magic
tech gf180mcuC
magscale 1 10
timestamp 1654786971
<< metal1 >>
rect 1120 18842 32816 18876
rect 1120 18790 4960 18842
rect 5012 18790 5064 18842
rect 5116 18790 5168 18842
rect 5220 18790 12900 18842
rect 12952 18790 13004 18842
rect 13056 18790 13108 18842
rect 13160 18790 20840 18842
rect 20892 18790 20944 18842
rect 20996 18790 21048 18842
rect 21100 18790 28780 18842
rect 28832 18790 28884 18842
rect 28936 18790 28988 18842
rect 29040 18790 32816 18842
rect 1120 18756 32816 18790
rect 1878 18618 1930 18630
rect 1878 18554 1930 18566
rect 6918 18618 6970 18630
rect 6918 18554 6970 18566
rect 16494 18618 16546 18630
rect 16494 18554 16546 18566
rect 21870 18618 21922 18630
rect 21870 18554 21922 18566
rect 23102 18618 23154 18630
rect 23102 18554 23154 18566
rect 25790 18618 25842 18630
rect 25790 18554 25842 18566
rect 3390 18506 3442 18518
rect 1530 18410 1542 18462
rect 1594 18410 1606 18462
rect 3390 18442 3442 18454
rect 6078 18506 6130 18518
rect 23998 18506 24050 18518
rect 6078 18442 6130 18454
rect 7142 18450 7194 18462
rect 2942 18394 2994 18406
rect 2942 18330 2994 18342
rect 3950 18394 4002 18406
rect 3950 18330 4002 18342
rect 4510 18394 4562 18406
rect 4510 18330 4562 18342
rect 6526 18394 6578 18406
rect 7142 18386 7194 18398
rect 9998 18450 10050 18462
rect 10154 18454 10166 18506
rect 10218 18454 10230 18506
rect 8698 18342 8710 18394
rect 8762 18342 8774 18394
rect 9998 18386 10050 18398
rect 11342 18450 11394 18462
rect 15822 18450 15874 18462
rect 15978 18454 15990 18506
rect 16042 18454 16054 18506
rect 6526 18330 6578 18342
rect 10154 18320 10166 18372
rect 10218 18320 10230 18372
rect 10602 18342 10614 18394
rect 10666 18342 10678 18394
rect 11162 18342 11174 18394
rect 11226 18342 11238 18394
rect 11342 18386 11394 18398
rect 11722 18380 11734 18432
rect 11786 18380 11798 18432
rect 13290 18398 13302 18450
rect 13354 18398 13366 18450
rect 14858 18342 14870 18394
rect 14922 18342 14934 18394
rect 15418 18380 15430 18432
rect 15482 18380 15494 18432
rect 17210 18410 17222 18462
rect 17274 18410 17286 18462
rect 17994 18454 18006 18506
rect 18058 18454 18070 18506
rect 15822 18386 15874 18398
rect 16606 18394 16658 18406
rect 15978 18320 15990 18372
rect 16042 18320 16054 18372
rect 16426 18342 16438 18394
rect 16490 18342 16502 18394
rect 18286 18394 18338 18406
rect 18622 18394 18674 18406
rect 19226 18398 19238 18450
rect 19290 18398 19302 18450
rect 21130 18410 21142 18462
rect 21194 18410 21206 18462
rect 22586 18410 22598 18462
rect 22650 18410 22662 18462
rect 23998 18442 24050 18454
rect 24558 18506 24610 18518
rect 28142 18506 28194 18518
rect 24558 18442 24610 18454
rect 27178 18410 27190 18462
rect 27242 18410 27254 18462
rect 28142 18442 28194 18454
rect 30718 18506 30770 18518
rect 30718 18442 30770 18454
rect 23774 18394 23826 18406
rect 16606 18330 16658 18342
rect 17994 18320 18006 18372
rect 18058 18320 18070 18372
rect 18442 18342 18454 18394
rect 18506 18342 18518 18394
rect 20570 18342 20582 18394
rect 20634 18342 20646 18394
rect 18286 18330 18338 18342
rect 18622 18330 18674 18342
rect 23774 18330 23826 18342
rect 25006 18394 25058 18406
rect 27626 18380 27638 18432
rect 27690 18380 27702 18432
rect 30494 18394 30546 18406
rect 25006 18330 25058 18342
rect 30494 18330 30546 18342
rect 32398 18394 32450 18406
rect 32398 18330 32450 18342
rect 2158 18282 2210 18294
rect 2158 18218 2210 18230
rect 2550 18282 2602 18294
rect 2550 18218 2602 18230
rect 2718 18282 2770 18294
rect 2718 18218 2770 18230
rect 3166 18282 3218 18294
rect 3166 18218 3218 18230
rect 4342 18282 4394 18294
rect 4342 18218 4394 18230
rect 6302 18282 6354 18294
rect 9326 18282 9378 18294
rect 7970 18230 7982 18282
rect 8034 18230 8046 18282
rect 6302 18218 6354 18230
rect 9326 18218 9378 18230
rect 9718 18282 9770 18294
rect 9718 18218 9770 18230
rect 10446 18282 10498 18294
rect 10446 18218 10498 18230
rect 10782 18282 10834 18294
rect 10782 18218 10834 18230
rect 11006 18282 11058 18294
rect 11006 18218 11058 18230
rect 12070 18282 12122 18294
rect 12070 18218 12122 18230
rect 12406 18282 12458 18294
rect 12406 18218 12458 18230
rect 12742 18282 12794 18294
rect 15094 18282 15146 18294
rect 14018 18230 14030 18282
rect 14082 18230 14094 18282
rect 12742 18218 12794 18230
rect 15094 18218 15146 18230
rect 17558 18282 17610 18294
rect 17558 18218 17610 18230
rect 17838 18282 17890 18294
rect 21478 18282 21530 18294
rect 19730 18230 19742 18282
rect 19794 18230 19806 18282
rect 17838 18218 17890 18230
rect 21478 18218 21530 18230
rect 21982 18282 22034 18294
rect 21982 18218 22034 18230
rect 22262 18282 22314 18294
rect 22262 18218 22314 18230
rect 22990 18282 23042 18294
rect 22990 18218 23042 18230
rect 23438 18282 23490 18294
rect 23438 18218 23490 18230
rect 23550 18282 23602 18294
rect 23550 18218 23602 18230
rect 25398 18282 25450 18294
rect 25398 18218 25450 18230
rect 25902 18282 25954 18294
rect 25902 18218 25954 18230
rect 26238 18282 26290 18294
rect 26238 18218 26290 18230
rect 26630 18282 26682 18294
rect 26630 18218 26682 18230
rect 26854 18282 26906 18294
rect 26854 18218 26906 18230
rect 27974 18282 28026 18294
rect 27974 18218 28026 18230
rect 29374 18282 29426 18294
rect 29374 18218 29426 18230
rect 29486 18282 29538 18294
rect 29486 18218 29538 18230
rect 30102 18282 30154 18294
rect 30102 18218 30154 18230
rect 31334 18282 31386 18294
rect 31334 18218 31386 18230
rect 31726 18282 31778 18294
rect 31726 18218 31778 18230
rect 32006 18282 32058 18294
rect 32006 18218 32058 18230
rect 1120 18058 32816 18092
rect 1120 18006 8930 18058
rect 8982 18006 9034 18058
rect 9086 18006 9138 18058
rect 9190 18006 16870 18058
rect 16922 18006 16974 18058
rect 17026 18006 17078 18058
rect 17130 18006 24810 18058
rect 24862 18006 24914 18058
rect 24966 18006 25018 18058
rect 25070 18006 32816 18058
rect 1120 17972 32816 18006
rect 1486 17834 1538 17846
rect 1486 17770 1538 17782
rect 5854 17834 5906 17846
rect 5854 17770 5906 17782
rect 10054 17834 10106 17846
rect 15430 17834 15482 17846
rect 11778 17782 11790 17834
rect 11842 17782 11854 17834
rect 10054 17770 10106 17782
rect 15430 17770 15482 17782
rect 16438 17834 16490 17846
rect 16438 17770 16490 17782
rect 17278 17834 17330 17846
rect 20582 17834 20634 17846
rect 32510 17834 32562 17846
rect 19506 17782 19518 17834
rect 19570 17782 19582 17834
rect 23202 17782 23214 17834
rect 23266 17782 23278 17834
rect 26114 17782 26126 17834
rect 26178 17782 26190 17834
rect 17278 17770 17330 17782
rect 20582 17770 20634 17782
rect 32510 17770 32562 17782
rect 2046 17722 2098 17734
rect 2538 17692 2550 17744
rect 2602 17692 2614 17744
rect 15822 17722 15874 17734
rect 2046 17658 2098 17670
rect 2382 17666 2434 17678
rect 6794 17670 6806 17722
rect 6858 17670 6870 17722
rect 6974 17666 7026 17678
rect 2382 17602 2434 17614
rect 3726 17610 3778 17622
rect 2538 17558 2550 17610
rect 2602 17558 2614 17610
rect 3726 17546 3778 17558
rect 6414 17610 6466 17622
rect 6974 17602 7026 17614
rect 7254 17666 7306 17678
rect 9482 17633 9494 17685
rect 9546 17633 9558 17685
rect 10950 17666 11002 17678
rect 12618 17670 12630 17722
rect 12682 17670 12694 17722
rect 7254 17602 7306 17614
rect 8094 17610 8146 17622
rect 6414 17546 6466 17558
rect 8922 17558 8934 17610
rect 8986 17558 8998 17610
rect 9762 17558 9774 17610
rect 9826 17558 9838 17610
rect 10378 17602 10390 17654
rect 10442 17602 10454 17654
rect 10782 17610 10834 17622
rect 10950 17602 11002 17614
rect 12854 17666 12906 17678
rect 14410 17670 14422 17722
rect 14474 17670 14486 17722
rect 14970 17633 14982 17685
rect 15034 17633 15046 17685
rect 15822 17658 15874 17670
rect 16102 17722 16154 17734
rect 17838 17722 17890 17734
rect 17658 17670 17670 17722
rect 17722 17670 17734 17722
rect 16102 17658 16154 17670
rect 17838 17658 17890 17670
rect 18062 17722 18114 17734
rect 18398 17722 18450 17734
rect 18218 17670 18230 17722
rect 18282 17670 18294 17722
rect 22094 17722 22146 17734
rect 18062 17658 18114 17670
rect 18398 17658 18450 17670
rect 12854 17602 12906 17614
rect 13694 17610 13746 17622
rect 8094 17546 8146 17558
rect 10782 17546 10834 17558
rect 13694 17546 13746 17558
rect 16830 17610 16882 17622
rect 20010 17614 20022 17666
rect 20074 17614 20086 17666
rect 18778 17558 18790 17610
rect 18842 17558 18854 17610
rect 20906 17602 20918 17654
rect 20970 17602 20982 17654
rect 21354 17633 21366 17685
rect 21418 17633 21430 17685
rect 22094 17658 22146 17670
rect 22374 17666 22426 17678
rect 27190 17666 27242 17678
rect 28746 17670 28758 17722
rect 28810 17670 28822 17722
rect 26730 17614 26742 17666
rect 26794 17614 26806 17666
rect 29094 17666 29146 17678
rect 22374 17602 22426 17614
rect 24042 17558 24054 17610
rect 24106 17558 24118 17610
rect 16830 17546 16882 17558
rect 1878 17498 1930 17510
rect 1878 17434 1930 17446
rect 2942 17498 2994 17510
rect 2942 17434 2994 17446
rect 3054 17498 3106 17510
rect 3054 17434 3106 17446
rect 3390 17498 3442 17510
rect 3390 17434 3442 17446
rect 3502 17498 3554 17510
rect 3502 17434 3554 17446
rect 5966 17498 6018 17510
rect 5966 17434 6018 17446
rect 6302 17498 6354 17510
rect 6302 17434 6354 17446
rect 6862 17498 6914 17510
rect 14970 17485 14982 17537
rect 15034 17485 15046 17537
rect 17726 17498 17778 17510
rect 6862 17434 6914 17446
rect 17726 17434 17778 17446
rect 21422 17498 21474 17510
rect 21422 17434 21474 17446
rect 21982 17498 22034 17510
rect 21982 17434 22034 17446
rect 24446 17498 24498 17510
rect 24714 17508 24726 17560
rect 24778 17508 24790 17560
rect 25274 17558 25286 17610
rect 25338 17558 25350 17610
rect 27190 17602 27242 17614
rect 28030 17610 28082 17622
rect 29094 17602 29146 17614
rect 29934 17610 29986 17622
rect 31322 17614 31334 17666
rect 31386 17614 31398 17666
rect 32062 17610 32114 17622
rect 28030 17546 28082 17558
rect 30762 17558 30774 17610
rect 30826 17558 30838 17610
rect 29934 17546 29986 17558
rect 32062 17546 32114 17558
rect 24446 17434 24498 17446
rect 30998 17498 31050 17510
rect 30998 17434 31050 17446
rect 1120 17274 32816 17308
rect 1120 17222 4960 17274
rect 5012 17222 5064 17274
rect 5116 17222 5168 17274
rect 5220 17222 12900 17274
rect 12952 17222 13004 17274
rect 13056 17222 13108 17274
rect 13160 17222 20840 17274
rect 20892 17222 20944 17274
rect 20996 17222 21048 17274
rect 21100 17222 28780 17274
rect 28832 17222 28884 17274
rect 28936 17222 28988 17274
rect 29040 17222 32816 17274
rect 1120 17188 32816 17222
rect 1878 17050 1930 17062
rect 1878 16986 1930 16998
rect 6022 17050 6074 17062
rect 12282 16998 12294 17050
rect 12346 16998 12358 17050
rect 15978 16998 15990 17050
rect 16042 16998 16054 17050
rect 6022 16986 6074 16998
rect 31322 16959 31334 17011
rect 31386 16959 31398 17011
rect 7534 16938 7586 16950
rect 1530 16842 1542 16894
rect 1594 16842 1606 16894
rect 2650 16830 2662 16882
rect 2714 16830 2726 16882
rect 6346 16842 6358 16894
rect 6410 16842 6422 16894
rect 6694 16882 6746 16894
rect 4286 16826 4338 16838
rect 3882 16774 3894 16826
rect 3946 16774 3958 16826
rect 8362 16886 8374 16938
rect 8426 16886 8438 16938
rect 7534 16874 7586 16886
rect 8598 16882 8650 16894
rect 10154 16886 10166 16938
rect 10218 16886 10230 16938
rect 6694 16818 6746 16830
rect 10714 16842 10726 16894
rect 10778 16842 10790 16894
rect 11610 16842 11622 16894
rect 11674 16842 11686 16894
rect 13302 16882 13354 16894
rect 14970 16886 14982 16938
rect 15034 16886 15046 16938
rect 8598 16818 8650 16830
rect 17210 16842 17222 16894
rect 17274 16842 17286 16894
rect 17838 16882 17890 16894
rect 17994 16886 18006 16938
rect 18058 16886 18070 16938
rect 18554 16886 18566 16938
rect 18618 16886 18630 16938
rect 24938 16886 24950 16938
rect 25002 16886 25014 16938
rect 26854 16882 26906 16894
rect 28410 16886 28422 16938
rect 28474 16886 28486 16938
rect 30874 16886 30886 16938
rect 30938 16886 30950 16938
rect 11946 16774 11958 16826
rect 12010 16774 12022 16826
rect 13302 16818 13354 16830
rect 20010 16830 20022 16882
rect 20074 16830 20086 16882
rect 15530 16774 15542 16826
rect 15594 16774 15606 16826
rect 17838 16818 17890 16830
rect 4286 16762 4338 16774
rect 17994 16752 18006 16804
rect 18058 16752 18070 16804
rect 20458 16774 20470 16826
rect 20522 16774 20534 16826
rect 22250 16812 22262 16864
rect 22314 16812 22326 16864
rect 23370 16830 23382 16882
rect 23434 16830 23446 16882
rect 26282 16830 26294 16882
rect 26346 16830 26358 16882
rect 29530 16830 29542 16882
rect 29594 16830 29606 16882
rect 24602 16774 24614 16826
rect 24666 16774 24678 16826
rect 26854 16818 26906 16830
rect 31210 16811 31222 16863
rect 31274 16811 31286 16863
rect 2046 16714 2098 16726
rect 4678 16714 4730 16726
rect 11062 16714 11114 16726
rect 3154 16662 3166 16714
rect 3218 16662 3230 16714
rect 9426 16662 9438 16714
rect 9490 16662 9502 16714
rect 2046 16650 2098 16662
rect 4678 16650 4730 16662
rect 11062 16650 11114 16662
rect 11286 16714 11338 16726
rect 12910 16714 12962 16726
rect 15262 16714 15314 16726
rect 11286 16650 11338 16662
rect 12350 16658 12402 16670
rect 12350 16594 12402 16606
rect 12574 16658 12626 16670
rect 14130 16662 14142 16714
rect 14194 16662 14206 16714
rect 16438 16714 16490 16726
rect 12910 16650 12962 16662
rect 15262 16650 15314 16662
rect 15934 16658 15986 16670
rect 12574 16594 12626 16606
rect 15934 16594 15986 16606
rect 16158 16658 16210 16670
rect 16438 16650 16490 16662
rect 16774 16714 16826 16726
rect 16774 16650 16826 16662
rect 17558 16714 17610 16726
rect 20302 16714 20354 16726
rect 19282 16662 19294 16714
rect 19346 16662 19358 16714
rect 17558 16650 17610 16662
rect 20302 16650 20354 16662
rect 20638 16714 20690 16726
rect 20638 16650 20690 16662
rect 21310 16714 21362 16726
rect 21310 16650 21362 16662
rect 21422 16714 21474 16726
rect 21422 16650 21474 16662
rect 21758 16714 21810 16726
rect 21758 16650 21810 16662
rect 21870 16714 21922 16726
rect 21870 16650 21922 16662
rect 22598 16714 22650 16726
rect 23874 16662 23886 16714
rect 23938 16662 23950 16714
rect 25778 16662 25790 16714
rect 25842 16662 25854 16714
rect 27682 16662 27694 16714
rect 27746 16662 27758 16714
rect 30034 16662 30046 16714
rect 30098 16662 30110 16714
rect 22598 16650 22650 16662
rect 16158 16594 16210 16606
rect 1120 16490 32816 16524
rect 1120 16438 8930 16490
rect 8982 16438 9034 16490
rect 9086 16438 9138 16490
rect 9190 16438 16870 16490
rect 16922 16438 16974 16490
rect 17026 16438 17078 16490
rect 17130 16438 24810 16490
rect 24862 16438 24914 16490
rect 24966 16438 25018 16490
rect 25070 16438 32816 16490
rect 1120 16404 32816 16438
rect 6638 16266 6690 16278
rect 3714 16214 3726 16266
rect 3778 16214 3790 16266
rect 6638 16202 6690 16214
rect 9830 16266 9882 16278
rect 9830 16202 9882 16214
rect 10110 16266 10162 16278
rect 10110 16202 10162 16214
rect 10222 16266 10274 16278
rect 10222 16202 10274 16214
rect 10558 16266 10610 16278
rect 10558 16202 10610 16214
rect 11006 16266 11058 16278
rect 15710 16266 15762 16278
rect 12114 16214 12126 16266
rect 12178 16214 12190 16266
rect 14858 16214 14870 16266
rect 14922 16214 14934 16266
rect 11006 16202 11058 16214
rect 15710 16202 15762 16214
rect 15822 16266 15874 16278
rect 15822 16202 15874 16214
rect 18734 16266 18786 16278
rect 18734 16202 18786 16214
rect 19294 16266 19346 16278
rect 21646 16266 21698 16278
rect 20402 16214 20414 16266
rect 20466 16214 20478 16266
rect 19294 16202 19346 16214
rect 21646 16202 21698 16214
rect 22654 16266 22706 16278
rect 22654 16202 22706 16214
rect 24110 16266 24162 16278
rect 24110 16202 24162 16214
rect 24502 16266 24554 16278
rect 24502 16202 24554 16214
rect 25230 16266 25282 16278
rect 25230 16202 25282 16214
rect 25566 16266 25618 16278
rect 25566 16202 25618 16214
rect 26126 16266 26178 16278
rect 28478 16266 28530 16278
rect 27234 16214 27246 16266
rect 27298 16214 27310 16266
rect 26126 16202 26178 16214
rect 28478 16202 28530 16214
rect 31502 16266 31554 16278
rect 31502 16202 31554 16214
rect 8878 16154 8930 16166
rect 1530 16034 1542 16086
rect 1594 16034 1606 16086
rect 2538 16065 2550 16117
rect 2602 16065 2614 16117
rect 4554 16102 4566 16154
rect 4618 16102 4630 16154
rect 2986 16046 2998 16098
rect 3050 16046 3062 16098
rect 4890 16065 4902 16117
rect 4954 16065 4966 16117
rect 7030 16098 7082 16110
rect 6750 16042 6802 16054
rect 11162 16124 11174 16176
rect 11226 16124 11238 16176
rect 11554 16102 11566 16154
rect 11618 16102 11630 16154
rect 11778 16102 11790 16154
rect 11842 16102 11854 16154
rect 14634 16102 14646 16154
rect 14698 16102 14710 16154
rect 8878 16090 8930 16102
rect 15598 16098 15650 16110
rect 16202 16102 16214 16154
rect 16266 16102 16278 16154
rect 16762 16124 16774 16176
rect 16826 16124 16838 16176
rect 17614 16154 17666 16166
rect 19070 16154 19122 16166
rect 7030 16034 7082 16046
rect 7870 16042 7922 16054
rect 6750 15978 6802 15990
rect 8698 15990 8710 16042
rect 8762 15990 8774 16042
rect 9482 16034 9494 16086
rect 9546 16034 9558 16086
rect 10670 16042 10722 16054
rect 13290 16046 13302 16098
rect 13354 16046 13366 16098
rect 13514 16046 13526 16098
rect 13578 16046 13590 16098
rect 11162 15990 11174 16042
rect 11226 15990 11238 16042
rect 15598 16034 15650 16046
rect 16606 16098 16658 16110
rect 16606 16034 16658 16046
rect 17390 16098 17442 16110
rect 17994 16102 18006 16154
rect 18058 16102 18070 16154
rect 17614 16090 17666 16102
rect 18342 16098 18394 16110
rect 16762 15990 16774 16042
rect 16826 15990 16838 16042
rect 17390 16034 17442 16046
rect 18342 16034 18394 16046
rect 18622 16098 18674 16110
rect 18622 16034 18674 16046
rect 18846 16098 18898 16110
rect 19070 16090 19122 16102
rect 21534 16154 21586 16166
rect 22250 16124 22262 16176
rect 22314 16124 22326 16176
rect 22810 16124 22822 16176
rect 22874 16124 22886 16176
rect 23370 16124 23382 16176
rect 23434 16124 23446 16176
rect 23774 16154 23826 16166
rect 28366 16154 28418 16166
rect 19898 16046 19910 16098
rect 19962 16046 19974 16098
rect 21534 16090 21586 16102
rect 22094 16098 22146 16110
rect 18846 16034 18898 16046
rect 21130 15990 21142 16042
rect 21194 15990 21206 16042
rect 21690 15990 21702 16042
rect 21754 15990 21766 16042
rect 22094 16034 22146 16046
rect 23214 16098 23266 16110
rect 25386 16102 25398 16154
rect 25450 16102 25462 16154
rect 25946 16102 25958 16154
rect 26010 16102 26022 16154
rect 26506 16102 26518 16154
rect 26570 16102 26582 16154
rect 23774 16090 23826 16102
rect 28086 16098 28138 16110
rect 22250 15990 22262 16042
rect 22314 15990 22326 16042
rect 22810 15990 22822 16042
rect 22874 15990 22886 16042
rect 23214 16034 23266 16046
rect 24782 16042 24834 16054
rect 23370 15990 23382 16042
rect 23434 15990 23446 16042
rect 28366 16090 28418 16102
rect 28870 16098 28922 16110
rect 28086 16034 28138 16046
rect 31098 16064 31110 16116
rect 31162 16064 31174 16116
rect 28870 16034 28922 16046
rect 29710 16042 29762 16054
rect 7870 15978 7922 15990
rect 10670 15978 10722 15990
rect 24782 15978 24834 15990
rect 30538 15990 30550 16042
rect 30602 15990 30614 16042
rect 29710 15978 29762 15990
rect 1878 15930 1930 15942
rect 1878 15866 1930 15878
rect 2494 15930 2546 15942
rect 2494 15866 2546 15878
rect 4958 15930 5010 15942
rect 26014 15930 26066 15942
rect 17546 15878 17558 15930
rect 17610 15878 17622 15930
rect 4958 15866 5010 15878
rect 26014 15866 26066 15878
rect 30774 15930 30826 15942
rect 30774 15866 30826 15878
rect 31614 15930 31666 15942
rect 31614 15866 31666 15878
rect 1120 15706 32816 15740
rect 1120 15654 4960 15706
rect 5012 15654 5064 15706
rect 5116 15654 5168 15706
rect 5220 15654 12900 15706
rect 12952 15654 13004 15706
rect 13056 15654 13108 15706
rect 13160 15654 20840 15706
rect 20892 15654 20944 15706
rect 20996 15654 21048 15706
rect 21100 15654 28780 15706
rect 28832 15654 28884 15706
rect 28936 15654 28988 15706
rect 29040 15654 32816 15706
rect 1120 15620 32816 15654
rect 18734 15538 18786 15550
rect 2270 15482 2322 15494
rect 2270 15418 2322 15430
rect 2382 15482 2434 15494
rect 2382 15418 2434 15430
rect 6470 15482 6522 15494
rect 6470 15418 6522 15430
rect 10670 15482 10722 15494
rect 10670 15418 10722 15430
rect 12506 15386 12518 15438
rect 12570 15386 12582 15438
rect 13738 15430 13750 15482
rect 13802 15430 13814 15482
rect 14366 15426 14418 15438
rect 14970 15430 14982 15482
rect 15034 15430 15046 15482
rect 16762 15430 16774 15482
rect 16826 15430 16838 15482
rect 17322 15430 17334 15482
rect 17386 15430 17398 15482
rect 18734 15474 18786 15486
rect 18958 15538 19010 15550
rect 18958 15474 19010 15486
rect 23942 15482 23994 15494
rect 5518 15370 5570 15382
rect 2874 15318 2886 15370
rect 2938 15318 2950 15370
rect 3222 15314 3274 15326
rect 4778 15318 4790 15370
rect 4842 15318 4854 15370
rect 5518 15306 5570 15318
rect 6694 15314 6746 15326
rect 3222 15250 3274 15262
rect 4062 15258 4114 15270
rect 2874 15184 2886 15236
rect 2938 15184 2950 15236
rect 6122 15244 6134 15296
rect 6186 15244 6198 15296
rect 8598 15314 8650 15326
rect 10266 15318 10278 15370
rect 10330 15318 10342 15370
rect 14366 15362 14418 15374
rect 14590 15370 14642 15382
rect 15754 15374 15766 15426
rect 15818 15374 15830 15426
rect 19786 15386 19798 15438
rect 19850 15386 19862 15438
rect 20526 15370 20578 15382
rect 6694 15250 6746 15262
rect 7534 15258 7586 15270
rect 4062 15194 4114 15206
rect 8250 15206 8262 15258
rect 8314 15206 8326 15258
rect 8598 15250 8650 15262
rect 10602 15243 10614 15295
rect 10666 15243 10678 15295
rect 12058 15250 12070 15302
rect 12122 15250 12134 15302
rect 12618 15274 12630 15326
rect 12682 15274 12694 15326
rect 14590 15306 14642 15318
rect 16158 15314 16210 15326
rect 13806 15258 13858 15270
rect 13402 15206 13414 15258
rect 13466 15206 13478 15258
rect 15194 15248 15206 15300
rect 15258 15248 15270 15300
rect 16158 15250 16210 15262
rect 16270 15314 16322 15326
rect 16270 15250 16322 15262
rect 17950 15314 18002 15326
rect 18106 15318 18118 15370
rect 18170 15318 18182 15370
rect 7534 15194 7586 15206
rect 13806 15194 13858 15206
rect 16718 15202 16770 15214
rect 16986 15206 16998 15258
rect 17050 15206 17062 15258
rect 17950 15250 18002 15262
rect 18554 15248 18566 15300
rect 18618 15248 18630 15300
rect 19674 15274 19686 15326
rect 19738 15274 19750 15326
rect 20078 15314 20130 15326
rect 20526 15306 20578 15318
rect 21198 15370 21250 15382
rect 22250 15374 22262 15426
rect 22314 15374 22326 15426
rect 23146 15384 23158 15436
rect 23210 15384 23222 15436
rect 23942 15418 23994 15430
rect 25722 15384 25734 15436
rect 25786 15384 25798 15436
rect 31322 15391 31334 15443
rect 31386 15391 31398 15443
rect 21198 15306 21250 15318
rect 22766 15370 22818 15382
rect 22766 15306 22818 15318
rect 24558 15370 24610 15382
rect 24558 15306 24610 15318
rect 25118 15370 25170 15382
rect 25566 15370 25618 15382
rect 30046 15370 30098 15382
rect 25118 15306 25170 15318
rect 25342 15314 25394 15326
rect 20078 15250 20130 15262
rect 21690 15248 21702 15300
rect 21754 15248 21766 15300
rect 1486 15146 1538 15158
rect 1486 15082 1538 15094
rect 1878 15146 1930 15158
rect 1878 15082 1930 15094
rect 2718 15146 2770 15158
rect 2718 15082 2770 15094
rect 5406 15146 5458 15158
rect 11398 15146 11450 15158
rect 9426 15094 9438 15146
rect 9490 15094 9502 15146
rect 5406 15082 5458 15094
rect 11398 15082 11450 15094
rect 11734 15146 11786 15158
rect 12462 15146 12514 15158
rect 11734 15082 11786 15094
rect 12238 15090 12290 15102
rect 15486 15146 15538 15158
rect 12462 15082 12514 15094
rect 14030 15090 14082 15102
rect 12238 15026 12290 15038
rect 15486 15082 15538 15094
rect 15710 15146 15762 15158
rect 15710 15082 15762 15094
rect 16494 15146 16546 15158
rect 18106 15184 18118 15236
rect 18170 15184 18182 15236
rect 22530 15206 22542 15258
rect 22594 15206 22606 15258
rect 23034 15242 23046 15294
rect 23098 15242 23110 15294
rect 23214 15258 23266 15270
rect 23214 15194 23266 15206
rect 24894 15258 24946 15270
rect 25566 15306 25618 15318
rect 26686 15314 26738 15326
rect 28746 15318 28758 15370
rect 28810 15318 28822 15370
rect 29206 15314 29258 15326
rect 25342 15250 25394 15262
rect 26014 15258 26066 15270
rect 27402 15262 27414 15314
rect 27466 15262 27478 15314
rect 24894 15194 24946 15206
rect 26506 15206 26518 15258
rect 26570 15206 26582 15258
rect 26686 15250 26738 15262
rect 27918 15258 27970 15270
rect 30874 15318 30886 15370
rect 30938 15318 30950 15370
rect 30046 15306 30098 15318
rect 29206 15250 29258 15262
rect 31210 15243 31222 15295
rect 31274 15243 31286 15295
rect 32330 15244 32342 15296
rect 32394 15244 32406 15296
rect 26014 15194 26066 15206
rect 27918 15194 27970 15206
rect 16718 15138 16770 15150
rect 17614 15146 17666 15158
rect 19854 15146 19906 15158
rect 21534 15146 21586 15158
rect 16494 15082 16546 15094
rect 17390 15090 17442 15102
rect 14030 15026 14082 15038
rect 19002 15094 19014 15146
rect 19066 15094 19078 15146
rect 20290 15094 20302 15146
rect 20354 15094 20366 15146
rect 23438 15146 23490 15158
rect 17614 15082 17666 15094
rect 19854 15082 19906 15094
rect 21534 15082 21586 15094
rect 21982 15090 22034 15102
rect 17390 15026 17442 15038
rect 21982 15026 22034 15038
rect 22206 15090 22258 15102
rect 23438 15082 23490 15094
rect 24334 15146 24386 15158
rect 26350 15146 26402 15158
rect 24334 15082 24386 15094
rect 25790 15090 25842 15102
rect 22206 15026 22258 15038
rect 26350 15082 26402 15094
rect 31838 15146 31890 15158
rect 31838 15082 31890 15094
rect 32006 15146 32058 15158
rect 32006 15082 32058 15094
rect 25790 15026 25842 15038
rect 1120 14922 32816 14956
rect 1120 14870 8930 14922
rect 8982 14870 9034 14922
rect 9086 14870 9138 14922
rect 9190 14870 16870 14922
rect 16922 14870 16974 14922
rect 17026 14870 17078 14922
rect 17130 14870 24810 14922
rect 24862 14870 24914 14922
rect 24966 14870 25018 14922
rect 25070 14870 32816 14922
rect 1120 14836 32816 14870
rect 12170 14728 12182 14780
rect 12234 14728 12246 14780
rect 19070 14754 19122 14766
rect 4678 14698 4730 14710
rect 4678 14634 4730 14646
rect 6862 14698 6914 14710
rect 13190 14698 13242 14710
rect 22206 14754 22258 14766
rect 8082 14646 8094 14698
rect 8146 14646 8158 14698
rect 6862 14634 6914 14646
rect 13190 14634 13242 14646
rect 14634 14612 14646 14664
rect 14698 14612 14710 14664
rect 16538 14646 16550 14698
rect 16602 14646 16614 14698
rect 19070 14690 19122 14702
rect 19294 14698 19346 14710
rect 20458 14646 20470 14698
rect 20522 14646 20534 14698
rect 21634 14646 21646 14698
rect 21698 14646 21710 14698
rect 22206 14690 22258 14702
rect 23886 14698 23938 14710
rect 19294 14634 19346 14646
rect 23886 14634 23938 14646
rect 26126 14698 26178 14710
rect 26126 14634 26178 14646
rect 26574 14698 26626 14710
rect 26574 14634 26626 14646
rect 27582 14698 27634 14710
rect 27582 14634 27634 14646
rect 27806 14698 27858 14710
rect 27806 14634 27858 14646
rect 27918 14698 27970 14710
rect 27918 14634 27970 14646
rect 28254 14698 28306 14710
rect 28254 14634 28306 14646
rect 28366 14698 28418 14710
rect 28366 14634 28418 14646
rect 31054 14698 31106 14710
rect 31054 14634 31106 14646
rect 31838 14698 31890 14710
rect 31838 14634 31890 14646
rect 1486 14586 1538 14598
rect 1486 14522 1538 14534
rect 2102 14530 2154 14542
rect 3770 14534 3782 14586
rect 3834 14534 3846 14586
rect 7254 14530 7306 14542
rect 8810 14534 8822 14586
rect 8874 14534 8886 14586
rect 2102 14466 2154 14478
rect 2942 14474 2994 14486
rect 4106 14472 4118 14524
rect 4170 14472 4182 14524
rect 5002 14466 5014 14518
rect 5066 14466 5078 14518
rect 6974 14474 7026 14486
rect 2942 14410 2994 14422
rect 9706 14496 9718 14548
rect 9770 14496 9782 14548
rect 10266 14534 10278 14586
rect 10330 14534 10342 14586
rect 10938 14556 10950 14608
rect 11002 14556 11014 14608
rect 11498 14556 11510 14608
rect 11562 14556 11574 14608
rect 14030 14586 14082 14598
rect 22430 14586 22482 14598
rect 26350 14586 26402 14598
rect 10446 14530 10498 14542
rect 7254 14466 7306 14478
rect 10446 14466 10498 14478
rect 10782 14530 10834 14542
rect 10782 14466 10834 14478
rect 11342 14530 11394 14542
rect 11834 14490 11846 14542
rect 11898 14490 11910 14542
rect 10938 14422 10950 14474
rect 11002 14422 11014 14474
rect 11342 14466 11394 14478
rect 12170 14466 12182 14518
rect 12234 14466 12246 14518
rect 12394 14490 12406 14542
rect 12458 14490 12470 14542
rect 12842 14534 12854 14586
rect 12906 14534 12918 14586
rect 13806 14530 13858 14542
rect 13626 14466 13638 14518
rect 13690 14466 13702 14518
rect 14030 14522 14082 14534
rect 14310 14530 14362 14542
rect 19742 14530 19794 14542
rect 19954 14534 19966 14586
rect 20018 14534 20030 14586
rect 21074 14534 21086 14586
rect 21138 14534 21150 14586
rect 21298 14534 21310 14586
rect 21362 14534 21374 14586
rect 13806 14466 13858 14478
rect 14746 14478 14758 14530
rect 14810 14478 14822 14530
rect 15530 14478 15542 14530
rect 15594 14478 15606 14530
rect 16090 14478 16102 14530
rect 16154 14478 16166 14530
rect 16314 14478 16326 14530
rect 16378 14478 16390 14530
rect 14310 14466 14362 14478
rect 17390 14474 17442 14486
rect 17658 14478 17670 14530
rect 17722 14478 17734 14530
rect 6974 14410 7026 14422
rect 17390 14410 17442 14422
rect 18622 14474 18674 14486
rect 18890 14466 18902 14518
rect 18954 14466 18966 14518
rect 22430 14522 22482 14534
rect 22654 14530 22706 14542
rect 23662 14530 23714 14542
rect 19742 14466 19794 14478
rect 20458 14466 20470 14518
rect 20522 14466 20534 14518
rect 22026 14458 22038 14510
rect 22090 14458 22102 14510
rect 22922 14478 22934 14530
rect 22986 14478 22998 14530
rect 24042 14484 24054 14536
rect 24106 14484 24118 14536
rect 25342 14530 25394 14542
rect 24378 14478 24390 14530
rect 24442 14478 24454 14530
rect 22654 14466 22706 14478
rect 23662 14466 23714 14478
rect 25342 14466 25394 14478
rect 25566 14530 25618 14542
rect 25946 14534 25958 14586
rect 26010 14534 26022 14586
rect 26730 14534 26742 14586
rect 26794 14534 26806 14586
rect 27402 14556 27414 14608
rect 27466 14556 27478 14608
rect 31726 14586 31778 14598
rect 26350 14522 26402 14534
rect 26910 14530 26962 14542
rect 25566 14466 25618 14478
rect 26910 14466 26962 14478
rect 27246 14530 27298 14542
rect 29306 14478 29318 14530
rect 29370 14478 29382 14530
rect 31726 14522 31778 14534
rect 27246 14466 27298 14478
rect 29934 14474 29986 14486
rect 1878 14362 1930 14374
rect 4218 14349 4230 14401
rect 4282 14349 4294 14401
rect 9382 14362 9434 14374
rect 1878 14298 1930 14310
rect 9382 14298 9434 14310
rect 10334 14362 10386 14374
rect 10334 14298 10386 14310
rect 11454 14362 11506 14374
rect 14074 14354 14086 14406
rect 14138 14354 14150 14406
rect 17882 14360 17894 14412
rect 17946 14360 17958 14412
rect 18622 14410 18674 14422
rect 18062 14362 18114 14374
rect 11454 14298 11506 14310
rect 18062 14298 18114 14310
rect 18398 14362 18450 14374
rect 19002 14356 19014 14408
rect 19066 14356 19078 14408
rect 23034 14372 23046 14424
rect 23098 14372 23110 14424
rect 30762 14422 30774 14474
rect 30826 14422 30838 14474
rect 29934 14410 29986 14422
rect 23326 14362 23378 14374
rect 18398 14298 18450 14310
rect 20234 14274 20246 14326
rect 20298 14274 20310 14326
rect 22586 14310 22598 14362
rect 22650 14310 22662 14362
rect 23930 14356 23942 14408
rect 23994 14356 24006 14408
rect 28702 14362 28754 14374
rect 25610 14310 25622 14362
rect 25674 14310 25686 14362
rect 23326 14298 23378 14310
rect 28702 14298 28754 14310
rect 28814 14362 28866 14374
rect 28814 14298 28866 14310
rect 31446 14362 31498 14374
rect 31446 14298 31498 14310
rect 1120 14138 32816 14172
rect 1120 14086 4960 14138
rect 5012 14086 5064 14138
rect 5116 14086 5168 14138
rect 5220 14086 12900 14138
rect 12952 14086 13004 14138
rect 13056 14086 13108 14138
rect 13160 14086 20840 14138
rect 20892 14086 20944 14138
rect 20996 14086 21048 14138
rect 21100 14086 28780 14138
rect 28832 14086 28884 14138
rect 28936 14086 28988 14138
rect 29040 14086 32816 14138
rect 1120 14052 32816 14086
rect 23214 13970 23266 13982
rect 5518 13914 5570 13926
rect 5518 13850 5570 13862
rect 6694 13914 6746 13926
rect 9494 13914 9546 13926
rect 11286 13914 11338 13926
rect 8138 13862 8150 13914
rect 8202 13862 8214 13914
rect 9818 13862 9830 13914
rect 9882 13862 9894 13914
rect 6694 13850 6746 13862
rect 9494 13850 9546 13862
rect 11286 13850 11338 13862
rect 15306 13816 15318 13868
rect 15370 13816 15382 13868
rect 22642 13862 22654 13914
rect 22706 13862 22718 13914
rect 23214 13906 23266 13918
rect 24558 13970 24610 13982
rect 24558 13906 24610 13918
rect 24782 13970 24834 13982
rect 24782 13906 24834 13918
rect 27526 13914 27578 13926
rect 22990 13858 23042 13870
rect 3502 13802 3554 13814
rect 12686 13802 12738 13814
rect 19574 13802 19626 13814
rect 20682 13806 20694 13858
rect 20746 13806 20758 13858
rect 22094 13802 22146 13814
rect 2158 13746 2210 13758
rect 2314 13750 2326 13802
rect 2378 13750 2390 13802
rect 4218 13750 4230 13802
rect 4282 13750 4294 13802
rect 2986 13694 2998 13746
rect 3050 13694 3062 13746
rect 3502 13738 3554 13750
rect 6346 13706 6358 13758
rect 6410 13706 6422 13758
rect 6906 13706 6918 13758
rect 6970 13706 6982 13758
rect 2158 13682 2210 13694
rect 5854 13690 5906 13702
rect 2314 13616 2326 13668
rect 2378 13616 2390 13668
rect 7242 13682 7254 13734
rect 7306 13682 7318 13734
rect 7466 13706 7478 13758
rect 7530 13706 7542 13758
rect 8430 13746 8482 13758
rect 8206 13690 8258 13702
rect 7802 13638 7814 13690
rect 7866 13638 7878 13690
rect 9930 13694 9942 13746
rect 9994 13694 10006 13746
rect 10154 13694 10166 13746
rect 10218 13694 10230 13746
rect 12394 13706 12406 13758
rect 12458 13706 12470 13758
rect 13626 13750 13638 13802
rect 13690 13750 13702 13802
rect 18330 13750 18342 13802
rect 18394 13750 18406 13802
rect 12686 13738 12738 13750
rect 8430 13682 8482 13694
rect 11790 13690 11842 13702
rect 5854 13626 5906 13638
rect 8206 13626 8258 13638
rect 11790 13626 11842 13638
rect 12238 13690 12290 13702
rect 14074 13694 14086 13746
rect 14138 13694 14150 13746
rect 14758 13690 14810 13702
rect 12238 13626 12290 13638
rect 13626 13616 13638 13668
rect 13690 13616 13702 13668
rect 1486 13578 1538 13590
rect 1486 13514 1538 13526
rect 1878 13578 1930 13590
rect 1878 13514 1930 13526
rect 4622 13578 4674 13590
rect 4622 13514 4674 13526
rect 4734 13578 4786 13590
rect 4734 13514 4786 13526
rect 5406 13578 5458 13590
rect 5406 13514 5458 13526
rect 5966 13578 6018 13590
rect 5966 13514 6018 13526
rect 9102 13578 9154 13590
rect 7130 13470 7142 13522
rect 7194 13470 7206 13522
rect 9102 13514 9154 13526
rect 10950 13578 11002 13590
rect 10950 13514 11002 13526
rect 11454 13578 11506 13590
rect 12126 13578 12178 13590
rect 11454 13514 11506 13526
rect 12014 13522 12066 13534
rect 12126 13514 12178 13526
rect 13470 13578 13522 13590
rect 14186 13582 14198 13634
rect 14250 13582 14262 13634
rect 14758 13626 14810 13638
rect 15262 13690 15314 13702
rect 15418 13688 15430 13740
rect 15482 13688 15494 13740
rect 15754 13694 15766 13746
rect 15818 13694 15830 13746
rect 16426 13694 16438 13746
rect 16490 13694 16502 13746
rect 17658 13694 17670 13746
rect 17722 13694 17734 13746
rect 18778 13706 18790 13758
rect 18842 13706 18854 13758
rect 19574 13738 19626 13750
rect 21310 13746 21362 13758
rect 21466 13750 21478 13802
rect 21530 13750 21542 13802
rect 27526 13850 27578 13862
rect 27806 13914 27858 13926
rect 27806 13850 27858 13862
rect 31110 13914 31162 13926
rect 31110 13850 31162 13862
rect 22990 13794 23042 13806
rect 30046 13802 30098 13814
rect 18958 13690 19010 13702
rect 17322 13638 17334 13690
rect 17386 13638 17398 13690
rect 15262 13626 15314 13638
rect 13470 13514 13522 13526
rect 15038 13578 15090 13590
rect 17770 13582 17782 13634
rect 17834 13582 17846 13634
rect 18330 13616 18342 13668
rect 18394 13616 18406 13668
rect 18958 13626 19010 13638
rect 19294 13690 19346 13702
rect 19294 13626 19346 13638
rect 20302 13690 20354 13702
rect 20302 13626 20354 13638
rect 20526 13690 20578 13702
rect 22094 13738 22146 13750
rect 23886 13746 23938 13758
rect 24042 13750 24054 13802
rect 24106 13750 24118 13802
rect 21310 13682 21362 13694
rect 21914 13682 21926 13734
rect 21978 13682 21990 13734
rect 22262 13690 22314 13702
rect 20526 13626 20578 13638
rect 23886 13682 23938 13694
rect 25062 13749 25114 13761
rect 25498 13750 25510 13802
rect 25562 13750 25574 13802
rect 26058 13706 26070 13758
rect 26122 13706 26134 13758
rect 26394 13706 26406 13758
rect 26458 13706 26470 13758
rect 29206 13746 29258 13758
rect 25062 13685 25114 13697
rect 26618 13682 26630 13734
rect 26682 13682 26694 13734
rect 30046 13738 30098 13750
rect 29206 13682 29258 13694
rect 22262 13626 22314 13638
rect 24042 13616 24054 13668
rect 24106 13616 24118 13668
rect 25498 13616 25510 13668
rect 25562 13616 25574 13668
rect 30762 13638 30774 13690
rect 30826 13638 30838 13690
rect 31434 13676 31446 13728
rect 31498 13676 31510 13728
rect 18174 13578 18226 13590
rect 17098 13526 17110 13578
rect 17162 13526 17174 13578
rect 15038 13514 15090 13526
rect 18174 13514 18226 13526
rect 19966 13578 20018 13590
rect 19114 13470 19126 13522
rect 19178 13470 19190 13522
rect 19966 13514 20018 13526
rect 20750 13578 20802 13590
rect 20750 13514 20802 13526
rect 21422 13578 21474 13590
rect 21422 13514 21474 13526
rect 23606 13578 23658 13590
rect 25342 13578 25394 13590
rect 24490 13526 24502 13578
rect 24554 13526 24566 13578
rect 23606 13514 23658 13526
rect 25342 13514 25394 13526
rect 25790 13578 25842 13590
rect 25790 13514 25842 13526
rect 27134 13578 27186 13590
rect 27134 13514 27186 13526
rect 27918 13578 27970 13590
rect 27918 13514 27970 13526
rect 28254 13578 28306 13590
rect 28254 13514 28306 13526
rect 28366 13578 28418 13590
rect 28366 13514 28418 13526
rect 12014 13458 12066 13470
rect 26394 13444 26406 13496
rect 26458 13444 26470 13496
rect 1120 13354 32816 13388
rect 1120 13302 8930 13354
rect 8982 13302 9034 13354
rect 9086 13302 9138 13354
rect 9190 13302 16870 13354
rect 16922 13302 16974 13354
rect 17026 13302 17078 13354
rect 17130 13302 24810 13354
rect 24862 13302 24914 13354
rect 24966 13302 25018 13354
rect 25070 13302 32816 13354
rect 1120 13268 32816 13302
rect 8654 13186 8706 13198
rect 1598 13130 1650 13142
rect 6638 13130 6690 13142
rect 3490 13078 3502 13130
rect 3554 13078 3566 13130
rect 1598 13066 1650 13078
rect 6638 13066 6690 13078
rect 6862 13130 6914 13142
rect 7578 13078 7590 13130
rect 7642 13078 7654 13130
rect 8654 13122 8706 13134
rect 8878 13130 8930 13142
rect 14746 13134 14758 13186
rect 14810 13134 14822 13186
rect 20470 13130 20522 13142
rect 6862 13066 6914 13078
rect 8878 13066 8930 13078
rect 16606 13074 16658 13086
rect 2438 13018 2490 13030
rect 2438 12954 2490 12966
rect 2662 12962 2714 12974
rect 4554 12966 4566 13018
rect 4618 12966 4630 13018
rect 7018 12988 7030 13040
rect 7082 12988 7094 13040
rect 7926 13018 7978 13030
rect 12058 13022 12070 13074
rect 12122 13022 12134 13074
rect 16158 13018 16210 13030
rect 1710 12906 1762 12918
rect 2090 12898 2102 12950
rect 2154 12898 2166 12950
rect 6246 12962 6298 12974
rect 2662 12898 2714 12910
rect 5406 12906 5458 12918
rect 4218 12854 4230 12906
rect 4282 12854 4294 12906
rect 8250 12966 8262 13018
rect 8314 12966 8326 13018
rect 10434 12966 10446 13018
rect 10498 12966 10510 13018
rect 7926 12954 7978 12966
rect 6246 12898 6298 12910
rect 9662 12906 9714 12918
rect 7018 12854 7030 12906
rect 7082 12854 7094 12906
rect 1710 12842 1762 12854
rect 5406 12842 5458 12854
rect 9662 12842 9714 12854
rect 10110 12906 10162 12918
rect 10938 12910 10950 12962
rect 11002 12910 11014 12962
rect 11386 12910 11398 12962
rect 11450 12910 11462 12962
rect 11946 12910 11958 12962
rect 12010 12910 12022 12962
rect 13290 12918 13302 12970
rect 13354 12918 13366 12970
rect 15990 12962 16042 12974
rect 10110 12842 10162 12854
rect 12630 12906 12682 12918
rect 13962 12898 13974 12950
rect 14026 12898 14038 12950
rect 14634 12910 14646 12962
rect 14698 12910 14710 12962
rect 14970 12909 14982 12961
rect 15034 12909 15046 12961
rect 20470 13066 20522 13078
rect 21030 13130 21082 13142
rect 21030 13066 21082 13078
rect 21646 13130 21698 13142
rect 22586 13134 22598 13186
rect 22650 13134 22662 13186
rect 24166 13130 24218 13142
rect 23818 13078 23830 13130
rect 23882 13078 23894 13130
rect 21646 13066 21698 13078
rect 24166 13066 24218 13078
rect 16606 13010 16658 13022
rect 18286 13018 18338 13030
rect 16158 12954 16210 12966
rect 16382 12962 16434 12974
rect 15990 12898 16042 12910
rect 17434 12928 17446 12980
rect 17498 12928 17510 12980
rect 18286 12954 18338 12966
rect 18510 13018 18562 13030
rect 21758 13018 21810 13030
rect 30494 13018 30546 13030
rect 19170 12966 19182 13018
rect 19234 12966 19246 13018
rect 19730 12966 19742 13018
rect 19794 12966 19806 13018
rect 20122 12966 20134 13018
rect 20186 12966 20198 13018
rect 18510 12954 18562 12966
rect 16382 12898 16434 12910
rect 17782 12906 17834 12918
rect 12630 12842 12682 12854
rect 17994 12898 18006 12950
rect 18058 12898 18070 12950
rect 20694 12906 20746 12918
rect 21354 12910 21366 12962
rect 21418 12910 21430 12962
rect 21758 12954 21810 12966
rect 22250 12922 22262 12974
rect 22314 12922 22326 12974
rect 13022 12794 13074 12806
rect 8586 12742 8598 12794
rect 8650 12742 8662 12794
rect 9874 12742 9886 12794
rect 9938 12742 9950 12794
rect 11498 12742 11510 12794
rect 11562 12742 11574 12794
rect 13022 12730 13074 12742
rect 13358 12794 13410 12806
rect 13358 12730 13410 12742
rect 13638 12794 13690 12806
rect 14522 12798 14534 12850
rect 14586 12798 14598 12850
rect 17782 12842 17834 12854
rect 22474 12898 22486 12950
rect 22538 12898 22550 12950
rect 22810 12922 22822 12974
rect 22874 12922 22886 12974
rect 23270 12962 23322 12974
rect 28534 12962 28586 12974
rect 30202 12966 30214 13018
rect 30266 12966 30278 13018
rect 22990 12906 23042 12918
rect 18330 12798 18342 12850
rect 18394 12798 18406 12850
rect 20694 12842 20746 12854
rect 23270 12898 23322 12910
rect 24490 12898 24502 12950
rect 24554 12898 24566 12950
rect 24782 12906 24834 12918
rect 25610 12910 25622 12962
rect 25674 12910 25686 12962
rect 22990 12842 23042 12854
rect 24782 12842 24834 12854
rect 26126 12906 26178 12918
rect 27178 12910 27190 12962
rect 27242 12910 27254 12962
rect 28030 12906 28082 12918
rect 26842 12854 26854 12906
rect 26906 12854 26918 12906
rect 26126 12842 26178 12854
rect 19406 12794 19458 12806
rect 27290 12804 27302 12856
rect 27354 12804 27366 12856
rect 30494 12954 30546 12966
rect 28534 12898 28586 12910
rect 29374 12906 29426 12918
rect 28030 12842 28082 12854
rect 29374 12842 29426 12854
rect 16090 12742 16102 12794
rect 16154 12742 16166 12794
rect 27582 12794 27634 12806
rect 13638 12730 13690 12742
rect 19406 12730 19458 12742
rect 23550 12738 23602 12750
rect 23550 12674 23602 12686
rect 23774 12738 23826 12750
rect 27582 12730 27634 12742
rect 27918 12794 27970 12806
rect 30762 12781 30774 12833
rect 30826 12781 30838 12833
rect 27918 12730 27970 12742
rect 23774 12674 23826 12686
rect 1120 12570 32816 12604
rect 1120 12518 4960 12570
rect 5012 12518 5064 12570
rect 5116 12518 5168 12570
rect 5220 12518 12900 12570
rect 12952 12518 13004 12570
rect 13056 12518 13108 12570
rect 13160 12518 20840 12570
rect 20892 12518 20944 12570
rect 20996 12518 21048 12570
rect 21100 12518 28780 12570
rect 28832 12518 28884 12570
rect 28936 12518 28988 12570
rect 29040 12518 32816 12570
rect 1120 12484 32816 12518
rect 7198 12346 7250 12358
rect 7198 12282 7250 12294
rect 17334 12346 17386 12358
rect 1598 12234 1650 12246
rect 3166 12234 3218 12246
rect 2314 12182 2326 12234
rect 2378 12182 2390 12234
rect 4230 12234 4282 12246
rect 1598 12170 1650 12182
rect 3166 12170 3218 12182
rect 4006 12178 4058 12190
rect 4230 12170 4282 12182
rect 5854 12234 5906 12246
rect 11162 12238 11174 12290
rect 11226 12238 11238 12290
rect 17334 12282 17386 12294
rect 20358 12346 20410 12358
rect 5854 12170 5906 12182
rect 12518 12234 12570 12246
rect 18218 12238 18230 12290
rect 18282 12238 18294 12290
rect 20358 12282 20410 12294
rect 22206 12346 22258 12358
rect 22206 12282 22258 12294
rect 22318 12346 22370 12358
rect 22318 12282 22370 12294
rect 23606 12346 23658 12358
rect 23606 12282 23658 12294
rect 24558 12346 24610 12358
rect 24558 12282 24610 12294
rect 26854 12346 26906 12358
rect 26854 12282 26906 12294
rect 32006 12346 32058 12358
rect 32006 12282 32058 12294
rect 20750 12234 20802 12246
rect 13402 12182 13414 12234
rect 13466 12182 13478 12234
rect 4006 12114 4058 12126
rect 4554 12108 4566 12160
rect 4618 12108 4630 12160
rect 6246 12122 6298 12134
rect 8810 12108 8822 12160
rect 8874 12108 8886 12160
rect 9482 12126 9494 12178
rect 9546 12126 9558 12178
rect 11610 12126 11622 12178
rect 11674 12126 11686 12178
rect 12518 12170 12570 12182
rect 17054 12178 17106 12190
rect 12170 12108 12182 12160
rect 12234 12108 12246 12160
rect 13738 12126 13750 12178
rect 13802 12126 13814 12178
rect 14366 12122 14418 12134
rect 6246 12058 6298 12070
rect 6458 12024 6470 12076
rect 6522 12024 6534 12076
rect 15082 12114 15094 12166
rect 15146 12114 15158 12166
rect 15306 12114 15318 12166
rect 15370 12114 15382 12166
rect 15642 12114 15654 12166
rect 15706 12114 15718 12166
rect 15866 12114 15878 12166
rect 15930 12114 15942 12166
rect 16202 12114 16214 12166
rect 16266 12114 16278 12166
rect 16426 12114 16438 12166
rect 16490 12114 16502 12166
rect 16718 12122 16770 12134
rect 1374 12010 1426 12022
rect 1374 11946 1426 11958
rect 2158 12010 2210 12022
rect 2158 11946 2210 11958
rect 5518 12010 5570 12022
rect 5518 11946 5570 11958
rect 7086 12010 7138 12022
rect 7086 11946 7138 11958
rect 9158 12010 9210 12022
rect 11722 12014 11734 12066
rect 11786 12014 11798 12066
rect 14366 12058 14418 12070
rect 16874 12070 16886 12122
rect 16938 12070 16950 12122
rect 17054 12114 17106 12126
rect 17950 12178 18002 12190
rect 27470 12234 27522 12246
rect 17950 12114 18002 12126
rect 18510 12122 18562 12134
rect 19002 12126 19014 12178
rect 19066 12126 19078 12178
rect 19338 12126 19350 12178
rect 19402 12126 19414 12178
rect 20750 12170 20802 12182
rect 23034 12138 23046 12190
rect 23098 12138 23110 12190
rect 20638 12122 20690 12134
rect 20010 12070 20022 12122
rect 20074 12070 20086 12122
rect 16718 12058 16770 12070
rect 18510 12058 18562 12070
rect 20638 12058 20690 12070
rect 22766 12122 22818 12134
rect 23370 12114 23382 12166
rect 23434 12114 23446 12166
rect 25050 12126 25062 12178
rect 25114 12126 25126 12178
rect 27470 12170 27522 12182
rect 29206 12178 29258 12190
rect 30762 12182 30774 12234
rect 30826 12182 30838 12234
rect 23930 12070 23942 12122
rect 23994 12070 24006 12122
rect 24490 12070 24502 12122
rect 24554 12070 24566 12122
rect 26618 12070 26630 12122
rect 26682 12070 26694 12122
rect 27178 12108 27190 12160
rect 27242 12108 27254 12160
rect 28310 12122 28362 12134
rect 28634 12108 28646 12160
rect 28698 12108 28710 12160
rect 29206 12114 29258 12126
rect 30046 12122 30098 12134
rect 22766 12058 22818 12070
rect 28310 12058 28362 12070
rect 32330 12108 32342 12160
rect 32394 12108 32406 12160
rect 30046 12058 30098 12070
rect 9158 11946 9210 11958
rect 12798 12010 12850 12022
rect 12798 11946 12850 11958
rect 17670 12010 17722 12022
rect 19014 12010 19066 12022
rect 15418 11876 15430 11928
rect 15482 11876 15494 11928
rect 16090 11902 16102 11954
rect 16154 11902 16166 11954
rect 17670 11946 17722 11958
rect 18286 11954 18338 11966
rect 19014 11946 19066 11958
rect 21534 12010 21586 12022
rect 21534 11946 21586 11958
rect 21926 12010 21978 12022
rect 21926 11946 21978 11958
rect 24670 12010 24722 12022
rect 31838 12010 31890 12022
rect 25778 11958 25790 12010
rect 25842 11958 25854 12010
rect 24670 11946 24722 11958
rect 31838 11946 31890 11958
rect 18286 11890 18338 11902
rect 23146 11876 23158 11928
rect 23210 11876 23222 11928
rect 1120 11786 32816 11820
rect 1120 11734 8930 11786
rect 8982 11734 9034 11786
rect 9086 11734 9138 11786
rect 9190 11734 16870 11786
rect 16922 11734 16974 11786
rect 17026 11734 17078 11786
rect 17130 11734 24810 11786
rect 24862 11734 24914 11786
rect 24966 11734 25018 11786
rect 25070 11734 32816 11786
rect 1120 11700 32816 11734
rect 2214 11562 2266 11574
rect 3266 11510 3278 11562
rect 3330 11510 3342 11562
rect 6234 11535 6246 11587
rect 6298 11535 6310 11587
rect 9326 11562 9378 11574
rect 8138 11510 8150 11562
rect 8202 11510 8214 11562
rect 2214 11498 2266 11510
rect 9326 11498 9378 11510
rect 9662 11562 9714 11574
rect 9662 11498 9714 11510
rect 10110 11562 10162 11574
rect 10110 11498 10162 11510
rect 10558 11562 10610 11574
rect 10558 11498 10610 11510
rect 10950 11562 11002 11574
rect 10950 11498 11002 11510
rect 12686 11562 12738 11574
rect 17390 11562 17442 11574
rect 16426 11510 16438 11562
rect 16490 11510 16502 11562
rect 12686 11498 12738 11510
rect 17390 11498 17442 11510
rect 17502 11562 17554 11574
rect 17502 11498 17554 11510
rect 18006 11562 18058 11574
rect 19674 11535 19686 11587
rect 19738 11535 19750 11587
rect 18006 11498 18058 11510
rect 9886 11450 9938 11462
rect 1866 11360 1878 11412
rect 1930 11360 1942 11412
rect 1598 11338 1650 11350
rect 2650 11342 2662 11394
rect 2714 11342 2726 11394
rect 4442 11361 4454 11413
rect 4506 11361 4518 11413
rect 5786 11342 5798 11394
rect 5850 11342 5862 11394
rect 6794 11342 6806 11394
rect 6858 11342 6870 11394
rect 7130 11348 7142 11400
rect 7194 11348 7206 11400
rect 11386 11420 11398 11472
rect 11450 11420 11462 11472
rect 8250 11342 8262 11394
rect 8314 11342 8326 11394
rect 9886 11386 9938 11398
rect 11230 11394 11282 11406
rect 11834 11398 11846 11450
rect 11898 11398 11910 11450
rect 13402 11444 13414 11496
rect 13466 11444 13478 11496
rect 13750 11450 13802 11462
rect 4106 11286 4118 11338
rect 4170 11286 4182 11338
rect 6010 11286 6022 11338
rect 6074 11286 6086 11338
rect 8026 11286 8038 11338
rect 8090 11286 8102 11338
rect 11230 11330 11282 11342
rect 12014 11394 12066 11406
rect 12954 11342 12966 11394
rect 13018 11342 13030 11394
rect 13750 11386 13802 11398
rect 15038 11450 15090 11462
rect 24054 11450 24106 11462
rect 15418 11398 15430 11450
rect 15482 11398 15494 11450
rect 15038 11386 15090 11398
rect 15642 11342 15654 11394
rect 15706 11342 15718 11394
rect 17782 11391 17834 11403
rect 11386 11286 11398 11338
rect 11450 11286 11462 11338
rect 12014 11330 12066 11342
rect 17782 11327 17834 11339
rect 18062 11394 18114 11406
rect 19226 11342 19238 11394
rect 19290 11342 19302 11394
rect 18062 11330 18114 11342
rect 18778 11286 18790 11338
rect 18842 11286 18854 11338
rect 21130 11330 21142 11382
rect 21194 11330 21206 11382
rect 21746 11342 21758 11394
rect 21810 11342 21822 11394
rect 24054 11386 24106 11398
rect 25286 11450 25338 11462
rect 26842 11398 26854 11450
rect 26906 11398 26918 11450
rect 25286 11386 25338 11398
rect 27290 11361 27302 11413
rect 27354 11361 27366 11413
rect 24726 11338 24778 11350
rect 1598 11274 1650 11286
rect 4510 11226 4562 11238
rect 7466 11230 7478 11282
rect 7530 11230 7542 11282
rect 24726 11274 24778 11286
rect 26574 11282 26626 11294
rect 4510 11162 4562 11174
rect 10222 11226 10274 11238
rect 10222 11162 10274 11174
rect 11902 11226 11954 11238
rect 11902 11162 11954 11174
rect 12574 11226 12626 11238
rect 14478 11226 14530 11238
rect 12574 11162 12626 11174
rect 14142 11170 14194 11182
rect 14478 11162 14530 11174
rect 14926 11226 14978 11238
rect 27402 11236 27414 11288
rect 27466 11236 27478 11288
rect 26574 11218 26626 11230
rect 14926 11162 14978 11174
rect 18286 11170 18338 11182
rect 14142 11106 14194 11118
rect 18286 11106 18338 11118
rect 1120 11002 32816 11036
rect 1120 10950 4960 11002
rect 5012 10950 5064 11002
rect 5116 10950 5168 11002
rect 5220 10950 12900 11002
rect 12952 10950 13004 11002
rect 13056 10950 13108 11002
rect 13160 10950 20840 11002
rect 20892 10950 20944 11002
rect 20996 10950 21048 11002
rect 21100 10950 28780 11002
rect 28832 10950 28884 11002
rect 28936 10950 28988 11002
rect 29040 10950 32816 11002
rect 1120 10916 32816 10950
rect 9662 10834 9714 10846
rect 8934 10778 8986 10790
rect 8934 10714 8986 10726
rect 9438 10778 9490 10790
rect 16942 10834 16994 10846
rect 9662 10770 9714 10782
rect 10782 10778 10834 10790
rect 9438 10714 9490 10726
rect 2270 10666 2322 10678
rect 10154 10668 10166 10720
rect 10218 10668 10230 10720
rect 10782 10714 10834 10726
rect 12014 10778 12066 10790
rect 15754 10726 15766 10778
rect 15818 10726 15830 10778
rect 16942 10770 16994 10782
rect 23998 10778 24050 10790
rect 12014 10714 12066 10726
rect 12842 10670 12854 10722
rect 12906 10670 12918 10722
rect 13738 10670 13750 10722
rect 13802 10670 13814 10722
rect 14298 10670 14310 10722
rect 14362 10670 14374 10722
rect 23998 10714 24050 10726
rect 24558 10778 24610 10790
rect 24558 10714 24610 10726
rect 25342 10778 25394 10790
rect 25342 10714 25394 10726
rect 20750 10666 20802 10678
rect 1430 10610 1482 10622
rect 4218 10614 4230 10666
rect 4282 10614 4294 10666
rect 2270 10602 2322 10614
rect 1430 10546 1482 10558
rect 2986 10502 2998 10554
rect 3050 10502 3062 10554
rect 3546 10535 3558 10587
rect 3610 10535 3622 10587
rect 5450 10546 5462 10598
rect 5514 10546 5526 10598
rect 5898 10546 5910 10598
rect 5962 10546 5974 10598
rect 9930 10570 9942 10622
rect 9994 10570 10006 10622
rect 10334 10610 10386 10622
rect 11386 10614 11398 10666
rect 11450 10614 11462 10666
rect 19786 10614 19798 10666
rect 19850 10614 19862 10666
rect 21870 10666 21922 10678
rect 8262 10554 8314 10566
rect 10334 10546 10386 10558
rect 12282 10544 12294 10596
rect 12346 10544 12358 10596
rect 12574 10554 12626 10566
rect 8262 10490 8314 10502
rect 11386 10480 11398 10532
rect 11450 10480 11462 10532
rect 11902 10498 11954 10510
rect 4846 10442 4898 10454
rect 4846 10378 4898 10390
rect 9102 10442 9154 10454
rect 10894 10442 10946 10454
rect 9102 10378 9154 10390
rect 10110 10386 10162 10398
rect 10894 10378 10946 10390
rect 11230 10442 11282 10454
rect 12574 10490 12626 10502
rect 13358 10554 13410 10566
rect 13570 10558 13582 10610
rect 13634 10558 13646 10610
rect 13358 10490 13410 10502
rect 13806 10554 13858 10566
rect 14410 10558 14422 10610
rect 14474 10558 14486 10610
rect 13806 10490 13858 10502
rect 15710 10554 15762 10566
rect 17334 10554 17386 10566
rect 16090 10502 16102 10554
rect 16154 10502 16166 10554
rect 15710 10490 15762 10502
rect 17334 10490 17386 10502
rect 18230 10554 18282 10566
rect 19002 10540 19014 10592
rect 19066 10540 19078 10592
rect 20010 10558 20022 10610
rect 20074 10558 20086 10610
rect 20750 10602 20802 10614
rect 21354 10570 21366 10622
rect 21418 10570 21430 10622
rect 21870 10602 21922 10614
rect 24110 10554 24162 10566
rect 11902 10434 11954 10446
rect 12798 10442 12850 10454
rect 11230 10378 11282 10390
rect 16606 10442 16658 10454
rect 17490 10446 17502 10498
rect 17554 10446 17566 10498
rect 18230 10490 18282 10502
rect 24110 10490 24162 10502
rect 24894 10554 24946 10566
rect 24894 10490 24946 10502
rect 25454 10554 25506 10566
rect 25454 10490 25506 10502
rect 25846 10554 25898 10566
rect 25846 10490 25898 10502
rect 27302 10554 27354 10566
rect 28074 10540 28086 10592
rect 28138 10540 28150 10592
rect 27302 10490 27354 10502
rect 12798 10378 12850 10390
rect 14758 10386 14810 10398
rect 10110 10322 10162 10334
rect 14758 10322 14810 10334
rect 15486 10386 15538 10398
rect 16606 10378 16658 10390
rect 18622 10442 18674 10454
rect 18622 10378 18674 10390
rect 19350 10442 19402 10454
rect 19350 10378 19402 10390
rect 21702 10442 21754 10454
rect 21702 10378 21754 10390
rect 23550 10442 23602 10454
rect 23550 10378 23602 10390
rect 24446 10442 24498 10454
rect 24446 10378 24498 10390
rect 25006 10442 25058 10454
rect 27750 10442 27802 10454
rect 25006 10378 25058 10390
rect 27134 10386 27186 10398
rect 15486 10322 15538 10334
rect 27750 10378 27802 10390
rect 27134 10322 27186 10334
rect 1120 10218 32816 10252
rect 1120 10166 8930 10218
rect 8982 10166 9034 10218
rect 9086 10166 9138 10218
rect 9190 10166 16870 10218
rect 16922 10166 16974 10218
rect 17026 10166 17078 10218
rect 17130 10166 24810 10218
rect 24862 10166 24914 10218
rect 24966 10166 25018 10218
rect 25070 10166 32816 10218
rect 1120 10132 32816 10166
rect 6458 10024 6470 10076
rect 6522 10024 6534 10076
rect 9662 10050 9714 10062
rect 4062 9994 4114 10006
rect 3042 9942 3054 9994
rect 3106 9942 3118 9994
rect 4062 9930 4114 9942
rect 4902 9994 4954 10006
rect 8710 9994 8762 10006
rect 4902 9930 4954 9942
rect 8094 9938 8146 9950
rect 5910 9882 5962 9894
rect 5562 9830 5574 9882
rect 5626 9830 5638 9882
rect 1530 9762 1542 9814
rect 1594 9762 1606 9814
rect 2538 9774 2550 9826
rect 2602 9774 2614 9826
rect 5910 9818 5962 9830
rect 6190 9882 6242 9894
rect 6190 9818 6242 9830
rect 6750 9882 6802 9894
rect 14926 10050 14978 10062
rect 9662 9986 9714 9998
rect 13526 9994 13578 10006
rect 12842 9942 12854 9994
rect 12906 9942 12918 9994
rect 14926 9986 14978 9998
rect 16046 9994 16098 10006
rect 8710 9930 8762 9942
rect 13526 9930 13578 9942
rect 15150 9938 15202 9950
rect 7186 9830 7198 9882
rect 7250 9830 7262 9882
rect 7410 9830 7422 9882
rect 7474 9830 7486 9882
rect 7746 9830 7758 9882
rect 7810 9830 7822 9882
rect 8094 9874 8146 9886
rect 9438 9882 9490 9894
rect 6750 9818 6802 9830
rect 8318 9826 8370 9838
rect 3882 9718 3894 9770
rect 3946 9718 3958 9770
rect 4554 9762 4566 9814
rect 4618 9762 4630 9814
rect 5070 9770 5122 9782
rect 6458 9762 6470 9814
rect 6522 9762 6534 9814
rect 10042 9830 10054 9882
rect 10106 9830 10118 9882
rect 11498 9830 11510 9882
rect 11562 9830 11574 9882
rect 12058 9852 12070 9904
rect 12122 9852 12134 9904
rect 12518 9882 12570 9894
rect 9438 9818 9490 9830
rect 11902 9826 11954 9838
rect 8318 9762 8370 9774
rect 14702 9882 14754 9894
rect 12518 9818 12570 9830
rect 13694 9826 13746 9838
rect 11902 9762 11954 9774
rect 14074 9803 14086 9855
rect 14138 9803 14150 9855
rect 16046 9930 16098 9942
rect 15150 9874 15202 9886
rect 20358 9882 20410 9894
rect 15418 9830 15430 9882
rect 15482 9830 15494 9882
rect 14702 9818 14754 9830
rect 15822 9826 15874 9838
rect 12058 9718 12070 9770
rect 12122 9718 12134 9770
rect 13694 9762 13746 9774
rect 14522 9754 14534 9806
rect 14586 9754 14598 9806
rect 16538 9792 16550 9844
rect 16602 9792 16614 9844
rect 24166 9882 24218 9894
rect 20358 9818 20410 9830
rect 15822 9762 15874 9774
rect 16886 9770 16938 9782
rect 17434 9762 17446 9814
rect 17498 9762 17510 9814
rect 17994 9762 18006 9814
rect 18058 9762 18070 9814
rect 21354 9786 21366 9838
rect 21418 9786 21430 9838
rect 21802 9786 21814 9838
rect 21866 9786 21878 9838
rect 24166 9818 24218 9830
rect 21030 9770 21082 9782
rect 5070 9706 5122 9718
rect 16886 9706 16938 9718
rect 21030 9706 21082 9718
rect 24838 9770 24890 9782
rect 24838 9706 24890 9718
rect 25230 9770 25282 9782
rect 25230 9706 25282 9718
rect 25454 9770 25506 9782
rect 25946 9774 25958 9826
rect 26010 9774 26022 9826
rect 25454 9706 25506 9718
rect 26574 9770 26626 9782
rect 27806 9770 27858 9782
rect 27290 9718 27302 9770
rect 27354 9718 27366 9770
rect 26574 9706 26626 9718
rect 27806 9706 27858 9718
rect 1878 9658 1930 9670
rect 11174 9658 11226 9670
rect 9594 9606 9606 9658
rect 9658 9606 9670 9658
rect 13918 9658 13970 9670
rect 27694 9658 27746 9670
rect 1878 9594 1930 9606
rect 11174 9594 11226 9606
rect 13470 9602 13522 9614
rect 14634 9606 14646 9658
rect 14698 9606 14710 9658
rect 15866 9606 15878 9658
rect 15930 9606 15942 9658
rect 13918 9594 13970 9606
rect 27694 9594 27746 9606
rect 13470 9538 13522 9550
rect 1120 9434 32816 9468
rect 1120 9382 4960 9434
rect 5012 9382 5064 9434
rect 5116 9382 5168 9434
rect 5220 9382 12900 9434
rect 12952 9382 13004 9434
rect 13056 9382 13108 9434
rect 13160 9382 20840 9434
rect 20892 9382 20944 9434
rect 20996 9382 21048 9434
rect 21100 9382 28780 9434
rect 28832 9382 28884 9434
rect 28936 9382 28988 9434
rect 29040 9382 32816 9434
rect 1120 9348 32816 9382
rect 13582 9266 13634 9278
rect 4118 9210 4170 9222
rect 10054 9210 10106 9222
rect 7578 9158 7590 9210
rect 7642 9158 7654 9210
rect 4118 9146 4170 9158
rect 10054 9146 10106 9158
rect 10278 9210 10330 9222
rect 10278 9146 10330 9158
rect 10502 9210 10554 9222
rect 11902 9210 11954 9222
rect 10502 9146 10554 9158
rect 1486 9098 1538 9110
rect 2718 9098 2770 9110
rect 3726 9098 3778 9110
rect 1486 9034 1538 9046
rect 1878 9042 1930 9054
rect 1598 8986 1650 8998
rect 3434 9046 3446 9098
rect 3498 9046 3510 9098
rect 2718 9034 2770 9046
rect 3726 9034 3778 9046
rect 4734 9098 4786 9110
rect 4734 9034 4786 9046
rect 6134 9098 6186 9110
rect 11722 9108 11734 9160
rect 11786 9108 11798 9160
rect 12618 9158 12630 9210
rect 12682 9158 12694 9210
rect 13582 9202 13634 9214
rect 19350 9210 19402 9222
rect 11902 9146 11954 9158
rect 19350 9146 19402 9158
rect 19630 9210 19682 9222
rect 19630 9146 19682 9158
rect 20358 9210 20410 9222
rect 20358 9146 20410 9158
rect 22262 9210 22314 9222
rect 13974 9098 14026 9110
rect 6134 9034 6186 9046
rect 8766 9042 8818 9054
rect 1878 8978 1930 8990
rect 4510 8986 4562 8998
rect 1598 8922 1650 8934
rect 5450 8967 5462 9019
rect 5514 8967 5526 9019
rect 7534 8986 7586 8998
rect 21578 9096 21590 9148
rect 21642 9096 21654 9148
rect 22262 9146 22314 9158
rect 23494 9210 23546 9222
rect 23494 9146 23546 9158
rect 32006 9210 32058 9222
rect 32006 9146 32058 9158
rect 26910 9098 26962 9110
rect 13974 9034 14026 9046
rect 4510 8922 4562 8934
rect 7914 8934 7926 8986
rect 7978 8934 7990 8986
rect 8138 8934 8150 8986
rect 8202 8934 8214 8986
rect 8766 8978 8818 8990
rect 11610 8982 11622 9034
rect 11674 8982 11686 9034
rect 14410 9002 14422 9054
rect 14474 9002 14486 9054
rect 14634 9002 14646 9054
rect 14698 9002 14710 9054
rect 14970 9002 14982 9054
rect 15034 9002 15046 9054
rect 12574 8986 12626 8998
rect 12170 8934 12182 8986
rect 12234 8934 12246 8986
rect 7534 8922 7586 8934
rect 12574 8922 12626 8934
rect 12798 8986 12850 8998
rect 12798 8922 12850 8934
rect 13358 8986 13410 8998
rect 15866 8978 15878 9030
rect 15930 8978 15942 9030
rect 16258 8990 16270 9042
rect 16322 8990 16334 9042
rect 19966 8986 20018 8998
rect 13358 8922 13410 8934
rect 20682 8972 20694 9024
rect 20746 8972 20758 9024
rect 21422 8986 21474 8998
rect 19966 8922 20018 8934
rect 21690 8982 21702 9034
rect 21754 8982 21766 9034
rect 23146 9002 23158 9054
rect 23210 9002 23222 9054
rect 26070 9042 26122 9054
rect 24166 8986 24218 8998
rect 27626 9046 27638 9098
rect 27690 9046 27702 9098
rect 26910 9034 26962 9046
rect 21422 8922 21474 8934
rect 25722 8934 25734 8986
rect 25786 8934 25798 8986
rect 26070 8978 26122 8990
rect 32330 8972 32342 9024
rect 32394 8972 32406 9024
rect 24166 8922 24218 8934
rect 8654 8874 8706 8886
rect 7310 8818 7362 8830
rect 7310 8754 7362 8766
rect 8542 8818 8594 8830
rect 8654 8810 8706 8822
rect 9102 8874 9154 8886
rect 9102 8810 9154 8822
rect 9214 8874 9266 8886
rect 10838 8874 10890 8886
rect 19742 8874 19794 8886
rect 9762 8822 9774 8874
rect 9826 8822 9838 8874
rect 18666 8822 18678 8874
rect 18730 8822 18742 8874
rect 9214 8810 9266 8822
rect 10838 8810 10890 8822
rect 14746 8766 14758 8818
rect 14810 8766 14822 8818
rect 19742 8810 19794 8822
rect 22654 8874 22706 8886
rect 31838 8874 31890 8886
rect 22654 8810 22706 8822
rect 25454 8818 25506 8830
rect 31838 8810 31890 8822
rect 8542 8754 8594 8766
rect 25454 8754 25506 8766
rect 1120 8650 32816 8684
rect 1120 8598 8930 8650
rect 8982 8598 9034 8650
rect 9086 8598 9138 8650
rect 9190 8598 16870 8650
rect 16922 8598 16974 8650
rect 17026 8598 17078 8650
rect 17130 8598 24810 8650
rect 24862 8598 24914 8650
rect 24966 8598 25018 8650
rect 25070 8598 32816 8650
rect 1120 8564 32816 8598
rect 8362 8456 8374 8508
rect 8426 8456 8438 8508
rect 1486 8426 1538 8438
rect 3210 8374 3222 8426
rect 3274 8374 3286 8426
rect 6346 8399 6358 8451
rect 6410 8399 6422 8451
rect 17278 8426 17330 8438
rect 1486 8362 1538 8374
rect 17278 8362 17330 8374
rect 18902 8426 18954 8438
rect 18902 8362 18954 8374
rect 20526 8426 20578 8438
rect 20526 8362 20578 8374
rect 20974 8426 21026 8438
rect 20974 8362 21026 8374
rect 24054 8426 24106 8438
rect 4734 8314 4786 8326
rect 3994 8262 4006 8314
rect 4058 8262 4070 8314
rect 2426 8206 2438 8258
rect 2490 8206 2502 8258
rect 3770 8206 3782 8258
rect 3834 8206 3846 8258
rect 4734 8250 4786 8262
rect 4958 8314 5010 8326
rect 4958 8250 5010 8262
rect 7422 8314 7474 8326
rect 12294 8314 12346 8326
rect 5898 8206 5910 8258
rect 5962 8206 5974 8258
rect 6638 8202 6690 8214
rect 7018 8206 7030 8258
rect 7082 8206 7094 8258
rect 7422 8250 7474 8262
rect 8138 8218 8150 8270
rect 8202 8218 8214 8270
rect 5450 8150 5462 8202
rect 5514 8150 5526 8202
rect 8474 8194 8486 8246
rect 8538 8194 8550 8246
rect 8698 8194 8710 8246
rect 8762 8194 8774 8246
rect 9370 8218 9382 8270
rect 9434 8218 9446 8270
rect 12294 8250 12346 8262
rect 16214 8314 16266 8326
rect 9930 8194 9942 8246
rect 9994 8194 10006 8246
rect 12966 8202 13018 8214
rect 1978 8094 1990 8146
rect 2042 8094 2054 8146
rect 6638 8138 6690 8150
rect 13290 8194 13302 8246
rect 13354 8194 13366 8246
rect 13794 8206 13806 8258
rect 13858 8206 13870 8258
rect 16214 8250 16266 8262
rect 17558 8314 17610 8326
rect 17558 8250 17610 8262
rect 17950 8314 18002 8326
rect 17950 8250 18002 8262
rect 18622 8314 18674 8326
rect 18622 8250 18674 8262
rect 19294 8314 19346 8326
rect 19294 8250 19346 8262
rect 19742 8314 19794 8326
rect 19742 8250 19794 8262
rect 19966 8314 20018 8326
rect 22026 8318 22038 8370
rect 22090 8318 22102 8370
rect 24054 8362 24106 8374
rect 19966 8250 20018 8262
rect 24334 8314 24386 8326
rect 16886 8202 16938 8214
rect 20794 8206 20806 8258
rect 20858 8206 20870 8258
rect 22362 8206 22374 8258
rect 22426 8206 22438 8258
rect 24334 8250 24386 8262
rect 25286 8314 25338 8326
rect 25286 8250 25338 8262
rect 26574 8314 26626 8326
rect 26574 8250 26626 8262
rect 26742 8314 26794 8326
rect 26742 8250 26794 8262
rect 12966 8138 13018 8150
rect 23706 8194 23718 8246
rect 23770 8194 23782 8246
rect 24602 8198 24614 8250
rect 24666 8198 24678 8250
rect 16886 8138 16938 8150
rect 4342 8090 4394 8102
rect 4342 8026 4394 8038
rect 7086 8090 7138 8102
rect 7086 8026 7138 8038
rect 18230 8090 18282 8102
rect 18230 8026 18282 8038
rect 19630 8090 19682 8102
rect 19630 8026 19682 8038
rect 20414 8090 20466 8102
rect 24490 8100 24502 8152
rect 24554 8100 24566 8152
rect 20414 8026 20466 8038
rect 1120 7866 32816 7900
rect 1120 7814 4960 7866
rect 5012 7814 5064 7866
rect 5116 7814 5168 7866
rect 5220 7814 12900 7866
rect 12952 7814 13004 7866
rect 13056 7814 13108 7866
rect 13160 7814 20840 7866
rect 20892 7814 20944 7866
rect 20996 7814 21048 7866
rect 21100 7814 28780 7866
rect 28832 7814 28884 7866
rect 28936 7814 28988 7866
rect 29040 7814 32816 7866
rect 1120 7780 32816 7814
rect 6862 7642 6914 7654
rect 3098 7590 3110 7642
rect 3162 7590 3174 7642
rect 6862 7578 6914 7590
rect 8934 7642 8986 7654
rect 8934 7578 8986 7590
rect 11622 7642 11674 7654
rect 11622 7578 11674 7590
rect 13750 7642 13802 7654
rect 13750 7578 13802 7590
rect 15430 7642 15482 7654
rect 15430 7578 15482 7590
rect 16102 7642 16154 7654
rect 16102 7578 16154 7590
rect 17446 7642 17498 7654
rect 6022 7530 6074 7542
rect 2986 7478 2998 7530
rect 3050 7478 3062 7530
rect 4062 7474 4114 7486
rect 2550 7418 2602 7430
rect 3770 7422 3782 7474
rect 3834 7422 3846 7474
rect 4062 7410 4114 7422
rect 4286 7474 4338 7486
rect 5674 7434 5686 7486
rect 5738 7434 5750 7486
rect 6022 7466 6074 7478
rect 4286 7410 4338 7422
rect 6346 7404 6358 7456
rect 6410 7404 6422 7456
rect 8586 7434 8598 7486
rect 8650 7434 8662 7486
rect 12506 7478 12518 7530
rect 12570 7478 12582 7530
rect 16874 7528 16886 7580
rect 16938 7528 16950 7580
rect 17446 7578 17498 7590
rect 18174 7642 18226 7654
rect 18174 7578 18226 7590
rect 18510 7642 18562 7654
rect 18510 7578 18562 7590
rect 19574 7642 19626 7654
rect 19574 7578 19626 7590
rect 20246 7642 20298 7654
rect 22766 7642 22818 7654
rect 20246 7578 20298 7590
rect 21914 7540 21926 7592
rect 21978 7540 21990 7592
rect 22766 7578 22818 7590
rect 25118 7586 25170 7598
rect 6794 7366 6806 7418
rect 6858 7366 6870 7418
rect 8026 7366 8038 7418
rect 8090 7366 8102 7418
rect 9482 7404 9494 7456
rect 9546 7404 9558 7456
rect 10490 7366 10502 7418
rect 10554 7366 10566 7418
rect 11050 7404 11062 7456
rect 11114 7404 11126 7456
rect 11946 7404 11958 7456
rect 12010 7404 12022 7456
rect 13402 7434 13414 7486
rect 13466 7434 13478 7486
rect 12798 7418 12850 7430
rect 2550 7354 2602 7366
rect 12506 7344 12518 7396
rect 12570 7344 12582 7396
rect 14410 7404 14422 7456
rect 14474 7404 14486 7456
rect 15082 7434 15094 7486
rect 15146 7434 15158 7486
rect 17770 7434 17782 7486
rect 17834 7434 17846 7486
rect 22418 7478 22430 7530
rect 22482 7478 22494 7530
rect 25118 7522 25170 7534
rect 25790 7586 25842 7598
rect 25790 7522 25842 7534
rect 26126 7530 26178 7542
rect 15710 7418 15762 7430
rect 12798 7354 12850 7366
rect 15710 7354 15762 7366
rect 17166 7418 17218 7430
rect 18106 7422 18118 7474
rect 18170 7422 18182 7474
rect 17166 7354 17218 7366
rect 18846 7418 18898 7430
rect 19226 7404 19238 7456
rect 19290 7404 19302 7456
rect 21690 7422 21702 7474
rect 21754 7422 21766 7474
rect 26126 7466 26178 7478
rect 22094 7418 22146 7430
rect 18846 7354 18898 7366
rect 23370 7404 23382 7456
rect 23434 7404 23446 7456
rect 23930 7366 23942 7418
rect 23994 7366 24006 7418
rect 25386 7366 25398 7418
rect 25450 7366 25462 7418
rect 22094 7354 22146 7366
rect 1486 7306 1538 7318
rect 1486 7242 1538 7254
rect 1598 7306 1650 7318
rect 4678 7306 4730 7318
rect 3210 7254 3222 7306
rect 3274 7254 3286 7306
rect 1598 7242 1650 7254
rect 4678 7242 4730 7254
rect 4958 7306 5010 7318
rect 4958 7242 5010 7254
rect 5350 7306 5402 7318
rect 5350 7242 5402 7254
rect 6974 7306 7026 7318
rect 6974 7242 7026 7254
rect 7422 7306 7474 7318
rect 7422 7242 7474 7254
rect 7646 7306 7698 7318
rect 7646 7242 7698 7254
rect 7870 7306 7922 7318
rect 7870 7242 7922 7254
rect 8206 7306 8258 7318
rect 8206 7242 8258 7254
rect 9158 7306 9210 7318
rect 9158 7242 9210 7254
rect 9774 7306 9826 7318
rect 9774 7242 9826 7254
rect 10334 7306 10386 7318
rect 10334 7242 10386 7254
rect 10670 7306 10722 7318
rect 10670 7242 10722 7254
rect 11398 7306 11450 7318
rect 11398 7242 11450 7254
rect 12350 7306 12402 7318
rect 12350 7242 12402 7254
rect 13918 7306 13970 7318
rect 13918 7242 13970 7254
rect 14758 7306 14810 7318
rect 14758 7242 14810 7254
rect 16942 7306 16994 7318
rect 16942 7242 16994 7254
rect 19854 7306 19906 7318
rect 19854 7242 19906 7254
rect 23046 7306 23098 7318
rect 23046 7242 23098 7254
rect 1120 7082 32816 7116
rect 1120 7030 8930 7082
rect 8982 7030 9034 7082
rect 9086 7030 9138 7082
rect 9190 7030 16870 7082
rect 16922 7030 16974 7082
rect 17026 7030 17078 7082
rect 17130 7030 24810 7082
rect 24862 7030 24914 7082
rect 24966 7030 25018 7082
rect 25070 7030 32816 7082
rect 1120 6996 32816 7030
rect 11902 6914 11954 6926
rect 2818 6806 2830 6858
rect 2882 6806 2894 6858
rect 7242 6831 7254 6883
rect 7306 6831 7318 6883
rect 12618 6862 12630 6914
rect 12682 6862 12694 6914
rect 11902 6850 11954 6862
rect 16830 6858 16882 6870
rect 15978 6806 15990 6858
rect 16042 6806 16054 6858
rect 4566 6746 4618 6758
rect 5450 6750 5462 6802
rect 5514 6750 5526 6802
rect 6234 6750 6246 6802
rect 6298 6750 6310 6802
rect 16830 6794 16882 6806
rect 19294 6858 19346 6870
rect 24334 6858 24386 6870
rect 23146 6806 23158 6858
rect 23210 6806 23222 6858
rect 19294 6794 19346 6806
rect 24334 6794 24386 6806
rect 6862 6746 6914 6758
rect 11678 6746 11730 6758
rect 6682 6694 6694 6746
rect 6746 6694 6758 6746
rect 11274 6694 11286 6746
rect 11338 6694 11350 6746
rect 24110 6746 24162 6758
rect 4566 6682 4618 6694
rect 1530 6626 1542 6678
rect 1594 6626 1606 6678
rect 1878 6634 1930 6646
rect 1878 6570 1930 6582
rect 2270 6634 2322 6646
rect 3434 6626 3446 6678
rect 3498 6626 3510 6678
rect 3726 6634 3778 6646
rect 5226 6638 5238 6690
rect 5290 6638 5302 6690
rect 6122 6638 6134 6690
rect 6186 6638 6198 6690
rect 6862 6682 6914 6694
rect 7690 6638 7702 6690
rect 7754 6638 7766 6690
rect 11678 6682 11730 6694
rect 2270 6570 2322 6582
rect 8138 6582 8150 6634
rect 8202 6582 8214 6634
rect 8810 6626 8822 6678
rect 8874 6626 8886 6678
rect 9930 6626 9942 6678
rect 9994 6626 10006 6678
rect 10334 6634 10386 6646
rect 10938 6630 10950 6682
rect 11002 6630 11014 6682
rect 12282 6626 12294 6678
rect 12346 6626 12358 6678
rect 12506 6626 12518 6678
rect 12570 6626 12582 6678
rect 12842 6626 12854 6678
rect 12906 6626 12918 6678
rect 13066 6650 13078 6702
rect 13130 6650 13142 6702
rect 13626 6626 13638 6678
rect 13690 6626 13702 6678
rect 17882 6656 17894 6708
rect 17946 6656 17958 6708
rect 18666 6656 18678 6708
rect 18730 6656 18742 6708
rect 20234 6650 20246 6702
rect 20298 6650 20310 6702
rect 18230 6634 18282 6646
rect 3726 6570 3778 6582
rect 2494 6522 2546 6534
rect 2494 6458 2546 6470
rect 3110 6522 3162 6534
rect 5674 6526 5686 6578
rect 5738 6526 5750 6578
rect 10334 6570 10386 6582
rect 3110 6458 3162 6470
rect 6750 6522 6802 6534
rect 6750 6458 6802 6470
rect 8486 6522 8538 6534
rect 8486 6458 8538 6470
rect 9606 6522 9658 6534
rect 9606 6458 9658 6470
rect 10670 6522 10722 6534
rect 10826 6532 10838 6584
rect 10890 6532 10902 6584
rect 18230 6570 18282 6582
rect 19686 6634 19738 6646
rect 20850 6638 20862 6690
rect 20914 6638 20926 6690
rect 24110 6682 24162 6694
rect 24558 6690 24610 6702
rect 24558 6626 24610 6638
rect 24714 6618 24726 6670
rect 24778 6618 24790 6670
rect 25274 6638 25286 6690
rect 25338 6638 25350 6690
rect 26282 6630 26294 6682
rect 26346 6630 26358 6682
rect 26954 6626 26966 6678
rect 27018 6626 27030 6678
rect 19686 6570 19738 6582
rect 16662 6522 16714 6534
rect 11610 6470 11622 6522
rect 11674 6470 11686 6522
rect 10670 6458 10722 6470
rect 16662 6458 16714 6470
rect 19014 6522 19066 6534
rect 19014 6458 19066 6470
rect 23830 6522 23882 6534
rect 25386 6532 25398 6584
rect 25450 6532 25462 6584
rect 25678 6522 25730 6534
rect 24042 6470 24054 6522
rect 24106 6470 24118 6522
rect 23830 6458 23882 6470
rect 25678 6458 25730 6470
rect 26014 6522 26066 6534
rect 26170 6532 26182 6584
rect 26234 6532 26246 6584
rect 26014 6458 26066 6470
rect 26630 6522 26682 6534
rect 26630 6458 26682 6470
rect 1120 6298 32816 6332
rect 1120 6246 4960 6298
rect 5012 6246 5064 6298
rect 5116 6246 5168 6298
rect 5220 6246 12900 6298
rect 12952 6246 13004 6298
rect 13056 6246 13108 6298
rect 13160 6246 20840 6298
rect 20892 6246 20944 6298
rect 20996 6246 21048 6298
rect 21100 6246 28780 6298
rect 28832 6246 28884 6298
rect 28936 6246 28988 6298
rect 29040 6246 32816 6298
rect 1120 6212 32816 6246
rect 4734 6074 4786 6086
rect 12070 6074 12122 6086
rect 2314 6022 2326 6074
rect 2378 6022 2390 6074
rect 5842 6022 5854 6074
rect 5906 6022 5918 6074
rect 6402 6022 6414 6074
rect 6466 6022 6478 6074
rect 4734 6010 4786 6022
rect 12070 6010 12122 6022
rect 12854 6074 12906 6086
rect 18566 6074 18618 6086
rect 14298 6022 14310 6074
rect 14362 6022 14374 6074
rect 12854 6010 12906 6022
rect 18566 6010 18618 6022
rect 21254 6074 21306 6086
rect 21254 6010 21306 6022
rect 22038 6074 22090 6086
rect 22038 6010 22090 6022
rect 3726 5962 3778 5974
rect 2762 5866 2774 5918
rect 2826 5866 2838 5918
rect 3726 5898 3778 5910
rect 3950 5962 4002 5974
rect 7422 5962 7474 5974
rect 3950 5898 4002 5910
rect 7198 5906 7250 5918
rect 1990 5850 2042 5862
rect 3098 5842 3110 5894
rect 3162 5842 3174 5894
rect 3322 5842 3334 5894
rect 3386 5842 3398 5894
rect 4330 5854 4342 5906
rect 4394 5854 4406 5906
rect 20414 5962 20466 5974
rect 7422 5898 7474 5910
rect 1990 5786 2042 5798
rect 4106 5750 4118 5802
rect 4170 5750 4182 5802
rect 6178 5798 6190 5850
rect 6242 5798 6254 5850
rect 7198 5842 7250 5854
rect 7578 5840 7590 5892
rect 7642 5840 7654 5892
rect 8586 5866 8598 5918
rect 8650 5866 8662 5918
rect 9034 5866 9046 5918
rect 9098 5866 9110 5918
rect 12506 5866 12518 5918
rect 12570 5866 12582 5918
rect 11398 5850 11450 5862
rect 8026 5798 8038 5850
rect 8090 5798 8102 5850
rect 13514 5836 13526 5888
rect 13578 5836 13590 5888
rect 14970 5866 14982 5918
rect 15034 5866 15046 5918
rect 20414 5898 20466 5910
rect 26462 5962 26514 5974
rect 26462 5898 26514 5910
rect 13862 5850 13914 5862
rect 11398 5786 11450 5798
rect 13862 5786 13914 5798
rect 14646 5850 14698 5862
rect 15530 5842 15542 5894
rect 15594 5842 15606 5894
rect 17894 5850 17946 5862
rect 14646 5786 14698 5798
rect 17894 5786 17946 5798
rect 18790 5850 18842 5862
rect 18790 5786 18842 5798
rect 19182 5850 19234 5862
rect 19182 5786 19234 5798
rect 19686 5850 19738 5862
rect 21578 5836 21590 5888
rect 21642 5836 21654 5888
rect 22710 5850 22762 5862
rect 19686 5786 19738 5798
rect 25050 5842 25062 5894
rect 25114 5842 25126 5894
rect 25498 5842 25510 5894
rect 25562 5842 25574 5894
rect 25846 5850 25898 5862
rect 22710 5786 22762 5798
rect 25846 5786 25898 5798
rect 1486 5738 1538 5750
rect 1486 5674 1538 5686
rect 1598 5738 1650 5750
rect 2494 5738 2546 5750
rect 1598 5674 1650 5686
rect 2270 5682 2322 5694
rect 2494 5674 2546 5686
rect 4846 5738 4898 5750
rect 2986 5630 2998 5682
rect 3050 5630 3062 5682
rect 4846 5674 4898 5686
rect 5406 5738 5458 5750
rect 5406 5674 5458 5686
rect 5518 5738 5570 5750
rect 7870 5738 7922 5750
rect 7130 5686 7142 5738
rect 7194 5686 7206 5738
rect 5518 5674 5570 5686
rect 7870 5674 7922 5686
rect 8206 5738 8258 5750
rect 8206 5674 8258 5686
rect 14142 5738 14194 5750
rect 26238 5738 26290 5750
rect 14142 5674 14194 5686
rect 14366 5682 14418 5694
rect 20010 5686 20022 5738
rect 20074 5686 20086 5738
rect 26238 5674 26290 5686
rect 2270 5618 2322 5630
rect 14366 5618 14418 5630
rect 1120 5514 32816 5548
rect 1120 5462 8930 5514
rect 8982 5462 9034 5514
rect 9086 5462 9138 5514
rect 9190 5462 16870 5514
rect 16922 5462 16974 5514
rect 17026 5462 17078 5514
rect 17130 5462 24810 5514
rect 24862 5462 24914 5514
rect 24966 5462 25018 5514
rect 25070 5462 32816 5514
rect 1120 5428 32816 5462
rect 2158 5346 2210 5358
rect 15374 5346 15426 5358
rect 2158 5282 2210 5294
rect 3334 5290 3386 5302
rect 3334 5226 3386 5238
rect 5294 5290 5346 5302
rect 5294 5226 5346 5238
rect 5854 5290 5906 5302
rect 6906 5238 6918 5290
rect 6970 5238 6982 5290
rect 8474 5238 8486 5290
rect 8538 5238 8550 5290
rect 15374 5282 15426 5294
rect 20582 5290 20634 5302
rect 5854 5226 5906 5238
rect 19966 5234 20018 5246
rect 3838 5178 3890 5190
rect 7086 5178 7138 5190
rect 1978 5090 1990 5142
rect 2042 5090 2054 5142
rect 2382 5122 2434 5134
rect 3434 5084 3446 5136
rect 3498 5084 3510 5136
rect 4498 5126 4510 5178
rect 4562 5126 4574 5178
rect 3838 5114 3890 5126
rect 7086 5114 7138 5126
rect 7310 5178 7362 5190
rect 12742 5178 12794 5190
rect 7690 5126 7702 5178
rect 7754 5126 7766 5178
rect 7310 5114 7362 5126
rect 8250 5070 8262 5122
rect 8314 5070 8326 5122
rect 9818 5082 9830 5134
rect 9882 5082 9894 5134
rect 12742 5114 12794 5126
rect 14534 5178 14586 5190
rect 14746 5172 14758 5224
rect 14810 5172 14822 5224
rect 15598 5178 15650 5190
rect 14534 5114 14586 5126
rect 16606 5178 16658 5190
rect 15598 5114 15650 5126
rect 16046 5122 16098 5134
rect 2382 5058 2434 5070
rect 10378 5058 10390 5110
rect 10442 5058 10454 5110
rect 15866 5058 15878 5110
rect 15930 5058 15942 5110
rect 16370 5070 16382 5122
rect 16434 5070 16446 5122
rect 16606 5114 16658 5126
rect 17726 5178 17778 5190
rect 17322 5070 17334 5122
rect 17386 5070 17398 5122
rect 17726 5114 17778 5126
rect 18174 5178 18226 5190
rect 20582 5226 20634 5238
rect 21186 5182 21198 5234
rect 21250 5182 21262 5234
rect 19966 5170 20018 5182
rect 21366 5178 21418 5190
rect 22810 5186 22822 5238
rect 22874 5186 22886 5238
rect 18174 5114 18226 5126
rect 18442 5078 18454 5130
rect 18506 5078 18518 5130
rect 18778 5070 18790 5122
rect 18842 5070 18854 5122
rect 21366 5114 21418 5126
rect 23046 5178 23098 5190
rect 23046 5114 23098 5126
rect 24726 5178 24778 5190
rect 24726 5114 24778 5126
rect 26014 5178 26066 5190
rect 26014 5114 26066 5126
rect 26238 5178 26290 5190
rect 26238 5114 26290 5126
rect 16046 5058 16098 5070
rect 25610 5058 25622 5110
rect 25674 5058 25686 5110
rect 31838 5066 31890 5078
rect 1486 4954 1538 4966
rect 2202 4948 2214 5000
rect 2266 4948 2278 5000
rect 3054 4954 3106 4966
rect 1486 4890 1538 4902
rect 1710 4898 1762 4910
rect 3054 4890 3106 4902
rect 3278 4954 3330 4966
rect 5070 4954 5122 4966
rect 4162 4902 4174 4954
rect 4226 4902 4238 4954
rect 4722 4902 4734 4954
rect 4786 4902 4798 4954
rect 5338 4952 5350 5004
rect 5402 4952 5414 5004
rect 5898 4952 5910 5004
rect 5962 4952 5974 5004
rect 6078 4954 6130 4966
rect 3278 4890 3330 4902
rect 5070 4890 5122 4902
rect 6078 4890 6130 4902
rect 6526 4954 6578 4966
rect 6526 4890 6578 4902
rect 6750 4954 6802 4966
rect 6750 4890 6802 4902
rect 13414 4954 13466 4966
rect 13414 4890 13466 4902
rect 13806 4954 13858 4966
rect 13806 4890 13858 4902
rect 14142 4954 14194 4966
rect 15642 4958 15654 5010
rect 15706 4958 15718 5010
rect 16650 4958 16662 5010
rect 16714 4958 16726 5010
rect 17434 4952 17446 5004
rect 17498 4952 17510 5004
rect 18330 4952 18342 5004
rect 18394 4952 18406 5004
rect 18890 4964 18902 5016
rect 18954 4964 18966 5016
rect 23438 5010 23490 5022
rect 19182 4954 19234 4966
rect 14142 4890 14194 4902
rect 19182 4890 19234 4902
rect 19518 4954 19570 4966
rect 19518 4890 19570 4902
rect 19630 4954 19682 4966
rect 21758 4954 21810 4966
rect 19630 4890 19682 4902
rect 20190 4898 20242 4910
rect 1710 4834 1762 4846
rect 21758 4890 21810 4902
rect 22094 4954 22146 4966
rect 32330 5058 32342 5110
rect 32394 5058 32406 5110
rect 23438 4946 23490 4958
rect 23774 4954 23826 4966
rect 25286 4954 25338 4966
rect 22094 4890 22146 4902
rect 24378 4902 24390 4954
rect 24442 4902 24454 4954
rect 26170 4952 26182 5004
rect 26234 4952 26246 5004
rect 31838 5002 31890 5014
rect 32006 4954 32058 4966
rect 23774 4890 23826 4902
rect 25286 4890 25338 4902
rect 32006 4890 32058 4902
rect 20190 4834 20242 4846
rect 1120 4730 32816 4764
rect 1120 4678 4960 4730
rect 5012 4678 5064 4730
rect 5116 4678 5168 4730
rect 5220 4678 12900 4730
rect 12952 4678 13004 4730
rect 13056 4678 13108 4730
rect 13160 4678 20840 4730
rect 20892 4678 20944 4730
rect 20996 4678 21048 4730
rect 21100 4678 28780 4730
rect 28832 4678 28884 4730
rect 28936 4678 28988 4730
rect 29040 4678 32816 4730
rect 1120 4644 32816 4678
rect 6862 4562 6914 4574
rect 3994 4490 4006 4542
rect 4058 4490 4070 4542
rect 5742 4506 5794 4518
rect 2202 4408 2214 4460
rect 2266 4408 2278 4460
rect 1934 4394 1986 4406
rect 2874 4404 2886 4456
rect 2938 4404 2950 4456
rect 6862 4498 6914 4510
rect 10390 4506 10442 4518
rect 5742 4442 5794 4454
rect 6234 4404 6246 4456
rect 6298 4404 6310 4456
rect 10390 4442 10442 4454
rect 11342 4506 11394 4518
rect 11342 4442 11394 4454
rect 12014 4506 12066 4518
rect 12014 4442 12066 4454
rect 12126 4506 12178 4518
rect 12798 4506 12850 4518
rect 12126 4442 12178 4454
rect 1710 4338 1762 4350
rect 7086 4394 7138 4406
rect 1934 4330 1986 4342
rect 1474 4230 1486 4282
rect 1538 4230 1550 4282
rect 1710 4274 1762 4286
rect 2158 4282 2210 4294
rect 2762 4286 2774 4338
rect 2826 4286 2838 4338
rect 3770 4298 3782 4350
rect 3834 4298 3846 4350
rect 4846 4338 4898 4350
rect 2158 4218 2210 4230
rect 3166 4282 3218 4294
rect 4106 4274 4118 4326
rect 4170 4274 4182 4326
rect 4510 4282 4562 4294
rect 7646 4394 7698 4406
rect 12506 4404 12518 4456
rect 12570 4404 12582 4456
rect 12798 4442 12850 4454
rect 19742 4506 19794 4518
rect 19742 4442 19794 4454
rect 21590 4506 21642 4518
rect 21590 4442 21642 4454
rect 14702 4394 14754 4406
rect 7086 4330 7138 4342
rect 7242 4306 7254 4358
rect 7306 4306 7318 4358
rect 7914 4342 7926 4394
rect 7978 4342 7990 4394
rect 7646 4330 7698 4342
rect 3166 4218 3218 4230
rect 3502 4226 3554 4238
rect 4666 4230 4678 4282
rect 4730 4230 4742 4282
rect 4846 4274 4898 4286
rect 5406 4282 5458 4294
rect 4510 4218 4562 4230
rect 5406 4218 5458 4230
rect 6414 4282 6466 4294
rect 8250 4286 8262 4338
rect 8314 4286 8326 4338
rect 9370 4268 9382 4320
rect 9434 4268 9446 4320
rect 10042 4298 10054 4350
rect 10106 4298 10118 4350
rect 10938 4294 10950 4346
rect 11002 4294 11014 4346
rect 10670 4282 10722 4294
rect 11274 4286 11286 4338
rect 11338 4286 11350 4338
rect 6414 4218 6466 4230
rect 10670 4218 10722 4230
rect 11678 4282 11730 4294
rect 12394 4286 12406 4338
rect 12458 4286 12470 4338
rect 14522 4298 14534 4350
rect 14586 4298 14598 4350
rect 19462 4394 19514 4406
rect 14702 4330 14754 4342
rect 11678 4218 11730 4230
rect 13246 4282 13298 4294
rect 13918 4282 13970 4294
rect 13402 4230 13414 4282
rect 13466 4230 13478 4282
rect 13246 4218 13298 4230
rect 13918 4218 13970 4230
rect 14142 4282 14194 4294
rect 15082 4274 15094 4326
rect 15146 4274 15158 4326
rect 15306 4298 15318 4350
rect 15370 4298 15382 4350
rect 21198 4394 21250 4406
rect 19462 4330 19514 4342
rect 15642 4274 15654 4326
rect 15706 4274 15718 4326
rect 15866 4274 15878 4326
rect 15930 4274 15942 4326
rect 16426 4274 16438 4326
rect 16490 4274 16502 4326
rect 20010 4294 20022 4346
rect 20074 4294 20086 4346
rect 20682 4298 20694 4350
rect 20746 4298 20758 4350
rect 21198 4330 21250 4342
rect 24602 4298 24614 4350
rect 24666 4298 24678 4350
rect 25162 4274 25174 4326
rect 25226 4274 25238 4326
rect 25790 4282 25842 4294
rect 14142 4218 14194 4230
rect 25790 4218 25842 4230
rect 3502 4162 3554 4174
rect 5630 4170 5682 4182
rect 2382 4114 2434 4126
rect 4218 4118 4230 4170
rect 4282 4118 4294 4170
rect 5630 4106 5682 4118
rect 6190 4170 6242 4182
rect 9718 4170 9770 4182
rect 6794 4118 6806 4170
rect 6858 4118 6870 4170
rect 6190 4106 6242 4118
rect 9718 4106 9770 4118
rect 10782 4170 10834 4182
rect 10782 4106 10834 4118
rect 13582 4170 13634 4182
rect 19854 4170 19906 4182
rect 18778 4118 18790 4170
rect 18842 4118 18854 4170
rect 13582 4106 13634 4118
rect 19854 4106 19906 4118
rect 20358 4170 20410 4182
rect 25398 4170 25450 4182
rect 22250 4118 22262 4170
rect 22314 4118 22326 4170
rect 20358 4106 20410 4118
rect 25398 4106 25450 4118
rect 26014 4170 26066 4182
rect 26014 4106 26066 4118
rect 2382 4050 2434 4062
rect 14298 4036 14310 4088
rect 14362 4036 14374 4088
rect 15418 4036 15430 4088
rect 15482 4036 15494 4088
rect 1120 3946 32816 3980
rect 1120 3894 8930 3946
rect 8982 3894 9034 3946
rect 9086 3894 9138 3946
rect 9190 3894 16870 3946
rect 16922 3894 16974 3946
rect 17026 3894 17078 3946
rect 17130 3894 24810 3946
rect 24862 3894 24914 3946
rect 24966 3894 25018 3946
rect 25070 3894 32816 3946
rect 1120 3860 32816 3894
rect 1866 3726 1878 3778
rect 1930 3726 1942 3778
rect 7578 3752 7590 3804
rect 7642 3752 7654 3804
rect 8362 3752 8374 3804
rect 8426 3752 8438 3804
rect 2774 3722 2826 3734
rect 12350 3722 12402 3734
rect 3322 3670 3334 3722
rect 3386 3670 3398 3722
rect 4778 3670 4790 3722
rect 4842 3670 4854 3722
rect 2774 3658 2826 3670
rect 12350 3658 12402 3670
rect 12742 3722 12794 3734
rect 15194 3726 15206 3778
rect 15258 3726 15270 3778
rect 16550 3722 16602 3734
rect 12742 3658 12794 3670
rect 14030 3666 14082 3678
rect 14578 3670 14590 3722
rect 14642 3670 14654 3722
rect 6078 3610 6130 3622
rect 1530 3514 1542 3566
rect 1594 3514 1606 3566
rect 1754 3514 1766 3566
rect 1818 3514 1830 3566
rect 2718 3554 2770 3566
rect 2090 3490 2102 3542
rect 2154 3490 2166 3542
rect 2718 3490 2770 3502
rect 2998 3554 3050 3566
rect 4330 3558 4342 3610
rect 4394 3558 4406 3610
rect 5786 3558 5798 3610
rect 5850 3558 5862 3610
rect 7870 3610 7922 3622
rect 4106 3502 4118 3554
rect 4170 3502 4182 3554
rect 5562 3502 5574 3554
rect 5626 3502 5638 3554
rect 6078 3546 6130 3558
rect 6682 3520 6694 3572
rect 6746 3520 6758 3572
rect 7354 3514 7366 3566
rect 7418 3514 7430 3566
rect 9326 3610 9378 3622
rect 9662 3610 9714 3622
rect 7870 3546 7922 3558
rect 2998 3490 3050 3502
rect 6302 3498 6354 3510
rect 6302 3434 6354 3446
rect 7030 3498 7082 3510
rect 7578 3490 7590 3542
rect 7642 3490 7654 3542
rect 8138 3514 8150 3566
rect 8202 3514 8214 3566
rect 8474 3490 8486 3542
rect 8538 3490 8550 3542
rect 8698 3514 8710 3566
rect 8762 3514 8774 3566
rect 9482 3558 9494 3610
rect 9546 3558 9558 3610
rect 9326 3546 9378 3558
rect 9662 3546 9714 3558
rect 10334 3610 10386 3622
rect 9930 3502 9942 3554
rect 9994 3502 10006 3554
rect 10334 3546 10386 3558
rect 11510 3610 11562 3622
rect 11722 3604 11734 3656
rect 11786 3604 11798 3656
rect 13470 3610 13522 3622
rect 11510 3546 11562 3558
rect 15934 3666 15986 3678
rect 14030 3602 14082 3614
rect 14198 3610 14250 3622
rect 13066 3502 13078 3554
rect 13130 3502 13142 3554
rect 13470 3546 13522 3558
rect 13750 3554 13802 3566
rect 25498 3695 25510 3747
rect 25562 3695 25574 3747
rect 16550 3658 16602 3670
rect 15934 3602 15986 3614
rect 20246 3610 20298 3622
rect 14198 3546 14250 3558
rect 13750 3490 13802 3502
rect 14970 3490 14982 3542
rect 15034 3490 15046 3542
rect 15306 3514 15318 3566
rect 15370 3514 15382 3566
rect 16158 3554 16210 3566
rect 15530 3490 15542 3542
rect 15594 3490 15606 3542
rect 17322 3514 17334 3566
rect 17386 3514 17398 3566
rect 17882 3514 17894 3566
rect 17946 3514 17958 3566
rect 24054 3610 24106 3622
rect 20246 3546 20298 3558
rect 21242 3514 21254 3566
rect 21306 3514 21318 3566
rect 16158 3490 16210 3502
rect 20918 3498 20970 3510
rect 21746 3502 21758 3554
rect 21810 3502 21822 3554
rect 24054 3546 24106 3558
rect 25834 3502 25846 3554
rect 25898 3502 25910 3554
rect 7030 3434 7082 3446
rect 2494 3386 2546 3398
rect 10042 3396 10054 3448
rect 10106 3396 10118 3448
rect 2494 3322 2546 3334
rect 10782 3386 10834 3398
rect 10782 3322 10834 3334
rect 11118 3386 11170 3398
rect 13178 3396 13190 3448
rect 13242 3396 13254 3448
rect 25610 3446 25622 3498
rect 25674 3446 25686 3498
rect 20918 3434 20970 3446
rect 11118 3322 11170 3334
rect 24726 3386 24778 3398
rect 24726 3322 24778 3334
rect 1120 3162 32816 3196
rect 1120 3110 4960 3162
rect 5012 3110 5064 3162
rect 5116 3110 5168 3162
rect 5220 3110 12900 3162
rect 12952 3110 13004 3162
rect 13056 3110 13108 3162
rect 13160 3110 20840 3162
rect 20892 3110 20944 3162
rect 20996 3110 21048 3162
rect 21100 3110 28780 3162
rect 28832 3110 28884 3162
rect 28936 3110 28988 3162
rect 29040 3110 32816 3162
rect 1120 3076 32816 3110
rect 20302 2938 20354 2950
rect 1486 2826 1538 2838
rect 7310 2826 7362 2838
rect 2650 2774 2662 2826
rect 2714 2774 2726 2826
rect 6346 2774 6358 2826
rect 6410 2774 6422 2826
rect 1486 2762 1538 2774
rect 2426 2718 2438 2770
rect 2490 2718 2502 2770
rect 4330 2718 4342 2770
rect 4394 2718 4406 2770
rect 4846 2714 4898 2726
rect 5898 2718 5910 2770
rect 5962 2718 5974 2770
rect 7310 2762 7362 2774
rect 8654 2826 8706 2838
rect 4666 2662 4678 2714
rect 4730 2662 4742 2714
rect 4846 2650 4898 2662
rect 7422 2714 7474 2726
rect 7578 2712 7590 2764
rect 7642 2712 7654 2764
rect 8654 2762 8706 2774
rect 9158 2826 9210 2838
rect 14186 2830 14198 2882
rect 14250 2830 14262 2882
rect 20302 2874 20354 2886
rect 24838 2938 24890 2950
rect 24838 2874 24890 2886
rect 9158 2762 9210 2774
rect 15206 2826 15258 2838
rect 8878 2714 8930 2726
rect 7422 2650 7474 2662
rect 3222 2602 3274 2614
rect 2102 2546 2154 2558
rect 3222 2538 3274 2550
rect 4510 2602 4562 2614
rect 7690 2606 7702 2658
rect 7754 2606 7766 2658
rect 8878 2650 8930 2662
rect 9830 2714 9882 2726
rect 12170 2706 12182 2758
rect 12234 2706 12246 2758
rect 12730 2706 12742 2758
rect 12794 2706 12806 2758
rect 14074 2718 14086 2770
rect 14138 2718 14150 2770
rect 15206 2762 15258 2774
rect 19630 2826 19682 2838
rect 18162 2718 18174 2770
rect 18226 2718 18238 2770
rect 19630 2762 19682 2774
rect 18666 2706 18678 2758
rect 18730 2706 18742 2758
rect 20570 2726 20582 2778
rect 20634 2726 20646 2778
rect 21242 2730 21254 2782
rect 21306 2730 21318 2782
rect 21802 2730 21814 2782
rect 21866 2730 21878 2782
rect 19406 2714 19458 2726
rect 9830 2650 9882 2662
rect 25386 2700 25398 2752
rect 25450 2700 25462 2752
rect 19406 2650 19458 2662
rect 8262 2602 8314 2614
rect 4510 2538 4562 2550
rect 5798 2546 5850 2558
rect 2102 2482 2154 2494
rect 5798 2482 5850 2494
rect 7198 2546 7250 2558
rect 8262 2538 8314 2550
rect 13246 2602 13298 2614
rect 13246 2538 13298 2550
rect 13470 2602 13522 2614
rect 19014 2602 19066 2614
rect 14858 2550 14870 2602
rect 14922 2550 14934 2602
rect 15866 2550 15878 2602
rect 15930 2550 15942 2602
rect 13470 2538 13522 2550
rect 19014 2538 19066 2550
rect 19966 2602 20018 2614
rect 19966 2538 20018 2550
rect 20414 2602 20466 2614
rect 25062 2602 25114 2614
rect 24154 2550 24166 2602
rect 24218 2550 24230 2602
rect 20414 2538 20466 2550
rect 25062 2538 25114 2550
rect 25678 2602 25730 2614
rect 25678 2538 25730 2550
rect 25902 2602 25954 2614
rect 25902 2538 25954 2550
rect 7198 2482 7250 2494
rect 1120 2378 32816 2412
rect 1120 2326 8930 2378
rect 8982 2326 9034 2378
rect 9086 2326 9138 2378
rect 9190 2326 16870 2378
rect 16922 2326 16974 2378
rect 17026 2326 17078 2378
rect 17130 2326 24810 2378
rect 24862 2326 24914 2378
rect 24966 2326 25018 2378
rect 25070 2326 32816 2378
rect 1120 2292 32816 2326
rect 4790 2154 4842 2166
rect 3994 2102 4006 2154
rect 4058 2102 4070 2154
rect 7690 2127 7702 2179
rect 7754 2127 7766 2179
rect 17278 2154 17330 2166
rect 2090 2046 2102 2098
rect 2154 2046 2166 2098
rect 4790 2090 4842 2102
rect 3334 2042 3386 2054
rect 5574 2042 5626 2054
rect 6346 2046 6358 2098
rect 6410 2046 6422 2098
rect 6906 2046 6918 2098
rect 6970 2046 6982 2098
rect 17278 2090 17330 2102
rect 23214 2154 23266 2166
rect 23214 2090 23266 2102
rect 24334 2154 24386 2166
rect 24334 2090 24386 2102
rect 32006 2154 32058 2166
rect 32006 2090 32058 2102
rect 4442 1990 4454 2042
rect 4506 1990 4518 2042
rect 3334 1978 3386 1990
rect 5574 1978 5626 1990
rect 12406 2042 12458 2054
rect 2438 1930 2490 1942
rect 6122 1934 6134 1986
rect 6186 1934 6198 1986
rect 7018 1934 7030 1986
rect 7082 1934 7094 1986
rect 8138 1934 8150 1986
rect 8202 1934 8214 1986
rect 7914 1878 7926 1930
rect 7978 1878 7990 1930
rect 9594 1922 9606 1974
rect 9658 1922 9670 1974
rect 10098 1934 10110 1986
rect 10162 1934 10174 1986
rect 12406 1978 12458 1990
rect 16214 2042 16266 2054
rect 16214 1978 16266 1990
rect 17950 2042 18002 2054
rect 21478 2042 21530 2054
rect 17950 1978 18002 1990
rect 13078 1930 13130 1942
rect 13290 1922 13302 1974
rect 13354 1922 13366 1974
rect 13850 1922 13862 1974
rect 13914 1922 13926 1974
rect 18330 1934 18342 1986
rect 18394 1934 18406 1986
rect 18554 1946 18566 1998
rect 18618 1946 18630 1998
rect 19114 1946 19126 1998
rect 19178 1946 19190 1998
rect 21478 1978 21530 1990
rect 22766 2042 22818 2054
rect 22150 1930 22202 1942
rect 22362 1934 22374 1986
rect 22426 1934 22438 1986
rect 22766 1978 22818 1990
rect 23102 2042 23154 2054
rect 23102 1978 23154 1990
rect 23774 2042 23826 2054
rect 23774 1978 23826 1990
rect 2438 1866 2490 1878
rect 6682 1822 6694 1874
rect 6746 1822 6758 1874
rect 13078 1866 13130 1878
rect 23370 1926 23382 1978
rect 23434 1926 23446 1978
rect 24042 1926 24054 1978
rect 24106 1926 24118 1978
rect 31838 1930 31890 1942
rect 22150 1866 22202 1878
rect 32330 1922 32342 1974
rect 32394 1922 32406 1974
rect 16886 1818 16938 1830
rect 16886 1754 16938 1766
rect 18286 1818 18338 1830
rect 22474 1816 22486 1868
rect 22538 1816 22550 1868
rect 23930 1816 23942 1868
rect 23994 1816 24006 1868
rect 31838 1866 31890 1878
rect 18286 1754 18338 1766
rect 1120 1594 32816 1628
rect 1120 1542 4960 1594
rect 5012 1542 5064 1594
rect 5116 1542 5168 1594
rect 5220 1542 12900 1594
rect 12952 1542 13004 1594
rect 13056 1542 13108 1594
rect 13160 1542 20840 1594
rect 20892 1542 20944 1594
rect 20996 1542 21048 1594
rect 21100 1542 28780 1594
rect 28832 1542 28884 1594
rect 28936 1542 28988 1594
rect 29040 1542 32816 1594
rect 1120 1508 32816 1542
rect 11566 1426 11618 1438
rect 4342 1370 4394 1382
rect 6750 1370 6802 1382
rect 7646 1370 7698 1382
rect 8822 1370 8874 1382
rect 6402 1318 6414 1370
rect 6466 1318 6478 1370
rect 6962 1318 6974 1370
rect 7026 1318 7038 1370
rect 7298 1318 7310 1370
rect 7362 1318 7374 1370
rect 7858 1318 7870 1370
rect 7922 1318 7934 1370
rect 4342 1306 4394 1318
rect 6750 1306 6802 1318
rect 7646 1306 7698 1318
rect 8822 1306 8874 1318
rect 9718 1370 9770 1382
rect 9718 1306 9770 1318
rect 10838 1370 10890 1382
rect 10838 1306 10890 1318
rect 11230 1370 11282 1382
rect 11566 1362 11618 1374
rect 14086 1370 14138 1382
rect 11230 1306 11282 1318
rect 14086 1306 14138 1318
rect 14814 1370 14866 1382
rect 14814 1306 14866 1318
rect 16438 1370 16490 1382
rect 16438 1306 16490 1318
rect 17558 1370 17610 1382
rect 17558 1306 17610 1318
rect 17782 1370 17834 1382
rect 17782 1306 17834 1318
rect 18454 1370 18506 1382
rect 18454 1306 18506 1318
rect 19126 1370 19178 1382
rect 19126 1306 19178 1318
rect 20022 1370 20074 1382
rect 20022 1306 20074 1318
rect 21758 1370 21810 1382
rect 21758 1306 21810 1318
rect 22374 1370 22426 1382
rect 13358 1258 13410 1270
rect 1530 1150 1542 1202
rect 1594 1150 1606 1202
rect 4666 1132 4678 1184
rect 4730 1132 4742 1184
rect 5786 1162 5798 1214
rect 5850 1162 5862 1214
rect 8474 1162 8486 1214
rect 8538 1162 8550 1214
rect 10042 1162 10054 1214
rect 10106 1162 10118 1214
rect 13358 1194 13410 1206
rect 16606 1258 16658 1270
rect 21914 1256 21926 1308
rect 21978 1256 21990 1308
rect 22374 1306 22426 1318
rect 23494 1370 23546 1382
rect 23494 1306 23546 1318
rect 25622 1370 25674 1382
rect 25622 1306 25674 1318
rect 16606 1194 16658 1206
rect 5518 1146 5570 1158
rect 5518 1082 5570 1094
rect 6078 1146 6130 1158
rect 6078 1082 6130 1094
rect 8094 1146 8146 1158
rect 10490 1132 10502 1184
rect 10554 1132 10566 1184
rect 17210 1162 17222 1214
rect 17274 1162 17286 1214
rect 18106 1162 18118 1214
rect 18170 1162 18182 1214
rect 18778 1162 18790 1214
rect 18842 1162 18854 1214
rect 21354 1162 21366 1214
rect 21418 1162 21430 1214
rect 11958 1146 12010 1158
rect 14478 1146 14530 1158
rect 8094 1082 8146 1094
rect 13738 1094 13750 1146
rect 13802 1094 13814 1146
rect 11958 1082 12010 1094
rect 2550 1034 2602 1046
rect 12114 1038 12126 1090
rect 12178 1038 12190 1090
rect 14478 1082 14530 1094
rect 15206 1146 15258 1158
rect 16046 1146 16098 1158
rect 15206 1082 15258 1094
rect 15418 1048 15430 1100
rect 15482 1048 15494 1100
rect 20346 1094 20358 1146
rect 20410 1094 20422 1146
rect 22026 1142 22038 1194
rect 22090 1142 22102 1194
rect 22698 1162 22710 1214
rect 22762 1162 22774 1214
rect 23146 1162 23158 1214
rect 23210 1162 23222 1214
rect 25946 1132 25958 1184
rect 26010 1132 26022 1184
rect 16046 1082 16098 1094
rect 2550 970 2602 982
rect 19518 1034 19570 1046
rect 19518 970 19570 982
rect 19742 1034 19794 1046
rect 19742 970 19794 982
rect 21030 1034 21082 1046
rect 21030 970 21082 982
rect 26238 1034 26290 1046
rect 26238 970 26290 982
rect 5786 900 5798 952
rect 5850 900 5862 952
rect 1120 810 32816 844
rect 1120 758 8930 810
rect 8982 758 9034 810
rect 9086 758 9138 810
rect 9190 758 16870 810
rect 16922 758 16974 810
rect 17026 758 17078 810
rect 17130 758 24810 810
rect 24862 758 24914 810
rect 24966 758 25018 810
rect 25070 758 32816 810
rect 1120 724 32816 758
rect 20122 534 20134 586
rect 20186 583 20198 586
rect 21018 583 21030 586
rect 20186 537 21030 583
rect 20186 534 20198 537
rect 21018 534 21030 537
rect 21082 534 21094 586
<< via1 >>
rect 4960 18790 5012 18842
rect 5064 18790 5116 18842
rect 5168 18790 5220 18842
rect 12900 18790 12952 18842
rect 13004 18790 13056 18842
rect 13108 18790 13160 18842
rect 20840 18790 20892 18842
rect 20944 18790 20996 18842
rect 21048 18790 21100 18842
rect 28780 18790 28832 18842
rect 28884 18790 28936 18842
rect 28988 18790 29040 18842
rect 1878 18566 1930 18618
rect 6918 18566 6970 18618
rect 16494 18566 16546 18618
rect 21870 18566 21922 18618
rect 23102 18566 23154 18618
rect 25790 18566 25842 18618
rect 1542 18410 1594 18462
rect 3390 18454 3442 18506
rect 6078 18454 6130 18506
rect 2942 18342 2994 18394
rect 3950 18342 4002 18394
rect 4510 18342 4562 18394
rect 6526 18342 6578 18394
rect 7142 18398 7194 18450
rect 10166 18454 10218 18506
rect 9998 18398 10050 18450
rect 8710 18342 8762 18394
rect 15990 18454 16042 18506
rect 11342 18398 11394 18450
rect 10166 18320 10218 18372
rect 10614 18342 10666 18394
rect 11174 18342 11226 18394
rect 11734 18380 11786 18432
rect 13302 18398 13354 18450
rect 14870 18342 14922 18394
rect 15430 18380 15482 18432
rect 15822 18398 15874 18450
rect 17222 18410 17274 18462
rect 18006 18454 18058 18506
rect 15990 18320 16042 18372
rect 16438 18342 16490 18394
rect 16606 18342 16658 18394
rect 19238 18398 19290 18450
rect 21142 18410 21194 18462
rect 22598 18410 22650 18462
rect 23998 18454 24050 18506
rect 24558 18454 24610 18506
rect 27190 18410 27242 18462
rect 28142 18454 28194 18506
rect 30718 18454 30770 18506
rect 18006 18320 18058 18372
rect 18286 18342 18338 18394
rect 18454 18342 18506 18394
rect 18622 18342 18674 18394
rect 20582 18342 20634 18394
rect 23774 18342 23826 18394
rect 25006 18342 25058 18394
rect 27638 18380 27690 18432
rect 30494 18342 30546 18394
rect 32398 18342 32450 18394
rect 2158 18230 2210 18282
rect 2550 18230 2602 18282
rect 2718 18230 2770 18282
rect 3166 18230 3218 18282
rect 4342 18230 4394 18282
rect 6302 18230 6354 18282
rect 7982 18230 8034 18282
rect 9326 18230 9378 18282
rect 9718 18230 9770 18282
rect 10446 18230 10498 18282
rect 10782 18230 10834 18282
rect 11006 18230 11058 18282
rect 12070 18230 12122 18282
rect 12406 18230 12458 18282
rect 12742 18230 12794 18282
rect 14030 18230 14082 18282
rect 15094 18230 15146 18282
rect 17558 18230 17610 18282
rect 17838 18230 17890 18282
rect 19742 18230 19794 18282
rect 21478 18230 21530 18282
rect 21982 18230 22034 18282
rect 22262 18230 22314 18282
rect 22990 18230 23042 18282
rect 23438 18230 23490 18282
rect 23550 18230 23602 18282
rect 25398 18230 25450 18282
rect 25902 18230 25954 18282
rect 26238 18230 26290 18282
rect 26630 18230 26682 18282
rect 26854 18230 26906 18282
rect 27974 18230 28026 18282
rect 29374 18230 29426 18282
rect 29486 18230 29538 18282
rect 30102 18230 30154 18282
rect 31334 18230 31386 18282
rect 31726 18230 31778 18282
rect 32006 18230 32058 18282
rect 8930 18006 8982 18058
rect 9034 18006 9086 18058
rect 9138 18006 9190 18058
rect 16870 18006 16922 18058
rect 16974 18006 17026 18058
rect 17078 18006 17130 18058
rect 24810 18006 24862 18058
rect 24914 18006 24966 18058
rect 25018 18006 25070 18058
rect 1486 17782 1538 17834
rect 5854 17782 5906 17834
rect 10054 17782 10106 17834
rect 11790 17782 11842 17834
rect 15430 17782 15482 17834
rect 16438 17782 16490 17834
rect 17278 17782 17330 17834
rect 19518 17782 19570 17834
rect 20582 17782 20634 17834
rect 23214 17782 23266 17834
rect 26126 17782 26178 17834
rect 32510 17782 32562 17834
rect 2046 17670 2098 17722
rect 2550 17692 2602 17744
rect 6806 17670 6858 17722
rect 2382 17614 2434 17666
rect 2550 17558 2602 17610
rect 3726 17558 3778 17610
rect 6414 17558 6466 17610
rect 6974 17614 7026 17666
rect 7254 17614 7306 17666
rect 9494 17633 9546 17685
rect 12630 17670 12682 17722
rect 8094 17558 8146 17610
rect 8934 17558 8986 17610
rect 9774 17558 9826 17610
rect 10390 17602 10442 17654
rect 10782 17558 10834 17610
rect 10950 17614 11002 17666
rect 14422 17670 14474 17722
rect 12854 17614 12906 17666
rect 14982 17633 15034 17685
rect 15822 17670 15874 17722
rect 16102 17670 16154 17722
rect 17670 17670 17722 17722
rect 17838 17670 17890 17722
rect 18062 17670 18114 17722
rect 18230 17670 18282 17722
rect 18398 17670 18450 17722
rect 13694 17558 13746 17610
rect 20022 17614 20074 17666
rect 16830 17558 16882 17610
rect 18790 17558 18842 17610
rect 20918 17602 20970 17654
rect 21366 17633 21418 17685
rect 22094 17670 22146 17722
rect 28758 17670 28810 17722
rect 22374 17614 22426 17666
rect 26742 17614 26794 17666
rect 27190 17614 27242 17666
rect 24054 17558 24106 17610
rect 1878 17446 1930 17498
rect 2942 17446 2994 17498
rect 3054 17446 3106 17498
rect 3390 17446 3442 17498
rect 3502 17446 3554 17498
rect 5966 17446 6018 17498
rect 6302 17446 6354 17498
rect 6862 17446 6914 17498
rect 14982 17485 15034 17537
rect 17726 17446 17778 17498
rect 21422 17446 21474 17498
rect 21982 17446 22034 17498
rect 24726 17508 24778 17560
rect 25286 17558 25338 17610
rect 28030 17558 28082 17610
rect 29094 17614 29146 17666
rect 31334 17614 31386 17666
rect 29934 17558 29986 17610
rect 30774 17558 30826 17610
rect 32062 17558 32114 17610
rect 24446 17446 24498 17498
rect 30998 17446 31050 17498
rect 4960 17222 5012 17274
rect 5064 17222 5116 17274
rect 5168 17222 5220 17274
rect 12900 17222 12952 17274
rect 13004 17222 13056 17274
rect 13108 17222 13160 17274
rect 20840 17222 20892 17274
rect 20944 17222 20996 17274
rect 21048 17222 21100 17274
rect 28780 17222 28832 17274
rect 28884 17222 28936 17274
rect 28988 17222 29040 17274
rect 1878 16998 1930 17050
rect 6022 16998 6074 17050
rect 12294 16998 12346 17050
rect 15990 16998 16042 17050
rect 31334 16959 31386 17011
rect 1542 16842 1594 16894
rect 2662 16830 2714 16882
rect 6358 16842 6410 16894
rect 3894 16774 3946 16826
rect 4286 16774 4338 16826
rect 6694 16830 6746 16882
rect 7534 16886 7586 16938
rect 8374 16886 8426 16938
rect 10166 16886 10218 16938
rect 8598 16830 8650 16882
rect 10726 16842 10778 16894
rect 11622 16842 11674 16894
rect 14982 16886 15034 16938
rect 13302 16830 13354 16882
rect 17222 16842 17274 16894
rect 18006 16886 18058 16938
rect 18566 16886 18618 16938
rect 24950 16886 25002 16938
rect 28422 16886 28474 16938
rect 30886 16886 30938 16938
rect 11958 16774 12010 16826
rect 17838 16830 17890 16882
rect 20022 16830 20074 16882
rect 15542 16774 15594 16826
rect 18006 16752 18058 16804
rect 20470 16774 20522 16826
rect 22262 16812 22314 16864
rect 23382 16830 23434 16882
rect 26294 16830 26346 16882
rect 26854 16830 26906 16882
rect 29542 16830 29594 16882
rect 24614 16774 24666 16826
rect 31222 16811 31274 16863
rect 2046 16662 2098 16714
rect 3166 16662 3218 16714
rect 4678 16662 4730 16714
rect 9438 16662 9490 16714
rect 11062 16662 11114 16714
rect 11286 16662 11338 16714
rect 12350 16606 12402 16658
rect 12574 16606 12626 16658
rect 12910 16662 12962 16714
rect 14142 16662 14194 16714
rect 15262 16662 15314 16714
rect 15934 16606 15986 16658
rect 16158 16606 16210 16658
rect 16438 16662 16490 16714
rect 16774 16662 16826 16714
rect 17558 16662 17610 16714
rect 19294 16662 19346 16714
rect 20302 16662 20354 16714
rect 20638 16662 20690 16714
rect 21310 16662 21362 16714
rect 21422 16662 21474 16714
rect 21758 16662 21810 16714
rect 21870 16662 21922 16714
rect 22598 16662 22650 16714
rect 23886 16662 23938 16714
rect 25790 16662 25842 16714
rect 27694 16662 27746 16714
rect 30046 16662 30098 16714
rect 8930 16438 8982 16490
rect 9034 16438 9086 16490
rect 9138 16438 9190 16490
rect 16870 16438 16922 16490
rect 16974 16438 17026 16490
rect 17078 16438 17130 16490
rect 24810 16438 24862 16490
rect 24914 16438 24966 16490
rect 25018 16438 25070 16490
rect 3726 16214 3778 16266
rect 6638 16214 6690 16266
rect 9830 16214 9882 16266
rect 10110 16214 10162 16266
rect 10222 16214 10274 16266
rect 10558 16214 10610 16266
rect 11006 16214 11058 16266
rect 12126 16214 12178 16266
rect 14870 16214 14922 16266
rect 15710 16214 15762 16266
rect 15822 16214 15874 16266
rect 18734 16214 18786 16266
rect 19294 16214 19346 16266
rect 20414 16214 20466 16266
rect 21646 16214 21698 16266
rect 22654 16214 22706 16266
rect 24110 16214 24162 16266
rect 24502 16214 24554 16266
rect 25230 16214 25282 16266
rect 25566 16214 25618 16266
rect 26126 16214 26178 16266
rect 27246 16214 27298 16266
rect 28478 16214 28530 16266
rect 31502 16214 31554 16266
rect 1542 16034 1594 16086
rect 2550 16065 2602 16117
rect 4566 16102 4618 16154
rect 2998 16046 3050 16098
rect 4902 16065 4954 16117
rect 6750 15990 6802 16042
rect 7030 16046 7082 16098
rect 8878 16102 8930 16154
rect 11174 16124 11226 16176
rect 11566 16102 11618 16154
rect 11790 16102 11842 16154
rect 14646 16102 14698 16154
rect 16214 16102 16266 16154
rect 16774 16124 16826 16176
rect 7870 15990 7922 16042
rect 8710 15990 8762 16042
rect 9494 16034 9546 16086
rect 13302 16046 13354 16098
rect 13526 16046 13578 16098
rect 15598 16046 15650 16098
rect 10670 15990 10722 16042
rect 11174 15990 11226 16042
rect 16606 16046 16658 16098
rect 17390 16046 17442 16098
rect 17614 16102 17666 16154
rect 18006 16102 18058 16154
rect 16774 15990 16826 16042
rect 18342 16046 18394 16098
rect 18622 16046 18674 16098
rect 18846 16046 18898 16098
rect 19070 16102 19122 16154
rect 21534 16102 21586 16154
rect 22262 16124 22314 16176
rect 22822 16124 22874 16176
rect 23382 16124 23434 16176
rect 19910 16046 19962 16098
rect 22094 16046 22146 16098
rect 21142 15990 21194 16042
rect 21702 15990 21754 16042
rect 23214 16046 23266 16098
rect 23774 16102 23826 16154
rect 25398 16102 25450 16154
rect 25958 16102 26010 16154
rect 26518 16102 26570 16154
rect 22262 15990 22314 16042
rect 22822 15990 22874 16042
rect 23382 15990 23434 16042
rect 24782 15990 24834 16042
rect 28086 16046 28138 16098
rect 28366 16102 28418 16154
rect 28870 16046 28922 16098
rect 31110 16064 31162 16116
rect 29710 15990 29762 16042
rect 30550 15990 30602 16042
rect 1878 15878 1930 15930
rect 2494 15878 2546 15930
rect 4958 15878 5010 15930
rect 17558 15878 17610 15930
rect 26014 15878 26066 15930
rect 30774 15878 30826 15930
rect 31614 15878 31666 15930
rect 4960 15654 5012 15706
rect 5064 15654 5116 15706
rect 5168 15654 5220 15706
rect 12900 15654 12952 15706
rect 13004 15654 13056 15706
rect 13108 15654 13160 15706
rect 20840 15654 20892 15706
rect 20944 15654 20996 15706
rect 21048 15654 21100 15706
rect 28780 15654 28832 15706
rect 28884 15654 28936 15706
rect 28988 15654 29040 15706
rect 2270 15430 2322 15482
rect 2382 15430 2434 15482
rect 6470 15430 6522 15482
rect 18734 15486 18786 15538
rect 10670 15430 10722 15482
rect 12518 15386 12570 15438
rect 13750 15430 13802 15482
rect 14982 15430 15034 15482
rect 16774 15430 16826 15482
rect 17334 15430 17386 15482
rect 18958 15486 19010 15538
rect 14366 15374 14418 15426
rect 2886 15318 2938 15370
rect 4790 15318 4842 15370
rect 5518 15318 5570 15370
rect 3222 15262 3274 15314
rect 2886 15184 2938 15236
rect 4062 15206 4114 15258
rect 6134 15244 6186 15296
rect 6694 15262 6746 15314
rect 10278 15318 10330 15370
rect 15766 15374 15818 15426
rect 19798 15386 19850 15438
rect 8598 15262 8650 15314
rect 7534 15206 7586 15258
rect 8262 15206 8314 15258
rect 10614 15243 10666 15295
rect 12070 15250 12122 15302
rect 12630 15274 12682 15326
rect 14590 15318 14642 15370
rect 13414 15206 13466 15258
rect 13806 15206 13858 15258
rect 15206 15248 15258 15300
rect 16158 15262 16210 15314
rect 16270 15262 16322 15314
rect 18118 15318 18170 15370
rect 17950 15262 18002 15314
rect 16998 15206 17050 15258
rect 18566 15248 18618 15300
rect 19686 15274 19738 15326
rect 20078 15262 20130 15314
rect 20526 15318 20578 15370
rect 22262 15374 22314 15426
rect 23158 15384 23210 15436
rect 23942 15430 23994 15482
rect 25734 15384 25786 15436
rect 31334 15391 31386 15443
rect 21198 15318 21250 15370
rect 22766 15318 22818 15370
rect 24558 15318 24610 15370
rect 25118 15318 25170 15370
rect 21702 15248 21754 15300
rect 1486 15094 1538 15146
rect 1878 15094 1930 15146
rect 2718 15094 2770 15146
rect 5406 15094 5458 15146
rect 9438 15094 9490 15146
rect 11398 15094 11450 15146
rect 11734 15094 11786 15146
rect 12238 15038 12290 15090
rect 12462 15094 12514 15146
rect 14030 15038 14082 15090
rect 15486 15094 15538 15146
rect 15710 15094 15762 15146
rect 16494 15094 16546 15146
rect 16718 15150 16770 15202
rect 18118 15184 18170 15236
rect 22542 15206 22594 15258
rect 23046 15242 23098 15294
rect 23214 15206 23266 15258
rect 24894 15206 24946 15258
rect 25342 15262 25394 15314
rect 25566 15318 25618 15370
rect 28758 15318 28810 15370
rect 26686 15262 26738 15314
rect 27414 15262 27466 15314
rect 26014 15206 26066 15258
rect 26518 15206 26570 15258
rect 27918 15206 27970 15258
rect 29206 15262 29258 15314
rect 30046 15318 30098 15370
rect 30886 15318 30938 15370
rect 31222 15243 31274 15295
rect 32342 15244 32394 15296
rect 17390 15038 17442 15090
rect 17614 15094 17666 15146
rect 19014 15094 19066 15146
rect 19854 15094 19906 15146
rect 20302 15094 20354 15146
rect 21534 15094 21586 15146
rect 21982 15038 22034 15090
rect 22206 15038 22258 15090
rect 23438 15094 23490 15146
rect 24334 15094 24386 15146
rect 25790 15038 25842 15090
rect 26350 15094 26402 15146
rect 31838 15094 31890 15146
rect 32006 15094 32058 15146
rect 8930 14870 8982 14922
rect 9034 14870 9086 14922
rect 9138 14870 9190 14922
rect 16870 14870 16922 14922
rect 16974 14870 17026 14922
rect 17078 14870 17130 14922
rect 24810 14870 24862 14922
rect 24914 14870 24966 14922
rect 25018 14870 25070 14922
rect 12182 14728 12234 14780
rect 4678 14646 4730 14698
rect 19070 14702 19122 14754
rect 6862 14646 6914 14698
rect 8094 14646 8146 14698
rect 13190 14646 13242 14698
rect 14646 14612 14698 14664
rect 16550 14646 16602 14698
rect 22206 14702 22258 14754
rect 19294 14646 19346 14698
rect 20470 14646 20522 14698
rect 21646 14646 21698 14698
rect 23886 14646 23938 14698
rect 26126 14646 26178 14698
rect 26574 14646 26626 14698
rect 27582 14646 27634 14698
rect 27806 14646 27858 14698
rect 27918 14646 27970 14698
rect 28254 14646 28306 14698
rect 28366 14646 28418 14698
rect 31054 14646 31106 14698
rect 31838 14646 31890 14698
rect 1486 14534 1538 14586
rect 3782 14534 3834 14586
rect 2102 14478 2154 14530
rect 8822 14534 8874 14586
rect 2942 14422 2994 14474
rect 4118 14472 4170 14524
rect 5014 14466 5066 14518
rect 6974 14422 7026 14474
rect 7254 14478 7306 14530
rect 9718 14496 9770 14548
rect 10278 14534 10330 14586
rect 10950 14556 11002 14608
rect 11510 14556 11562 14608
rect 10446 14478 10498 14530
rect 10782 14478 10834 14530
rect 11342 14478 11394 14530
rect 11846 14490 11898 14542
rect 10950 14422 11002 14474
rect 12182 14466 12234 14518
rect 12406 14490 12458 14542
rect 12854 14534 12906 14586
rect 13638 14466 13690 14518
rect 13806 14478 13858 14530
rect 14030 14534 14082 14586
rect 19966 14534 20018 14586
rect 21086 14534 21138 14586
rect 21310 14534 21362 14586
rect 22430 14534 22482 14586
rect 14310 14478 14362 14530
rect 14758 14478 14810 14530
rect 15542 14478 15594 14530
rect 16102 14478 16154 14530
rect 16326 14478 16378 14530
rect 17670 14478 17722 14530
rect 17390 14422 17442 14474
rect 18622 14422 18674 14474
rect 18902 14466 18954 14518
rect 19742 14478 19794 14530
rect 20470 14466 20522 14518
rect 22038 14458 22090 14510
rect 22654 14478 22706 14530
rect 22934 14478 22986 14530
rect 23662 14478 23714 14530
rect 24054 14484 24106 14536
rect 24390 14478 24442 14530
rect 25342 14478 25394 14530
rect 25958 14534 26010 14586
rect 26350 14534 26402 14586
rect 26742 14534 26794 14586
rect 27414 14556 27466 14608
rect 25566 14478 25618 14530
rect 26910 14478 26962 14530
rect 31726 14534 31778 14586
rect 27246 14478 27298 14530
rect 29318 14478 29370 14530
rect 1878 14310 1930 14362
rect 4230 14349 4282 14401
rect 9382 14310 9434 14362
rect 10334 14310 10386 14362
rect 11454 14310 11506 14362
rect 14086 14354 14138 14406
rect 17894 14360 17946 14412
rect 18062 14310 18114 14362
rect 18398 14310 18450 14362
rect 19014 14356 19066 14408
rect 23046 14372 23098 14424
rect 29934 14422 29986 14474
rect 30774 14422 30826 14474
rect 20246 14274 20298 14326
rect 22598 14310 22650 14362
rect 23326 14310 23378 14362
rect 23942 14356 23994 14408
rect 25622 14310 25674 14362
rect 28702 14310 28754 14362
rect 28814 14310 28866 14362
rect 31446 14310 31498 14362
rect 4960 14086 5012 14138
rect 5064 14086 5116 14138
rect 5168 14086 5220 14138
rect 12900 14086 12952 14138
rect 13004 14086 13056 14138
rect 13108 14086 13160 14138
rect 20840 14086 20892 14138
rect 20944 14086 20996 14138
rect 21048 14086 21100 14138
rect 28780 14086 28832 14138
rect 28884 14086 28936 14138
rect 28988 14086 29040 14138
rect 5518 13862 5570 13914
rect 23214 13918 23266 13970
rect 6694 13862 6746 13914
rect 8150 13862 8202 13914
rect 9494 13862 9546 13914
rect 9830 13862 9882 13914
rect 11286 13862 11338 13914
rect 15318 13816 15370 13868
rect 22654 13862 22706 13914
rect 24558 13918 24610 13970
rect 24782 13918 24834 13970
rect 20694 13806 20746 13858
rect 2326 13750 2378 13802
rect 3502 13750 3554 13802
rect 4230 13750 4282 13802
rect 2158 13694 2210 13746
rect 2998 13694 3050 13746
rect 6358 13706 6410 13758
rect 6918 13706 6970 13758
rect 2326 13616 2378 13668
rect 5854 13638 5906 13690
rect 7254 13682 7306 13734
rect 7478 13706 7530 13758
rect 7814 13638 7866 13690
rect 8206 13638 8258 13690
rect 8430 13694 8482 13746
rect 9942 13694 9994 13746
rect 10166 13694 10218 13746
rect 12406 13706 12458 13758
rect 12686 13750 12738 13802
rect 13638 13750 13690 13802
rect 18342 13750 18394 13802
rect 11790 13638 11842 13690
rect 14086 13694 14138 13746
rect 12238 13638 12290 13690
rect 13638 13616 13690 13668
rect 14758 13638 14810 13690
rect 1486 13526 1538 13578
rect 1878 13526 1930 13578
rect 4622 13526 4674 13578
rect 4734 13526 4786 13578
rect 5406 13526 5458 13578
rect 5966 13526 6018 13578
rect 9102 13526 9154 13578
rect 7142 13470 7194 13522
rect 10950 13526 11002 13578
rect 11454 13526 11506 13578
rect 12014 13470 12066 13522
rect 12126 13526 12178 13578
rect 14198 13582 14250 13634
rect 15262 13638 15314 13690
rect 15430 13688 15482 13740
rect 15766 13694 15818 13746
rect 16438 13694 16490 13746
rect 17670 13694 17722 13746
rect 18790 13706 18842 13758
rect 19574 13750 19626 13802
rect 21478 13750 21530 13802
rect 22094 13750 22146 13802
rect 22990 13806 23042 13858
rect 27526 13862 27578 13914
rect 27806 13862 27858 13914
rect 31110 13862 31162 13914
rect 17334 13638 17386 13690
rect 13470 13526 13522 13578
rect 17782 13582 17834 13634
rect 18342 13616 18394 13668
rect 18958 13638 19010 13690
rect 19294 13638 19346 13690
rect 20302 13638 20354 13690
rect 20526 13638 20578 13690
rect 21310 13694 21362 13746
rect 24054 13750 24106 13802
rect 21926 13682 21978 13734
rect 22262 13638 22314 13690
rect 23886 13694 23938 13746
rect 25510 13750 25562 13802
rect 25062 13697 25114 13749
rect 26070 13706 26122 13758
rect 26406 13706 26458 13758
rect 26630 13682 26682 13734
rect 29206 13694 29258 13746
rect 30046 13750 30098 13802
rect 24054 13616 24106 13668
rect 25510 13616 25562 13668
rect 30774 13638 30826 13690
rect 31446 13676 31498 13728
rect 15038 13526 15090 13578
rect 17110 13526 17162 13578
rect 18174 13526 18226 13578
rect 19966 13526 20018 13578
rect 19126 13470 19178 13522
rect 20750 13526 20802 13578
rect 21422 13526 21474 13578
rect 23606 13526 23658 13578
rect 24502 13526 24554 13578
rect 25342 13526 25394 13578
rect 25790 13526 25842 13578
rect 27134 13526 27186 13578
rect 27918 13526 27970 13578
rect 28254 13526 28306 13578
rect 28366 13526 28418 13578
rect 26406 13444 26458 13496
rect 8930 13302 8982 13354
rect 9034 13302 9086 13354
rect 9138 13302 9190 13354
rect 16870 13302 16922 13354
rect 16974 13302 17026 13354
rect 17078 13302 17130 13354
rect 24810 13302 24862 13354
rect 24914 13302 24966 13354
rect 25018 13302 25070 13354
rect 1598 13078 1650 13130
rect 3502 13078 3554 13130
rect 6638 13078 6690 13130
rect 8654 13134 8706 13186
rect 6862 13078 6914 13130
rect 7590 13078 7642 13130
rect 14758 13134 14810 13186
rect 8878 13078 8930 13130
rect 2438 12966 2490 13018
rect 4566 12966 4618 13018
rect 7030 12988 7082 13040
rect 12070 13022 12122 13074
rect 1710 12854 1762 12906
rect 2102 12898 2154 12950
rect 2662 12910 2714 12962
rect 4230 12854 4282 12906
rect 5406 12854 5458 12906
rect 6246 12910 6298 12962
rect 7926 12966 7978 13018
rect 8262 12966 8314 13018
rect 10446 12966 10498 13018
rect 7030 12854 7082 12906
rect 9662 12854 9714 12906
rect 10950 12910 11002 12962
rect 11398 12910 11450 12962
rect 11958 12910 12010 12962
rect 13302 12918 13354 12970
rect 10110 12854 10162 12906
rect 12630 12854 12682 12906
rect 13974 12898 14026 12950
rect 14646 12910 14698 12962
rect 14982 12909 15034 12961
rect 15990 12910 16042 12962
rect 16158 12966 16210 13018
rect 16606 13022 16658 13074
rect 20470 13078 20522 13130
rect 21030 13078 21082 13130
rect 22598 13134 22650 13186
rect 21646 13078 21698 13130
rect 23830 13078 23882 13130
rect 24166 13078 24218 13130
rect 16382 12910 16434 12962
rect 17446 12928 17498 12980
rect 18286 12966 18338 13018
rect 18510 12966 18562 13018
rect 19182 12966 19234 13018
rect 19742 12966 19794 13018
rect 20134 12966 20186 13018
rect 21758 12966 21810 13018
rect 17782 12854 17834 12906
rect 18006 12898 18058 12950
rect 21366 12910 21418 12962
rect 22262 12922 22314 12974
rect 8598 12742 8650 12794
rect 9886 12742 9938 12794
rect 11510 12742 11562 12794
rect 13022 12742 13074 12794
rect 13358 12742 13410 12794
rect 14534 12798 14586 12850
rect 20694 12854 20746 12906
rect 22486 12898 22538 12950
rect 22822 12922 22874 12974
rect 30214 12966 30266 13018
rect 30494 12966 30546 13018
rect 18342 12798 18394 12850
rect 22990 12854 23042 12906
rect 23270 12910 23322 12962
rect 24502 12898 24554 12950
rect 25622 12910 25674 12962
rect 24782 12854 24834 12906
rect 27190 12910 27242 12962
rect 26126 12854 26178 12906
rect 26854 12854 26906 12906
rect 27302 12804 27354 12856
rect 28030 12854 28082 12906
rect 28534 12910 28586 12962
rect 29374 12854 29426 12906
rect 13638 12742 13690 12794
rect 16102 12742 16154 12794
rect 19406 12742 19458 12794
rect 23550 12686 23602 12738
rect 23774 12686 23826 12738
rect 27582 12742 27634 12794
rect 27918 12742 27970 12794
rect 30774 12781 30826 12833
rect 4960 12518 5012 12570
rect 5064 12518 5116 12570
rect 5168 12518 5220 12570
rect 12900 12518 12952 12570
rect 13004 12518 13056 12570
rect 13108 12518 13160 12570
rect 20840 12518 20892 12570
rect 20944 12518 20996 12570
rect 21048 12518 21100 12570
rect 28780 12518 28832 12570
rect 28884 12518 28936 12570
rect 28988 12518 29040 12570
rect 7198 12294 7250 12346
rect 17334 12294 17386 12346
rect 1598 12182 1650 12234
rect 2326 12182 2378 12234
rect 3166 12182 3218 12234
rect 4006 12126 4058 12178
rect 4230 12182 4282 12234
rect 11174 12238 11226 12290
rect 20358 12294 20410 12346
rect 5854 12182 5906 12234
rect 18230 12238 18282 12290
rect 22206 12294 22258 12346
rect 22318 12294 22370 12346
rect 23606 12294 23658 12346
rect 24558 12294 24610 12346
rect 26854 12294 26906 12346
rect 32006 12294 32058 12346
rect 12518 12182 12570 12234
rect 13414 12182 13466 12234
rect 4566 12108 4618 12160
rect 6246 12070 6298 12122
rect 8822 12108 8874 12160
rect 9494 12126 9546 12178
rect 11622 12126 11674 12178
rect 12182 12108 12234 12160
rect 13750 12126 13802 12178
rect 6470 12024 6522 12076
rect 14366 12070 14418 12122
rect 15094 12114 15146 12166
rect 15318 12114 15370 12166
rect 15654 12114 15706 12166
rect 15878 12114 15930 12166
rect 16214 12114 16266 12166
rect 16438 12114 16490 12166
rect 17054 12126 17106 12178
rect 1374 11958 1426 12010
rect 2158 11958 2210 12010
rect 5518 11958 5570 12010
rect 7086 11958 7138 12010
rect 11734 12014 11786 12066
rect 16718 12070 16770 12122
rect 16886 12070 16938 12122
rect 20750 12182 20802 12234
rect 17950 12126 18002 12178
rect 19014 12126 19066 12178
rect 19350 12126 19402 12178
rect 23046 12138 23098 12190
rect 27470 12182 27522 12234
rect 18510 12070 18562 12122
rect 20022 12070 20074 12122
rect 20638 12070 20690 12122
rect 22766 12070 22818 12122
rect 23382 12114 23434 12166
rect 25062 12126 25114 12178
rect 30774 12182 30826 12234
rect 23942 12070 23994 12122
rect 24502 12070 24554 12122
rect 26630 12070 26682 12122
rect 27190 12108 27242 12160
rect 28310 12070 28362 12122
rect 28646 12108 28698 12160
rect 29206 12126 29258 12178
rect 30046 12070 30098 12122
rect 32342 12108 32394 12160
rect 9158 11958 9210 12010
rect 12798 11958 12850 12010
rect 17670 11958 17722 12010
rect 15430 11876 15482 11928
rect 16102 11902 16154 11954
rect 18286 11902 18338 11954
rect 19014 11958 19066 12010
rect 21534 11958 21586 12010
rect 21926 11958 21978 12010
rect 24670 11958 24722 12010
rect 25790 11958 25842 12010
rect 31838 11958 31890 12010
rect 23158 11876 23210 11928
rect 8930 11734 8982 11786
rect 9034 11734 9086 11786
rect 9138 11734 9190 11786
rect 16870 11734 16922 11786
rect 16974 11734 17026 11786
rect 17078 11734 17130 11786
rect 24810 11734 24862 11786
rect 24914 11734 24966 11786
rect 25018 11734 25070 11786
rect 2214 11510 2266 11562
rect 3278 11510 3330 11562
rect 6246 11535 6298 11587
rect 8150 11510 8202 11562
rect 9326 11510 9378 11562
rect 9662 11510 9714 11562
rect 10110 11510 10162 11562
rect 10558 11510 10610 11562
rect 10950 11510 11002 11562
rect 12686 11510 12738 11562
rect 16438 11510 16490 11562
rect 17390 11510 17442 11562
rect 17502 11510 17554 11562
rect 18006 11510 18058 11562
rect 19686 11535 19738 11587
rect 1878 11360 1930 11412
rect 2662 11342 2714 11394
rect 4454 11361 4506 11413
rect 5798 11342 5850 11394
rect 6806 11342 6858 11394
rect 7142 11348 7194 11400
rect 9886 11398 9938 11450
rect 11398 11420 11450 11472
rect 8262 11342 8314 11394
rect 11846 11398 11898 11450
rect 13414 11444 13466 11496
rect 11230 11342 11282 11394
rect 1598 11286 1650 11338
rect 4118 11286 4170 11338
rect 6022 11286 6074 11338
rect 8038 11286 8090 11338
rect 13750 11398 13802 11450
rect 12014 11342 12066 11394
rect 12966 11342 13018 11394
rect 15038 11398 15090 11450
rect 15430 11398 15482 11450
rect 15654 11342 15706 11394
rect 11398 11286 11450 11338
rect 17782 11339 17834 11391
rect 24054 11398 24106 11450
rect 18062 11342 18114 11394
rect 19238 11342 19290 11394
rect 18790 11286 18842 11338
rect 21142 11330 21194 11382
rect 21758 11342 21810 11394
rect 25286 11398 25338 11450
rect 26854 11398 26906 11450
rect 27302 11361 27354 11413
rect 24726 11286 24778 11338
rect 7478 11230 7530 11282
rect 4510 11174 4562 11226
rect 10222 11174 10274 11226
rect 11902 11174 11954 11226
rect 12574 11174 12626 11226
rect 14142 11118 14194 11170
rect 14478 11174 14530 11226
rect 14926 11174 14978 11226
rect 26574 11230 26626 11282
rect 27414 11236 27466 11288
rect 18286 11118 18338 11170
rect 4960 10950 5012 11002
rect 5064 10950 5116 11002
rect 5168 10950 5220 11002
rect 12900 10950 12952 11002
rect 13004 10950 13056 11002
rect 13108 10950 13160 11002
rect 20840 10950 20892 11002
rect 20944 10950 20996 11002
rect 21048 10950 21100 11002
rect 28780 10950 28832 11002
rect 28884 10950 28936 11002
rect 28988 10950 29040 11002
rect 8934 10726 8986 10778
rect 9438 10726 9490 10778
rect 9662 10782 9714 10834
rect 10782 10726 10834 10778
rect 10166 10668 10218 10720
rect 16942 10782 16994 10834
rect 12014 10726 12066 10778
rect 15766 10726 15818 10778
rect 23998 10726 24050 10778
rect 12854 10670 12906 10722
rect 13750 10670 13802 10722
rect 14310 10670 14362 10722
rect 24558 10726 24610 10778
rect 25342 10726 25394 10778
rect 1430 10558 1482 10610
rect 2270 10614 2322 10666
rect 4230 10614 4282 10666
rect 2998 10502 3050 10554
rect 3558 10535 3610 10587
rect 5462 10546 5514 10598
rect 5910 10546 5962 10598
rect 9942 10570 9994 10622
rect 11398 10614 11450 10666
rect 19798 10614 19850 10666
rect 20750 10614 20802 10666
rect 8262 10502 8314 10554
rect 10334 10558 10386 10610
rect 12294 10544 12346 10596
rect 11398 10480 11450 10532
rect 4846 10390 4898 10442
rect 9102 10390 9154 10442
rect 10110 10334 10162 10386
rect 10894 10390 10946 10442
rect 11230 10390 11282 10442
rect 11902 10446 11954 10498
rect 12574 10502 12626 10554
rect 13582 10558 13634 10610
rect 13358 10502 13410 10554
rect 14422 10558 14474 10610
rect 13806 10502 13858 10554
rect 15710 10502 15762 10554
rect 16102 10502 16154 10554
rect 17334 10502 17386 10554
rect 18230 10502 18282 10554
rect 19014 10540 19066 10592
rect 20022 10558 20074 10610
rect 21366 10570 21418 10622
rect 21870 10614 21922 10666
rect 12798 10390 12850 10442
rect 17502 10446 17554 10498
rect 24110 10502 24162 10554
rect 24894 10502 24946 10554
rect 25454 10502 25506 10554
rect 25846 10502 25898 10554
rect 27302 10502 27354 10554
rect 28086 10540 28138 10592
rect 14758 10334 14810 10386
rect 15486 10334 15538 10386
rect 16606 10390 16658 10442
rect 18622 10390 18674 10442
rect 19350 10390 19402 10442
rect 21702 10390 21754 10442
rect 23550 10390 23602 10442
rect 24446 10390 24498 10442
rect 25006 10390 25058 10442
rect 27134 10334 27186 10386
rect 27750 10390 27802 10442
rect 8930 10166 8982 10218
rect 9034 10166 9086 10218
rect 9138 10166 9190 10218
rect 16870 10166 16922 10218
rect 16974 10166 17026 10218
rect 17078 10166 17130 10218
rect 24810 10166 24862 10218
rect 24914 10166 24966 10218
rect 25018 10166 25070 10218
rect 6470 10024 6522 10076
rect 3054 9942 3106 9994
rect 4062 9942 4114 9994
rect 4902 9942 4954 9994
rect 5574 9830 5626 9882
rect 5910 9830 5962 9882
rect 1542 9762 1594 9814
rect 2550 9774 2602 9826
rect 6190 9830 6242 9882
rect 8094 9886 8146 9938
rect 8710 9942 8762 9994
rect 9662 9998 9714 10050
rect 12854 9942 12906 9994
rect 13526 9942 13578 9994
rect 14926 9998 14978 10050
rect 6750 9830 6802 9882
rect 7198 9830 7250 9882
rect 7422 9830 7474 9882
rect 7758 9830 7810 9882
rect 3894 9718 3946 9770
rect 4566 9762 4618 9814
rect 5070 9718 5122 9770
rect 6470 9762 6522 9814
rect 8318 9774 8370 9826
rect 9438 9830 9490 9882
rect 10054 9830 10106 9882
rect 11510 9830 11562 9882
rect 12070 9852 12122 9904
rect 11902 9774 11954 9826
rect 12518 9830 12570 9882
rect 13694 9774 13746 9826
rect 14086 9803 14138 9855
rect 14702 9830 14754 9882
rect 15150 9886 15202 9938
rect 16046 9942 16098 9994
rect 15430 9830 15482 9882
rect 12070 9718 12122 9770
rect 14534 9754 14586 9806
rect 15822 9774 15874 9826
rect 16550 9792 16602 9844
rect 20358 9830 20410 9882
rect 16886 9718 16938 9770
rect 17446 9762 17498 9814
rect 18006 9762 18058 9814
rect 21366 9786 21418 9838
rect 21814 9786 21866 9838
rect 24166 9830 24218 9882
rect 21030 9718 21082 9770
rect 24838 9718 24890 9770
rect 25230 9718 25282 9770
rect 25958 9774 26010 9826
rect 25454 9718 25506 9770
rect 26574 9718 26626 9770
rect 27302 9718 27354 9770
rect 27806 9718 27858 9770
rect 1878 9606 1930 9658
rect 9606 9606 9658 9658
rect 11174 9606 11226 9658
rect 13470 9550 13522 9602
rect 13918 9606 13970 9658
rect 14646 9606 14698 9658
rect 15878 9606 15930 9658
rect 27694 9606 27746 9658
rect 4960 9382 5012 9434
rect 5064 9382 5116 9434
rect 5168 9382 5220 9434
rect 12900 9382 12952 9434
rect 13004 9382 13056 9434
rect 13108 9382 13160 9434
rect 20840 9382 20892 9434
rect 20944 9382 20996 9434
rect 21048 9382 21100 9434
rect 28780 9382 28832 9434
rect 28884 9382 28936 9434
rect 28988 9382 29040 9434
rect 4118 9158 4170 9210
rect 7590 9158 7642 9210
rect 10054 9158 10106 9210
rect 10278 9158 10330 9210
rect 10502 9158 10554 9210
rect 13582 9214 13634 9266
rect 1486 9046 1538 9098
rect 1598 8934 1650 8986
rect 1878 8990 1930 9042
rect 2718 9046 2770 9098
rect 3446 9046 3498 9098
rect 3726 9046 3778 9098
rect 4734 9046 4786 9098
rect 11734 9108 11786 9160
rect 11902 9158 11954 9210
rect 12630 9158 12682 9210
rect 19350 9158 19402 9210
rect 19630 9158 19682 9210
rect 20358 9158 20410 9210
rect 22262 9158 22314 9210
rect 6134 9046 6186 9098
rect 4510 8934 4562 8986
rect 5462 8967 5514 9019
rect 8766 8990 8818 9042
rect 13974 9046 14026 9098
rect 21590 9096 21642 9148
rect 23494 9158 23546 9210
rect 32006 9158 32058 9210
rect 7534 8934 7586 8986
rect 7926 8934 7978 8986
rect 8150 8934 8202 8986
rect 11622 8982 11674 9034
rect 14422 9002 14474 9054
rect 14646 9002 14698 9054
rect 14982 9002 15034 9054
rect 12182 8934 12234 8986
rect 12574 8934 12626 8986
rect 12798 8934 12850 8986
rect 13358 8934 13410 8986
rect 15878 8978 15930 9030
rect 16270 8990 16322 9042
rect 19966 8934 20018 8986
rect 20694 8972 20746 9024
rect 21422 8934 21474 8986
rect 21702 8982 21754 9034
rect 23158 9002 23210 9054
rect 26070 8990 26122 9042
rect 26910 9046 26962 9098
rect 27638 9046 27690 9098
rect 24166 8934 24218 8986
rect 25734 8934 25786 8986
rect 32342 8972 32394 9024
rect 7310 8766 7362 8818
rect 8542 8766 8594 8818
rect 8654 8822 8706 8874
rect 9102 8822 9154 8874
rect 9214 8822 9266 8874
rect 9774 8822 9826 8874
rect 10838 8822 10890 8874
rect 18678 8822 18730 8874
rect 19742 8822 19794 8874
rect 14758 8766 14810 8818
rect 22654 8822 22706 8874
rect 25454 8766 25506 8818
rect 31838 8822 31890 8874
rect 8930 8598 8982 8650
rect 9034 8598 9086 8650
rect 9138 8598 9190 8650
rect 16870 8598 16922 8650
rect 16974 8598 17026 8650
rect 17078 8598 17130 8650
rect 24810 8598 24862 8650
rect 24914 8598 24966 8650
rect 25018 8598 25070 8650
rect 8374 8456 8426 8508
rect 1486 8374 1538 8426
rect 3222 8374 3274 8426
rect 6358 8399 6410 8451
rect 17278 8374 17330 8426
rect 18902 8374 18954 8426
rect 20526 8374 20578 8426
rect 20974 8374 21026 8426
rect 24054 8374 24106 8426
rect 4006 8262 4058 8314
rect 4734 8262 4786 8314
rect 2438 8206 2490 8258
rect 3782 8206 3834 8258
rect 4958 8262 5010 8314
rect 7422 8262 7474 8314
rect 5910 8206 5962 8258
rect 7030 8206 7082 8258
rect 8150 8218 8202 8270
rect 5462 8150 5514 8202
rect 6638 8150 6690 8202
rect 8486 8194 8538 8246
rect 8710 8194 8762 8246
rect 9382 8218 9434 8270
rect 12294 8262 12346 8314
rect 16214 8262 16266 8314
rect 9942 8194 9994 8246
rect 1990 8094 2042 8146
rect 12966 8150 13018 8202
rect 13302 8194 13354 8246
rect 13806 8206 13858 8258
rect 17558 8262 17610 8314
rect 17950 8262 18002 8314
rect 18622 8262 18674 8314
rect 19294 8262 19346 8314
rect 19742 8262 19794 8314
rect 22038 8318 22090 8370
rect 19966 8262 20018 8314
rect 24334 8262 24386 8314
rect 20806 8206 20858 8258
rect 22374 8206 22426 8258
rect 25286 8262 25338 8314
rect 26574 8262 26626 8314
rect 26742 8262 26794 8314
rect 16886 8150 16938 8202
rect 23718 8194 23770 8246
rect 24614 8198 24666 8250
rect 4342 8038 4394 8090
rect 7086 8038 7138 8090
rect 18230 8038 18282 8090
rect 19630 8038 19682 8090
rect 24502 8100 24554 8152
rect 20414 8038 20466 8090
rect 4960 7814 5012 7866
rect 5064 7814 5116 7866
rect 5168 7814 5220 7866
rect 12900 7814 12952 7866
rect 13004 7814 13056 7866
rect 13108 7814 13160 7866
rect 20840 7814 20892 7866
rect 20944 7814 20996 7866
rect 21048 7814 21100 7866
rect 28780 7814 28832 7866
rect 28884 7814 28936 7866
rect 28988 7814 29040 7866
rect 3110 7590 3162 7642
rect 6862 7590 6914 7642
rect 8934 7590 8986 7642
rect 11622 7590 11674 7642
rect 13750 7590 13802 7642
rect 15430 7590 15482 7642
rect 16102 7590 16154 7642
rect 17446 7590 17498 7642
rect 2998 7478 3050 7530
rect 3782 7422 3834 7474
rect 4062 7422 4114 7474
rect 2550 7366 2602 7418
rect 4286 7422 4338 7474
rect 5686 7434 5738 7486
rect 6022 7478 6074 7530
rect 6358 7404 6410 7456
rect 8598 7434 8650 7486
rect 12518 7478 12570 7530
rect 16886 7528 16938 7580
rect 18174 7590 18226 7642
rect 18510 7590 18562 7642
rect 19574 7590 19626 7642
rect 20246 7590 20298 7642
rect 21926 7540 21978 7592
rect 22766 7590 22818 7642
rect 25118 7534 25170 7586
rect 6806 7366 6858 7418
rect 8038 7366 8090 7418
rect 9494 7404 9546 7456
rect 10502 7366 10554 7418
rect 11062 7404 11114 7456
rect 11958 7404 12010 7456
rect 13414 7434 13466 7486
rect 12518 7344 12570 7396
rect 12798 7366 12850 7418
rect 14422 7404 14474 7456
rect 15094 7434 15146 7486
rect 17782 7434 17834 7486
rect 22430 7478 22482 7530
rect 25790 7534 25842 7586
rect 26126 7478 26178 7530
rect 15710 7366 15762 7418
rect 18118 7422 18170 7474
rect 17166 7366 17218 7418
rect 18846 7366 18898 7418
rect 19238 7404 19290 7456
rect 21702 7422 21754 7474
rect 22094 7366 22146 7418
rect 23382 7404 23434 7456
rect 23942 7366 23994 7418
rect 25398 7366 25450 7418
rect 1486 7254 1538 7306
rect 1598 7254 1650 7306
rect 3222 7254 3274 7306
rect 4678 7254 4730 7306
rect 4958 7254 5010 7306
rect 5350 7254 5402 7306
rect 6974 7254 7026 7306
rect 7422 7254 7474 7306
rect 7646 7254 7698 7306
rect 7870 7254 7922 7306
rect 8206 7254 8258 7306
rect 9158 7254 9210 7306
rect 9774 7254 9826 7306
rect 10334 7254 10386 7306
rect 10670 7254 10722 7306
rect 11398 7254 11450 7306
rect 12350 7254 12402 7306
rect 13918 7254 13970 7306
rect 14758 7254 14810 7306
rect 16942 7254 16994 7306
rect 19854 7254 19906 7306
rect 23046 7254 23098 7306
rect 8930 7030 8982 7082
rect 9034 7030 9086 7082
rect 9138 7030 9190 7082
rect 16870 7030 16922 7082
rect 16974 7030 17026 7082
rect 17078 7030 17130 7082
rect 24810 7030 24862 7082
rect 24914 7030 24966 7082
rect 25018 7030 25070 7082
rect 2830 6806 2882 6858
rect 7254 6831 7306 6883
rect 11902 6862 11954 6914
rect 12630 6862 12682 6914
rect 15990 6806 16042 6858
rect 16830 6806 16882 6858
rect 5462 6750 5514 6802
rect 6246 6750 6298 6802
rect 19294 6806 19346 6858
rect 23158 6806 23210 6858
rect 24334 6806 24386 6858
rect 4566 6694 4618 6746
rect 6694 6694 6746 6746
rect 6862 6694 6914 6746
rect 11286 6694 11338 6746
rect 11678 6694 11730 6746
rect 1542 6626 1594 6678
rect 1878 6582 1930 6634
rect 2270 6582 2322 6634
rect 3446 6626 3498 6678
rect 5238 6638 5290 6690
rect 6134 6638 6186 6690
rect 7702 6638 7754 6690
rect 3726 6582 3778 6634
rect 8150 6582 8202 6634
rect 8822 6626 8874 6678
rect 9942 6626 9994 6678
rect 10334 6582 10386 6634
rect 10950 6630 11002 6682
rect 12294 6626 12346 6678
rect 12518 6626 12570 6678
rect 12854 6626 12906 6678
rect 13078 6650 13130 6702
rect 13638 6626 13690 6678
rect 17894 6656 17946 6708
rect 18678 6656 18730 6708
rect 20246 6650 20298 6702
rect 24110 6694 24162 6746
rect 2494 6470 2546 6522
rect 5686 6526 5738 6578
rect 3110 6470 3162 6522
rect 6750 6470 6802 6522
rect 8486 6470 8538 6522
rect 9606 6470 9658 6522
rect 10838 6532 10890 6584
rect 18230 6582 18282 6634
rect 20862 6638 20914 6690
rect 24558 6638 24610 6690
rect 19686 6582 19738 6634
rect 24726 6618 24778 6670
rect 25286 6638 25338 6690
rect 26294 6630 26346 6682
rect 26966 6626 27018 6678
rect 10670 6470 10722 6522
rect 11622 6470 11674 6522
rect 16662 6470 16714 6522
rect 19014 6470 19066 6522
rect 25398 6532 25450 6584
rect 23830 6470 23882 6522
rect 24054 6470 24106 6522
rect 25678 6470 25730 6522
rect 26182 6532 26234 6584
rect 26014 6470 26066 6522
rect 26630 6470 26682 6522
rect 4960 6246 5012 6298
rect 5064 6246 5116 6298
rect 5168 6246 5220 6298
rect 12900 6246 12952 6298
rect 13004 6246 13056 6298
rect 13108 6246 13160 6298
rect 20840 6246 20892 6298
rect 20944 6246 20996 6298
rect 21048 6246 21100 6298
rect 28780 6246 28832 6298
rect 28884 6246 28936 6298
rect 28988 6246 29040 6298
rect 2326 6022 2378 6074
rect 4734 6022 4786 6074
rect 5854 6022 5906 6074
rect 6414 6022 6466 6074
rect 12070 6022 12122 6074
rect 12854 6022 12906 6074
rect 14310 6022 14362 6074
rect 18566 6022 18618 6074
rect 21254 6022 21306 6074
rect 22038 6022 22090 6074
rect 2774 5866 2826 5918
rect 3726 5910 3778 5962
rect 3950 5910 4002 5962
rect 1990 5798 2042 5850
rect 3110 5842 3162 5894
rect 3334 5842 3386 5894
rect 4342 5854 4394 5906
rect 7198 5854 7250 5906
rect 7422 5910 7474 5962
rect 4118 5750 4170 5802
rect 6190 5798 6242 5850
rect 7590 5840 7642 5892
rect 8598 5866 8650 5918
rect 9046 5866 9098 5918
rect 12518 5866 12570 5918
rect 8038 5798 8090 5850
rect 11398 5798 11450 5850
rect 13526 5836 13578 5888
rect 14982 5866 15034 5918
rect 20414 5910 20466 5962
rect 26462 5910 26514 5962
rect 13862 5798 13914 5850
rect 14646 5798 14698 5850
rect 15542 5842 15594 5894
rect 17894 5798 17946 5850
rect 18790 5798 18842 5850
rect 19182 5798 19234 5850
rect 19686 5798 19738 5850
rect 21590 5836 21642 5888
rect 22710 5798 22762 5850
rect 25062 5842 25114 5894
rect 25510 5842 25562 5894
rect 25846 5798 25898 5850
rect 1486 5686 1538 5738
rect 1598 5686 1650 5738
rect 2270 5630 2322 5682
rect 2494 5686 2546 5738
rect 4846 5686 4898 5738
rect 2998 5630 3050 5682
rect 5406 5686 5458 5738
rect 5518 5686 5570 5738
rect 7142 5686 7194 5738
rect 7870 5686 7922 5738
rect 8206 5686 8258 5738
rect 14142 5686 14194 5738
rect 20022 5686 20074 5738
rect 26238 5686 26290 5738
rect 14366 5630 14418 5682
rect 8930 5462 8982 5514
rect 9034 5462 9086 5514
rect 9138 5462 9190 5514
rect 16870 5462 16922 5514
rect 16974 5462 17026 5514
rect 17078 5462 17130 5514
rect 24810 5462 24862 5514
rect 24914 5462 24966 5514
rect 25018 5462 25070 5514
rect 2158 5294 2210 5346
rect 3334 5238 3386 5290
rect 5294 5238 5346 5290
rect 15374 5294 15426 5346
rect 5854 5238 5906 5290
rect 6918 5238 6970 5290
rect 8486 5238 8538 5290
rect 1990 5090 2042 5142
rect 2382 5070 2434 5122
rect 3446 5084 3498 5136
rect 3838 5126 3890 5178
rect 4510 5126 4562 5178
rect 7086 5126 7138 5178
rect 7310 5126 7362 5178
rect 7702 5126 7754 5178
rect 8262 5070 8314 5122
rect 9830 5082 9882 5134
rect 12742 5126 12794 5178
rect 14534 5126 14586 5178
rect 14758 5172 14810 5224
rect 15598 5126 15650 5178
rect 16606 5126 16658 5178
rect 10390 5058 10442 5110
rect 15878 5058 15930 5110
rect 16046 5070 16098 5122
rect 16382 5070 16434 5122
rect 17726 5126 17778 5178
rect 17334 5070 17386 5122
rect 18174 5126 18226 5178
rect 19966 5182 20018 5234
rect 20582 5238 20634 5290
rect 21198 5182 21250 5234
rect 22822 5186 22874 5238
rect 18454 5078 18506 5130
rect 21366 5126 21418 5178
rect 18790 5070 18842 5122
rect 23046 5126 23098 5178
rect 24726 5126 24778 5178
rect 26014 5126 26066 5178
rect 26238 5126 26290 5178
rect 25622 5058 25674 5110
rect 1486 4902 1538 4954
rect 2214 4948 2266 5000
rect 1710 4846 1762 4898
rect 3054 4902 3106 4954
rect 3278 4902 3330 4954
rect 4174 4902 4226 4954
rect 4734 4902 4786 4954
rect 5070 4902 5122 4954
rect 5350 4952 5402 5004
rect 5910 4952 5962 5004
rect 6078 4902 6130 4954
rect 6526 4902 6578 4954
rect 6750 4902 6802 4954
rect 13414 4902 13466 4954
rect 13806 4902 13858 4954
rect 15654 4958 15706 5010
rect 16662 4958 16714 5010
rect 14142 4902 14194 4954
rect 17446 4952 17498 5004
rect 18342 4952 18394 5004
rect 18902 4964 18954 5016
rect 19182 4902 19234 4954
rect 19518 4902 19570 4954
rect 19630 4902 19682 4954
rect 20190 4846 20242 4898
rect 21758 4902 21810 4954
rect 22094 4902 22146 4954
rect 23438 4958 23490 5010
rect 31838 5014 31890 5066
rect 32342 5058 32394 5110
rect 23774 4902 23826 4954
rect 24390 4902 24442 4954
rect 25286 4902 25338 4954
rect 26182 4952 26234 5004
rect 32006 4902 32058 4954
rect 4960 4678 5012 4730
rect 5064 4678 5116 4730
rect 5168 4678 5220 4730
rect 12900 4678 12952 4730
rect 13004 4678 13056 4730
rect 13108 4678 13160 4730
rect 20840 4678 20892 4730
rect 20944 4678 20996 4730
rect 21048 4678 21100 4730
rect 28780 4678 28832 4730
rect 28884 4678 28936 4730
rect 28988 4678 29040 4730
rect 4006 4490 4058 4542
rect 2214 4408 2266 4460
rect 2886 4404 2938 4456
rect 5742 4454 5794 4506
rect 6862 4510 6914 4562
rect 6246 4404 6298 4456
rect 10390 4454 10442 4506
rect 11342 4454 11394 4506
rect 12014 4454 12066 4506
rect 12126 4454 12178 4506
rect 1710 4286 1762 4338
rect 1934 4342 1986 4394
rect 1486 4230 1538 4282
rect 2774 4286 2826 4338
rect 3782 4298 3834 4350
rect 2158 4230 2210 4282
rect 3166 4230 3218 4282
rect 4118 4274 4170 4326
rect 4846 4286 4898 4338
rect 7086 4342 7138 4394
rect 12518 4404 12570 4456
rect 12798 4454 12850 4506
rect 19742 4454 19794 4506
rect 21590 4454 21642 4506
rect 7254 4306 7306 4358
rect 7646 4342 7698 4394
rect 7926 4342 7978 4394
rect 3502 4174 3554 4226
rect 4510 4230 4562 4282
rect 4678 4230 4730 4282
rect 5406 4230 5458 4282
rect 8262 4286 8314 4338
rect 6414 4230 6466 4282
rect 9382 4268 9434 4320
rect 10054 4298 10106 4350
rect 10950 4294 11002 4346
rect 11286 4286 11338 4338
rect 10670 4230 10722 4282
rect 12406 4286 12458 4338
rect 14534 4298 14586 4350
rect 14702 4342 14754 4394
rect 11678 4230 11730 4282
rect 13246 4230 13298 4282
rect 13414 4230 13466 4282
rect 13918 4230 13970 4282
rect 14142 4230 14194 4282
rect 15094 4274 15146 4326
rect 15318 4298 15370 4350
rect 19462 4342 19514 4394
rect 15654 4274 15706 4326
rect 15878 4274 15930 4326
rect 16438 4274 16490 4326
rect 20022 4294 20074 4346
rect 20694 4298 20746 4350
rect 21198 4342 21250 4394
rect 24614 4298 24666 4350
rect 25174 4274 25226 4326
rect 25790 4230 25842 4282
rect 4230 4118 4282 4170
rect 5630 4118 5682 4170
rect 2382 4062 2434 4114
rect 6190 4118 6242 4170
rect 6806 4118 6858 4170
rect 9718 4118 9770 4170
rect 10782 4118 10834 4170
rect 13582 4118 13634 4170
rect 18790 4118 18842 4170
rect 19854 4118 19906 4170
rect 20358 4118 20410 4170
rect 22262 4118 22314 4170
rect 25398 4118 25450 4170
rect 26014 4118 26066 4170
rect 14310 4036 14362 4088
rect 15430 4036 15482 4088
rect 8930 3894 8982 3946
rect 9034 3894 9086 3946
rect 9138 3894 9190 3946
rect 16870 3894 16922 3946
rect 16974 3894 17026 3946
rect 17078 3894 17130 3946
rect 24810 3894 24862 3946
rect 24914 3894 24966 3946
rect 25018 3894 25070 3946
rect 1878 3726 1930 3778
rect 7590 3752 7642 3804
rect 8374 3752 8426 3804
rect 2774 3670 2826 3722
rect 3334 3670 3386 3722
rect 4790 3670 4842 3722
rect 12350 3670 12402 3722
rect 15206 3726 15258 3778
rect 12742 3670 12794 3722
rect 14590 3670 14642 3722
rect 1542 3514 1594 3566
rect 1766 3514 1818 3566
rect 2102 3490 2154 3542
rect 2718 3502 2770 3554
rect 4342 3558 4394 3610
rect 5798 3558 5850 3610
rect 6078 3558 6130 3610
rect 2998 3502 3050 3554
rect 4118 3502 4170 3554
rect 5574 3502 5626 3554
rect 6694 3520 6746 3572
rect 7366 3514 7418 3566
rect 7870 3558 7922 3610
rect 6302 3446 6354 3498
rect 7030 3446 7082 3498
rect 7590 3490 7642 3542
rect 8150 3514 8202 3566
rect 8486 3490 8538 3542
rect 8710 3514 8762 3566
rect 9326 3558 9378 3610
rect 9494 3558 9546 3610
rect 9662 3558 9714 3610
rect 10334 3558 10386 3610
rect 9942 3502 9994 3554
rect 11510 3558 11562 3610
rect 11734 3604 11786 3656
rect 13470 3558 13522 3610
rect 14030 3614 14082 3666
rect 13078 3502 13130 3554
rect 13750 3502 13802 3554
rect 14198 3558 14250 3610
rect 15934 3614 15986 3666
rect 16550 3670 16602 3722
rect 25510 3695 25562 3747
rect 14982 3490 15034 3542
rect 15318 3514 15370 3566
rect 15542 3490 15594 3542
rect 16158 3502 16210 3554
rect 17334 3514 17386 3566
rect 17894 3514 17946 3566
rect 20246 3558 20298 3610
rect 21254 3514 21306 3566
rect 24054 3558 24106 3610
rect 21758 3502 21810 3554
rect 25846 3502 25898 3554
rect 10054 3396 10106 3448
rect 2494 3334 2546 3386
rect 10782 3334 10834 3386
rect 13190 3396 13242 3448
rect 20918 3446 20970 3498
rect 25622 3446 25674 3498
rect 11118 3334 11170 3386
rect 24726 3334 24778 3386
rect 4960 3110 5012 3162
rect 5064 3110 5116 3162
rect 5168 3110 5220 3162
rect 12900 3110 12952 3162
rect 13004 3110 13056 3162
rect 13108 3110 13160 3162
rect 20840 3110 20892 3162
rect 20944 3110 20996 3162
rect 21048 3110 21100 3162
rect 28780 3110 28832 3162
rect 28884 3110 28936 3162
rect 28988 3110 29040 3162
rect 20302 2886 20354 2938
rect 1486 2774 1538 2826
rect 2662 2774 2714 2826
rect 6358 2774 6410 2826
rect 7310 2774 7362 2826
rect 2438 2718 2490 2770
rect 4342 2718 4394 2770
rect 5910 2718 5962 2770
rect 8654 2774 8706 2826
rect 4678 2662 4730 2714
rect 4846 2662 4898 2714
rect 7422 2662 7474 2714
rect 7590 2712 7642 2764
rect 14198 2830 14250 2882
rect 24838 2886 24890 2938
rect 9158 2774 9210 2826
rect 15206 2774 15258 2826
rect 8878 2662 8930 2714
rect 2102 2494 2154 2546
rect 3222 2550 3274 2602
rect 7702 2606 7754 2658
rect 9830 2662 9882 2714
rect 12182 2706 12234 2758
rect 12742 2706 12794 2758
rect 14086 2718 14138 2770
rect 19630 2774 19682 2826
rect 18174 2718 18226 2770
rect 18678 2706 18730 2758
rect 20582 2726 20634 2778
rect 21254 2730 21306 2782
rect 21814 2730 21866 2782
rect 19406 2662 19458 2714
rect 25398 2700 25450 2752
rect 4510 2550 4562 2602
rect 5798 2494 5850 2546
rect 7198 2494 7250 2546
rect 8262 2550 8314 2602
rect 13246 2550 13298 2602
rect 13470 2550 13522 2602
rect 14870 2550 14922 2602
rect 15878 2550 15930 2602
rect 19014 2550 19066 2602
rect 19966 2550 20018 2602
rect 20414 2550 20466 2602
rect 24166 2550 24218 2602
rect 25062 2550 25114 2602
rect 25678 2550 25730 2602
rect 25902 2550 25954 2602
rect 8930 2326 8982 2378
rect 9034 2326 9086 2378
rect 9138 2326 9190 2378
rect 16870 2326 16922 2378
rect 16974 2326 17026 2378
rect 17078 2326 17130 2378
rect 24810 2326 24862 2378
rect 24914 2326 24966 2378
rect 25018 2326 25070 2378
rect 4006 2102 4058 2154
rect 4790 2102 4842 2154
rect 7702 2127 7754 2179
rect 2102 2046 2154 2098
rect 17278 2102 17330 2154
rect 6358 2046 6410 2098
rect 6918 2046 6970 2098
rect 23214 2102 23266 2154
rect 24334 2102 24386 2154
rect 32006 2102 32058 2154
rect 3334 1990 3386 2042
rect 4454 1990 4506 2042
rect 5574 1990 5626 2042
rect 12406 1990 12458 2042
rect 6134 1934 6186 1986
rect 7030 1934 7082 1986
rect 8150 1934 8202 1986
rect 2438 1878 2490 1930
rect 7926 1878 7978 1930
rect 9606 1922 9658 1974
rect 10110 1934 10162 1986
rect 16214 1990 16266 2042
rect 17950 1990 18002 2042
rect 13078 1878 13130 1930
rect 13302 1922 13354 1974
rect 13862 1922 13914 1974
rect 18342 1934 18394 1986
rect 18566 1946 18618 1998
rect 19126 1946 19178 1998
rect 21478 1990 21530 2042
rect 22766 1990 22818 2042
rect 22374 1934 22426 1986
rect 23102 1990 23154 2042
rect 23774 1990 23826 2042
rect 6694 1822 6746 1874
rect 22150 1878 22202 1930
rect 23382 1926 23434 1978
rect 24054 1926 24106 1978
rect 31838 1878 31890 1930
rect 32342 1922 32394 1974
rect 16886 1766 16938 1818
rect 18286 1766 18338 1818
rect 22486 1816 22538 1868
rect 23942 1816 23994 1868
rect 4960 1542 5012 1594
rect 5064 1542 5116 1594
rect 5168 1542 5220 1594
rect 12900 1542 12952 1594
rect 13004 1542 13056 1594
rect 13108 1542 13160 1594
rect 20840 1542 20892 1594
rect 20944 1542 20996 1594
rect 21048 1542 21100 1594
rect 28780 1542 28832 1594
rect 28884 1542 28936 1594
rect 28988 1542 29040 1594
rect 4342 1318 4394 1370
rect 6414 1318 6466 1370
rect 6750 1318 6802 1370
rect 6974 1318 7026 1370
rect 7310 1318 7362 1370
rect 7646 1318 7698 1370
rect 7870 1318 7922 1370
rect 8822 1318 8874 1370
rect 9718 1318 9770 1370
rect 10838 1318 10890 1370
rect 11230 1318 11282 1370
rect 11566 1374 11618 1426
rect 14086 1318 14138 1370
rect 14814 1318 14866 1370
rect 16438 1318 16490 1370
rect 17558 1318 17610 1370
rect 17782 1318 17834 1370
rect 18454 1318 18506 1370
rect 19126 1318 19178 1370
rect 20022 1318 20074 1370
rect 21758 1318 21810 1370
rect 22374 1318 22426 1370
rect 1542 1150 1594 1202
rect 4678 1132 4730 1184
rect 5798 1162 5850 1214
rect 8486 1162 8538 1214
rect 10054 1162 10106 1214
rect 13358 1206 13410 1258
rect 16606 1206 16658 1258
rect 21926 1256 21978 1308
rect 23494 1318 23546 1370
rect 25622 1318 25674 1370
rect 5518 1094 5570 1146
rect 6078 1094 6130 1146
rect 8094 1094 8146 1146
rect 10502 1132 10554 1184
rect 17222 1162 17274 1214
rect 18118 1162 18170 1214
rect 18790 1162 18842 1214
rect 21366 1162 21418 1214
rect 11958 1094 12010 1146
rect 13750 1094 13802 1146
rect 14478 1094 14530 1146
rect 12126 1038 12178 1090
rect 15206 1094 15258 1146
rect 15430 1048 15482 1100
rect 16046 1094 16098 1146
rect 20358 1094 20410 1146
rect 22038 1142 22090 1194
rect 22710 1162 22762 1214
rect 23158 1162 23210 1214
rect 25958 1132 26010 1184
rect 2550 982 2602 1034
rect 19518 982 19570 1034
rect 19742 982 19794 1034
rect 21030 982 21082 1034
rect 26238 982 26290 1034
rect 5798 900 5850 952
rect 8930 758 8982 810
rect 9034 758 9086 810
rect 9138 758 9190 810
rect 16870 758 16922 810
rect 16974 758 17026 810
rect 17078 758 17130 810
rect 24810 758 24862 810
rect 24914 758 24966 810
rect 25018 758 25070 810
rect 20134 534 20186 586
rect 21030 534 21082 586
<< metal2 >>
rect 1176 19200 1288 20000
rect 3752 19200 3864 20000
rect 6328 19200 6440 20000
rect 9016 19200 9128 20000
rect 11592 19200 11704 20000
rect 14168 19200 14280 20000
rect 16856 19200 16968 20000
rect 19432 19200 19544 20000
rect 22120 19200 22232 20000
rect 24696 19200 24808 20000
rect 27272 19200 27384 20000
rect 29960 19200 30072 20000
rect 32536 19200 32648 20000
rect 1204 18508 1260 19200
rect 1204 18442 1260 18452
rect 1428 19068 1484 19078
rect 1428 18396 1484 19012
rect 1876 18620 1932 18630
rect 1876 18526 1932 18564
rect 1540 18508 1596 18518
rect 1540 18410 1542 18452
rect 1594 18410 1596 18452
rect 3388 18508 3444 18518
rect 3388 18414 3444 18452
rect 1540 18398 1596 18410
rect 1428 17846 1484 18340
rect 2940 18396 2996 18406
rect 3780 18396 3836 19200
rect 4958 18844 5222 18854
rect 5014 18788 5062 18844
rect 5118 18788 5166 18844
rect 4958 18778 5222 18788
rect 6076 18508 6132 18518
rect 6356 18508 6412 19200
rect 6916 18620 6972 18630
rect 6916 18618 7420 18620
rect 6916 18566 6918 18618
rect 6970 18566 7420 18618
rect 6916 18564 7420 18566
rect 6916 18554 6972 18564
rect 6076 18506 6524 18508
rect 6076 18454 6078 18506
rect 6130 18454 6524 18506
rect 6076 18452 6524 18454
rect 6076 18442 6132 18452
rect 6468 18406 6524 18452
rect 7140 18450 7196 18462
rect 3892 18396 4004 18406
rect 3780 18340 3892 18396
rect 3948 18394 4004 18396
rect 3948 18342 3950 18394
rect 4002 18342 4004 18394
rect 3948 18340 4004 18342
rect 2940 18302 2996 18340
rect 3892 18330 4004 18340
rect 4508 18396 4564 18406
rect 6468 18394 6580 18406
rect 6468 18342 6526 18394
rect 6578 18342 6580 18394
rect 6468 18340 6580 18342
rect 1652 18284 1708 18294
rect 2156 18284 2212 18294
rect 1428 17834 1540 17846
rect 1428 17782 1486 17834
rect 1538 17782 1540 17834
rect 1428 17780 1540 17782
rect 1484 17770 1540 17780
rect 1652 17276 1708 18228
rect 2100 18282 2212 18284
rect 2100 18230 2158 18282
rect 2210 18230 2212 18282
rect 2100 18218 2212 18230
rect 2548 18282 2604 18294
rect 2548 18230 2550 18282
rect 2602 18230 2604 18282
rect 2100 18060 2156 18218
rect 2548 18172 2604 18230
rect 2716 18284 2772 18294
rect 2716 18190 2772 18228
rect 3164 18282 3220 18294
rect 3164 18230 3166 18282
rect 3218 18230 3220 18282
rect 3892 18264 3948 18330
rect 4508 18302 4564 18340
rect 6524 18330 6580 18340
rect 7140 18398 7142 18450
rect 7194 18398 7196 18450
rect 4340 18284 4396 18294
rect 2548 18106 2604 18116
rect 2100 17994 2156 18004
rect 3164 18060 3220 18230
rect 4340 18190 4396 18228
rect 6300 18284 6356 18294
rect 6300 18190 6356 18228
rect 3164 17994 3220 18004
rect 2660 17836 2716 17846
rect 2548 17780 2660 17836
rect 2548 17744 2604 17780
rect 2660 17770 2716 17780
rect 3724 17836 3780 17846
rect 2044 17724 2100 17734
rect 1540 17220 1708 17276
rect 1764 17722 2100 17724
rect 1764 17670 2046 17722
rect 2098 17670 2100 17722
rect 2548 17692 2550 17744
rect 2602 17692 2604 17744
rect 2548 17680 2604 17692
rect 1764 17668 2100 17670
rect 1540 16940 1596 17220
rect 1540 16842 1542 16884
rect 1594 16842 1596 16884
rect 1540 16808 1596 16842
rect 1428 16716 1484 16726
rect 1764 16716 1820 17668
rect 2044 17658 2100 17668
rect 2380 17666 2436 17678
rect 2380 17614 2382 17666
rect 2434 17614 2436 17666
rect 1876 17500 1932 17510
rect 1876 17406 1932 17444
rect 2380 17276 2436 17614
rect 2548 17612 2604 17622
rect 2548 17518 2604 17556
rect 3724 17612 3780 17780
rect 3724 17518 3780 17556
rect 5852 17836 5908 17846
rect 2940 17500 2996 17510
rect 1876 17220 2436 17276
rect 2660 17498 2996 17500
rect 2660 17446 2942 17498
rect 2994 17446 2996 17498
rect 2660 17444 2996 17446
rect 1876 17050 1932 17220
rect 1876 16998 1878 17050
rect 1930 16998 1932 17050
rect 1876 16986 1932 16998
rect 2660 16882 2716 17444
rect 2940 17434 2996 17444
rect 3052 17498 3108 17510
rect 3052 17446 3054 17498
rect 3106 17446 3108 17498
rect 3052 16940 3108 17446
rect 3388 17500 3444 17510
rect 3388 17406 3444 17444
rect 3500 17498 3556 17510
rect 3500 17446 3502 17498
rect 3554 17446 3556 17498
rect 3500 17052 3556 17446
rect 4958 17276 5222 17286
rect 5014 17220 5062 17276
rect 5118 17220 5166 17276
rect 4958 17210 5222 17220
rect 5852 17052 5908 17780
rect 7140 17836 7196 18398
rect 7140 17770 7196 17780
rect 6804 17724 6860 17734
rect 6804 17630 6860 17668
rect 6972 17666 7028 17678
rect 6412 17612 6468 17622
rect 6972 17614 6974 17666
rect 7026 17614 7028 17666
rect 6972 17612 7028 17614
rect 7252 17666 7308 17678
rect 7252 17614 7254 17666
rect 7306 17614 7308 17666
rect 7252 17612 7308 17614
rect 6972 17556 7196 17612
rect 6412 17518 6468 17556
rect 5964 17500 6020 17510
rect 5964 17406 6020 17444
rect 6300 17498 6356 17510
rect 6300 17446 6302 17498
rect 6354 17446 6356 17498
rect 6300 17276 6356 17446
rect 6300 17210 6356 17220
rect 6692 17500 6748 17510
rect 6020 17052 6076 17062
rect 5852 17050 6076 17052
rect 5852 16998 6022 17050
rect 6074 16998 6076 17050
rect 5852 16996 6076 16998
rect 3500 16986 3556 16996
rect 6020 16986 6076 16996
rect 6356 17052 6412 17062
rect 2660 16830 2662 16882
rect 2714 16830 2716 16882
rect 2660 16818 2716 16830
rect 2996 16884 3108 16940
rect 6356 16894 6412 16996
rect 1428 15158 1484 16660
rect 1540 16660 1820 16716
rect 2044 16716 2100 16726
rect 1540 16086 1596 16660
rect 2044 16622 2100 16660
rect 2996 16380 3052 16884
rect 6356 16842 6358 16894
rect 6410 16842 6412 16894
rect 3892 16828 3948 16838
rect 4284 16828 4340 16838
rect 6356 16830 6412 16842
rect 6692 16882 6748 17444
rect 6860 17500 6916 17510
rect 6860 17498 6972 17500
rect 6860 17446 6862 17498
rect 6914 17446 6972 17498
rect 6860 17434 6972 17446
rect 6916 17276 6972 17434
rect 6916 17210 6972 17220
rect 6692 16830 6694 16882
rect 6746 16830 6748 16882
rect 3892 16826 4340 16828
rect 3892 16774 3894 16826
rect 3946 16774 4286 16826
rect 4338 16774 4340 16826
rect 6692 16818 6748 16830
rect 3892 16772 4340 16774
rect 3164 16716 3220 16726
rect 3164 16622 3220 16660
rect 3724 16716 3780 16726
rect 2436 16324 3052 16380
rect 2436 16156 2492 16324
rect 1540 16034 1542 16086
rect 1594 16034 1596 16086
rect 1540 15596 1596 16034
rect 2380 16100 2492 16156
rect 2548 16156 2604 16166
rect 1876 15932 1932 15942
rect 1540 15530 1596 15540
rect 1764 15930 1932 15932
rect 1764 15878 1878 15930
rect 1930 15878 1932 15930
rect 1764 15876 1932 15878
rect 1428 15146 1540 15158
rect 1428 15094 1486 15146
rect 1538 15094 1540 15146
rect 1428 15082 1540 15094
rect 1428 15036 1484 15082
rect 1204 14980 1484 15036
rect 1204 14364 1260 14980
rect 1484 14588 1540 14598
rect 1204 14298 1260 14308
rect 1316 14586 1540 14588
rect 1316 14534 1486 14586
rect 1538 14534 1540 14586
rect 1316 14532 1540 14534
rect 1204 13468 1260 13478
rect 1204 11228 1260 13412
rect 1316 13132 1372 14532
rect 1484 14522 1540 14532
rect 1596 13692 1652 13702
rect 1484 13580 1540 13590
rect 1316 12236 1372 13076
rect 1316 12170 1372 12180
rect 1428 13578 1540 13580
rect 1428 13526 1486 13578
rect 1538 13526 1540 13578
rect 1428 13514 1540 13526
rect 1428 12022 1484 13514
rect 1596 13130 1652 13636
rect 1764 13244 1820 15876
rect 1876 15866 1932 15876
rect 2268 15820 2324 15830
rect 2268 15482 2324 15764
rect 2268 15430 2270 15482
rect 2322 15430 2324 15482
rect 2268 15418 2324 15430
rect 2380 15482 2436 16100
rect 2548 16065 2550 16100
rect 2602 16065 2604 16100
rect 2548 16053 2604 16065
rect 2996 16098 3052 16324
rect 3724 16266 3780 16660
rect 3724 16214 3726 16266
rect 3778 16214 3780 16266
rect 3724 16202 3780 16214
rect 2996 16046 2998 16098
rect 3050 16046 3052 16098
rect 2996 16034 3052 16046
rect 2492 15932 2548 15942
rect 2492 15930 3052 15932
rect 2492 15878 2494 15930
rect 2546 15878 3052 15930
rect 2492 15876 3052 15878
rect 2492 15866 2548 15876
rect 2380 15430 2382 15482
rect 2434 15430 2436 15482
rect 2380 15418 2436 15430
rect 2884 15372 2940 15410
rect 2884 15306 2940 15316
rect 2884 15236 2940 15248
rect 2884 15184 2886 15236
rect 2938 15184 2940 15236
rect 1876 15148 1932 15158
rect 2100 15148 2156 15158
rect 2716 15148 2772 15158
rect 1876 15146 2044 15148
rect 1876 15094 1878 15146
rect 1930 15094 2044 15146
rect 1876 15092 2044 15094
rect 1876 15082 1932 15092
rect 1876 14362 1932 14374
rect 1876 14310 1878 14362
rect 1930 14310 1932 14362
rect 1876 13804 1932 14310
rect 1988 14252 2044 15092
rect 2100 14530 2156 15092
rect 2100 14478 2102 14530
rect 2154 14478 2156 14530
rect 2100 14466 2156 14478
rect 2548 15146 2772 15148
rect 2548 15094 2718 15146
rect 2770 15094 2772 15146
rect 2548 15092 2772 15094
rect 2548 14476 2604 15092
rect 2716 15082 2772 15092
rect 2884 14924 2940 15184
rect 2884 14858 2940 14868
rect 2996 14700 3052 15876
rect 3220 15372 3276 15382
rect 3220 15314 3276 15316
rect 2324 14420 2604 14476
rect 2772 14644 3052 14700
rect 3108 15260 3164 15270
rect 3220 15262 3222 15314
rect 3274 15262 3276 15314
rect 3220 15250 3276 15262
rect 1988 14196 2212 14252
rect 1876 13738 1932 13748
rect 2156 13746 2212 14196
rect 2156 13694 2158 13746
rect 2210 13694 2212 13746
rect 2324 13802 2380 14420
rect 2324 13750 2326 13802
rect 2378 13750 2380 13802
rect 2324 13738 2380 13750
rect 2156 13682 2212 13694
rect 2324 13668 2380 13680
rect 2324 13616 2326 13668
rect 2378 13616 2380 13668
rect 1764 13178 1820 13188
rect 1876 13578 1932 13590
rect 1876 13526 1878 13578
rect 1930 13526 1932 13578
rect 1596 13078 1598 13130
rect 1650 13078 1652 13130
rect 1596 13066 1652 13078
rect 1708 12908 1764 12918
rect 1708 12814 1764 12852
rect 1876 12460 1932 13526
rect 2324 13580 2380 13616
rect 1876 12394 1932 12404
rect 2100 12950 2156 12962
rect 2100 12898 2102 12950
rect 2154 12898 2156 12950
rect 1596 12236 1652 12246
rect 2100 12236 2156 12898
rect 2324 12460 2380 13524
rect 2436 13020 2492 13030
rect 2436 12926 2492 12964
rect 2660 12962 2716 12974
rect 2660 12910 2662 12962
rect 2714 12910 2716 12962
rect 2660 12908 2716 12910
rect 2660 12842 2716 12852
rect 2324 12404 2492 12460
rect 2324 12236 2380 12246
rect 2100 12180 2324 12236
rect 1596 12142 1652 12180
rect 2324 12104 2380 12180
rect 1372 12010 1484 12022
rect 1372 11958 1374 12010
rect 1426 11958 1484 12010
rect 1372 11956 1484 11958
rect 1876 12012 1932 12022
rect 1372 11900 1428 11956
rect 1372 11834 1428 11844
rect 1876 11412 1932 11956
rect 2156 12012 2212 12022
rect 2436 12012 2492 12404
rect 2156 12010 2492 12012
rect 2156 11958 2158 12010
rect 2210 11958 2492 12010
rect 2156 11956 2492 11958
rect 2156 11946 2212 11956
rect 2212 11676 2268 11686
rect 2212 11562 2268 11620
rect 2660 11676 2716 11686
rect 2212 11510 2214 11562
rect 2266 11510 2268 11562
rect 2212 11498 2268 11510
rect 2324 11564 2380 11574
rect 1876 11360 1878 11412
rect 1930 11360 1932 11412
rect 1596 11340 1652 11350
rect 1876 11348 1932 11360
rect 1540 11338 1652 11340
rect 1540 11286 1598 11338
rect 1650 11286 1652 11338
rect 1540 11274 1652 11286
rect 1204 11172 1484 11228
rect 1428 10610 1484 11172
rect 1428 10558 1430 10610
rect 1482 10558 1484 10610
rect 1428 10546 1484 10558
rect 1540 9996 1596 11274
rect 2324 10678 2380 11508
rect 2660 11394 2716 11620
rect 2660 11342 2662 11394
rect 2714 11342 2716 11394
rect 2660 11330 2716 11342
rect 2772 11228 2828 14644
rect 3108 14588 3164 15204
rect 3892 14700 3948 16772
rect 4284 16762 4340 16772
rect 4676 16714 4732 16726
rect 4676 16662 4678 16714
rect 4730 16662 4732 16714
rect 4564 16156 4620 16166
rect 4676 16156 4732 16662
rect 4564 16154 4732 16156
rect 4564 16102 4566 16154
rect 4618 16102 4732 16154
rect 4564 16100 4732 16102
rect 4900 16716 4956 16726
rect 4900 16117 4956 16660
rect 4564 16090 4620 16100
rect 4900 16065 4902 16117
rect 4954 16065 4956 16117
rect 4900 16053 4956 16065
rect 6636 16268 6692 16278
rect 4956 15932 5012 15942
rect 4788 15930 5012 15932
rect 4788 15878 4958 15930
rect 5010 15878 5012 15930
rect 4788 15876 5012 15878
rect 4788 15370 4844 15876
rect 4956 15866 5012 15876
rect 6636 15820 6692 16212
rect 7028 16098 7084 16110
rect 6748 16044 6804 16054
rect 7028 16046 7030 16098
rect 7082 16046 7084 16098
rect 7028 16044 7084 16046
rect 6748 16042 7084 16044
rect 6748 15990 6750 16042
rect 6802 15990 7084 16042
rect 6748 15988 7084 15990
rect 6748 15978 6804 15988
rect 6636 15764 6748 15820
rect 4958 15708 5222 15718
rect 5014 15652 5062 15708
rect 5118 15652 5166 15708
rect 4958 15642 5222 15652
rect 6468 15484 6524 15494
rect 6468 15390 6524 15428
rect 4788 15318 4790 15370
rect 4842 15318 4844 15370
rect 4788 15306 4844 15318
rect 5516 15372 5572 15382
rect 5516 15278 5572 15316
rect 6692 15314 6748 15764
rect 7140 15596 7196 17556
rect 7252 17546 7308 17556
rect 7364 15708 7420 18564
rect 8708 18394 8764 18406
rect 8708 18342 8710 18394
rect 8762 18342 8764 18394
rect 7980 18284 8036 18294
rect 7924 18282 8036 18284
rect 7924 18230 7982 18282
rect 8034 18230 8036 18282
rect 7924 18218 8036 18230
rect 7924 17724 7980 18218
rect 8708 17836 8764 18342
rect 9044 18284 9100 19200
rect 11172 18732 11228 18742
rect 9996 18620 10052 18630
rect 9996 18450 10052 18564
rect 9996 18398 9998 18450
rect 10050 18398 10052 18450
rect 10164 18508 10220 18546
rect 10164 18442 10220 18452
rect 9996 18386 10052 18398
rect 10612 18394 10668 18406
rect 10164 18372 10220 18384
rect 10164 18320 10166 18372
rect 10218 18320 10220 18372
rect 9044 18218 9100 18228
rect 9268 18284 9380 18294
rect 9716 18284 9772 18294
rect 9324 18282 9380 18284
rect 9324 18230 9326 18282
rect 9378 18230 9380 18282
rect 9324 18228 9380 18230
rect 9268 18218 9380 18228
rect 9604 18282 9772 18284
rect 9604 18230 9718 18282
rect 9770 18230 9772 18282
rect 9604 18228 9772 18230
rect 8928 18060 9192 18070
rect 8984 18004 9032 18060
rect 9088 18004 9136 18060
rect 8928 17994 9192 18004
rect 8708 17770 8764 17780
rect 7532 16940 7588 16950
rect 7924 16940 7980 17668
rect 9492 17724 9548 17734
rect 9492 17633 9494 17668
rect 9546 17633 9548 17668
rect 8092 17610 8148 17622
rect 8092 17558 8094 17610
rect 8146 17558 8148 17610
rect 8092 17164 8148 17558
rect 8092 17098 8148 17108
rect 8372 17612 8428 17622
rect 7532 16938 7980 16940
rect 7532 16886 7534 16938
rect 7586 16886 7980 16938
rect 7532 16884 7980 16886
rect 8372 16938 8428 17556
rect 8932 17612 8988 17622
rect 9492 17621 9548 17633
rect 8932 17518 8988 17556
rect 8372 16886 8374 16938
rect 8426 16886 8428 16938
rect 7532 16874 7588 16884
rect 8372 16874 8428 16886
rect 8596 17276 8652 17286
rect 8596 16882 8652 17220
rect 8596 16830 8598 16882
rect 8650 16830 8652 16882
rect 8596 16818 8652 16830
rect 9436 17164 9492 17174
rect 9436 16714 9492 17108
rect 9436 16662 9438 16714
rect 9490 16662 9492 16714
rect 9436 16650 9492 16662
rect 8928 16492 9192 16502
rect 8984 16436 9032 16492
rect 9088 16436 9136 16492
rect 8928 16426 9192 16436
rect 8876 16156 8932 16166
rect 7868 16044 7924 16054
rect 7868 16042 7980 16044
rect 7868 15990 7870 16042
rect 7922 15990 7980 16042
rect 7868 15978 7980 15990
rect 7364 15642 7420 15652
rect 7140 15530 7196 15540
rect 6132 15296 6188 15308
rect 4060 15260 4116 15270
rect 4060 15166 4116 15204
rect 6132 15260 6134 15296
rect 6186 15260 6188 15296
rect 6692 15262 6694 15314
rect 6746 15262 6748 15314
rect 6692 15250 6748 15262
rect 6916 15372 6972 15382
rect 6132 15194 6188 15204
rect 5404 15148 5460 15158
rect 5404 15054 5460 15092
rect 6916 14710 6972 15316
rect 7532 15260 7588 15270
rect 7532 15166 7588 15204
rect 7924 15260 7980 15978
rect 8708 16042 8764 16054
rect 8708 15990 8710 16042
rect 8762 15990 8764 16042
rect 8708 15484 8764 15990
rect 8876 15932 8932 16100
rect 8876 15866 8932 15876
rect 9492 16086 9548 16098
rect 9492 16034 9494 16086
rect 9546 16034 9548 16086
rect 8596 15372 8652 15382
rect 8596 15314 8652 15316
rect 7924 15194 7980 15204
rect 8260 15258 8316 15270
rect 8260 15206 8262 15258
rect 8314 15206 8316 15258
rect 8596 15262 8598 15314
rect 8650 15262 8652 15314
rect 8596 15250 8652 15262
rect 4676 14700 4732 14710
rect 6860 14700 6972 14710
rect 2940 14532 3164 14588
rect 3780 14698 4732 14700
rect 3780 14646 4678 14698
rect 4730 14646 4732 14698
rect 3780 14644 4732 14646
rect 3780 14586 3836 14644
rect 4676 14634 4732 14644
rect 6692 14698 6972 14700
rect 6692 14646 6862 14698
rect 6914 14646 6972 14698
rect 6692 14644 6972 14646
rect 8092 15148 8148 15158
rect 8092 14698 8148 15092
rect 8092 14646 8094 14698
rect 8146 14646 8148 14698
rect 3780 14534 3782 14586
rect 3834 14534 3836 14586
rect 2940 14474 2996 14532
rect 3780 14522 3836 14534
rect 4116 14524 4172 14536
rect 2940 14422 2942 14474
rect 2994 14422 2996 14474
rect 2940 14410 2996 14422
rect 4116 14472 4118 14524
rect 4170 14472 4172 14524
rect 3500 14364 3556 14374
rect 3500 13802 3556 14308
rect 2996 13746 3052 13758
rect 2996 13694 2998 13746
rect 3050 13694 3052 13746
rect 2996 13692 3052 13694
rect 2996 13626 3052 13636
rect 3500 13750 3502 13802
rect 3554 13750 3556 13802
rect 3500 13130 3556 13750
rect 3500 13078 3502 13130
rect 3554 13078 3556 13130
rect 3500 13066 3556 13078
rect 4004 13580 4060 13590
rect 3164 12796 3220 12806
rect 3164 12234 3220 12740
rect 3164 12182 3166 12234
rect 3218 12182 3220 12234
rect 3164 12170 3220 12182
rect 4004 12178 4060 13524
rect 4116 12796 4172 14472
rect 5012 14518 5068 14530
rect 5012 14466 5014 14518
rect 5066 14466 5068 14518
rect 4228 14401 4284 14413
rect 4228 14349 4230 14401
rect 4282 14349 4284 14401
rect 4228 13802 4284 14349
rect 5012 14364 5068 14466
rect 5012 14298 5068 14308
rect 5516 14252 5572 14262
rect 4958 14140 5222 14150
rect 5014 14084 5062 14140
rect 5118 14084 5166 14140
rect 4958 14074 5222 14084
rect 5516 13914 5572 14196
rect 5516 13862 5518 13914
rect 5570 13862 5572 13914
rect 5516 13850 5572 13862
rect 6244 14252 6300 14262
rect 4228 13750 4230 13802
rect 4282 13750 4284 13802
rect 4228 13738 4284 13750
rect 5852 13692 5908 13702
rect 5852 13598 5908 13636
rect 4620 13578 4676 13590
rect 4620 13526 4622 13578
rect 4674 13526 4676 13578
rect 4620 13468 4676 13526
rect 4620 13402 4676 13412
rect 4732 13578 4788 13590
rect 4732 13526 4734 13578
rect 4786 13526 4788 13578
rect 4564 13020 4620 13030
rect 4732 13020 4788 13526
rect 5404 13580 5460 13590
rect 5404 13486 5460 13524
rect 5964 13580 6020 13590
rect 5964 13486 6020 13524
rect 4564 12926 4620 12964
rect 4676 12964 4788 13020
rect 4116 12730 4172 12740
rect 4228 12906 4284 12918
rect 4228 12854 4230 12906
rect 4282 12854 4284 12906
rect 4004 12126 4006 12178
rect 4058 12126 4060 12178
rect 4228 12236 4284 12854
rect 4228 12142 4284 12180
rect 4564 12160 4620 12172
rect 4004 12114 4060 12126
rect 4564 12108 4566 12160
rect 4618 12108 4620 12160
rect 3276 11564 3332 11574
rect 3276 11470 3332 11508
rect 4564 11564 4620 12108
rect 4676 11676 4732 12964
rect 6244 12962 6300 14196
rect 6356 13916 6412 13926
rect 6356 13758 6412 13860
rect 6692 13914 6748 14644
rect 6860 14634 6916 14644
rect 8092 14634 8148 14646
rect 7252 14530 7308 14542
rect 6972 14476 7028 14486
rect 7252 14478 7254 14530
rect 7306 14478 7308 14530
rect 7252 14476 7308 14478
rect 6972 14474 7308 14476
rect 6972 14422 6974 14474
rect 7026 14422 7308 14474
rect 6972 14420 7308 14422
rect 6972 14410 7028 14420
rect 8260 14364 8316 15206
rect 8260 14298 8316 14308
rect 8596 14924 8652 14934
rect 8036 14140 8092 14150
rect 6692 13862 6694 13914
rect 6746 13862 6748 13914
rect 6692 13850 6748 13862
rect 7476 14028 7532 14038
rect 6356 13706 6358 13758
rect 6410 13706 6412 13758
rect 6356 13694 6412 13706
rect 6916 13804 6972 13814
rect 6916 13706 6918 13748
rect 6970 13706 6972 13748
rect 7476 13758 7532 13972
rect 6916 13694 6972 13706
rect 7252 13734 7308 13746
rect 7252 13692 7254 13734
rect 7306 13692 7308 13734
rect 7476 13706 7478 13758
rect 7530 13706 7532 13758
rect 7476 13694 7532 13706
rect 7252 13626 7308 13636
rect 7812 13690 7868 13702
rect 7812 13638 7814 13690
rect 7866 13638 7868 13690
rect 7140 13580 7196 13590
rect 7140 13522 7196 13524
rect 7140 13470 7142 13522
rect 7194 13470 7196 13522
rect 7140 13458 7196 13470
rect 7812 13356 7868 13638
rect 7476 13300 7868 13356
rect 6860 13244 6916 13254
rect 6636 13132 6692 13142
rect 6636 13038 6692 13076
rect 6860 13130 6916 13188
rect 6860 13078 6862 13130
rect 6914 13078 6916 13130
rect 6860 13066 6916 13078
rect 7028 13132 7084 13142
rect 7028 13040 7084 13076
rect 7028 12988 7030 13040
rect 7082 12988 7084 13040
rect 7028 12976 7084 12988
rect 5404 12906 5460 12918
rect 5404 12854 5406 12906
rect 5458 12854 5460 12906
rect 6244 12910 6246 12962
rect 6298 12910 6300 12962
rect 6244 12898 6300 12910
rect 7028 12908 7084 12918
rect 7476 12908 7532 13300
rect 7588 13132 7644 13142
rect 7588 13038 7644 13076
rect 7028 12906 7532 12908
rect 5404 12796 5460 12854
rect 7028 12854 7030 12906
rect 7082 12854 7532 12906
rect 7028 12852 7532 12854
rect 7924 13018 7980 13030
rect 7924 12966 7926 13018
rect 7978 12966 7980 13018
rect 7028 12842 7084 12852
rect 5404 12730 5460 12740
rect 4958 12572 5222 12582
rect 5014 12516 5062 12572
rect 5118 12516 5166 12572
rect 4958 12506 5222 12516
rect 6468 12460 6524 12470
rect 6244 12348 6300 12358
rect 5852 12236 5908 12246
rect 5852 12142 5908 12180
rect 6244 12122 6300 12292
rect 6244 12070 6246 12122
rect 6298 12070 6300 12122
rect 6244 12058 6300 12070
rect 6468 12076 6524 12404
rect 7196 12348 7252 12358
rect 7196 12254 7252 12292
rect 6468 12024 6470 12076
rect 6522 12024 6524 12076
rect 5516 12012 5572 12022
rect 6468 12012 6524 12024
rect 7084 12012 7140 12022
rect 5516 11918 5572 11956
rect 7028 11956 7084 12012
rect 4676 11610 4732 11620
rect 7028 11880 7140 11956
rect 7924 12012 7980 12966
rect 8036 12168 8092 14084
rect 8148 13916 8204 13926
rect 8148 13822 8204 13860
rect 8428 13804 8484 13814
rect 8428 13746 8484 13748
rect 8204 13692 8260 13702
rect 8428 13694 8430 13746
rect 8482 13694 8484 13746
rect 8428 13682 8484 13694
rect 8596 13692 8652 14868
rect 8708 14588 8764 15428
rect 9492 15158 9548 16034
rect 9436 15148 9548 15158
rect 9492 15092 9548 15148
rect 9436 15054 9492 15092
rect 8928 14924 9192 14934
rect 8984 14868 9032 14924
rect 9088 14868 9136 14924
rect 8928 14858 9192 14868
rect 9604 14812 9660 18228
rect 9716 18218 9772 18228
rect 10164 18284 10220 18320
rect 10612 18342 10614 18394
rect 10666 18342 10668 18394
rect 10164 18218 10220 18228
rect 10444 18284 10500 18294
rect 10612 18284 10668 18342
rect 11172 18394 11228 18676
rect 11172 18342 11174 18394
rect 11226 18342 11228 18394
rect 11340 18620 11396 18630
rect 11340 18450 11396 18564
rect 11620 18508 11676 19200
rect 12898 18844 13162 18854
rect 12954 18788 13002 18844
rect 13058 18788 13106 18844
rect 12898 18778 13162 18788
rect 11620 18452 11788 18508
rect 11340 18398 11342 18450
rect 11394 18398 11396 18450
rect 11340 18386 11396 18398
rect 11732 18432 11788 18452
rect 11732 18396 11734 18432
rect 11786 18396 11788 18432
rect 13300 18450 13356 18462
rect 11172 18330 11228 18342
rect 11732 18330 11788 18340
rect 12516 18396 12572 18406
rect 10444 18282 10556 18284
rect 10444 18230 10446 18282
rect 10498 18230 10556 18282
rect 10444 18218 10556 18230
rect 10052 17836 10108 17846
rect 10052 17742 10108 17780
rect 10388 17654 10444 17666
rect 9772 17612 9828 17622
rect 10388 17612 10390 17654
rect 10442 17612 10444 17654
rect 9772 17610 9996 17612
rect 9772 17558 9774 17610
rect 9826 17558 9996 17610
rect 9772 17556 9996 17558
rect 9772 17546 9828 17556
rect 9828 17388 9884 17398
rect 9828 16266 9884 17332
rect 9940 17164 9996 17556
rect 10500 17612 10556 18218
rect 10612 18060 10668 18228
rect 10780 18284 10836 18294
rect 11004 18284 11060 18294
rect 10780 18190 10836 18228
rect 10948 18282 11060 18284
rect 10948 18230 11006 18282
rect 11058 18230 11060 18282
rect 10948 18218 11060 18230
rect 12068 18284 12124 18294
rect 12068 18282 12236 18284
rect 12068 18230 12070 18282
rect 12122 18230 12236 18282
rect 12068 18228 12236 18230
rect 12068 18218 12124 18228
rect 10948 18172 11004 18218
rect 10948 18106 11004 18116
rect 11172 18172 11228 18182
rect 10612 17994 10668 18004
rect 10948 17666 11004 17678
rect 10612 17612 10668 17622
rect 10500 17556 10612 17612
rect 10388 17546 10444 17556
rect 10612 17546 10668 17556
rect 10780 17612 10836 17622
rect 10780 17518 10836 17556
rect 10948 17614 10950 17666
rect 11002 17614 11004 17666
rect 10948 17388 11004 17614
rect 10276 17332 11004 17388
rect 11060 17500 11116 17510
rect 9940 17108 10220 17164
rect 10164 16938 10220 17108
rect 10164 16886 10166 16938
rect 10218 16886 10220 16938
rect 10164 16874 10220 16886
rect 9828 16214 9830 16266
rect 9882 16214 9884 16266
rect 9828 16202 9884 16214
rect 10108 16492 10164 16502
rect 10108 16266 10164 16436
rect 10276 16278 10332 17332
rect 10724 17164 10780 17174
rect 10612 16940 10668 16950
rect 10612 16278 10668 16884
rect 10724 16894 10780 17108
rect 10724 16842 10726 16894
rect 10778 16842 10780 16894
rect 11060 16884 11116 17444
rect 10724 16830 10780 16842
rect 10108 16214 10110 16266
rect 10162 16214 10164 16266
rect 10108 16202 10164 16214
rect 10220 16266 10332 16278
rect 10220 16214 10222 16266
rect 10274 16214 10332 16266
rect 10220 16212 10332 16214
rect 10556 16266 10668 16278
rect 10556 16214 10558 16266
rect 10610 16214 10668 16266
rect 10556 16212 10668 16214
rect 10836 16828 11116 16884
rect 10220 16202 10276 16212
rect 10556 16202 10612 16212
rect 10668 16044 10724 16054
rect 10836 16044 10892 16828
rect 11060 16716 11116 16726
rect 11172 16716 11228 18116
rect 11788 17836 11844 17846
rect 11788 17742 11844 17780
rect 11508 17612 11564 17622
rect 11060 16714 11228 16716
rect 11060 16662 11062 16714
rect 11114 16662 11228 16714
rect 11060 16660 11228 16662
rect 11284 16940 11340 16950
rect 11284 16714 11340 16884
rect 11284 16662 11286 16714
rect 11338 16662 11340 16714
rect 11060 16650 11116 16660
rect 11284 16650 11340 16662
rect 11396 16828 11452 16838
rect 11004 16268 11060 16278
rect 11004 16174 11060 16212
rect 11172 16268 11228 16278
rect 11172 16176 11228 16212
rect 11172 16124 11174 16176
rect 11226 16124 11228 16176
rect 11172 16112 11228 16124
rect 10668 16042 10892 16044
rect 10668 15990 10670 16042
rect 10722 15990 10892 16042
rect 10668 15988 10892 15990
rect 11172 16044 11228 16054
rect 11396 16044 11452 16772
rect 11508 16716 11564 17556
rect 11620 17052 11676 17062
rect 11620 16894 11676 16996
rect 11620 16842 11622 16894
rect 11674 16842 11676 16894
rect 11620 16830 11676 16842
rect 11956 16828 12012 16838
rect 11956 16734 12012 16772
rect 11620 16716 11676 16726
rect 11508 16660 11620 16716
rect 11620 16166 11676 16660
rect 12180 16492 12236 18228
rect 12404 18282 12460 18294
rect 12404 18230 12406 18282
rect 12458 18230 12460 18282
rect 12404 18172 12460 18230
rect 12404 18106 12460 18116
rect 12516 17500 12572 18340
rect 13300 18398 13302 18450
rect 13354 18398 13356 18450
rect 13300 18396 13356 18398
rect 13300 18330 13356 18340
rect 14196 18396 14252 19200
rect 15988 18956 16044 18966
rect 15652 18732 15708 18742
rect 15428 18432 15484 18444
rect 14196 18330 14252 18340
rect 14868 18394 14924 18406
rect 14868 18342 14870 18394
rect 14922 18342 14924 18394
rect 12740 18282 12796 18294
rect 12740 18230 12742 18282
rect 12794 18230 12796 18282
rect 12628 17724 12684 17734
rect 12740 17724 12796 18230
rect 14028 18282 14084 18294
rect 14028 18230 14030 18282
rect 14082 18230 14084 18282
rect 14028 17836 14084 18230
rect 14028 17770 14084 17780
rect 14420 18172 14476 18182
rect 12628 17722 12796 17724
rect 12628 17670 12630 17722
rect 12682 17670 12796 17722
rect 14420 17722 14476 18116
rect 14868 17836 14924 18342
rect 15316 18396 15372 18406
rect 15428 18396 15430 18432
rect 15372 18380 15430 18396
rect 15482 18380 15484 18432
rect 15372 18340 15484 18380
rect 15092 18284 15148 18294
rect 15092 18190 15148 18228
rect 14868 17770 14924 17780
rect 12628 17668 12796 17670
rect 12628 17658 12684 17668
rect 12852 17666 12908 17678
rect 12852 17614 12854 17666
rect 12906 17614 12908 17666
rect 14420 17670 14422 17722
rect 14474 17670 14476 17722
rect 14420 17658 14476 17670
rect 14980 17724 15036 17734
rect 14980 17633 14982 17668
rect 15034 17633 15036 17668
rect 12852 17500 12908 17614
rect 13692 17612 13748 17622
rect 14980 17621 15036 17633
rect 15316 17668 15372 18340
rect 15428 17836 15484 17846
rect 15428 17742 15484 17780
rect 15316 17612 15484 17668
rect 13692 17610 13804 17612
rect 13692 17558 13694 17610
rect 13746 17558 13804 17610
rect 13692 17546 13804 17558
rect 12516 17444 12796 17500
rect 12292 17052 12348 17062
rect 12292 16958 12348 16996
rect 12348 16658 12404 16670
rect 12348 16606 12350 16658
rect 12402 16614 12404 16658
rect 12572 16658 12628 16670
rect 12402 16606 12460 16614
rect 12348 16604 12460 16606
rect 12348 16548 12404 16604
rect 12404 16538 12460 16548
rect 12572 16606 12574 16658
rect 12626 16606 12628 16658
rect 12180 16436 12348 16492
rect 12124 16268 12180 16278
rect 12124 16174 12180 16212
rect 11564 16156 11676 16166
rect 11564 16154 11620 16156
rect 11564 16102 11566 16154
rect 11618 16102 11620 16154
rect 11564 16100 11620 16102
rect 11564 16090 11676 16100
rect 11172 16042 11452 16044
rect 11172 15990 11174 16042
rect 11226 15990 11452 16042
rect 11620 16024 11676 16090
rect 11788 16156 11844 16166
rect 11788 16062 11844 16100
rect 11172 15988 11452 15990
rect 10668 15978 10724 15988
rect 11172 15978 11228 15988
rect 10668 15484 10724 15494
rect 10276 15482 10724 15484
rect 10276 15430 10670 15482
rect 10722 15430 10724 15482
rect 10276 15428 10724 15430
rect 10276 15370 10332 15428
rect 10668 15418 10724 15428
rect 10276 15318 10278 15370
rect 10330 15318 10332 15370
rect 10276 15306 10332 15318
rect 12292 15372 12348 16436
rect 12572 16268 12628 16606
rect 12572 16202 12628 16212
rect 12628 15708 12684 15718
rect 12516 15484 12572 15494
rect 12516 15386 12518 15428
rect 12570 15386 12572 15428
rect 12516 15374 12572 15386
rect 12292 15316 12404 15372
rect 10612 15295 10668 15307
rect 10612 15260 10614 15295
rect 10666 15260 10668 15295
rect 12068 15302 12124 15314
rect 10612 15194 10668 15204
rect 11060 15260 11116 15270
rect 9604 14746 9660 14756
rect 10052 14700 10108 14710
rect 10948 14700 11004 14710
rect 8820 14588 8876 14598
rect 8708 14586 9772 14588
rect 8708 14534 8822 14586
rect 8874 14548 9772 14586
rect 8874 14534 9718 14548
rect 8708 14532 9718 14534
rect 8820 14522 8876 14532
rect 9716 14496 9718 14532
rect 9770 14496 9772 14548
rect 9716 14484 9772 14496
rect 9380 14364 9436 14374
rect 9380 14270 9436 14308
rect 10052 14140 10108 14644
rect 10276 14644 10668 14700
rect 10276 14586 10332 14644
rect 10276 14534 10278 14586
rect 10330 14534 10332 14586
rect 10276 14522 10332 14534
rect 10444 14530 10500 14542
rect 10052 14074 10108 14084
rect 10164 14476 10220 14486
rect 9828 14028 9884 14038
rect 9492 13916 9548 13926
rect 9492 13822 9548 13860
rect 9828 13914 9884 13972
rect 9828 13862 9830 13914
rect 9882 13862 9884 13914
rect 9828 13850 9884 13862
rect 8204 13598 8260 13636
rect 8596 13468 8652 13636
rect 9940 13746 9996 13758
rect 9940 13694 9942 13746
rect 9994 13694 9996 13746
rect 9940 13692 9996 13694
rect 10164 13746 10220 14420
rect 10444 14478 10446 14530
rect 10498 14478 10500 14530
rect 10332 14364 10388 14374
rect 10164 13694 10166 13746
rect 10218 13694 10220 13746
rect 10164 13682 10220 13694
rect 10276 14362 10388 14364
rect 10276 14310 10334 14362
rect 10386 14310 10388 14362
rect 10276 14298 10388 14310
rect 9940 13626 9996 13636
rect 9044 13580 9156 13590
rect 9100 13578 9156 13580
rect 9100 13526 9102 13578
rect 9154 13526 9156 13578
rect 9100 13524 9156 13526
rect 9044 13514 9156 13524
rect 8540 13412 8652 13468
rect 8260 13356 8316 13366
rect 8540 13356 8596 13412
rect 8260 13018 8316 13300
rect 8260 12966 8262 13018
rect 8314 12966 8316 13018
rect 8260 12348 8316 12966
rect 8484 13300 8596 13356
rect 8928 13356 9192 13366
rect 8984 13300 9032 13356
rect 9088 13300 9136 13356
rect 8484 12796 8540 13300
rect 8928 13290 9192 13300
rect 8652 13244 8708 13254
rect 8652 13186 8708 13188
rect 8652 13134 8654 13186
rect 8706 13134 8708 13186
rect 8652 13122 8708 13134
rect 8876 13132 8932 13142
rect 8876 13038 8932 13076
rect 9660 12906 9716 12918
rect 10108 12908 10164 12918
rect 9660 12854 9662 12906
rect 9714 12854 9716 12906
rect 8596 12796 8652 12806
rect 8484 12794 8652 12796
rect 8484 12742 8598 12794
rect 8650 12742 8652 12794
rect 8484 12740 8652 12742
rect 9660 12796 9716 12854
rect 10052 12852 10108 12908
rect 10052 12814 10164 12852
rect 9884 12796 9940 12806
rect 9660 12740 9884 12796
rect 8596 12730 8652 12740
rect 8260 12282 8316 12292
rect 9492 12178 9548 12190
rect 8036 12112 8316 12168
rect 8820 12160 8876 12172
rect 8820 12124 8822 12160
rect 8874 12124 8876 12160
rect 7924 11946 7980 11956
rect 4564 11498 4620 11508
rect 6244 11587 6300 11599
rect 6244 11535 6246 11587
rect 6298 11535 6300 11587
rect 2268 10666 2380 10678
rect 2268 10614 2270 10666
rect 2322 10614 2380 10666
rect 2268 10612 2380 10614
rect 2436 11172 2828 11228
rect 3108 11452 3164 11462
rect 2268 10602 2324 10612
rect 1428 9940 1540 9996
rect 1316 9324 1372 9334
rect 1316 8428 1372 9268
rect 1428 9110 1484 9940
rect 1540 9930 1596 9940
rect 1540 9814 1596 9826
rect 1540 9762 1542 9814
rect 1594 9762 1596 9814
rect 1540 9324 1596 9762
rect 1540 9258 1596 9268
rect 1876 9658 1932 9670
rect 1876 9606 1878 9658
rect 1930 9606 1932 9658
rect 1876 9324 1932 9606
rect 1876 9258 1932 9268
rect 1428 9098 1540 9110
rect 1428 9046 1486 9098
rect 1538 9046 1540 9098
rect 1428 9044 1540 9046
rect 1876 9044 1932 9054
rect 1484 9034 1540 9044
rect 1596 9042 1932 9044
rect 1596 8990 1878 9042
rect 1930 8990 1932 9042
rect 1596 8988 1932 8990
rect 1596 8986 1652 8988
rect 1596 8934 1598 8986
rect 1650 8934 1652 8986
rect 1876 8978 1932 8988
rect 1596 8922 1652 8934
rect 1484 8428 1540 8438
rect 1316 8426 1540 8428
rect 1316 8374 1486 8426
rect 1538 8374 1540 8426
rect 1316 8372 1540 8374
rect 1484 8362 1540 8372
rect 2436 8258 2492 11172
rect 2996 10556 3052 10566
rect 2996 10462 3052 10500
rect 3108 10006 3164 11396
rect 4452 11452 4508 11462
rect 6244 11452 6300 11535
rect 4452 11361 4454 11396
rect 4506 11361 4508 11396
rect 4116 11338 4172 11350
rect 4452 11349 4508 11361
rect 5796 11394 5852 11406
rect 4116 11286 4118 11338
rect 4170 11286 4172 11338
rect 4116 11228 4172 11286
rect 5796 11342 5798 11394
rect 5850 11342 5852 11394
rect 6244 11386 6300 11396
rect 6804 11452 6860 11462
rect 6804 11394 6860 11396
rect 5796 11340 5852 11342
rect 5796 11274 5852 11284
rect 6020 11338 6076 11350
rect 6020 11286 6022 11338
rect 6074 11286 6076 11338
rect 6804 11342 6806 11394
rect 6858 11342 6860 11394
rect 6804 11330 6860 11342
rect 4508 11228 4564 11238
rect 4116 11226 4564 11228
rect 4116 11174 4510 11226
rect 4562 11174 4564 11226
rect 4116 11172 4564 11174
rect 4508 11162 4564 11172
rect 4958 11004 5222 11014
rect 5014 10948 5062 11004
rect 5118 10948 5166 11004
rect 4958 10938 5222 10948
rect 2548 9996 2604 10006
rect 3052 9996 3164 10006
rect 2548 9826 2604 9940
rect 2548 9774 2550 9826
rect 2602 9774 2604 9826
rect 2548 9762 2604 9774
rect 2772 9994 3164 9996
rect 2772 9942 3054 9994
rect 3106 9942 3164 9994
rect 2772 9940 3164 9942
rect 3556 10668 3612 10678
rect 3556 10587 3612 10612
rect 3556 10535 3558 10587
rect 3610 10535 3612 10587
rect 4228 10668 4284 10678
rect 4228 10574 4284 10612
rect 5460 10598 5516 10610
rect 2772 9110 2828 9940
rect 3052 9930 3108 9940
rect 2716 9098 2828 9110
rect 2716 9046 2718 9098
rect 2770 9046 2828 9098
rect 2716 9044 2828 9046
rect 3444 9100 3500 9110
rect 3556 9100 3612 10535
rect 4788 10556 4844 10566
rect 4788 10454 4844 10500
rect 5460 10546 5462 10598
rect 5514 10546 5516 10598
rect 4788 10442 4900 10454
rect 4788 10390 4846 10442
rect 4898 10390 4900 10442
rect 4788 10378 4900 10390
rect 5460 10444 5516 10546
rect 4060 9996 4116 10006
rect 4060 9902 4116 9940
rect 4564 9814 4620 9826
rect 3892 9770 3948 9782
rect 3892 9718 3894 9770
rect 3946 9718 3948 9770
rect 3892 9212 3948 9718
rect 4564 9762 4566 9814
rect 4618 9762 4620 9814
rect 4564 9660 4620 9762
rect 4564 9594 4620 9604
rect 4788 9772 4844 10378
rect 5460 10220 5516 10388
rect 5460 10154 5516 10164
rect 5908 10598 5964 10610
rect 5908 10546 5910 10598
rect 5962 10546 5964 10598
rect 4900 10108 4956 10118
rect 4900 9994 4956 10052
rect 5908 10108 5964 10546
rect 5908 10042 5964 10052
rect 4900 9942 4902 9994
rect 4954 9942 4956 9994
rect 4900 9930 4956 9942
rect 5572 9884 5628 9894
rect 5460 9882 5628 9884
rect 5460 9830 5574 9882
rect 5626 9830 5628 9882
rect 5460 9828 5628 9830
rect 4116 9212 4172 9222
rect 3892 9210 4172 9212
rect 3892 9158 4118 9210
rect 4170 9158 4172 9210
rect 3892 9156 4172 9158
rect 4116 9146 4172 9156
rect 4788 9110 4844 9716
rect 5068 9772 5124 9782
rect 5068 9678 5124 9716
rect 4958 9436 5222 9446
rect 5014 9380 5062 9436
rect 5118 9380 5166 9436
rect 4958 9370 5222 9380
rect 3724 9100 3780 9110
rect 3556 9098 3780 9100
rect 3556 9046 3726 9098
rect 3778 9046 3780 9098
rect 3556 9044 3780 9046
rect 2716 9034 2772 9044
rect 3444 9006 3500 9044
rect 3724 9034 3780 9044
rect 4564 9100 4620 9110
rect 4732 9100 4844 9110
rect 4620 9098 4844 9100
rect 4620 9046 4734 9098
rect 4786 9046 4844 9098
rect 4620 9044 4844 9046
rect 4564 8998 4620 9044
rect 4732 9034 4788 9044
rect 4508 8986 4620 8998
rect 4508 8934 4510 8986
rect 4562 8934 4620 8986
rect 4508 8932 4620 8934
rect 5460 9019 5516 9828
rect 5572 9818 5628 9828
rect 5908 9884 5964 9894
rect 5908 9790 5964 9828
rect 6020 9100 6076 11286
rect 7028 10668 7084 11880
rect 7140 11676 7196 11686
rect 7140 11400 7196 11620
rect 8148 11562 8204 11574
rect 8148 11510 8150 11562
rect 8202 11510 8204 11562
rect 7140 11348 7142 11400
rect 7194 11348 7196 11400
rect 7140 11336 7196 11348
rect 7252 11452 7308 11462
rect 7028 10602 7084 10612
rect 7252 10108 7308 11396
rect 8036 11338 8092 11350
rect 6468 10076 6524 10088
rect 6468 10024 6470 10076
rect 6522 10024 6524 10076
rect 6468 9996 6524 10024
rect 6468 9930 6524 9940
rect 7252 9894 7308 10052
rect 7476 11282 7532 11294
rect 7476 11230 7478 11282
rect 7530 11230 7532 11282
rect 7476 9996 7532 11230
rect 8036 11286 8038 11338
rect 8090 11286 8092 11338
rect 8036 11228 8092 11286
rect 8036 11162 8092 11172
rect 8148 11116 8204 11510
rect 8260 11394 8316 12112
rect 8260 11342 8262 11394
rect 8314 11342 8316 11394
rect 8260 11330 8316 11342
rect 8708 12068 8820 12124
rect 8708 11340 8764 12068
rect 8820 12058 8876 12068
rect 9492 12126 9494 12178
rect 9546 12126 9548 12178
rect 9156 12012 9212 12022
rect 9492 12012 9548 12126
rect 9156 12010 9324 12012
rect 9156 11958 9158 12010
rect 9210 11958 9324 12010
rect 9156 11956 9324 11958
rect 9156 11946 9212 11956
rect 9268 11900 9324 11956
rect 9492 11946 9548 11956
rect 9268 11834 9324 11844
rect 8928 11788 9192 11798
rect 8984 11732 9032 11788
rect 9088 11732 9136 11788
rect 8928 11722 9192 11732
rect 9324 11676 9380 11686
rect 9324 11562 9380 11620
rect 9716 11574 9772 12740
rect 9884 12702 9940 12740
rect 10052 12124 10108 12814
rect 10052 11900 10108 12068
rect 9324 11510 9326 11562
rect 9378 11510 9380 11562
rect 9324 11498 9380 11510
rect 9660 11564 9772 11574
rect 9660 11562 9716 11564
rect 9660 11510 9662 11562
rect 9714 11510 9716 11562
rect 9660 11508 9716 11510
rect 9660 11498 9772 11508
rect 9716 11432 9772 11498
rect 9884 11844 10108 11900
rect 10276 12236 10332 14298
rect 10444 14028 10500 14478
rect 10444 13972 10556 14028
rect 10500 13804 10556 13972
rect 10500 13468 10556 13748
rect 10612 13580 10668 14644
rect 10948 14608 11004 14644
rect 10948 14556 10950 14608
rect 11002 14556 11004 14608
rect 10948 14544 11004 14556
rect 10780 14530 10836 14542
rect 10780 14478 10782 14530
rect 10834 14478 10836 14530
rect 10780 14476 10836 14478
rect 10780 14410 10836 14420
rect 10948 14476 11004 14486
rect 11060 14476 11116 15204
rect 12068 15260 12070 15302
rect 12122 15260 12124 15302
rect 12068 15194 12124 15204
rect 11396 15146 11452 15158
rect 11396 15094 11398 15146
rect 11450 15094 11452 15146
rect 11396 15036 11452 15094
rect 11396 14970 11452 14980
rect 11732 15146 11788 15158
rect 11732 15094 11734 15146
rect 11786 15094 11788 15146
rect 11732 15036 11788 15094
rect 12236 15148 12292 15168
rect 12236 15090 12292 15092
rect 12236 15038 12238 15090
rect 12290 15038 12292 15090
rect 12236 15036 12292 15038
rect 11508 14924 11564 14934
rect 10948 14474 11116 14476
rect 10948 14422 10950 14474
rect 11002 14422 11116 14474
rect 10948 14420 11116 14422
rect 11172 14700 11228 14710
rect 10948 14410 11004 14420
rect 10948 13580 11004 13590
rect 10612 13578 11004 13580
rect 10612 13526 10950 13578
rect 11002 13526 11004 13578
rect 10612 13524 11004 13526
rect 10500 13412 10668 13468
rect 10444 13020 10500 13030
rect 10444 12926 10500 12964
rect 9884 11450 9940 11844
rect 10276 11788 10332 12180
rect 10612 12124 10668 13412
rect 10948 12962 11004 13524
rect 10948 12910 10950 12962
rect 11002 12910 11004 12962
rect 10948 12908 11004 12910
rect 10612 12058 10668 12068
rect 10836 12852 11004 12908
rect 10500 12012 10556 12022
rect 10276 11732 10444 11788
rect 10052 11564 10164 11574
rect 10108 11562 10164 11564
rect 10108 11510 10110 11562
rect 10162 11510 10164 11562
rect 10108 11508 10164 11510
rect 10052 11498 10164 11508
rect 9884 11398 9886 11450
rect 9938 11398 9940 11450
rect 9884 11386 9940 11398
rect 10276 11452 10332 11462
rect 9436 11340 9492 11350
rect 8764 11284 8988 11340
rect 8708 11208 8764 11284
rect 8148 11050 8204 11060
rect 8932 10778 8988 11284
rect 8932 10726 8934 10778
rect 8986 10726 8988 10778
rect 8932 10714 8988 10726
rect 9436 10780 9492 11284
rect 10276 11238 10332 11396
rect 10388 11340 10444 11732
rect 10500 11574 10556 11956
rect 10500 11562 10612 11574
rect 10500 11510 10558 11562
rect 10610 11510 10612 11562
rect 10500 11508 10612 11510
rect 10556 11498 10612 11508
rect 10836 11452 10892 12852
rect 11172 12290 11228 14644
rect 11508 14608 11564 14868
rect 11508 14556 11510 14608
rect 11562 14556 11564 14608
rect 11508 14544 11564 14556
rect 11340 14530 11396 14542
rect 11340 14478 11342 14530
rect 11394 14478 11396 14530
rect 11340 14476 11396 14478
rect 11340 14410 11396 14420
rect 11732 14476 11788 14980
rect 12068 14980 12292 15036
rect 11844 14812 11900 14822
rect 11844 14542 11900 14756
rect 11844 14490 11846 14542
rect 11898 14490 11900 14542
rect 11844 14478 11900 14490
rect 11732 14410 11788 14420
rect 11452 14364 11508 14374
rect 11452 14362 11676 14364
rect 11452 14310 11454 14362
rect 11506 14310 11676 14362
rect 11452 14308 11676 14310
rect 11452 14298 11508 14308
rect 11284 14140 11340 14150
rect 11284 13914 11340 14084
rect 11284 13862 11286 13914
rect 11338 13862 11340 13914
rect 11284 13850 11340 13862
rect 11508 14140 11564 14150
rect 11508 13804 11564 14084
rect 11508 13738 11564 13748
rect 11620 13692 11676 14308
rect 12068 14252 12124 14980
rect 12348 14924 12404 15316
rect 12628 15326 12684 15652
rect 12628 15274 12630 15326
rect 12682 15274 12684 15326
rect 12628 15262 12684 15274
rect 12460 15148 12516 15158
rect 12460 15146 12684 15148
rect 12460 15094 12462 15146
rect 12514 15094 12684 15146
rect 12460 15092 12684 15094
rect 12460 15082 12516 15092
rect 12628 15036 12684 15092
rect 12628 14970 12684 14980
rect 12292 14868 12404 14924
rect 12180 14812 12236 14822
rect 12180 14728 12182 14756
rect 12234 14728 12236 14756
rect 12180 14716 12236 14728
rect 12012 14196 12124 14252
rect 12180 14518 12236 14530
rect 12180 14476 12182 14518
rect 12234 14476 12236 14518
rect 11788 13692 11844 13702
rect 11620 13690 11844 13692
rect 11620 13638 11790 13690
rect 11842 13638 11844 13690
rect 11620 13636 11844 13638
rect 11788 13626 11844 13636
rect 11396 13580 11508 13590
rect 11452 13578 11508 13580
rect 11452 13526 11454 13578
rect 11506 13526 11508 13578
rect 11452 13524 11508 13526
rect 11396 13514 11508 13524
rect 12012 13522 12068 14196
rect 12180 13742 12236 14420
rect 12292 14364 12348 14868
rect 12404 14700 12460 14710
rect 12404 14542 12460 14644
rect 12404 14490 12406 14542
rect 12458 14490 12460 14542
rect 12404 14478 12460 14490
rect 12516 14476 12572 14486
rect 12292 14308 12460 14364
rect 12404 13758 12460 14308
rect 12180 13690 12292 13742
rect 12404 13706 12406 13758
rect 12458 13706 12460 13758
rect 12404 13694 12460 13706
rect 12180 13686 12238 13690
rect 12236 13638 12238 13686
rect 12290 13638 12292 13690
rect 12236 13626 12292 13638
rect 12012 13470 12014 13522
rect 12066 13470 12068 13522
rect 12124 13580 12180 13590
rect 12124 13486 12180 13524
rect 12012 13468 12068 13470
rect 12012 13402 12068 13412
rect 11508 13356 11564 13366
rect 11396 13020 11452 13030
rect 11396 12962 11452 12964
rect 11396 12910 11398 12962
rect 11450 12910 11452 12962
rect 11396 12898 11452 12910
rect 11172 12238 11174 12290
rect 11226 12238 11228 12290
rect 11172 12226 11228 12238
rect 11508 12794 11564 13300
rect 12068 13074 12124 13086
rect 12068 13022 12070 13074
rect 12122 13022 12124 13074
rect 11956 12962 12012 12974
rect 11956 12910 11958 12962
rect 12010 12910 12012 12962
rect 11956 12908 12012 12910
rect 11956 12842 12012 12852
rect 11508 12742 11510 12794
rect 11562 12742 11564 12794
rect 11508 11676 11564 12742
rect 12068 12796 12124 13022
rect 11732 12460 11788 12470
rect 11620 12178 11676 12190
rect 11620 12126 11622 12178
rect 11674 12126 11676 12178
rect 11620 12124 11676 12126
rect 11620 12058 11676 12068
rect 11732 12066 11788 12404
rect 11732 12014 11734 12066
rect 11786 12014 11788 12066
rect 11732 12002 11788 12014
rect 12068 11900 12124 12740
rect 12292 12796 12348 12806
rect 12180 12160 12236 12172
rect 12180 12108 12182 12160
rect 12234 12108 12236 12160
rect 12180 12012 12236 12108
rect 12180 11946 12236 11956
rect 12068 11834 12124 11844
rect 11508 11610 11564 11620
rect 11844 11788 11900 11798
rect 10948 11564 11004 11574
rect 10948 11470 11004 11508
rect 11396 11564 11452 11574
rect 11396 11472 11452 11508
rect 10836 11386 10892 11396
rect 11060 11452 11116 11462
rect 11396 11420 11398 11472
rect 11450 11420 11452 11472
rect 11396 11408 11452 11420
rect 11620 11564 11676 11574
rect 10388 11284 10556 11340
rect 9660 11228 9716 11238
rect 9660 10834 9716 11172
rect 10220 11226 10332 11238
rect 10220 11174 10222 11226
rect 10274 11174 10332 11226
rect 10220 11172 10332 11174
rect 10220 11162 10276 11172
rect 9660 10782 9662 10834
rect 9714 10782 9716 10834
rect 9436 10778 9548 10780
rect 9436 10726 9438 10778
rect 9490 10726 9548 10778
rect 9660 10770 9716 10782
rect 9940 11004 9996 11014
rect 9436 10714 9548 10726
rect 8260 10556 8316 10566
rect 8260 10462 8316 10500
rect 9100 10444 9156 10482
rect 9156 10388 9324 10444
rect 9100 10378 9156 10388
rect 8928 10220 9192 10230
rect 8984 10164 9032 10220
rect 9088 10164 9136 10220
rect 8928 10154 9192 10164
rect 7476 9894 7532 9940
rect 8092 10108 8148 10118
rect 8092 9938 8148 10052
rect 6188 9884 6244 9894
rect 6748 9884 6804 9894
rect 6188 9882 6300 9884
rect 6188 9830 6190 9882
rect 6242 9830 6300 9882
rect 6188 9818 6300 9830
rect 6748 9882 6860 9884
rect 6748 9830 6750 9882
rect 6802 9830 6860 9882
rect 6132 9100 6188 9110
rect 6020 9098 6188 9100
rect 6020 9046 6134 9098
rect 6186 9046 6188 9098
rect 6020 9044 6188 9046
rect 5460 8967 5462 9019
rect 5514 8967 5516 9019
rect 4508 8922 4564 8932
rect 2436 8206 2438 8258
rect 2490 8206 2492 8258
rect 2436 8194 2492 8206
rect 3220 8426 3276 8438
rect 3220 8374 3222 8426
rect 3274 8374 3276 8426
rect 1988 8146 2044 8158
rect 1316 8092 1372 8102
rect 1204 6972 1260 6982
rect 868 2604 924 2614
rect 1204 2604 1260 6916
rect 1316 6748 1372 8036
rect 1988 8094 1990 8146
rect 2042 8094 2044 8146
rect 1484 7306 1540 7318
rect 1484 7254 1486 7306
rect 1538 7254 1540 7306
rect 1484 7084 1540 7254
rect 1484 7018 1540 7028
rect 1596 7306 1652 7318
rect 1596 7254 1598 7306
rect 1650 7254 1652 7306
rect 1596 6860 1652 7254
rect 1988 6972 2044 8094
rect 2884 7700 3164 7756
rect 2548 7418 2604 7430
rect 2548 7366 2550 7418
rect 2602 7366 2604 7418
rect 2436 7084 2492 7094
rect 1988 6906 2044 6916
rect 2268 6972 2324 6982
rect 1596 6804 1708 6860
rect 1316 6692 1596 6748
rect 1540 6678 1596 6692
rect 1540 6626 1542 6678
rect 1594 6626 1596 6678
rect 1540 5896 1596 6626
rect 1652 6524 1708 6804
rect 1876 6636 1932 6646
rect 2268 6636 2324 6916
rect 1876 6634 2324 6636
rect 1876 6582 1878 6634
rect 1930 6582 2270 6634
rect 2322 6582 2324 6634
rect 1876 6580 2324 6582
rect 1876 6570 1932 6580
rect 2268 6570 2324 6580
rect 2436 6534 2492 7028
rect 2548 6748 2604 7366
rect 2884 6870 2940 7700
rect 3108 7642 3164 7700
rect 3108 7590 3110 7642
rect 3162 7590 3164 7642
rect 3108 7578 3164 7590
rect 2828 6858 2940 6870
rect 2828 6806 2830 6858
rect 2882 6806 2940 6858
rect 2828 6804 2940 6806
rect 2996 7530 3052 7542
rect 2996 7478 2998 7530
rect 3050 7478 3052 7530
rect 3220 7488 3276 8374
rect 4004 8314 4060 8326
rect 3780 8258 3836 8270
rect 3780 8206 3782 8258
rect 3834 8206 3836 8258
rect 3780 7644 3836 8206
rect 4004 8262 4006 8314
rect 4058 8262 4060 8314
rect 4004 7644 4060 8262
rect 4732 8316 4788 8326
rect 4956 8316 5012 8326
rect 4732 8314 4956 8316
rect 4732 8262 4734 8314
rect 4786 8262 4956 8314
rect 4732 8260 4956 8262
rect 4732 8250 4788 8260
rect 4956 8222 5012 8260
rect 5460 8202 5516 8967
rect 6132 8540 6188 9044
rect 6244 8764 6300 9818
rect 6468 9814 6524 9826
rect 6748 9818 6860 9830
rect 7196 9882 7308 9894
rect 7196 9830 7198 9882
rect 7250 9830 7308 9882
rect 7196 9828 7308 9830
rect 7420 9882 7532 9894
rect 7420 9830 7422 9882
rect 7474 9830 7532 9882
rect 7420 9828 7532 9830
rect 7756 9884 7812 9894
rect 8092 9886 8094 9938
rect 8146 9886 8148 9938
rect 8092 9874 8148 9886
rect 8316 9996 8372 10006
rect 7196 9818 7252 9828
rect 7420 9818 7476 9828
rect 6468 9762 6470 9814
rect 6522 9762 6524 9814
rect 6468 8988 6524 9762
rect 6468 8922 6524 8932
rect 6356 8764 6412 8774
rect 6244 8708 6356 8764
rect 6132 8474 6188 8484
rect 6356 8451 6412 8708
rect 6356 8399 6358 8451
rect 6410 8399 6412 8451
rect 6356 8387 6412 8399
rect 5460 8150 5462 8202
rect 5514 8150 5516 8202
rect 5908 8316 5964 8326
rect 5908 8258 5964 8260
rect 5908 8206 5910 8258
rect 5962 8206 5964 8258
rect 5908 8194 5964 8206
rect 6636 8204 6692 8214
rect 6580 8202 6692 8204
rect 4340 8092 4396 8102
rect 4340 7998 4396 8036
rect 4958 7868 5222 7878
rect 5014 7812 5062 7868
rect 5118 7812 5166 7868
rect 4958 7802 5222 7812
rect 4452 7756 4508 7766
rect 3780 7588 3948 7644
rect 4004 7588 4340 7644
rect 2828 6794 2884 6804
rect 2548 6692 2716 6748
rect 2436 6522 2548 6534
rect 2436 6470 2494 6522
rect 2546 6470 2548 6522
rect 2436 6468 2548 6470
rect 1652 6458 1708 6468
rect 2492 6458 2548 6468
rect 2324 6076 2380 6086
rect 2324 5982 2380 6020
rect 1316 5840 1596 5896
rect 1988 5850 2044 5862
rect 1316 2828 1372 5840
rect 1988 5798 1990 5850
rect 2042 5798 2044 5850
rect 1484 5740 1540 5750
rect 1484 5646 1540 5684
rect 1596 5738 1652 5750
rect 1596 5686 1598 5738
rect 1650 5686 1652 5738
rect 1484 5516 1540 5526
rect 1484 4954 1540 5460
rect 1596 5124 1652 5686
rect 1988 5740 2044 5798
rect 2492 5740 2548 5750
rect 1988 5292 2044 5684
rect 2268 5682 2324 5694
rect 2268 5630 2270 5682
rect 2322 5630 2324 5682
rect 2492 5646 2548 5684
rect 2156 5404 2212 5414
rect 2156 5346 2212 5348
rect 2156 5294 2158 5346
rect 2210 5294 2212 5346
rect 2156 5282 2212 5294
rect 1988 5142 2044 5236
rect 2268 5180 2324 5630
rect 1596 5068 1932 5124
rect 1988 5090 1990 5142
rect 2042 5090 2044 5142
rect 1988 5078 2044 5090
rect 2100 5124 2324 5180
rect 2548 5404 2604 5414
rect 1484 4902 1486 4954
rect 1538 4902 1540 4954
rect 1484 4890 1540 4902
rect 1708 4898 1764 4910
rect 1708 4846 1710 4898
rect 1762 4846 1764 4898
rect 1708 4620 1764 4846
rect 1708 4554 1764 4564
rect 1876 4406 1932 5068
rect 2100 4620 2156 5124
rect 2380 5122 2436 5134
rect 2380 5070 2382 5122
rect 2434 5070 2436 5122
rect 2212 5000 2268 5012
rect 2212 4948 2214 5000
rect 2266 4948 2268 5000
rect 2212 4732 2268 4948
rect 2380 4956 2436 5070
rect 2380 4890 2436 4900
rect 2548 4732 2604 5348
rect 2212 4666 2268 4676
rect 2324 4676 2604 4732
rect 2100 4554 2156 4564
rect 2212 4508 2268 4518
rect 2212 4408 2214 4452
rect 2266 4408 2268 4452
rect 1876 4394 1988 4406
rect 2212 4396 2268 4408
rect 1708 4338 1764 4350
rect 1876 4342 1934 4394
rect 1986 4342 1988 4394
rect 1876 4340 1988 4342
rect 1484 4284 1540 4294
rect 1484 4190 1540 4228
rect 1708 4286 1710 4338
rect 1762 4286 1764 4338
rect 1932 4330 1988 4340
rect 1708 4172 1764 4286
rect 2156 4284 2212 4294
rect 2324 4284 2380 4676
rect 2156 4282 2380 4284
rect 2156 4230 2158 4282
rect 2210 4230 2380 4282
rect 2156 4228 2380 4230
rect 2548 4508 2604 4518
rect 2156 4218 2212 4228
rect 1708 4106 1764 4116
rect 2380 4114 2436 4126
rect 1540 4060 1596 4070
rect 1540 3566 1596 4004
rect 2380 4062 2382 4114
rect 2434 4062 2436 4114
rect 1876 3778 1932 3790
rect 1540 3514 1542 3566
rect 1594 3514 1596 3566
rect 1540 3502 1596 3514
rect 1764 3724 1820 3734
rect 1764 3566 1820 3668
rect 1764 3514 1766 3566
rect 1818 3514 1820 3566
rect 1764 3276 1820 3514
rect 1876 3726 1878 3778
rect 1930 3726 1932 3778
rect 1876 3500 1932 3726
rect 2380 3724 2436 4062
rect 2380 3658 2436 3668
rect 2548 3612 2604 4452
rect 2660 3724 2716 6692
rect 2772 6076 2828 6086
rect 2772 5918 2828 6020
rect 2772 5866 2774 5918
rect 2826 5866 2828 5918
rect 2772 5854 2828 5866
rect 2996 5682 3052 7478
rect 3108 7432 3276 7488
rect 3892 7488 3948 7588
rect 3780 7474 3836 7486
rect 3108 7084 3164 7432
rect 3780 7422 3782 7474
rect 3834 7422 3836 7474
rect 3892 7474 4116 7488
rect 3892 7432 4062 7474
rect 3220 7308 3276 7318
rect 3220 7214 3276 7252
rect 3108 7018 3164 7028
rect 3780 6972 3836 7422
rect 4060 7422 4062 7432
rect 4114 7422 4116 7474
rect 4060 7420 4116 7422
rect 4060 7344 4116 7364
rect 4284 7474 4340 7588
rect 4284 7422 4286 7474
rect 4338 7422 4340 7474
rect 4284 6972 4340 7422
rect 3780 6916 4172 6972
rect 4284 6916 4396 6972
rect 4004 6748 4060 6758
rect 3444 6678 3500 6690
rect 3444 6636 3446 6678
rect 3498 6636 3500 6678
rect 3444 6570 3500 6580
rect 3724 6636 3780 6646
rect 3724 6542 3780 6580
rect 3108 6524 3164 6534
rect 3108 6522 3276 6524
rect 3108 6470 3110 6522
rect 3162 6470 3276 6522
rect 3108 6468 3276 6470
rect 3108 6458 3164 6468
rect 2996 5630 2998 5682
rect 3050 5630 3052 5682
rect 2996 5618 3052 5630
rect 3108 5894 3164 5906
rect 3108 5842 3110 5894
rect 3162 5842 3164 5894
rect 2996 5292 3052 5302
rect 2884 5068 2940 5078
rect 2884 4456 2940 5012
rect 2996 4966 3052 5236
rect 3108 5124 3164 5842
rect 3220 5292 3276 6468
rect 4004 5974 4060 6692
rect 3724 5964 3780 5974
rect 3556 5962 3780 5964
rect 3556 5910 3726 5962
rect 3778 5910 3780 5962
rect 3556 5908 3780 5910
rect 3220 5226 3276 5236
rect 3332 5894 3388 5906
rect 3332 5842 3334 5894
rect 3386 5842 3388 5894
rect 3332 5290 3388 5842
rect 3332 5238 3334 5290
rect 3386 5238 3388 5290
rect 3332 5226 3388 5238
rect 3444 5740 3500 5750
rect 3444 5136 3500 5684
rect 3108 5068 3220 5124
rect 3444 5084 3446 5136
rect 3498 5084 3500 5136
rect 3444 5072 3500 5084
rect 2996 4954 3108 4966
rect 2996 4902 3054 4954
rect 3106 4902 3108 4954
rect 2996 4900 3108 4902
rect 3052 4890 3108 4900
rect 3164 4742 3220 5068
rect 3276 4956 3332 4966
rect 3276 4954 3388 4956
rect 3276 4902 3278 4954
rect 3330 4902 3388 4954
rect 3276 4890 3388 4902
rect 2772 4396 2828 4406
rect 2884 4404 2886 4456
rect 2938 4404 2940 4456
rect 2884 4392 2940 4404
rect 2996 4732 3052 4742
rect 3164 4732 3276 4742
rect 3164 4676 3220 4732
rect 2772 4338 2828 4340
rect 2772 4286 2774 4338
rect 2826 4286 2828 4338
rect 2772 4274 2828 4286
rect 2996 3836 3052 4676
rect 3220 4666 3276 4676
rect 3332 4620 3388 4890
rect 3332 4554 3388 4564
rect 3556 4620 3612 5908
rect 3724 5898 3780 5908
rect 3948 5962 4060 5974
rect 3948 5910 3950 5962
rect 4002 5910 4060 5962
rect 3948 5908 4060 5910
rect 4116 6636 4172 6916
rect 3948 5898 4004 5908
rect 4116 5802 4172 6580
rect 4340 6412 4396 6916
rect 4452 6748 4508 7700
rect 4676 7308 4732 7318
rect 4452 6682 4508 6692
rect 4564 7306 4732 7308
rect 4564 7254 4678 7306
rect 4730 7254 4732 7306
rect 4564 7252 4732 7254
rect 4564 6746 4620 7252
rect 4676 7242 4732 7252
rect 4956 7306 5012 7318
rect 4956 7254 4958 7306
rect 5010 7254 5012 7306
rect 4956 7196 5012 7254
rect 4956 7130 5012 7140
rect 5348 7306 5404 7318
rect 5348 7254 5350 7306
rect 5402 7254 5404 7306
rect 5348 6860 5404 7254
rect 5460 7308 5516 8150
rect 6580 8150 6638 8202
rect 6690 8150 6692 8202
rect 6580 8138 6692 8150
rect 5684 7644 5740 7654
rect 5684 7486 5740 7588
rect 6580 7644 6636 8138
rect 6804 8092 6860 9818
rect 7756 9790 7812 9828
rect 8316 9826 8372 9940
rect 8708 9996 8764 10006
rect 8708 9902 8764 9940
rect 8316 9774 8318 9826
rect 8370 9774 8372 9826
rect 8316 9762 8372 9774
rect 8820 9772 8876 9782
rect 8260 9548 8316 9558
rect 8820 9548 8876 9716
rect 8036 9324 8092 9334
rect 7588 9212 7644 9222
rect 7588 9118 7644 9156
rect 7532 8988 7588 8998
rect 7532 8894 7588 8932
rect 7924 8988 7980 8998
rect 7924 8894 7980 8932
rect 7308 8818 7364 8830
rect 7308 8766 7310 8818
rect 7362 8766 7364 8818
rect 7308 8764 7364 8766
rect 7308 8698 7364 8708
rect 7420 8540 7476 8550
rect 7028 8316 7084 8326
rect 7028 8258 7084 8260
rect 7028 8206 7030 8258
rect 7082 8206 7084 8258
rect 7420 8314 7476 8484
rect 7420 8262 7422 8314
rect 7474 8262 7476 8314
rect 7420 8250 7476 8262
rect 7028 8194 7084 8206
rect 7084 8092 7140 8102
rect 6804 8090 7140 8092
rect 6804 8038 7086 8090
rect 7138 8038 7140 8090
rect 6804 8036 7140 8038
rect 7084 8026 7140 8036
rect 6804 7756 6860 7766
rect 6804 7654 6860 7700
rect 6804 7642 6916 7654
rect 6804 7590 6862 7642
rect 6914 7590 6916 7642
rect 6804 7588 6916 7590
rect 6580 7578 6636 7588
rect 6860 7578 6916 7588
rect 5684 7434 5686 7486
rect 5738 7434 5740 7486
rect 6020 7532 6076 7542
rect 6020 7438 6076 7476
rect 6692 7532 6748 7542
rect 6356 7456 6412 7468
rect 5684 7422 5740 7434
rect 5460 7242 5516 7252
rect 6356 7404 6358 7456
rect 6410 7404 6412 7456
rect 6356 7196 6412 7404
rect 6356 7130 6412 7140
rect 6468 7420 6524 7430
rect 6244 6860 6300 6870
rect 5348 6794 5404 6804
rect 5460 6802 5516 6814
rect 4564 6694 4566 6746
rect 4618 6694 4620 6746
rect 5460 6750 5462 6802
rect 5514 6750 5516 6802
rect 4564 6682 4620 6694
rect 5236 6690 5292 6702
rect 5236 6638 5238 6690
rect 5290 6638 5292 6690
rect 5236 6524 5292 6638
rect 5236 6458 5292 6468
rect 4340 6346 4396 6356
rect 4958 6300 5222 6310
rect 5014 6244 5062 6300
rect 5118 6244 5166 6300
rect 5460 6300 5516 6750
rect 6244 6802 6300 6804
rect 6244 6750 6246 6802
rect 6298 6750 6300 6802
rect 6244 6738 6300 6750
rect 6132 6690 6188 6702
rect 5684 6636 5740 6646
rect 5684 6578 5740 6580
rect 5684 6526 5686 6578
rect 5738 6526 5740 6578
rect 6132 6638 6134 6690
rect 6186 6638 6188 6690
rect 6132 6636 6188 6638
rect 6132 6570 6188 6580
rect 5684 6514 5740 6526
rect 6188 6412 6244 6422
rect 5460 6244 5908 6300
rect 4958 6234 5222 6244
rect 4732 6076 4788 6086
rect 4732 5982 4788 6020
rect 5852 6074 5908 6244
rect 5852 6022 5854 6074
rect 5906 6022 5908 6074
rect 5852 6010 5908 6022
rect 4116 5750 4118 5802
rect 4170 5750 4172 5802
rect 4116 5738 4172 5750
rect 4340 5906 4396 5918
rect 4340 5854 4342 5906
rect 4394 5854 4396 5906
rect 3836 5180 3892 5190
rect 3836 5086 3892 5124
rect 3556 4462 3612 4564
rect 3332 4406 3612 4462
rect 3668 4956 3724 4966
rect 4172 4956 4228 4966
rect 2772 3724 2828 3734
rect 2660 3722 2828 3724
rect 2660 3670 2774 3722
rect 2826 3670 2828 3722
rect 2660 3668 2828 3670
rect 2772 3658 2828 3668
rect 2548 3568 2716 3612
rect 2548 3556 2772 3568
rect 2660 3554 2772 3556
rect 1876 3434 1932 3444
rect 2100 3542 2156 3554
rect 2100 3490 2102 3542
rect 2154 3490 2156 3542
rect 2660 3512 2718 3554
rect 1764 3220 2044 3276
rect 1484 2828 1540 2838
rect 1316 2826 1540 2828
rect 1316 2774 1486 2826
rect 1538 2774 1540 2826
rect 1316 2772 1540 2774
rect 1484 2762 1540 2772
rect 1204 2548 1596 2604
rect 868 700 924 2548
rect 1540 1202 1596 2548
rect 1988 2380 2044 3220
rect 2100 2546 2156 3490
rect 2436 3500 2492 3510
rect 2716 3502 2718 3512
rect 2770 3502 2772 3554
rect 2492 3444 2548 3500
rect 2716 3490 2772 3502
rect 2996 3554 3052 3780
rect 3164 4282 3220 4294
rect 3164 4230 3166 4282
rect 3218 4230 3220 4282
rect 3164 3724 3220 4230
rect 3332 4060 3388 4406
rect 3500 4226 3556 4238
rect 3500 4174 3502 4226
rect 3554 4174 3556 4226
rect 3500 4172 3556 4174
rect 3500 4116 3612 4172
rect 3332 3994 3388 4004
rect 3332 3724 3388 3734
rect 3556 3724 3612 4116
rect 3668 4060 3724 4900
rect 4004 4954 4228 4956
rect 4004 4902 4174 4954
rect 4226 4902 4228 4954
rect 4004 4900 4228 4902
rect 4004 4732 4060 4900
rect 4172 4890 4228 4900
rect 3892 4676 4060 4732
rect 3780 4396 3836 4406
rect 3780 4298 3782 4340
rect 3834 4298 3836 4340
rect 3780 4286 3836 4298
rect 3892 4172 3948 4676
rect 4004 4542 4060 4554
rect 4004 4508 4006 4542
rect 4058 4508 4060 4542
rect 4004 4442 4060 4452
rect 4116 4326 4172 4338
rect 4116 4274 4118 4326
rect 4170 4274 4172 4326
rect 3892 4116 4060 4172
rect 3668 4004 3948 4060
rect 3164 3722 3612 3724
rect 3164 3670 3334 3722
rect 3386 3670 3612 3722
rect 3164 3668 3612 3670
rect 3332 3658 3388 3668
rect 2996 3502 2998 3554
rect 3050 3502 3052 3554
rect 2996 3490 3052 3502
rect 2436 3434 2548 3444
rect 2492 3386 2548 3434
rect 2492 3334 2494 3386
rect 2546 3334 2548 3386
rect 2492 3322 2548 3334
rect 2660 2826 2716 2838
rect 2100 2494 2102 2546
rect 2154 2494 2156 2546
rect 2100 2482 2156 2494
rect 2436 2770 2492 2782
rect 2436 2718 2438 2770
rect 2490 2718 2492 2770
rect 1988 2324 2156 2380
rect 2100 2098 2156 2324
rect 2100 2046 2102 2098
rect 2154 2046 2156 2098
rect 2100 2034 2156 2046
rect 2436 1932 2492 2718
rect 2660 2774 2662 2826
rect 2714 2774 2716 2826
rect 2660 2492 2716 2774
rect 3220 2604 3276 2614
rect 3220 2510 3276 2548
rect 2660 2426 2716 2436
rect 3332 2380 3388 2390
rect 3332 2042 3388 2324
rect 3892 2156 3948 4004
rect 4004 2380 4060 4116
rect 4116 3836 4172 4274
rect 4228 4172 4284 4182
rect 4340 4172 4396 5854
rect 6188 5850 6244 6356
rect 6468 6086 6524 7364
rect 6692 6746 6748 7476
rect 6804 7418 6860 7430
rect 6804 7366 6806 7418
rect 6858 7366 6860 7418
rect 6804 6972 6860 7366
rect 7252 7420 7308 7430
rect 6972 7306 7028 7318
rect 6972 7254 6974 7306
rect 7026 7254 7028 7306
rect 6972 7084 7028 7254
rect 6972 7018 7028 7028
rect 6804 6906 6860 6916
rect 7252 6883 7308 7364
rect 8036 7418 8092 9268
rect 8148 9212 8204 9222
rect 8148 8986 8204 9156
rect 8148 8934 8150 8986
rect 8202 8934 8204 8986
rect 8148 8922 8204 8934
rect 8260 8876 8316 9492
rect 8764 9492 8876 9548
rect 8764 9042 8820 9492
rect 9268 9100 9324 10388
rect 9492 10220 9548 10714
rect 9940 10622 9996 10948
rect 10332 10892 10388 10902
rect 9940 10570 9942 10622
rect 9994 10570 9996 10622
rect 10164 10720 10220 10732
rect 10164 10668 10166 10720
rect 10218 10668 10220 10720
rect 10164 10602 10220 10612
rect 10332 10610 10388 10836
rect 9940 10558 9996 10570
rect 10332 10558 10334 10610
rect 10386 10558 10388 10610
rect 10332 10546 10388 10558
rect 10108 10388 10164 10398
rect 10108 10386 10220 10388
rect 10108 10334 10110 10386
rect 10162 10334 10220 10386
rect 10108 10322 10220 10334
rect 10052 10220 10108 10230
rect 9492 10164 9716 10220
rect 9660 10050 9716 10164
rect 9660 9998 9662 10050
rect 9714 9998 9716 10050
rect 9660 9986 9716 9998
rect 9436 9884 9492 9894
rect 9436 9790 9492 9828
rect 10052 9882 10108 10164
rect 10164 9996 10220 10322
rect 10164 9930 10220 9940
rect 10276 10108 10332 10118
rect 10052 9830 10054 9882
rect 10106 9830 10108 9882
rect 10052 9818 10108 9830
rect 10164 9772 10220 9782
rect 9604 9660 9660 9670
rect 9604 9566 9660 9604
rect 10052 9212 10108 9222
rect 10164 9212 10220 9716
rect 10052 9210 10220 9212
rect 10052 9158 10054 9210
rect 10106 9158 10220 9210
rect 10052 9156 10220 9158
rect 10276 9210 10332 10052
rect 10276 9158 10278 9210
rect 10330 9158 10332 9210
rect 10052 9146 10108 9156
rect 9268 9044 9436 9100
rect 8148 8764 8204 8774
rect 8148 8270 8204 8708
rect 8148 8218 8150 8270
rect 8202 8218 8204 8270
rect 8260 8316 8316 8820
rect 8372 8988 8428 8998
rect 8764 8990 8766 9042
rect 8818 8990 8820 9042
rect 8764 8978 8820 8990
rect 8372 8508 8428 8932
rect 8540 8876 8596 8896
rect 8540 8818 8596 8820
rect 8540 8766 8542 8818
rect 8594 8766 8596 8818
rect 8540 8764 8596 8766
rect 8372 8456 8374 8508
rect 8426 8456 8428 8508
rect 8372 8444 8428 8456
rect 8484 8708 8596 8764
rect 8652 8874 8708 8886
rect 8652 8822 8654 8874
rect 8706 8822 8708 8874
rect 8484 8428 8540 8708
rect 8652 8652 8708 8822
rect 9100 8876 9156 8886
rect 9100 8782 9156 8820
rect 9212 8876 9268 8886
rect 9212 8874 9324 8876
rect 9212 8822 9214 8874
rect 9266 8822 9324 8874
rect 9212 8810 9324 8822
rect 8484 8362 8540 8372
rect 8596 8596 8708 8652
rect 8928 8652 9192 8662
rect 8984 8596 9032 8652
rect 9088 8596 9136 8652
rect 8260 8260 8428 8316
rect 8148 8206 8204 8218
rect 8372 8204 8428 8260
rect 8484 8246 8540 8258
rect 8484 8204 8486 8246
rect 8372 8194 8486 8204
rect 8538 8194 8540 8246
rect 8372 8148 8540 8194
rect 8596 7486 8652 8596
rect 8928 8586 9192 8596
rect 9268 8652 9324 8810
rect 9268 8586 9324 8596
rect 9380 8270 9436 9044
rect 9772 8874 9828 8886
rect 9772 8822 9774 8874
rect 9826 8822 9828 8874
rect 9772 8652 9828 8822
rect 9772 8586 9828 8596
rect 10276 8540 10332 9158
rect 10500 9210 10556 11284
rect 11060 11004 11116 11396
rect 10780 10948 11116 11004
rect 11228 11394 11284 11406
rect 11228 11342 11230 11394
rect 11282 11342 11284 11394
rect 10780 10778 10836 10948
rect 11228 10892 11284 11342
rect 11396 11340 11452 11350
rect 11396 11246 11452 11284
rect 11508 11228 11564 11238
rect 10780 10726 10782 10778
rect 10834 10726 10836 10778
rect 10780 10108 10836 10726
rect 11060 10836 11284 10892
rect 11396 10892 11452 10902
rect 10892 10444 10948 10454
rect 10892 10350 10948 10388
rect 10780 10042 10836 10052
rect 11060 9996 11116 10836
rect 11396 10666 11452 10836
rect 11396 10614 11398 10666
rect 11450 10614 11452 10666
rect 11396 10602 11452 10614
rect 11396 10532 11452 10544
rect 11396 10480 11398 10532
rect 11450 10480 11452 10532
rect 11228 10442 11284 10454
rect 11228 10390 11230 10442
rect 11282 10390 11284 10442
rect 11228 10108 11284 10390
rect 11396 10444 11452 10480
rect 11508 10444 11564 11172
rect 11396 10388 11564 10444
rect 11228 10042 11284 10052
rect 11620 10108 11676 11508
rect 11844 11450 11900 11732
rect 11844 11398 11846 11450
rect 11898 11398 11900 11450
rect 11844 11386 11900 11398
rect 12012 11394 12068 11406
rect 12012 11342 12014 11394
rect 12066 11342 12068 11394
rect 12012 11340 12068 11342
rect 12012 11274 12068 11284
rect 11900 11228 11956 11238
rect 11844 11226 11956 11228
rect 11844 11174 11902 11226
rect 11954 11174 11956 11226
rect 11844 11162 11956 11174
rect 11844 10780 11900 11162
rect 11732 10724 11900 10780
rect 12012 10780 12068 10790
rect 12292 10780 12348 12740
rect 12516 12236 12572 14420
rect 12740 13814 12796 17444
rect 12852 17434 12908 17444
rect 12898 17276 13162 17286
rect 12954 17220 13002 17276
rect 13058 17220 13106 17276
rect 12898 17210 13162 17220
rect 13300 16940 13356 16950
rect 13300 16882 13356 16884
rect 13300 16830 13302 16882
rect 13354 16830 13356 16882
rect 13300 16818 13356 16830
rect 12908 16716 12964 16726
rect 12908 16622 12964 16660
rect 13748 16380 13804 17546
rect 14980 17537 15036 17549
rect 14980 17485 14982 17537
rect 15034 17485 15036 17537
rect 13748 16314 13804 16324
rect 14140 16940 14196 16950
rect 14140 16714 14196 16884
rect 14980 16938 15036 17485
rect 14980 16886 14982 16938
rect 15034 16886 15036 16938
rect 14980 16874 15036 16886
rect 15092 17500 15148 17510
rect 15092 16716 15148 17444
rect 15428 16828 15484 17612
rect 15428 16762 15484 16772
rect 15540 16826 15596 16838
rect 15540 16774 15542 16826
rect 15594 16774 15596 16826
rect 14140 16662 14142 16714
rect 14194 16662 14196 16714
rect 14140 16380 14196 16662
rect 14140 16314 14196 16324
rect 14868 16660 15148 16716
rect 15260 16716 15316 16726
rect 15260 16714 15372 16716
rect 15260 16662 15262 16714
rect 15314 16662 15372 16714
rect 14868 16604 14924 16660
rect 15260 16650 15372 16662
rect 14868 16266 14924 16548
rect 14868 16214 14870 16266
rect 14922 16214 14924 16266
rect 14868 16202 14924 16214
rect 14644 16154 14700 16166
rect 13300 16098 13356 16110
rect 13300 16046 13302 16098
rect 13354 16046 13356 16098
rect 12898 15708 13162 15718
rect 12954 15652 13002 15708
rect 13058 15652 13106 15708
rect 12898 15642 13162 15652
rect 13300 14812 13356 16046
rect 13524 16098 13580 16110
rect 13524 16046 13526 16098
rect 13578 16046 13580 16098
rect 13412 15258 13468 15270
rect 13412 15206 13414 15258
rect 13466 15206 13468 15258
rect 13412 15148 13468 15206
rect 13412 15082 13468 15092
rect 13300 14746 13356 14756
rect 13188 14700 13244 14710
rect 13188 14606 13244 14644
rect 12852 14586 12908 14598
rect 12852 14534 12854 14586
rect 12906 14534 12908 14586
rect 12852 14476 12908 14534
rect 12852 14410 12908 14420
rect 13524 14364 13580 16046
rect 14644 16102 14646 16154
rect 14698 16102 14700 16154
rect 13748 15596 13804 15606
rect 13748 15482 13804 15540
rect 14644 15596 14700 16102
rect 14644 15530 14700 15540
rect 14980 16156 15036 16166
rect 13748 15430 13750 15482
rect 13802 15430 13804 15482
rect 13748 15418 13804 15430
rect 14364 15484 14420 15494
rect 14980 15484 15036 16100
rect 14364 15426 14420 15428
rect 14364 15374 14366 15426
rect 14418 15374 14420 15426
rect 14756 15482 15036 15484
rect 14756 15430 14982 15482
rect 15034 15430 15036 15482
rect 14756 15428 15036 15430
rect 14364 15362 14420 15374
rect 14588 15372 14644 15382
rect 14588 15278 14644 15316
rect 13804 15260 13860 15270
rect 13804 15166 13860 15204
rect 13636 15148 13692 15158
rect 14756 15148 14812 15428
rect 14980 15418 15036 15428
rect 15092 15820 15148 15830
rect 13636 14700 13692 15092
rect 14028 15090 14084 15102
rect 14028 15038 14030 15090
rect 14082 15038 14084 15090
rect 14028 14812 14084 15038
rect 14028 14746 14084 14756
rect 14644 15092 14812 15148
rect 14308 14700 14364 14710
rect 13636 14644 13860 14700
rect 13804 14530 13860 14644
rect 14028 14588 14084 14598
rect 13524 14298 13580 14308
rect 13636 14518 13692 14530
rect 13636 14466 13638 14518
rect 13690 14466 13692 14518
rect 12898 14140 13162 14150
rect 13636 14140 13692 14466
rect 12954 14084 13002 14140
rect 13058 14084 13106 14140
rect 12898 14074 13162 14084
rect 13412 14084 13692 14140
rect 13804 14478 13806 14530
rect 13858 14478 13860 14530
rect 12684 13802 12796 13814
rect 12684 13750 12686 13802
rect 12738 13750 12796 13802
rect 12684 13748 12796 13750
rect 13412 13804 13468 14084
rect 13804 14028 13860 14478
rect 12684 13738 12740 13748
rect 13412 13738 13468 13748
rect 13524 13972 13860 14028
rect 13972 14586 14084 14588
rect 13972 14534 14030 14586
rect 14082 14534 14084 14586
rect 13972 14522 14084 14534
rect 14308 14530 14364 14644
rect 14644 14664 14700 15092
rect 14644 14612 14646 14664
rect 14698 14612 14700 14664
rect 14644 14600 14700 14612
rect 13524 13590 13580 13972
rect 13636 13804 13692 13842
rect 13636 13738 13692 13748
rect 13972 13748 14028 14522
rect 14308 14478 14310 14530
rect 14362 14478 14364 14530
rect 14756 14530 14812 14542
rect 14084 14406 14140 14418
rect 14084 14364 14086 14406
rect 14138 14364 14140 14406
rect 14084 14298 14140 14308
rect 14084 13748 14140 13758
rect 13972 13746 14140 13748
rect 13972 13694 14086 13746
rect 14138 13694 14140 13746
rect 13972 13692 14140 13694
rect 13468 13580 13580 13590
rect 13412 13578 13580 13580
rect 13412 13526 13470 13578
rect 13522 13526 13580 13578
rect 13412 13524 13580 13526
rect 13636 13668 13692 13680
rect 13636 13616 13638 13668
rect 13690 13616 13692 13668
rect 13412 13514 13524 13524
rect 13300 13356 13356 13366
rect 13300 12970 13356 13300
rect 13300 12918 13302 12970
rect 13354 12918 13356 12970
rect 12628 12906 12684 12918
rect 13300 12906 13356 12918
rect 12628 12854 12630 12906
rect 12682 12854 12684 12906
rect 12628 12460 12684 12854
rect 13020 12796 13076 12834
rect 13412 12806 13468 13514
rect 13636 13244 13692 13616
rect 13636 13178 13692 13188
rect 13972 12950 14028 12962
rect 13972 12898 13974 12950
rect 14026 12898 14028 12950
rect 13020 12730 13076 12740
rect 13356 12794 13468 12806
rect 13356 12742 13358 12794
rect 13410 12742 13468 12794
rect 13356 12740 13468 12742
rect 13636 12794 13692 12806
rect 13636 12742 13638 12794
rect 13690 12742 13692 12794
rect 13356 12730 13412 12740
rect 13636 12684 13692 12742
rect 13524 12628 13636 12684
rect 12898 12572 13162 12582
rect 12954 12516 13002 12572
rect 13058 12516 13106 12572
rect 12898 12506 13162 12516
rect 12628 12394 12684 12404
rect 12516 12142 12572 12180
rect 13412 12234 13468 12246
rect 13412 12182 13414 12234
rect 13466 12182 13468 12234
rect 12796 12010 12852 12022
rect 12796 11958 12798 12010
rect 12850 11958 12852 12010
rect 12796 11900 12852 11958
rect 12796 11834 12852 11844
rect 12740 11676 12796 11686
rect 13412 11676 13468 12182
rect 12740 11574 12796 11620
rect 13300 11620 13468 11676
rect 12684 11562 12796 11574
rect 12684 11510 12686 11562
rect 12738 11510 12796 11562
rect 12684 11508 12796 11510
rect 12964 11564 13020 11574
rect 12684 11498 12740 11508
rect 12964 11394 13020 11508
rect 12012 10778 12348 10780
rect 12012 10726 12014 10778
rect 12066 10726 12348 10778
rect 12012 10724 12348 10726
rect 12404 11340 12460 11350
rect 12964 11342 12966 11394
rect 13018 11342 13020 11394
rect 13300 11452 13356 11620
rect 13524 11564 13580 12628
rect 13636 12618 13692 12628
rect 13748 12796 13804 12806
rect 13972 12796 14028 12898
rect 13804 12740 14028 12796
rect 13748 12178 13804 12740
rect 14084 12572 14140 13692
rect 14196 13634 14252 13646
rect 14196 13582 14198 13634
rect 14250 13582 14252 13634
rect 14196 13244 14252 13582
rect 14196 13020 14252 13188
rect 14196 12954 14252 12964
rect 14308 12908 14364 14478
rect 14532 14476 14588 14486
rect 14532 13580 14588 14420
rect 14532 13514 14588 13524
rect 14756 14478 14758 14530
rect 14810 14478 14812 14530
rect 14756 13690 14812 14478
rect 15092 14028 15148 15764
rect 15316 15372 15372 16650
rect 15540 16268 15596 16774
rect 15652 16380 15708 18676
rect 15820 18508 15876 18518
rect 15820 18450 15876 18452
rect 15820 18398 15822 18450
rect 15874 18398 15876 18450
rect 15988 18506 16044 18900
rect 16548 18732 16604 18742
rect 16548 18630 16604 18676
rect 16492 18618 16604 18630
rect 16492 18566 16494 18618
rect 16546 18566 16604 18618
rect 16492 18564 16604 18566
rect 16492 18554 16548 18564
rect 15988 18454 15990 18506
rect 16042 18454 16044 18506
rect 15988 18442 16044 18454
rect 16884 18508 16940 19200
rect 18004 18620 18060 18630
rect 16884 18462 17276 18508
rect 16884 18452 17222 18462
rect 15820 18386 15876 18398
rect 16436 18396 16492 18434
rect 17220 18410 17222 18452
rect 17274 18410 17276 18462
rect 18004 18506 18060 18564
rect 18004 18454 18006 18506
rect 18058 18454 18060 18506
rect 18004 18442 18060 18454
rect 19236 18620 19292 18630
rect 19236 18450 19292 18564
rect 15988 18372 16044 18384
rect 15988 18320 15990 18372
rect 16042 18320 16044 18372
rect 16436 18330 16492 18340
rect 16604 18396 16660 18406
rect 15820 17724 15932 17734
rect 15820 17722 15876 17724
rect 15820 17670 15822 17722
rect 15874 17670 15876 17722
rect 15820 17668 15876 17670
rect 15820 17658 15932 17668
rect 15988 17050 16044 18320
rect 16604 18302 16660 18340
rect 16212 18284 16268 18294
rect 16100 17724 16156 17734
rect 16100 17630 16156 17668
rect 16212 17500 16268 18228
rect 16436 18172 16492 18182
rect 16212 17434 16268 17444
rect 16324 18060 16380 18070
rect 15988 16998 15990 17050
rect 16042 16998 16044 17050
rect 15988 16986 16044 16998
rect 16324 16716 16380 18004
rect 16436 17834 16492 18116
rect 16868 18060 17132 18070
rect 16924 18004 16972 18060
rect 17028 18004 17076 18060
rect 16868 17994 17132 18004
rect 16436 17782 16438 17834
rect 16490 17782 16492 17834
rect 16436 17770 16492 17782
rect 17220 17846 17276 18410
rect 18228 18396 18340 18406
rect 18004 18372 18060 18384
rect 18004 18320 18006 18372
rect 18058 18320 18060 18372
rect 18284 18394 18340 18396
rect 18284 18342 18286 18394
rect 18338 18342 18340 18394
rect 18284 18340 18340 18342
rect 18228 18330 18340 18340
rect 18452 18394 18508 18406
rect 18452 18342 18454 18394
rect 18506 18342 18508 18394
rect 17556 18284 17612 18294
rect 17836 18284 17892 18294
rect 17556 18282 17892 18284
rect 17556 18230 17558 18282
rect 17610 18230 17838 18282
rect 17890 18230 17892 18282
rect 17556 18228 17892 18230
rect 17556 18218 17612 18228
rect 17836 18218 17892 18228
rect 18004 18172 18060 18320
rect 18452 18172 18508 18342
rect 18620 18396 18676 18406
rect 18620 18302 18676 18340
rect 19236 18398 19238 18450
rect 19290 18398 19292 18450
rect 19460 18508 19516 19200
rect 21868 18956 21924 18966
rect 20838 18844 21102 18854
rect 20894 18788 20942 18844
rect 20998 18788 21046 18844
rect 20838 18778 21102 18788
rect 21868 18618 21924 18900
rect 22148 18732 22204 19200
rect 22148 18676 22652 18732
rect 21868 18566 21870 18618
rect 21922 18566 21924 18618
rect 21868 18554 21924 18566
rect 19460 18442 19516 18452
rect 21140 18508 21196 18518
rect 21140 18410 21142 18452
rect 21194 18410 21196 18452
rect 18060 18116 18508 18172
rect 18004 18106 18060 18116
rect 17220 17834 17332 17846
rect 17220 17782 17278 17834
rect 17330 17782 17332 17834
rect 17220 17780 17332 17782
rect 17276 17770 17332 17780
rect 17668 17724 17724 17734
rect 17444 17722 17724 17724
rect 17444 17670 17670 17722
rect 17722 17670 17724 17722
rect 17444 17668 17724 17670
rect 16828 17612 16884 17622
rect 16828 17610 16940 17612
rect 16828 17558 16830 17610
rect 16882 17558 16940 17610
rect 16828 17546 16940 17558
rect 16772 17052 16828 17062
rect 16772 16884 16828 16996
rect 16660 16828 16828 16884
rect 16436 16716 16492 16726
rect 16324 16714 16492 16716
rect 15932 16658 15988 16670
rect 15932 16606 15934 16658
rect 15986 16606 15988 16658
rect 15652 16324 15764 16380
rect 15428 16212 15596 16268
rect 15708 16266 15764 16324
rect 15708 16214 15710 16266
rect 15762 16214 15764 16266
rect 15428 15820 15484 16212
rect 15708 16202 15764 16214
rect 15820 16268 15876 16278
rect 15820 16174 15876 16212
rect 15932 16156 15988 16606
rect 16156 16658 16212 16670
rect 16324 16662 16438 16714
rect 16490 16662 16492 16714
rect 16324 16660 16492 16662
rect 16156 16606 16158 16658
rect 16210 16606 16212 16658
rect 16436 16650 16492 16660
rect 16156 16380 16212 16606
rect 15596 16098 15652 16110
rect 15596 16046 15598 16098
rect 15650 16046 15652 16098
rect 15932 16090 15988 16100
rect 16100 16324 16212 16380
rect 16660 16380 16716 16828
rect 16772 16716 16828 16726
rect 16884 16716 16940 17546
rect 17220 16940 17276 16950
rect 17220 16842 17222 16884
rect 17274 16842 17276 16884
rect 17220 16830 17276 16842
rect 16828 16660 16940 16716
rect 16772 16622 16828 16660
rect 17444 16604 17500 17668
rect 17668 17658 17724 17668
rect 17836 17724 17892 17734
rect 18060 17724 18116 17734
rect 17836 17722 18116 17724
rect 17836 17670 17838 17722
rect 17890 17670 18062 17722
rect 18114 17670 18116 17722
rect 17836 17668 18116 17670
rect 17836 17658 17892 17668
rect 18060 17658 18116 17668
rect 18228 17722 18284 18116
rect 18228 17670 18230 17722
rect 18282 17670 18284 17722
rect 18228 17658 18284 17670
rect 18396 17724 18452 17734
rect 18396 17630 18452 17668
rect 18788 17612 18844 17622
rect 18564 17556 18788 17612
rect 17724 17500 17836 17510
rect 17724 17498 17780 17500
rect 17724 17446 17726 17498
rect 17778 17446 17780 17498
rect 17724 17444 17780 17446
rect 17724 17434 17836 17444
rect 17836 17276 17892 17286
rect 17836 16882 17892 17220
rect 17836 16830 17838 16882
rect 17890 16830 17892 16882
rect 18004 16940 18060 16978
rect 18004 16874 18060 16884
rect 18564 16938 18620 17556
rect 18788 17518 18844 17556
rect 19236 17500 19292 18398
rect 20580 18394 20636 18406
rect 21140 18398 21196 18410
rect 22596 18508 22652 18676
rect 23100 18620 23156 18630
rect 23100 18526 23156 18564
rect 22596 18410 22598 18452
rect 22650 18410 22652 18452
rect 23996 18508 24052 18518
rect 23996 18414 24052 18452
rect 24556 18508 24612 18518
rect 24724 18508 24780 19200
rect 26740 18956 26796 18966
rect 25788 18732 25844 18742
rect 25788 18618 25844 18676
rect 25788 18566 25790 18618
rect 25842 18566 25844 18618
rect 25788 18554 25844 18566
rect 24556 18506 25004 18508
rect 24556 18454 24558 18506
rect 24610 18454 25004 18506
rect 24556 18452 25004 18454
rect 24556 18442 24612 18452
rect 20580 18342 20582 18394
rect 20634 18342 20636 18394
rect 22596 18376 22652 18410
rect 24948 18406 25004 18452
rect 23772 18396 23828 18406
rect 19740 18282 19796 18294
rect 19740 18230 19742 18282
rect 19794 18230 19796 18282
rect 19516 17836 19572 17846
rect 19516 17742 19572 17780
rect 19740 17836 19796 18230
rect 20020 18284 20076 18294
rect 19740 17770 19796 17780
rect 19908 18172 19964 18182
rect 19236 17434 19292 17444
rect 18564 16886 18566 16938
rect 18618 16886 18620 16938
rect 17836 16818 17892 16830
rect 18004 16804 18060 16816
rect 18004 16752 18006 16804
rect 18058 16752 18060 16804
rect 17556 16716 17612 16726
rect 17556 16622 17612 16660
rect 17220 16548 17500 16604
rect 16868 16492 17132 16502
rect 16924 16436 16972 16492
rect 17028 16436 17076 16492
rect 16868 16426 17132 16436
rect 16660 16324 16828 16380
rect 15596 15932 15652 16046
rect 16100 15932 16156 16324
rect 16772 16176 16828 16324
rect 15596 15876 16156 15932
rect 15428 15754 15484 15764
rect 15204 15300 15260 15312
rect 15316 15306 15372 15316
rect 15652 15596 15708 15606
rect 15204 15248 15206 15300
rect 15258 15248 15260 15300
rect 15204 15148 15260 15248
rect 15652 15260 15708 15540
rect 16100 15484 16156 15876
rect 16212 16154 16268 16166
rect 16212 16102 16214 16154
rect 16266 16102 16268 16154
rect 16772 16124 16774 16176
rect 16826 16124 16828 16176
rect 16772 16112 16828 16124
rect 16212 15820 16268 16102
rect 16212 15596 16268 15764
rect 16212 15530 16268 15540
rect 16604 16098 16660 16110
rect 16604 16046 16606 16098
rect 16658 16046 16660 16098
rect 15764 15426 15820 15438
rect 15764 15374 15766 15426
rect 15818 15374 15820 15426
rect 16100 15418 16156 15428
rect 16324 15484 16380 15494
rect 15764 15372 15820 15374
rect 16324 15372 16380 15428
rect 15764 15316 15932 15372
rect 15876 15260 15932 15316
rect 16156 15314 16212 15326
rect 16156 15262 16158 15314
rect 16210 15262 16212 15314
rect 16156 15260 16212 15262
rect 15876 15204 16212 15260
rect 16268 15316 16380 15372
rect 16268 15314 16324 15316
rect 16268 15262 16270 15314
rect 16322 15262 16324 15314
rect 16268 15250 16324 15262
rect 15652 15158 15708 15204
rect 15484 15147 15540 15158
rect 15204 15082 15260 15092
rect 15428 15146 15540 15147
rect 15428 15094 15486 15146
rect 15538 15094 15540 15146
rect 15428 15082 15540 15094
rect 15652 15146 15764 15158
rect 16492 15147 16548 15158
rect 15652 15094 15710 15146
rect 15762 15094 15764 15146
rect 15652 15091 15764 15094
rect 15092 13962 15148 13972
rect 15204 14476 15260 14486
rect 14756 13638 14758 13690
rect 14810 13638 14812 13690
rect 14756 13580 14812 13638
rect 15204 13804 15260 14420
rect 15316 14364 15372 14374
rect 15428 14364 15484 15082
rect 15540 14924 15596 14934
rect 15540 14530 15596 14868
rect 15708 14700 15764 15091
rect 16436 15146 16548 15147
rect 16436 15094 16494 15146
rect 16546 15094 16548 15146
rect 16436 15082 16548 15094
rect 16324 15036 16380 15046
rect 15708 14644 16268 14700
rect 15540 14478 15542 14530
rect 15594 14478 15596 14530
rect 16100 14530 16156 14542
rect 16100 14520 16102 14530
rect 15540 14466 15596 14478
rect 15652 14478 16102 14520
rect 16154 14478 16156 14530
rect 15652 14464 16156 14478
rect 15652 14364 15708 14464
rect 15428 14308 15708 14364
rect 15316 13868 15372 14308
rect 15316 13816 15318 13868
rect 15370 13816 15372 13868
rect 15316 13804 15372 13816
rect 15204 13702 15260 13748
rect 15428 13740 15484 13752
rect 15204 13690 15316 13702
rect 15204 13638 15262 13690
rect 15314 13638 15316 13690
rect 15204 13636 15316 13638
rect 15260 13626 15316 13636
rect 15428 13692 15430 13740
rect 15482 13692 15484 13740
rect 15428 13626 15484 13636
rect 14756 13514 14812 13524
rect 15036 13580 15092 13590
rect 15036 13486 15092 13524
rect 15540 13468 15596 14308
rect 16100 14028 16156 14038
rect 15988 13804 16044 13814
rect 15764 13746 15820 13758
rect 15764 13694 15766 13746
rect 15818 13694 15820 13746
rect 15316 13412 15596 13468
rect 15652 13468 15708 13478
rect 14756 13356 14812 13366
rect 14644 13244 14700 13254
rect 14644 12962 14700 13188
rect 14756 13186 14812 13300
rect 14756 13134 14758 13186
rect 14810 13134 14812 13186
rect 14756 13122 14812 13134
rect 14644 12910 14646 12962
rect 14698 12910 14700 12962
rect 14308 12842 14364 12852
rect 14532 12850 14588 12862
rect 14532 12798 14534 12850
rect 14586 12798 14588 12850
rect 14532 12796 14588 12798
rect 14532 12730 14588 12740
rect 14084 12506 14140 12516
rect 13748 12126 13750 12178
rect 13802 12126 13804 12178
rect 13748 12114 13804 12126
rect 14364 12124 14476 12134
rect 14364 12122 14420 12124
rect 14364 12070 14366 12122
rect 14418 12070 14420 12122
rect 14364 12068 14420 12070
rect 14364 12058 14476 12068
rect 13300 11386 13356 11396
rect 13412 11496 13468 11508
rect 13524 11498 13580 11508
rect 14308 11564 14364 11574
rect 13412 11444 13414 11496
rect 13466 11444 13468 11496
rect 12964 11330 13020 11342
rect 11732 10220 11788 10724
rect 12012 10714 12068 10724
rect 12292 10596 12348 10608
rect 12292 10544 12294 10596
rect 12346 10544 12348 10596
rect 11732 10154 11788 10164
rect 11900 10498 11956 10510
rect 11900 10446 11902 10498
rect 11954 10446 11956 10498
rect 11620 10042 11676 10052
rect 11900 10108 11956 10446
rect 11900 10042 11956 10052
rect 11060 9930 11116 9940
rect 12068 9904 12236 9940
rect 11508 9882 11564 9894
rect 11508 9830 11510 9882
rect 11562 9830 11564 9882
rect 11508 9772 11564 9830
rect 11508 9706 11564 9716
rect 11732 9884 11788 9894
rect 12068 9852 12070 9904
rect 12122 9884 12236 9904
rect 12122 9852 12124 9884
rect 12068 9840 12124 9852
rect 11172 9658 11228 9670
rect 11172 9606 11174 9658
rect 11226 9606 11228 9658
rect 11172 9548 11228 9606
rect 11172 9482 11228 9492
rect 10500 9158 10502 9210
rect 10554 9158 10556 9210
rect 10500 9146 10556 9158
rect 11732 9160 11788 9828
rect 11900 9826 11956 9838
rect 11900 9774 11902 9826
rect 11954 9774 11956 9826
rect 11900 9660 11956 9774
rect 11900 9594 11956 9604
rect 12068 9770 12124 9782
rect 12068 9718 12070 9770
rect 12122 9718 12124 9770
rect 11732 9108 11734 9160
rect 11786 9108 11788 9160
rect 11900 9324 11956 9334
rect 11900 9210 11956 9268
rect 11900 9158 11902 9210
rect 11954 9158 11956 9210
rect 11900 9146 11956 9158
rect 11732 9096 11788 9108
rect 11620 9034 11676 9046
rect 11620 8988 11622 9034
rect 11674 8988 11676 9034
rect 12068 8988 12124 9718
rect 12180 9548 12236 9884
rect 12292 9884 12348 10544
rect 12292 9818 12348 9828
rect 12180 9482 12236 9492
rect 12292 9660 12348 9670
rect 12404 9660 12460 11284
rect 12572 11228 12628 11238
rect 12572 11134 12628 11172
rect 13300 11228 13356 11238
rect 12898 11004 13162 11014
rect 12954 10948 13002 11004
rect 13058 10948 13106 11004
rect 12898 10938 13162 10948
rect 13300 11004 13356 11172
rect 13300 10938 13356 10948
rect 13412 10892 13468 11444
rect 13748 11450 13804 11462
rect 13748 11398 13750 11450
rect 13802 11398 13804 11450
rect 13412 10826 13468 10836
rect 13580 11116 13636 11126
rect 12852 10780 12908 10790
rect 12852 10722 12908 10724
rect 12852 10670 12854 10722
rect 12906 10670 12908 10722
rect 12852 10658 12908 10670
rect 13580 10610 13636 11060
rect 13748 10722 13804 11398
rect 13748 10670 13750 10722
rect 13802 10670 13804 10722
rect 14140 11170 14196 11182
rect 14140 11118 14142 11170
rect 14194 11118 14196 11170
rect 14140 10780 14196 11118
rect 14308 11004 14364 11508
rect 14644 11452 14700 12910
rect 14980 12961 15036 12973
rect 14980 12909 14982 12961
rect 15034 12909 15036 12961
rect 14980 12348 15036 12909
rect 15316 12908 15372 13412
rect 15316 12842 15372 12852
rect 15540 13132 15596 13142
rect 15540 12908 15596 13076
rect 15540 12842 15596 12852
rect 15540 12684 15596 12694
rect 14980 12292 15260 12348
rect 15092 12166 15148 12178
rect 15092 12114 15094 12166
rect 15146 12114 15148 12166
rect 15092 11676 15148 12114
rect 15092 11610 15148 11620
rect 15036 11452 15092 11462
rect 14644 11450 15092 11452
rect 14644 11398 15038 11450
rect 15090 11398 15092 11450
rect 14644 11396 15092 11398
rect 15036 11386 15092 11396
rect 14476 11228 14532 11238
rect 14476 11134 14532 11172
rect 14924 11226 14980 11238
rect 14924 11174 14926 11226
rect 14978 11174 14980 11226
rect 14924 11004 14980 11174
rect 14308 10948 14980 11004
rect 14140 10714 14196 10724
rect 14308 10780 14364 10790
rect 14308 10722 14364 10724
rect 13748 10658 13804 10670
rect 14308 10670 14310 10722
rect 14362 10670 14364 10722
rect 14308 10658 14364 10670
rect 12572 10556 12628 10566
rect 12572 10462 12628 10500
rect 13356 10556 13412 10566
rect 13580 10558 13582 10610
rect 13634 10558 13636 10610
rect 14420 10610 14476 10948
rect 15204 10892 15260 12292
rect 14980 10836 15260 10892
rect 15316 12166 15372 12178
rect 15316 12114 15318 12166
rect 15370 12114 15372 12166
rect 15316 11340 15372 12114
rect 15428 11928 15484 11940
rect 15428 11876 15430 11928
rect 15482 11876 15484 11928
rect 15428 11450 15484 11876
rect 15540 11564 15596 12628
rect 15652 12572 15708 13412
rect 15764 12796 15820 13694
rect 15988 12962 16044 13748
rect 16100 13468 16156 13972
rect 16100 13402 16156 13412
rect 16212 13244 16268 14644
rect 16324 14530 16380 14980
rect 16324 14478 16326 14530
rect 16378 14478 16380 14530
rect 16324 14466 16380 14478
rect 16436 14364 16492 15082
rect 16604 15036 16660 16046
rect 16772 16044 16828 16054
rect 16772 15950 16828 15988
rect 16772 15820 16828 15830
rect 16772 15482 16828 15764
rect 16772 15430 16774 15482
rect 16826 15430 16828 15482
rect 16772 15418 16828 15430
rect 16996 15596 17052 15606
rect 16996 15258 17052 15540
rect 17220 15484 17276 16548
rect 17780 16380 17836 16390
rect 18004 16380 18060 16752
rect 18564 16716 18620 16886
rect 19908 16828 19964 18116
rect 20020 17666 20076 18228
rect 20580 17834 20636 18342
rect 24948 18394 25060 18406
rect 24948 18342 25006 18394
rect 25058 18342 25060 18394
rect 24948 18340 25060 18342
rect 23772 18302 23828 18340
rect 25004 18330 25060 18340
rect 26628 18396 26684 18406
rect 21476 18284 21532 18294
rect 21980 18284 22036 18294
rect 21476 18282 21756 18284
rect 21476 18230 21478 18282
rect 21530 18230 21756 18282
rect 21476 18228 21756 18230
rect 21476 18218 21532 18228
rect 20580 17782 20582 17834
rect 20634 17782 20636 17834
rect 20580 17770 20636 17782
rect 21364 17836 21420 17846
rect 21364 17685 21420 17780
rect 20020 17614 20022 17666
rect 20074 17614 20076 17666
rect 20020 17602 20076 17614
rect 20916 17654 20972 17666
rect 20916 17612 20918 17654
rect 20970 17612 20972 17654
rect 21364 17633 21366 17685
rect 21418 17633 21420 17685
rect 21364 17621 21420 17633
rect 20916 17546 20972 17556
rect 21420 17500 21476 17510
rect 21252 17498 21476 17500
rect 21252 17446 21422 17498
rect 21474 17446 21476 17498
rect 21252 17444 21476 17446
rect 20838 17276 21102 17286
rect 20894 17220 20942 17276
rect 20998 17220 21046 17276
rect 20838 17210 21102 17220
rect 19684 16772 19964 16828
rect 20020 16882 20076 16894
rect 21252 16884 21308 17444
rect 21420 17434 21476 17444
rect 20020 16830 20022 16882
rect 20074 16830 20076 16882
rect 20020 16828 20076 16830
rect 18564 16650 18620 16660
rect 19292 16714 19348 16726
rect 19292 16662 19294 16714
rect 19346 16662 19348 16714
rect 19292 16604 19348 16662
rect 19292 16538 19348 16548
rect 19460 16492 19516 16502
rect 17612 16156 17668 16166
rect 17388 16098 17444 16110
rect 17388 16046 17390 16098
rect 17442 16046 17444 16098
rect 17612 16062 17668 16100
rect 17388 15820 17444 16046
rect 17388 15754 17444 15764
rect 17556 15930 17612 15942
rect 17556 15878 17558 15930
rect 17610 15878 17612 15930
rect 17556 15820 17612 15878
rect 17556 15754 17612 15764
rect 17780 15708 17836 16324
rect 17892 16324 18060 16380
rect 18620 16380 18676 16390
rect 17892 16156 17948 16324
rect 17892 16090 17948 16100
rect 18004 16154 18060 16166
rect 18004 16102 18006 16154
rect 18058 16102 18060 16154
rect 18004 16044 18060 16102
rect 18340 16156 18396 16166
rect 18340 16098 18396 16100
rect 18340 16046 18342 16098
rect 18394 16046 18396 16098
rect 18340 16034 18396 16046
rect 18620 16098 18676 16324
rect 19292 16380 19348 16390
rect 18732 16268 18844 16278
rect 18732 16266 18788 16268
rect 18732 16214 18734 16266
rect 18786 16214 18788 16266
rect 18732 16212 18788 16214
rect 18732 16202 18844 16212
rect 19292 16266 19348 16324
rect 19292 16214 19294 16266
rect 19346 16214 19348 16266
rect 19292 16202 19348 16214
rect 19068 16156 19124 16166
rect 19068 16154 19180 16156
rect 18620 16046 18622 16098
rect 18674 16046 18676 16098
rect 18004 15978 18060 15988
rect 17780 15652 18004 15708
rect 17332 15484 17388 15494
rect 17220 15482 17388 15484
rect 17220 15430 17334 15482
rect 17386 15430 17388 15482
rect 17220 15428 17388 15430
rect 17332 15418 17388 15428
rect 16604 14970 16660 14980
rect 16716 15202 16772 15214
rect 16716 15150 16718 15202
rect 16770 15150 16772 15202
rect 16996 15206 16998 15258
rect 17050 15206 17052 15258
rect 17948 15314 18004 15652
rect 18620 15596 18676 16046
rect 18844 16098 18900 16110
rect 18844 16046 18846 16098
rect 18898 16046 18900 16098
rect 19068 16102 19070 16154
rect 19122 16102 19180 16154
rect 19068 16090 19180 16102
rect 18620 15530 18676 15540
rect 18732 15820 18788 15830
rect 18732 15538 18788 15764
rect 18732 15486 18734 15538
rect 18786 15486 18788 15538
rect 18732 15474 18788 15486
rect 17948 15262 17950 15314
rect 18002 15262 18004 15314
rect 18116 15372 18172 15410
rect 18116 15306 18172 15316
rect 17948 15250 18004 15262
rect 18564 15300 18620 15312
rect 18564 15260 18566 15300
rect 18618 15260 18620 15300
rect 16996 15194 17052 15206
rect 18116 15236 18172 15248
rect 16324 14308 16492 14364
rect 16548 14698 16604 14710
rect 16716 14700 16772 15150
rect 17220 15148 17276 15158
rect 17612 15148 17668 15186
rect 16868 14924 17132 14934
rect 16924 14868 16972 14924
rect 17028 14868 17076 14924
rect 16868 14858 17132 14868
rect 16548 14646 16550 14698
rect 16602 14646 16604 14698
rect 16324 13580 16380 14308
rect 16548 14028 16604 14646
rect 16548 13962 16604 13972
rect 16660 14644 16772 14700
rect 16324 13514 16380 13524
rect 16436 13746 16492 13758
rect 16436 13694 16438 13746
rect 16490 13694 16492 13746
rect 16436 13468 16492 13694
rect 16436 13402 16492 13412
rect 16660 13244 16716 14644
rect 17220 13692 17276 15092
rect 17388 15090 17444 15102
rect 17388 15038 17390 15090
rect 17442 15038 17444 15090
rect 17612 15082 17668 15092
rect 18116 15184 18118 15236
rect 18170 15184 18172 15236
rect 18564 15194 18620 15204
rect 17388 14700 17444 15038
rect 17388 14634 17444 14644
rect 17556 14812 17612 14822
rect 17388 14476 17444 14486
rect 17388 13916 17444 14420
rect 17388 13850 17444 13860
rect 17332 13692 17388 13702
rect 17220 13690 17388 13692
rect 17220 13638 17334 13690
rect 17386 13638 17388 13690
rect 17220 13636 17388 13638
rect 17108 13580 17164 13590
rect 17108 13486 17164 13524
rect 16868 13356 17132 13366
rect 16924 13300 16972 13356
rect 17028 13300 17076 13356
rect 16868 13290 17132 13300
rect 16212 13188 16604 13244
rect 16660 13188 16828 13244
rect 16548 13132 16604 13188
rect 16548 13076 16660 13132
rect 16604 13074 16660 13076
rect 15988 12910 15990 12962
rect 16042 12910 16044 12962
rect 16156 13020 16212 13030
rect 16604 13022 16606 13074
rect 16658 13022 16660 13074
rect 16156 13018 16268 13020
rect 16156 12966 16158 13018
rect 16210 12966 16268 13018
rect 16604 13010 16660 13022
rect 16156 12954 16268 12966
rect 15988 12898 16044 12910
rect 16100 12796 16156 12806
rect 15764 12794 16156 12796
rect 15764 12742 16102 12794
rect 16154 12742 16156 12794
rect 15764 12740 16156 12742
rect 16100 12730 16156 12740
rect 16212 12684 16268 12954
rect 16380 12962 16436 12974
rect 16380 12910 16382 12962
rect 16434 12910 16436 12962
rect 16380 12908 16436 12910
rect 16380 12842 16436 12852
rect 16772 12796 16828 13188
rect 16212 12618 16268 12628
rect 16660 12740 16828 12796
rect 16996 12908 17052 12918
rect 15652 12516 16156 12572
rect 15652 12166 15708 12178
rect 15652 12124 15654 12166
rect 15706 12124 15708 12166
rect 15652 12058 15708 12068
rect 15876 12166 15932 12178
rect 15876 12114 15878 12166
rect 15930 12114 15932 12166
rect 15876 11564 15932 12114
rect 15540 11508 15820 11564
rect 15428 11398 15430 11450
rect 15482 11398 15484 11450
rect 15428 11386 15484 11398
rect 15652 11396 15708 11406
rect 15540 11394 15708 11396
rect 13356 10554 13468 10556
rect 13356 10502 13358 10554
rect 13410 10502 13468 10554
rect 13580 10546 13636 10558
rect 13804 10556 13860 10566
rect 13356 10490 13468 10502
rect 12796 10444 12852 10454
rect 12796 10350 12852 10388
rect 12852 10220 12908 10230
rect 12852 9996 12908 10164
rect 12852 9902 12908 9940
rect 12516 9884 12572 9894
rect 12516 9790 12572 9828
rect 13412 9884 13468 10490
rect 13804 10462 13860 10500
rect 14420 10558 14422 10610
rect 14474 10558 14476 10610
rect 13692 10332 13748 10342
rect 13524 9994 13580 10006
rect 13524 9942 13526 9994
rect 13578 9942 13580 9994
rect 13524 9884 13580 9942
rect 13524 9828 13636 9884
rect 13412 9818 13468 9828
rect 12348 9604 12460 9660
rect 12292 9100 12348 9604
rect 13468 9602 13524 9614
rect 12180 8988 12236 8998
rect 12068 8986 12236 8988
rect 12068 8934 12182 8986
rect 12234 8934 12236 8986
rect 12068 8932 12236 8934
rect 11620 8922 11676 8932
rect 12180 8922 12236 8932
rect 10276 8474 10332 8484
rect 10836 8874 10892 8886
rect 10836 8822 10838 8874
rect 10890 8822 10892 8874
rect 8708 8246 8764 8258
rect 8708 8204 8710 8246
rect 8762 8204 8764 8246
rect 8708 8138 8764 8148
rect 9380 8218 9382 8270
rect 9434 8218 9436 8270
rect 8932 7644 8988 7654
rect 8932 7550 8988 7588
rect 8596 7434 8598 7486
rect 8650 7434 8652 7486
rect 8596 7422 8652 7434
rect 8036 7366 8038 7418
rect 8090 7366 8092 7418
rect 8036 7354 8092 7366
rect 7028 6860 7084 6870
rect 6916 6804 7028 6860
rect 7252 6831 7254 6883
rect 7306 6831 7308 6883
rect 7252 6819 7308 6831
rect 7420 7306 7476 7318
rect 7420 7254 7422 7306
rect 7474 7254 7476 7306
rect 7420 6860 7476 7254
rect 7644 7308 7700 7318
rect 7644 7214 7700 7252
rect 7868 7308 7924 7318
rect 8204 7308 8260 7318
rect 7868 7306 7980 7308
rect 7868 7254 7870 7306
rect 7922 7254 7980 7306
rect 7868 7242 7980 7254
rect 6916 6758 6972 6804
rect 7028 6794 7084 6804
rect 7420 6794 7476 6804
rect 7924 6860 7980 7242
rect 8204 7214 8260 7252
rect 9156 7308 9212 7318
rect 9156 7214 9212 7252
rect 8928 7084 9192 7094
rect 8984 7028 9032 7084
rect 9088 7028 9136 7084
rect 8928 7018 9192 7028
rect 7924 6794 7980 6804
rect 6692 6694 6694 6746
rect 6746 6694 6748 6746
rect 6692 6682 6748 6694
rect 6860 6746 6972 6758
rect 6860 6694 6862 6746
rect 6914 6694 6972 6746
rect 8148 6748 8204 6758
rect 6860 6692 6972 6694
rect 6860 6682 6916 6692
rect 7700 6690 7756 6702
rect 7700 6638 7702 6690
rect 7754 6638 7756 6690
rect 7700 6636 7756 6638
rect 6748 6524 6860 6534
rect 6748 6522 6804 6524
rect 6748 6470 6750 6522
rect 6802 6470 6804 6522
rect 6748 6468 6804 6470
rect 6748 6458 6860 6468
rect 7700 6300 7756 6580
rect 8148 6634 8204 6692
rect 8820 6678 8876 6690
rect 8148 6582 8150 6634
rect 8202 6582 8204 6634
rect 7700 6234 7756 6244
rect 8036 6524 8092 6534
rect 6412 6074 6524 6086
rect 6412 6022 6414 6074
rect 6466 6022 6524 6074
rect 6412 6020 6524 6022
rect 6412 6010 6468 6020
rect 7420 5964 7476 5974
rect 7196 5906 7252 5918
rect 7196 5896 7198 5906
rect 6188 5798 6190 5850
rect 6242 5798 6244 5850
rect 4844 5738 4900 5750
rect 4844 5686 4846 5738
rect 4898 5686 4900 5738
rect 4844 5684 4900 5686
rect 4508 5628 4900 5684
rect 5404 5738 5460 5750
rect 5404 5686 5406 5738
rect 5458 5686 5460 5738
rect 4508 5180 4564 5628
rect 4676 5516 4732 5526
rect 4676 5180 4732 5460
rect 5404 5404 5460 5686
rect 5404 5338 5460 5348
rect 5516 5738 5572 5750
rect 5516 5686 5518 5738
rect 5570 5686 5572 5738
rect 4508 5086 4564 5124
rect 4620 5068 4732 5124
rect 4788 5292 4844 5302
rect 5292 5292 5348 5302
rect 4452 4732 4508 4742
rect 4620 4732 4676 5068
rect 4788 4966 4844 5236
rect 5012 5290 5348 5292
rect 5012 5238 5294 5290
rect 5346 5238 5348 5290
rect 5012 5236 5348 5238
rect 5012 5124 5068 5236
rect 5292 5226 5348 5236
rect 4900 5068 5068 5124
rect 5516 5180 5572 5686
rect 5908 5516 5964 5526
rect 5908 5302 5964 5460
rect 5852 5290 5964 5302
rect 5852 5238 5854 5290
rect 5906 5238 5964 5290
rect 5852 5236 5964 5238
rect 6188 5292 6244 5798
rect 7028 5854 7198 5896
rect 7250 5854 7252 5906
rect 7420 5870 7476 5908
rect 7588 5892 7644 5904
rect 7028 5840 7252 5854
rect 7588 5840 7590 5892
rect 7642 5840 7644 5892
rect 5852 5226 5908 5236
rect 6188 5226 6244 5236
rect 6916 5292 6972 5302
rect 6916 5198 6972 5236
rect 5516 5114 5572 5124
rect 7028 5190 7084 5840
rect 7140 5740 7196 5750
rect 7140 5646 7196 5684
rect 7028 5178 7140 5190
rect 7028 5126 7086 5178
rect 7138 5126 7140 5178
rect 7028 5114 7140 5126
rect 7308 5180 7364 5190
rect 4900 5002 4956 5012
rect 5348 5004 5404 5016
rect 4732 4954 4844 4966
rect 4732 4902 4734 4954
rect 4786 4902 4844 4954
rect 4732 4900 4844 4902
rect 5068 4956 5124 4966
rect 4732 4890 4788 4900
rect 5068 4862 5124 4900
rect 5348 4952 5350 5004
rect 5402 4952 5404 5004
rect 4788 4732 4844 4742
rect 4958 4732 5222 4742
rect 4620 4676 4732 4732
rect 4452 4294 4508 4676
rect 4452 4282 4564 4294
rect 4452 4230 4510 4282
rect 4562 4230 4564 4282
rect 4452 4228 4564 4230
rect 4508 4218 4564 4228
rect 4676 4282 4732 4676
rect 4844 4676 4900 4732
rect 4788 4666 4900 4676
rect 5014 4676 5062 4732
rect 5118 4676 5166 4732
rect 4958 4666 5222 4676
rect 4676 4230 4678 4282
rect 4730 4230 4732 4282
rect 4228 4170 4396 4172
rect 4228 4118 4230 4170
rect 4282 4118 4396 4170
rect 4228 4116 4396 4118
rect 4228 4106 4284 4116
rect 4116 3770 4172 3780
rect 4340 3836 4396 3846
rect 4340 3610 4396 3780
rect 4116 3554 4172 3566
rect 4116 3502 4118 3554
rect 4170 3502 4172 3554
rect 4340 3558 4342 3610
rect 4394 3558 4396 3610
rect 4340 3546 4396 3558
rect 4116 3500 4172 3502
rect 4116 3434 4172 3444
rect 4676 3387 4732 4230
rect 4844 4338 4900 4666
rect 5348 4620 5404 4952
rect 5908 5004 5964 5016
rect 5908 4956 5910 5004
rect 5962 4956 5964 5004
rect 5908 4890 5964 4900
rect 6076 4954 6132 4966
rect 6076 4902 6078 4954
rect 6130 4902 6132 4954
rect 6076 4844 6132 4902
rect 6076 4778 6132 4788
rect 6524 4954 6580 4966
rect 6524 4902 6526 4954
rect 6578 4902 6580 4954
rect 5348 4554 5404 4564
rect 6524 4620 6580 4902
rect 6748 4956 6804 4966
rect 7028 4956 7084 5114
rect 7308 5086 7364 5124
rect 6748 4862 6804 4900
rect 6860 4900 7084 4956
rect 6580 4564 6636 4620
rect 6524 4554 6636 4564
rect 5740 4508 5796 4518
rect 6244 4508 6300 4518
rect 5740 4506 5852 4508
rect 5740 4454 5742 4506
rect 5794 4454 5852 4506
rect 5740 4442 5852 4454
rect 4844 4286 4846 4338
rect 4898 4286 4900 4338
rect 4844 3948 4900 4286
rect 5404 4284 5460 4294
rect 5236 4282 5460 4284
rect 5236 4230 5406 4282
rect 5458 4230 5460 4282
rect 5236 4228 5460 4230
rect 4844 3892 4956 3948
rect 4788 3724 4844 3734
rect 4788 3630 4844 3668
rect 4900 3612 4956 3892
rect 4900 3546 4956 3556
rect 5236 3387 5292 4228
rect 5404 4218 5460 4228
rect 5628 4172 5684 4182
rect 5572 4170 5684 4172
rect 5572 4118 5630 4170
rect 5682 4118 5684 4170
rect 5572 4106 5684 4118
rect 5572 3836 5628 4106
rect 5796 3948 5852 4442
rect 6244 4404 6246 4452
rect 6298 4404 6300 4452
rect 6244 4392 6300 4404
rect 6412 4282 6468 4294
rect 6412 4230 6414 4282
rect 6466 4230 6468 4282
rect 6188 4172 6244 4182
rect 6188 4170 6300 4172
rect 6188 4118 6190 4170
rect 6242 4118 6300 4170
rect 6188 4106 6300 4118
rect 6244 4060 6300 4106
rect 6244 3994 6300 4004
rect 5796 3882 5852 3892
rect 4004 2314 4060 2324
rect 4228 3331 4732 3387
rect 4788 3331 5292 3387
rect 5460 3780 5628 3836
rect 6412 3836 6468 4230
rect 4004 2156 4060 2166
rect 3892 2154 4060 2156
rect 3892 2102 4006 2154
rect 4058 2102 4060 2154
rect 3892 2100 4060 2102
rect 4004 2090 4060 2100
rect 3332 1990 3334 2042
rect 3386 1990 3388 2042
rect 3332 1978 3388 1990
rect 2436 1800 2492 1876
rect 1540 1150 1542 1202
rect 1594 1150 1596 1202
rect 1540 1138 1596 1150
rect 2548 1596 2604 1606
rect 2548 1034 2604 1540
rect 4228 1372 4284 3331
rect 4340 2828 4396 2838
rect 4340 2770 4396 2772
rect 4340 2718 4342 2770
rect 4394 2718 4396 2770
rect 4788 2726 4844 3331
rect 5348 3276 5404 3286
rect 4958 3164 5222 3174
rect 5014 3108 5062 3164
rect 5118 3108 5166 3164
rect 4958 3098 5222 3108
rect 5348 2828 5404 3220
rect 5460 2940 5516 3780
rect 6412 3770 6468 3780
rect 5796 3610 5852 3622
rect 5572 3554 5628 3566
rect 5572 3502 5574 3554
rect 5626 3502 5628 3554
rect 5572 3052 5628 3502
rect 5796 3558 5798 3610
rect 5850 3558 5852 3610
rect 5796 3276 5852 3558
rect 6076 3612 6132 3622
rect 6076 3518 6132 3556
rect 6300 3500 6356 3538
rect 6300 3434 6356 3444
rect 6580 3387 6636 4554
rect 6860 4562 6916 4900
rect 6860 4510 6862 4562
rect 6914 4510 6916 4562
rect 6860 4508 6916 4510
rect 6860 4432 6916 4452
rect 7252 4620 7308 4630
rect 7588 4620 7644 5840
rect 8036 5850 8092 6468
rect 8148 6412 8204 6582
rect 8596 6636 8652 6646
rect 8484 6524 8540 6534
rect 8484 6430 8540 6468
rect 8148 6346 8204 6356
rect 8036 5798 8038 5850
rect 8090 5798 8092 5850
rect 7868 5740 7924 5750
rect 7812 5738 7924 5740
rect 7812 5686 7870 5738
rect 7922 5686 7924 5738
rect 7812 5674 7924 5686
rect 7700 5178 7756 5190
rect 7700 5126 7702 5178
rect 7754 5126 7756 5178
rect 7700 4844 7756 5126
rect 7812 5180 7868 5674
rect 7812 5114 7868 5124
rect 8036 5068 8092 5798
rect 8372 5964 8428 5974
rect 8204 5740 8260 5750
rect 8036 5002 8092 5012
rect 8148 5738 8260 5740
rect 8148 5686 8206 5738
rect 8258 5686 8260 5738
rect 8148 5674 8260 5686
rect 7700 4778 7756 4788
rect 7924 4844 7980 4854
rect 7308 4564 7644 4620
rect 7084 4396 7140 4406
rect 7084 4302 7140 4340
rect 7252 4358 7308 4564
rect 7252 4306 7254 4358
rect 7306 4306 7308 4358
rect 7252 4294 7308 4306
rect 7364 4396 7420 4406
rect 6804 4172 6860 4182
rect 6804 4078 6860 4116
rect 7252 3948 7308 3958
rect 6916 3836 6972 3846
rect 6692 3724 6748 3734
rect 6692 3572 6748 3668
rect 6692 3520 6694 3572
rect 6746 3520 6748 3572
rect 6692 3508 6748 3520
rect 6580 3331 6748 3387
rect 5796 3210 5852 3220
rect 6356 3276 6412 3286
rect 5572 2996 5964 3052
rect 5460 2884 5628 2940
rect 5348 2762 5404 2772
rect 4340 2706 4396 2718
rect 4676 2714 4732 2726
rect 4676 2662 4678 2714
rect 4730 2662 4732 2714
rect 4508 2604 4620 2614
rect 4508 2602 4564 2604
rect 4508 2550 4510 2602
rect 4562 2550 4564 2602
rect 4508 2548 4564 2550
rect 4508 2538 4620 2548
rect 4452 2044 4508 2054
rect 4676 2044 4732 2662
rect 4788 2716 4900 2726
rect 4844 2714 4900 2716
rect 4844 2662 4846 2714
rect 4898 2662 4900 2714
rect 4844 2660 4900 2662
rect 4788 2650 4900 2660
rect 4788 2584 4844 2650
rect 5572 2604 5628 2884
rect 5460 2548 5628 2604
rect 5796 2828 5852 2838
rect 4788 2156 4844 2166
rect 4788 2062 4844 2100
rect 5460 2156 5516 2548
rect 5796 2546 5852 2772
rect 5796 2494 5798 2546
rect 5850 2494 5852 2546
rect 5796 2482 5852 2494
rect 5908 2770 5964 2996
rect 5908 2718 5910 2770
rect 5962 2718 5964 2770
rect 5460 2090 5516 2100
rect 5572 2380 5628 2390
rect 4452 2042 4732 2044
rect 4452 1990 4454 2042
rect 4506 1990 4732 2042
rect 4452 1988 4732 1990
rect 5572 2042 5628 2324
rect 5572 1990 5574 2042
rect 5626 1990 5628 2042
rect 4452 1820 4508 1988
rect 4452 1754 4508 1764
rect 4958 1596 5222 1606
rect 5014 1540 5062 1596
rect 5118 1540 5166 1596
rect 4958 1530 5222 1540
rect 4340 1372 4396 1382
rect 4228 1370 4396 1372
rect 4228 1318 4342 1370
rect 4394 1318 4396 1370
rect 4228 1316 4396 1318
rect 4340 1306 4396 1316
rect 4676 1184 4732 1196
rect 4676 1148 4678 1184
rect 4730 1148 4732 1184
rect 5572 1158 5628 1990
rect 4676 1082 4732 1092
rect 5516 1146 5628 1158
rect 5796 1932 5852 1942
rect 5796 1214 5852 1876
rect 5796 1162 5798 1214
rect 5850 1162 5852 1214
rect 5796 1150 5852 1162
rect 5516 1094 5518 1146
rect 5570 1094 5628 1146
rect 5516 1092 5628 1094
rect 5516 1082 5572 1092
rect 5908 1036 5964 2718
rect 6356 2826 6412 3220
rect 6356 2774 6358 2826
rect 6410 2774 6412 2826
rect 6356 2268 6412 2774
rect 6356 2202 6412 2212
rect 6356 2098 6412 2110
rect 6356 2046 6358 2098
rect 6410 2046 6412 2098
rect 6132 1986 6188 1998
rect 6132 1934 6134 1986
rect 6186 1934 6188 1986
rect 6132 1932 6188 1934
rect 6132 1866 6188 1876
rect 6356 1382 6412 2046
rect 6692 1874 6748 3331
rect 6916 2828 6972 3780
rect 7028 3500 7084 3510
rect 7028 3406 7084 3444
rect 7140 3164 7196 3174
rect 7140 2828 7196 3108
rect 7252 3052 7308 3892
rect 7364 3566 7420 4340
rect 7588 4396 7700 4406
rect 7644 4394 7700 4396
rect 7644 4342 7646 4394
rect 7698 4342 7700 4394
rect 7644 4340 7700 4342
rect 7588 4330 7700 4340
rect 7924 4394 7980 4788
rect 8148 4844 8204 5674
rect 8148 4778 8204 4788
rect 8260 5516 8316 5526
rect 8260 5122 8316 5460
rect 8372 5292 8428 5908
rect 8596 5918 8652 6580
rect 8596 5866 8598 5918
rect 8650 5866 8652 5918
rect 8820 6626 8822 6678
rect 8874 6626 8876 6678
rect 8820 6188 8876 6626
rect 9380 6636 9436 8218
rect 9940 8246 9996 8258
rect 9940 8194 9942 8246
rect 9994 8194 9996 8246
rect 9940 7644 9996 8194
rect 9940 7578 9996 7588
rect 9380 6570 9436 6580
rect 9492 7456 9548 7468
rect 9492 7404 9494 7456
rect 9546 7404 9548 7456
rect 9492 7308 9548 7404
rect 10500 7418 10556 7430
rect 10500 7366 10502 7418
rect 10554 7366 10556 7418
rect 9772 7308 9828 7318
rect 9492 7306 9828 7308
rect 9492 7254 9774 7306
rect 9826 7254 9828 7306
rect 9492 7252 9828 7254
rect 8820 5964 8876 6132
rect 8820 5898 8876 5908
rect 9044 6524 9100 6534
rect 9044 5918 9100 6468
rect 8596 5854 8652 5866
rect 9044 5866 9046 5918
rect 9098 5866 9100 5918
rect 9044 5854 9100 5866
rect 9492 5740 9548 7252
rect 9772 7242 9828 7252
rect 10332 7308 10388 7318
rect 10332 7306 10444 7308
rect 10332 7254 10334 7306
rect 10386 7254 10444 7306
rect 10332 7242 10444 7254
rect 10388 7196 10444 7242
rect 10388 7130 10444 7140
rect 9940 6678 9996 6690
rect 9828 6636 9884 6646
rect 9604 6524 9660 6534
rect 9604 6430 9660 6468
rect 8596 5684 9548 5740
rect 8484 5292 8540 5302
rect 8372 5236 8484 5292
rect 8484 5160 8540 5236
rect 8260 5070 8262 5122
rect 8314 5070 8316 5122
rect 7924 4342 7926 4394
rect 7978 4342 7980 4394
rect 7924 4330 7980 4342
rect 8260 4338 8316 5070
rect 8260 4286 8262 4338
rect 8314 4286 8316 4338
rect 8260 4274 8316 4286
rect 7588 4172 7644 4182
rect 7588 3804 7644 4116
rect 7588 3752 7590 3804
rect 7642 3752 7644 3804
rect 7588 3740 7644 3752
rect 8372 3948 8428 3958
rect 8372 3804 8428 3892
rect 8372 3752 8374 3804
rect 8426 3752 8428 3804
rect 8372 3740 8428 3752
rect 7364 3514 7366 3566
rect 7418 3514 7420 3566
rect 7364 3502 7420 3514
rect 7476 3612 7532 3622
rect 7868 3612 7924 3622
rect 7476 3164 7532 3556
rect 7812 3610 8204 3612
rect 7812 3558 7870 3610
rect 7922 3566 8204 3610
rect 7922 3558 8150 3566
rect 7812 3556 8150 3558
rect 7588 3542 7644 3554
rect 7588 3490 7590 3542
rect 7642 3490 7644 3542
rect 7588 3388 7644 3490
rect 7588 3322 7644 3332
rect 7812 3546 7924 3556
rect 7812 3164 7868 3546
rect 8148 3514 8150 3556
rect 8202 3514 8204 3566
rect 8148 3502 8204 3514
rect 8484 3542 8540 3554
rect 8484 3490 8486 3542
rect 8538 3490 8540 3542
rect 7476 3108 7644 3164
rect 7252 2996 7532 3052
rect 7308 2828 7364 2838
rect 7140 2826 7364 2828
rect 7140 2774 7310 2826
rect 7362 2774 7364 2826
rect 7140 2772 7364 2774
rect 6692 1822 6694 1874
rect 6746 1822 6748 1874
rect 6692 1810 6748 1822
rect 6804 2716 6860 2726
rect 6804 2044 6860 2660
rect 6916 2098 6972 2772
rect 7308 2762 7364 2772
rect 7476 2726 7532 2996
rect 6916 2046 6918 2098
rect 6970 2046 6972 2098
rect 6916 2034 6972 2046
rect 7028 2716 7084 2726
rect 6804 1382 6860 1988
rect 7028 1986 7084 2660
rect 7420 2714 7532 2726
rect 7420 2662 7422 2714
rect 7474 2662 7532 2714
rect 7420 2660 7532 2662
rect 7588 2764 7644 3108
rect 7812 3098 7868 3108
rect 8260 3388 8316 3398
rect 8484 3388 8540 3490
rect 8316 3332 8540 3388
rect 7588 2712 7590 2764
rect 7642 2712 7644 2764
rect 7420 2650 7476 2660
rect 7196 2546 7252 2558
rect 7196 2494 7198 2546
rect 7250 2494 7252 2546
rect 7196 2492 7252 2494
rect 7196 2426 7252 2436
rect 7028 1934 7030 1986
rect 7082 1934 7084 1986
rect 7028 1922 7084 1934
rect 7252 2268 7308 2278
rect 6356 1372 6468 1382
rect 6132 1370 6468 1372
rect 6132 1318 6414 1370
rect 6466 1318 6468 1370
rect 6132 1316 6468 1318
rect 6132 1158 6188 1316
rect 6412 1306 6468 1316
rect 6748 1370 6860 1382
rect 6748 1318 6750 1370
rect 6802 1318 6860 1370
rect 6748 1316 6860 1318
rect 6972 1820 7028 1830
rect 6972 1370 7028 1764
rect 6972 1318 6974 1370
rect 7026 1318 7028 1370
rect 6748 1306 6804 1316
rect 6972 1306 7028 1318
rect 7252 1382 7308 2212
rect 7588 1382 7644 2712
rect 7700 2658 7756 2670
rect 7700 2606 7702 2658
rect 7754 2606 7756 2658
rect 7700 2604 7756 2606
rect 7700 2538 7756 2548
rect 8260 2602 8316 3332
rect 8596 3052 8652 5684
rect 8928 5516 9192 5526
rect 8984 5460 9032 5516
rect 9088 5460 9136 5516
rect 8928 5450 9192 5460
rect 8708 5292 8764 5302
rect 8708 3566 8764 5236
rect 9828 5134 9884 6580
rect 9940 6626 9942 6678
rect 9994 6626 9996 6678
rect 9940 6524 9996 6626
rect 10332 6636 10388 6646
rect 10332 6542 10388 6580
rect 9940 6458 9996 6468
rect 10500 6412 10556 7366
rect 10668 7306 10724 7318
rect 10668 7254 10670 7306
rect 10722 7254 10724 7306
rect 10668 7084 10724 7254
rect 10836 7308 10892 8822
rect 12292 8764 12348 9044
rect 12516 9548 12572 9558
rect 12516 8998 12572 9492
rect 13468 9550 13470 9602
rect 13522 9550 13524 9602
rect 13468 9548 13524 9550
rect 13468 9482 13524 9492
rect 12898 9436 13162 9446
rect 12954 9380 13002 9436
rect 13058 9380 13106 9436
rect 12898 9370 13162 9380
rect 13580 9324 13636 9828
rect 13692 9826 13748 10276
rect 13692 9774 13694 9826
rect 13746 9774 13748 9826
rect 14084 9996 14140 10006
rect 14084 9855 14140 9940
rect 14084 9803 14086 9855
rect 14138 9803 14140 9855
rect 14084 9791 14140 9803
rect 13692 9762 13748 9774
rect 13916 9660 13972 9670
rect 13916 9566 13972 9604
rect 14420 9548 14476 10558
rect 14756 10780 14812 10790
rect 14756 10556 14812 10724
rect 14756 10386 14812 10500
rect 14756 10334 14758 10386
rect 14810 10334 14812 10386
rect 14756 10322 14812 10334
rect 14868 10444 14924 10454
rect 14868 10118 14924 10388
rect 14980 10332 15036 10836
rect 15148 10332 15204 10342
rect 14980 10276 15148 10332
rect 14868 10108 14980 10118
rect 14868 10052 14924 10108
rect 14924 10050 14980 10052
rect 14924 9998 14926 10050
rect 14978 9998 14980 10050
rect 14924 9986 14980 9998
rect 15148 9938 15204 10276
rect 14700 9884 14756 9894
rect 14980 9884 15036 9894
rect 14700 9882 14924 9884
rect 14700 9830 14702 9882
rect 14754 9830 14924 9882
rect 14700 9828 14924 9830
rect 14700 9818 14756 9828
rect 14420 9482 14476 9492
rect 14532 9806 14588 9818
rect 14532 9772 14534 9806
rect 14586 9772 14588 9806
rect 13580 9266 13636 9268
rect 12628 9212 12684 9222
rect 12628 9118 12684 9156
rect 13188 9212 13244 9222
rect 13580 9214 13582 9266
rect 13634 9214 13636 9266
rect 13580 9192 13636 9214
rect 12180 8708 12348 8764
rect 12404 8988 12460 8998
rect 12516 8986 12628 8998
rect 12516 8934 12574 8986
rect 12626 8934 12628 8986
rect 12516 8932 12628 8934
rect 12180 8204 12236 8708
rect 12292 8316 12348 8326
rect 12292 8222 12348 8260
rect 12180 8138 12236 8148
rect 11620 7756 11676 7766
rect 11620 7642 11676 7700
rect 11620 7590 11622 7642
rect 11674 7590 11676 7642
rect 11620 7578 11676 7590
rect 12404 7532 12460 8932
rect 12572 8922 12628 8932
rect 12796 8988 12852 8998
rect 12796 8894 12852 8932
rect 12964 8652 13020 8662
rect 12964 8202 13020 8596
rect 13188 8428 13244 9156
rect 13972 9100 14028 9110
rect 13972 9006 14028 9044
rect 14420 9100 14476 9110
rect 14420 9002 14422 9044
rect 14474 9002 14476 9044
rect 13356 8988 13412 8998
rect 14420 8990 14476 9002
rect 13356 8894 13412 8932
rect 13188 8372 13468 8428
rect 12964 8150 12966 8202
rect 13018 8150 13020 8202
rect 12964 8138 13020 8150
rect 13300 8246 13356 8258
rect 13300 8194 13302 8246
rect 13354 8194 13356 8246
rect 12898 7868 13162 7878
rect 12954 7812 13002 7868
rect 13058 7812 13106 7868
rect 12898 7802 13162 7812
rect 12516 7532 12572 7542
rect 12404 7530 12572 7532
rect 12404 7478 12518 7530
rect 12570 7478 12572 7530
rect 12404 7476 12572 7478
rect 10836 7242 10892 7252
rect 11060 7456 11116 7468
rect 11060 7404 11062 7456
rect 11114 7404 11116 7456
rect 10668 7018 10724 7028
rect 10836 6972 10892 6982
rect 10836 6584 10892 6916
rect 10500 6346 10556 6356
rect 10668 6522 10724 6534
rect 10668 6470 10670 6522
rect 10722 6470 10724 6522
rect 10836 6532 10838 6584
rect 10890 6532 10892 6584
rect 10836 6520 10892 6532
rect 10948 6682 11004 6694
rect 10948 6630 10950 6682
rect 11002 6630 11004 6682
rect 10668 6076 10724 6470
rect 10668 6010 10724 6020
rect 10948 5628 11004 6630
rect 10948 5562 11004 5572
rect 9828 5082 9830 5134
rect 9882 5082 9884 5134
rect 9828 5070 9884 5082
rect 10388 5110 10444 5122
rect 10388 5058 10390 5110
rect 10442 5058 10444 5110
rect 10052 4620 10108 4630
rect 9940 4508 9996 4518
rect 9380 4320 9436 4332
rect 9380 4268 9382 4320
rect 9434 4268 9436 4320
rect 9380 4060 9436 4268
rect 9716 4172 9772 4182
rect 9716 4170 9884 4172
rect 9716 4118 9718 4170
rect 9770 4118 9884 4170
rect 9716 4116 9884 4118
rect 9716 4106 9772 4116
rect 9380 3994 9436 4004
rect 8928 3948 9192 3958
rect 8984 3892 9032 3948
rect 9088 3892 9136 3948
rect 8928 3882 9192 3892
rect 9492 3836 9548 3846
rect 8708 3514 8710 3566
rect 8762 3514 8764 3566
rect 9268 3612 9380 3622
rect 9324 3610 9380 3612
rect 9324 3558 9326 3610
rect 9378 3558 9380 3610
rect 9324 3556 9380 3558
rect 9268 3546 9380 3556
rect 9492 3610 9548 3780
rect 9492 3558 9494 3610
rect 9546 3558 9548 3610
rect 8708 3502 8764 3514
rect 8260 2550 8262 2602
rect 8314 2550 8316 2602
rect 7700 2179 7756 2191
rect 7700 2127 7702 2179
rect 7754 2127 7756 2179
rect 7700 1932 7756 2127
rect 7700 1866 7756 1876
rect 7924 2044 7980 2054
rect 7924 1930 7980 1988
rect 7924 1878 7926 1930
rect 7978 1878 7980 1930
rect 7924 1866 7980 1878
rect 8148 1986 8204 1998
rect 8148 1934 8150 1986
rect 8202 1934 8204 1986
rect 8148 1820 8204 1934
rect 8148 1754 8204 1764
rect 7252 1370 7364 1382
rect 7252 1318 7310 1370
rect 7362 1318 7364 1370
rect 7252 1316 7364 1318
rect 7588 1370 7700 1382
rect 7588 1318 7646 1370
rect 7698 1318 7700 1370
rect 7588 1316 7700 1318
rect 7308 1306 7364 1316
rect 7644 1306 7700 1316
rect 7868 1372 7924 1382
rect 8260 1372 8316 2550
rect 7868 1370 8316 1372
rect 7868 1318 7870 1370
rect 7922 1318 8316 1370
rect 7868 1316 8316 1318
rect 8372 2996 8652 3052
rect 9492 3388 9548 3558
rect 9660 3612 9716 3622
rect 9660 3387 9716 3556
rect 7868 1306 7924 1316
rect 6076 1146 6188 1158
rect 6076 1094 6078 1146
rect 6130 1094 6188 1146
rect 6076 1092 6188 1094
rect 8092 1148 8148 1158
rect 6076 1082 6132 1092
rect 8092 1054 8148 1092
rect 2548 982 2550 1034
rect 2602 982 2604 1034
rect 2548 970 2604 982
rect 5796 980 5964 1036
rect 8372 1036 8428 2996
rect 8652 2828 8708 2838
rect 8652 2734 8708 2772
rect 9156 2828 9212 2838
rect 9156 2734 9212 2772
rect 8876 2716 8932 2726
rect 8876 2622 8932 2660
rect 8928 2380 9192 2390
rect 8984 2324 9032 2380
rect 9088 2324 9136 2380
rect 8928 2314 9192 2324
rect 9492 2156 9548 3332
rect 9604 3331 9716 3387
rect 9604 2828 9660 3331
rect 9604 2762 9660 2772
rect 9828 2714 9884 4116
rect 9940 3554 9996 4452
rect 10052 4350 10108 4564
rect 10388 4506 10444 5058
rect 10388 4454 10390 4506
rect 10442 4454 10444 4506
rect 10388 4442 10444 4454
rect 10948 4508 11004 4518
rect 11060 4508 11116 7404
rect 11956 7456 12012 7468
rect 12516 7466 12572 7476
rect 11956 7420 11958 7456
rect 12010 7420 12012 7456
rect 12796 7420 12852 7430
rect 11956 7354 12012 7364
rect 12516 7396 12572 7408
rect 12516 7344 12518 7396
rect 12570 7344 12572 7396
rect 11396 7306 11452 7318
rect 11396 7254 11398 7306
rect 11450 7254 11452 7306
rect 11284 7196 11340 7206
rect 11284 6746 11340 7140
rect 11284 6694 11286 6746
rect 11338 6694 11340 6746
rect 11284 6682 11340 6694
rect 11396 5850 11452 7254
rect 12348 7306 12404 7318
rect 12348 7254 12350 7306
rect 12402 7254 12404 7306
rect 11900 7084 11956 7094
rect 11900 6914 11956 7028
rect 11900 6862 11902 6914
rect 11954 6862 11956 6914
rect 12348 6972 12404 7254
rect 12516 7308 12572 7344
rect 12796 7326 12852 7364
rect 12516 7242 12572 7252
rect 13300 7308 13356 8194
rect 13412 7486 13468 8372
rect 13804 8258 13860 8270
rect 13804 8206 13806 8258
rect 13858 8206 13860 8258
rect 13804 8204 13860 8206
rect 13748 8148 13860 8204
rect 14532 8204 14588 9716
rect 14644 9660 14700 9670
rect 14644 9566 14700 9604
rect 14756 9548 14812 9558
rect 14644 9100 14700 9110
rect 14644 9002 14646 9044
rect 14698 9002 14700 9044
rect 14644 8990 14700 9002
rect 14756 8818 14812 9492
rect 14756 8766 14758 8818
rect 14810 8766 14812 8818
rect 14756 8754 14812 8766
rect 14868 8652 14924 9828
rect 15148 9886 15150 9938
rect 15202 9886 15204 9938
rect 15148 9874 15204 9886
rect 14980 9054 15036 9828
rect 14980 9002 14982 9054
rect 15034 9002 15036 9054
rect 15316 9772 15372 11284
rect 15540 11342 15654 11394
rect 15706 11342 15708 11394
rect 15540 11340 15708 11342
rect 15540 10780 15596 11340
rect 15652 11330 15708 11340
rect 15764 11004 15820 11508
rect 15876 11498 15932 11508
rect 15988 12124 16044 12134
rect 15540 10714 15596 10724
rect 15652 10948 15820 11004
rect 15652 10566 15708 10948
rect 15764 10780 15820 10790
rect 15764 10778 15932 10780
rect 15764 10726 15766 10778
rect 15818 10726 15932 10778
rect 15764 10724 15932 10726
rect 15764 10714 15820 10724
rect 15484 10556 15540 10566
rect 15652 10554 15764 10566
rect 15652 10502 15710 10554
rect 15762 10502 15764 10554
rect 15652 10500 15764 10502
rect 15484 10386 15540 10500
rect 15708 10490 15764 10500
rect 15484 10334 15486 10386
rect 15538 10334 15540 10386
rect 15484 10220 15540 10334
rect 15484 10154 15540 10164
rect 15876 10108 15932 10724
rect 15652 10052 15932 10108
rect 15316 9100 15372 9716
rect 15428 9882 15484 9894
rect 15428 9830 15430 9882
rect 15482 9830 15484 9882
rect 15428 9548 15484 9830
rect 15428 9482 15484 9492
rect 15316 9034 15372 9044
rect 14980 8990 15036 9002
rect 14868 8586 14924 8596
rect 13748 7642 13804 8148
rect 14532 8138 14588 8148
rect 13748 7590 13750 7642
rect 13802 7590 13804 7642
rect 13748 7578 13804 7590
rect 15428 7644 15484 7654
rect 15428 7550 15484 7588
rect 13412 7434 13414 7486
rect 13466 7434 13468 7486
rect 15092 7532 15148 7542
rect 13412 7422 13468 7434
rect 14420 7456 14476 7468
rect 14420 7404 14422 7456
rect 14474 7404 14476 7456
rect 15092 7434 15094 7476
rect 15146 7434 15148 7476
rect 15092 7422 15148 7434
rect 15652 7430 15708 10052
rect 15988 10006 16044 12068
rect 16100 11954 16156 12516
rect 16100 11902 16102 11954
rect 16154 11902 16156 11954
rect 16212 12166 16268 12178
rect 16212 12114 16214 12166
rect 16266 12114 16268 12166
rect 16212 12012 16268 12114
rect 16436 12166 16492 12178
rect 16436 12124 16438 12166
rect 16490 12124 16492 12166
rect 16660 12134 16716 12740
rect 16996 12348 17052 12852
rect 17332 12572 17388 13636
rect 17556 13468 17612 14756
rect 17668 14700 17724 14710
rect 17668 14530 17724 14644
rect 18116 14700 18172 15184
rect 18844 15148 18900 16046
rect 18956 15596 19012 15606
rect 18956 15538 19012 15540
rect 18956 15486 18958 15538
rect 19010 15486 19012 15538
rect 18956 15474 19012 15486
rect 18116 14634 18172 14644
rect 18788 15092 18900 15148
rect 19012 15148 19068 15158
rect 19124 15148 19180 16090
rect 19012 15146 19180 15148
rect 19012 15094 19014 15146
rect 19066 15094 19180 15146
rect 19012 15092 19180 15094
rect 17668 14478 17670 14530
rect 17722 14478 17724 14530
rect 17668 14466 17724 14478
rect 18620 14476 18676 14486
rect 17892 14412 17948 14424
rect 17892 14360 17894 14412
rect 17946 14360 17948 14412
rect 18620 14382 18676 14420
rect 18060 14364 18116 14374
rect 17780 13916 17836 13926
rect 17668 13746 17724 13758
rect 17668 13694 17670 13746
rect 17722 13694 17724 13746
rect 17668 13692 17724 13694
rect 17668 13626 17724 13636
rect 17780 13634 17836 13860
rect 17892 13804 17948 14360
rect 17892 13738 17948 13748
rect 18004 14362 18116 14364
rect 18004 14310 18062 14362
rect 18114 14310 18116 14362
rect 18004 14298 18116 14310
rect 18396 14364 18452 14374
rect 17780 13582 17782 13634
rect 17834 13582 17836 13634
rect 17780 13570 17836 13582
rect 17332 12506 17388 12516
rect 17444 13244 17500 13254
rect 17444 12980 17500 13188
rect 17444 12928 17446 12980
rect 17498 12928 17500 12980
rect 17332 12348 17388 12358
rect 17444 12348 17500 12928
rect 17556 12796 17612 13412
rect 17892 13356 17948 13366
rect 17892 13020 17948 13300
rect 18004 13132 18060 14298
rect 18396 14270 18452 14308
rect 18788 14252 18844 15092
rect 19012 15082 19068 15092
rect 19460 14924 19516 16436
rect 19068 14868 19516 14924
rect 19572 15596 19628 15606
rect 19572 15148 19628 15540
rect 19684 15326 19740 16772
rect 20020 16762 20076 16772
rect 20468 16828 20524 16838
rect 20916 16828 21308 16884
rect 21700 16884 21756 18228
rect 21980 18282 22204 18284
rect 21980 18230 21982 18282
rect 22034 18230 22204 18282
rect 21980 18228 22204 18230
rect 21980 18218 22036 18228
rect 22036 18060 22092 18070
rect 22036 17734 22092 18004
rect 22148 17948 22204 18228
rect 22260 18282 22316 18294
rect 22260 18230 22262 18282
rect 22314 18230 22316 18282
rect 22260 18172 22316 18230
rect 22988 18284 23044 18294
rect 23436 18284 23492 18294
rect 22988 18190 23044 18228
rect 23380 18282 23492 18284
rect 23380 18230 23438 18282
rect 23490 18230 23492 18282
rect 23380 18218 23492 18230
rect 23548 18284 23604 18294
rect 25396 18284 25452 18294
rect 25900 18284 25956 18294
rect 26236 18284 26292 18294
rect 26628 18284 26684 18340
rect 23548 18282 23660 18284
rect 23548 18230 23550 18282
rect 23602 18230 23660 18282
rect 23548 18218 23660 18230
rect 25396 18282 25564 18284
rect 25396 18230 25398 18282
rect 25450 18230 25564 18282
rect 25396 18228 25564 18230
rect 25396 18218 25452 18228
rect 22260 18106 22316 18116
rect 22148 17892 22428 17948
rect 22036 17722 22148 17734
rect 22036 17670 22094 17722
rect 22146 17670 22148 17722
rect 22036 17668 22148 17670
rect 22092 17658 22148 17668
rect 22372 17666 22428 17892
rect 23212 17836 23268 17846
rect 23212 17742 23268 17780
rect 22372 17614 22374 17666
rect 22426 17614 22428 17666
rect 22372 17602 22428 17614
rect 21980 17498 22036 17510
rect 21980 17446 21982 17498
rect 22034 17446 22036 17498
rect 21980 17052 22036 17446
rect 21980 16986 22036 16996
rect 21700 16828 21924 16884
rect 23380 16882 23436 18218
rect 20468 16826 20580 16828
rect 20468 16774 20470 16826
rect 20522 16774 20580 16826
rect 20468 16762 20580 16774
rect 20300 16716 20356 16726
rect 20132 16714 20356 16716
rect 20132 16662 20302 16714
rect 20354 16662 20356 16714
rect 20132 16660 20356 16662
rect 19908 16268 19964 16278
rect 19908 16098 19964 16212
rect 19908 16046 19910 16098
rect 19962 16046 19964 16098
rect 19908 16034 19964 16046
rect 20132 15820 20188 16660
rect 20300 16650 20356 16660
rect 20524 16716 20580 16762
rect 20412 16604 20468 16614
rect 20412 16266 20468 16548
rect 20412 16214 20414 16266
rect 20466 16214 20468 16266
rect 20412 16202 20468 16214
rect 20524 16156 20580 16660
rect 20636 16714 20692 16726
rect 20636 16662 20638 16714
rect 20690 16662 20692 16714
rect 20636 16380 20692 16662
rect 20636 16314 20692 16324
rect 20524 16100 20636 16156
rect 20076 15764 20188 15820
rect 19796 15708 19852 15718
rect 19796 15438 19852 15652
rect 19796 15386 19798 15438
rect 19850 15386 19852 15438
rect 19796 15374 19852 15386
rect 19684 15274 19686 15326
rect 19738 15274 19740 15326
rect 19684 15262 19740 15274
rect 20076 15314 20132 15764
rect 20580 15596 20636 16100
rect 20916 16044 20972 16828
rect 21308 16716 21364 16726
rect 21308 16622 21364 16660
rect 21420 16714 21476 16726
rect 21420 16662 21422 16714
rect 21474 16662 21476 16714
rect 21420 16492 21476 16662
rect 21028 16436 21476 16492
rect 21756 16714 21812 16726
rect 21756 16662 21758 16714
rect 21810 16662 21812 16714
rect 21756 16492 21812 16662
rect 21868 16714 21924 16828
rect 22260 16864 22316 16876
rect 22260 16828 22262 16864
rect 22314 16828 22316 16864
rect 23380 16830 23382 16882
rect 23434 16830 23436 16882
rect 23380 16818 23436 16830
rect 23604 16940 23660 18218
rect 24808 18060 25072 18070
rect 24864 18004 24912 18060
rect 24968 18004 25016 18060
rect 24808 17994 25072 18004
rect 22260 16762 22316 16772
rect 21868 16662 21870 16714
rect 21922 16662 21924 16714
rect 21868 16650 21924 16662
rect 22596 16714 22652 16726
rect 22596 16662 22598 16714
rect 22650 16662 22652 16714
rect 22596 16604 22652 16662
rect 22596 16538 22652 16548
rect 21028 16268 21084 16436
rect 21756 16426 21812 16436
rect 22652 16380 22708 16390
rect 21028 16202 21084 16212
rect 21252 16324 21700 16380
rect 21140 16044 21196 16054
rect 20916 16042 21196 16044
rect 20916 15990 21142 16042
rect 21194 15990 21196 16042
rect 20916 15988 21196 15990
rect 21140 15978 21196 15988
rect 20838 15708 21102 15718
rect 20894 15652 20942 15708
rect 20998 15652 21046 15708
rect 20838 15642 21102 15652
rect 21252 15606 21308 16324
rect 21644 16266 21700 16324
rect 23604 16380 23660 16884
rect 24052 17610 24108 17622
rect 24052 17558 24054 17610
rect 24106 17558 24108 17610
rect 23884 16716 23940 16726
rect 23884 16622 23940 16660
rect 24052 16604 24108 17558
rect 24724 17612 24780 17622
rect 24444 17500 24500 17510
rect 24388 17498 24500 17500
rect 24388 17446 24446 17498
rect 24498 17446 24500 17498
rect 24724 17508 24726 17556
rect 24778 17508 24780 17556
rect 25284 17612 25340 17622
rect 25284 17518 25340 17556
rect 24724 17496 24780 17508
rect 24388 17434 24500 17446
rect 24388 16716 24444 17434
rect 24388 16650 24444 16660
rect 24500 16996 24780 17052
rect 23604 16324 23996 16380
rect 21644 16214 21646 16266
rect 21698 16214 21700 16266
rect 21644 16202 21700 16214
rect 21812 16268 21868 16278
rect 20580 15382 20636 15540
rect 20076 15262 20078 15314
rect 20130 15262 20132 15314
rect 20524 15370 20636 15382
rect 20524 15318 20526 15370
rect 20578 15318 20636 15370
rect 20524 15316 20636 15318
rect 21196 15596 21308 15606
rect 21252 15540 21308 15596
rect 21532 16156 21588 16166
rect 21532 15596 21588 16100
rect 21700 16044 21756 16054
rect 21812 16044 21868 16212
rect 22260 16268 22316 16278
rect 22260 16176 22316 16212
rect 22652 16266 22708 16324
rect 22652 16214 22654 16266
rect 22706 16214 22708 16266
rect 22652 16202 22708 16214
rect 22820 16268 22876 16278
rect 22260 16124 22262 16176
rect 22314 16124 22316 16176
rect 22260 16112 22316 16124
rect 22820 16176 22876 16212
rect 22820 16124 22822 16176
rect 22874 16124 22876 16176
rect 22820 16112 22876 16124
rect 23380 16268 23436 16278
rect 23380 16176 23436 16212
rect 23380 16124 23382 16176
rect 23434 16124 23436 16176
rect 23380 16112 23436 16124
rect 23772 16156 23828 16166
rect 21700 16042 21868 16044
rect 21700 15990 21702 16042
rect 21754 15990 21868 16042
rect 21700 15988 21868 15990
rect 22092 16098 22148 16110
rect 22092 16046 22094 16098
rect 22146 16046 22148 16098
rect 23212 16098 23268 16110
rect 21700 15978 21756 15988
rect 22092 15596 22148 16046
rect 22260 16044 22316 16054
rect 22820 16044 22876 16054
rect 23212 16046 23214 16098
rect 23266 16046 23268 16098
rect 23772 16062 23828 16100
rect 23212 16044 23268 16046
rect 22260 16042 22540 16044
rect 22260 15990 22262 16042
rect 22314 15990 22540 16042
rect 22260 15988 22540 15990
rect 22260 15978 22316 15988
rect 21196 15370 21252 15540
rect 21532 15530 21588 15540
rect 22036 15540 22148 15596
rect 22372 15596 22428 15606
rect 21700 15484 21756 15494
rect 21196 15318 21198 15370
rect 21250 15318 21252 15370
rect 20524 15306 20580 15316
rect 21196 15306 21252 15318
rect 21364 15372 21420 15382
rect 20076 15250 20132 15262
rect 19068 14754 19124 14868
rect 19068 14702 19070 14754
rect 19122 14702 19124 14754
rect 19068 14690 19124 14702
rect 19292 14700 19348 14710
rect 19292 14606 19348 14644
rect 19572 14700 19628 15092
rect 19852 15146 19908 15158
rect 19852 15094 19854 15146
rect 19906 15094 19908 15146
rect 19852 14924 19908 15094
rect 20300 15148 20356 15158
rect 20300 15146 20412 15148
rect 20300 15094 20302 15146
rect 20354 15094 20412 15146
rect 20300 15082 20412 15094
rect 19852 14858 19908 14868
rect 20244 14812 20300 14822
rect 19572 14644 19964 14700
rect 18676 14196 18844 14252
rect 18900 14518 18956 14530
rect 18900 14466 18902 14518
rect 18954 14466 18956 14518
rect 18900 14252 18956 14466
rect 18340 13804 18396 13814
rect 18340 13802 18508 13804
rect 18340 13750 18342 13802
rect 18394 13750 18508 13802
rect 18340 13748 18508 13750
rect 18340 13738 18396 13748
rect 18340 13668 18396 13680
rect 18340 13616 18342 13668
rect 18394 13616 18396 13668
rect 18172 13578 18228 13590
rect 18172 13526 18174 13578
rect 18226 13526 18228 13578
rect 18172 13356 18228 13526
rect 18172 13290 18228 13300
rect 18340 13244 18396 13616
rect 18452 13356 18508 13748
rect 18452 13290 18508 13300
rect 18340 13178 18396 13188
rect 18564 13244 18620 13254
rect 18116 13132 18172 13142
rect 18004 13076 18116 13132
rect 17892 12964 18060 13020
rect 18004 12950 18060 12964
rect 17780 12908 17836 12918
rect 17780 12814 17836 12852
rect 18004 12898 18006 12950
rect 18058 12898 18060 12950
rect 17556 12730 17612 12740
rect 18004 12684 18060 12898
rect 18116 12684 18172 13076
rect 18564 13030 18620 13188
rect 18284 13020 18340 13030
rect 18228 13018 18340 13020
rect 18228 12966 18286 13018
rect 18338 12966 18340 13018
rect 18228 12954 18340 12966
rect 18508 13018 18620 13030
rect 18508 12966 18510 13018
rect 18562 12966 18620 13018
rect 18508 12964 18620 12966
rect 18228 12908 18284 12954
rect 18228 12842 18284 12852
rect 18340 12850 18396 12862
rect 18340 12798 18342 12850
rect 18394 12798 18396 12850
rect 18340 12796 18396 12798
rect 18340 12730 18396 12740
rect 18116 12628 18284 12684
rect 18004 12618 18060 12628
rect 16996 12292 17108 12348
rect 17052 12178 17108 12292
rect 17332 12346 17500 12348
rect 17332 12294 17334 12346
rect 17386 12294 17500 12346
rect 17332 12292 17500 12294
rect 17332 12282 17388 12292
rect 18228 12290 18284 12628
rect 16660 12122 16772 12134
rect 16660 12070 16718 12122
rect 16770 12070 16772 12122
rect 16660 12068 16772 12070
rect 16436 12058 16492 12068
rect 16716 12058 16772 12068
rect 16884 12122 16940 12134
rect 16884 12070 16886 12122
rect 16938 12070 16940 12122
rect 16212 11946 16268 11956
rect 16884 12012 16940 12070
rect 17052 12126 17054 12178
rect 17106 12126 17108 12178
rect 17052 12012 17108 12126
rect 17892 12236 17948 12246
rect 18228 12238 18230 12290
rect 18282 12238 18284 12290
rect 18228 12226 18284 12238
rect 17948 12180 18004 12190
rect 17892 12178 18004 12180
rect 17892 12126 17950 12178
rect 18002 12126 18004 12178
rect 17892 12124 18004 12126
rect 17780 12068 18004 12124
rect 18508 12124 18564 12964
rect 18676 12348 18732 14196
rect 18900 14186 18956 14196
rect 19012 14408 19068 14420
rect 19012 14356 19014 14408
rect 19066 14356 19068 14408
rect 19012 14140 19068 14356
rect 19012 14074 19068 14084
rect 19124 14364 19180 14374
rect 18788 13804 18844 13814
rect 18788 13706 18790 13748
rect 18842 13706 18844 13748
rect 18788 13694 18844 13706
rect 18956 13692 19012 13702
rect 18900 13690 19012 13692
rect 18900 13638 18958 13690
rect 19010 13638 19012 13690
rect 18900 13626 19012 13638
rect 18900 13244 18956 13626
rect 19124 13522 19180 14308
rect 19572 13802 19628 14644
rect 19908 14598 19964 14644
rect 19908 14586 20020 14598
rect 19740 14530 19796 14542
rect 19908 14534 19966 14586
rect 20018 14534 20020 14586
rect 19908 14532 20020 14534
rect 19740 14478 19742 14530
rect 19794 14478 19796 14530
rect 19964 14522 20020 14532
rect 19740 14028 19796 14478
rect 20244 14326 20300 14756
rect 20356 14700 20412 15082
rect 20692 15036 20748 15046
rect 20468 14700 20524 14710
rect 20356 14698 20524 14700
rect 20356 14646 20470 14698
rect 20522 14646 20524 14698
rect 20356 14644 20524 14646
rect 20468 14634 20524 14644
rect 20580 14700 20636 14710
rect 20244 14274 20246 14326
rect 20298 14274 20300 14326
rect 20244 14252 20300 14274
rect 20244 14186 20300 14196
rect 20468 14518 20524 14530
rect 20468 14476 20470 14518
rect 20522 14476 20524 14518
rect 20468 14252 20524 14420
rect 20468 14186 20524 14196
rect 19572 13750 19574 13802
rect 19626 13750 19628 13802
rect 19572 13738 19628 13750
rect 19684 13972 19796 14028
rect 19292 13692 19348 13702
rect 19124 13470 19126 13522
rect 19178 13470 19180 13522
rect 19124 13458 19180 13470
rect 19236 13690 19516 13692
rect 19236 13638 19294 13690
rect 19346 13638 19516 13690
rect 19236 13636 19516 13638
rect 19236 13626 19348 13636
rect 19236 13356 19292 13626
rect 19460 13580 19516 13636
rect 19684 13580 19740 13972
rect 20580 13916 20636 14644
rect 20356 13860 20636 13916
rect 20356 13702 20412 13860
rect 20692 13858 20748 14980
rect 21084 15036 21140 15046
rect 21084 14586 21140 14980
rect 21084 14534 21086 14586
rect 21138 14534 21140 14586
rect 21084 14522 21140 14534
rect 21252 15036 21308 15046
rect 21252 14598 21308 14980
rect 21364 14924 21420 15316
rect 21700 15300 21756 15428
rect 21700 15248 21702 15300
rect 21754 15248 21756 15300
rect 21532 15148 21588 15186
rect 21532 15082 21588 15092
rect 21700 15147 21756 15248
rect 22036 15260 22092 15540
rect 22260 15426 22316 15438
rect 22260 15374 22262 15426
rect 22314 15374 22316 15426
rect 22260 15372 22316 15374
rect 22372 15372 22428 15540
rect 22484 15484 22540 15988
rect 22820 16042 22988 16044
rect 22820 15990 22822 16042
rect 22874 15990 22988 16042
rect 22820 15988 22988 15990
rect 22820 15978 22876 15988
rect 22484 15428 22708 15484
rect 22260 15316 22428 15372
rect 22036 15194 22092 15204
rect 21700 15091 21868 15147
rect 21364 14868 21532 14924
rect 21252 14586 21364 14598
rect 21252 14534 21310 14586
rect 21362 14534 21364 14586
rect 21252 14522 21364 14534
rect 21252 14364 21308 14522
rect 21252 14298 21308 14308
rect 20838 14140 21102 14150
rect 21476 14140 21532 14868
rect 21644 14700 21700 14710
rect 21644 14606 21700 14644
rect 21812 14588 21868 15091
rect 21980 15090 22036 15102
rect 21980 15038 21982 15090
rect 22034 15038 22036 15090
rect 21980 14812 22036 15038
rect 21980 14746 22036 14756
rect 22204 15090 22260 15102
rect 22204 15038 22206 15090
rect 22258 15038 22260 15090
rect 22204 14754 22260 15038
rect 22372 14812 22428 15316
rect 22204 14702 22206 14754
rect 22258 14702 22260 14754
rect 22204 14700 22260 14702
rect 22204 14624 22260 14644
rect 22316 14756 22428 14812
rect 22540 15258 22596 15270
rect 22540 15206 22542 15258
rect 22594 15206 22596 15258
rect 21812 14532 22092 14588
rect 22036 14510 22092 14532
rect 21700 14476 21756 14486
rect 21756 14420 21868 14476
rect 21700 14410 21756 14420
rect 20894 14084 20942 14140
rect 20998 14084 21046 14140
rect 20838 14074 21102 14084
rect 21308 14084 21532 14140
rect 21700 14140 21756 14150
rect 20692 13806 20694 13858
rect 20746 13806 20748 13858
rect 20692 13794 20748 13806
rect 21308 13746 21364 14084
rect 20300 13690 20412 13702
rect 20300 13638 20302 13690
rect 20354 13638 20412 13690
rect 20300 13636 20412 13638
rect 20524 13692 20580 13702
rect 21308 13694 21310 13746
rect 21362 13694 21364 13746
rect 21476 13804 21532 13814
rect 21700 13804 21756 14084
rect 21476 13802 21756 13804
rect 21476 13750 21478 13802
rect 21530 13750 21756 13802
rect 21476 13748 21756 13750
rect 21476 13738 21532 13748
rect 21308 13682 21364 13694
rect 21812 13692 21868 14420
rect 22036 14458 22038 14510
rect 22090 14458 22092 14510
rect 22036 14252 22092 14458
rect 22316 14364 22372 14756
rect 22428 14588 22484 14598
rect 22428 14494 22484 14532
rect 22540 14374 22596 15206
rect 22652 15148 22708 15428
rect 22764 15372 22820 15382
rect 22764 15278 22820 15316
rect 22652 15092 22876 15148
rect 22652 14532 22708 14542
rect 22652 14530 22764 14532
rect 22652 14478 22654 14530
rect 22706 14478 22764 14530
rect 22652 14466 22764 14478
rect 22316 14308 22428 14364
rect 22540 14362 22652 14374
rect 22540 14310 22598 14362
rect 22650 14310 22652 14362
rect 22540 14308 22652 14310
rect 22036 14186 22092 14196
rect 22092 13802 22148 13814
rect 22092 13750 22094 13802
rect 22146 13750 22148 13802
rect 20300 13626 20356 13636
rect 20524 13598 20580 13636
rect 21588 13636 21868 13692
rect 21924 13734 21980 13746
rect 21924 13682 21926 13734
rect 21978 13682 21980 13734
rect 22092 13702 22148 13750
rect 19460 13524 19740 13580
rect 19964 13580 20020 13590
rect 20748 13580 20804 13590
rect 21420 13580 21476 13590
rect 19964 13578 20076 13580
rect 19964 13526 19966 13578
rect 20018 13526 20076 13578
rect 19964 13514 20076 13526
rect 18900 13178 18956 13188
rect 19012 13300 19292 13356
rect 19012 12908 19068 13300
rect 19348 13244 19404 13254
rect 19180 13188 19348 13244
rect 19180 13020 19236 13188
rect 19348 13178 19404 13188
rect 19180 12926 19236 12964
rect 19740 13020 19796 13030
rect 20020 13020 20076 13514
rect 20748 13486 20804 13524
rect 21364 13578 21476 13580
rect 21364 13526 21422 13578
rect 21474 13526 21476 13578
rect 21364 13514 21476 13526
rect 21364 13468 21420 13514
rect 21364 13402 21420 13412
rect 20468 13244 20524 13254
rect 20468 13130 20524 13188
rect 21364 13244 21420 13254
rect 20468 13078 20470 13130
rect 20522 13078 20524 13130
rect 20468 13066 20524 13078
rect 21028 13132 21084 13142
rect 21028 13038 21084 13076
rect 20132 13020 20188 13030
rect 20020 13018 20188 13020
rect 20020 12966 20134 13018
rect 20186 12966 20188 13018
rect 20020 12964 20188 12966
rect 19740 12926 19796 12964
rect 18676 12282 18732 12292
rect 18900 12852 19068 12908
rect 17668 12012 17724 12022
rect 17052 11956 17276 12012
rect 16884 11946 16940 11956
rect 16100 11890 16156 11902
rect 16868 11788 17132 11798
rect 16924 11732 16972 11788
rect 17028 11732 17076 11788
rect 16868 11722 17132 11732
rect 16436 11562 16492 11574
rect 16436 11510 16438 11562
rect 16490 11510 16492 11562
rect 16436 11340 16492 11510
rect 16436 11274 16492 11284
rect 16940 11340 16996 11350
rect 16940 10834 16996 11284
rect 17220 11228 17276 11956
rect 17668 11918 17724 11956
rect 17388 11676 17444 11686
rect 17388 11562 17444 11620
rect 17388 11510 17390 11562
rect 17442 11510 17444 11562
rect 17388 11498 17444 11510
rect 17500 11564 17556 11574
rect 17500 11470 17556 11508
rect 17780 11391 17836 12068
rect 18284 12012 18340 12032
rect 18508 12030 18564 12068
rect 18284 11954 18340 11956
rect 18284 11902 18286 11954
rect 18338 11902 18340 11954
rect 18004 11676 18060 11686
rect 18004 11562 18060 11620
rect 18004 11510 18006 11562
rect 18058 11510 18060 11562
rect 18004 11498 18060 11510
rect 17780 11339 17782 11391
rect 17834 11339 17836 11391
rect 17220 11172 17500 11228
rect 16940 10782 16942 10834
rect 16994 10782 16996 10834
rect 16940 10770 16996 10782
rect 16100 10556 16156 10566
rect 17332 10556 17388 10566
rect 16100 10554 16268 10556
rect 16100 10502 16102 10554
rect 16154 10502 16268 10554
rect 16100 10500 16268 10502
rect 16100 10490 16156 10500
rect 15988 9994 16100 10006
rect 15988 9942 16046 9994
rect 16098 9942 16100 9994
rect 15988 9930 16100 9942
rect 15988 9884 16044 9930
rect 15820 9828 15876 9838
rect 15764 9826 15876 9828
rect 15764 9774 15822 9826
rect 15874 9774 15876 9826
rect 15988 9818 16044 9828
rect 15764 9772 15876 9774
rect 15820 9762 15876 9772
rect 15764 9706 15820 9716
rect 15876 9660 15932 9670
rect 16212 9660 16268 10500
rect 17444 10556 17500 11172
rect 17444 10500 17556 10556
rect 17332 10462 17388 10500
rect 17500 10498 17556 10500
rect 16604 10444 16660 10454
rect 16548 10442 16660 10444
rect 16548 10390 16606 10442
rect 16658 10390 16660 10442
rect 17500 10446 17502 10498
rect 17554 10446 17556 10498
rect 17500 10434 17556 10446
rect 17780 10444 17836 11339
rect 18060 11396 18116 11406
rect 18284 11396 18340 11902
rect 18900 11564 18956 12852
rect 19404 12796 19460 12806
rect 19348 12794 19460 12796
rect 19348 12742 19406 12794
rect 19458 12742 19460 12794
rect 19348 12730 19460 12742
rect 19124 12348 19180 12358
rect 19348 12348 19404 12730
rect 19180 12292 19404 12348
rect 19908 12460 19964 12470
rect 19012 12236 19068 12246
rect 19012 12178 19068 12180
rect 19012 12126 19014 12178
rect 19066 12126 19068 12178
rect 19012 12114 19068 12126
rect 19012 12012 19068 12022
rect 19124 12012 19180 12292
rect 19460 12236 19516 12246
rect 19012 12010 19180 12012
rect 19012 11958 19014 12010
rect 19066 11958 19180 12010
rect 19012 11956 19180 11958
rect 19348 12178 19404 12190
rect 19348 12126 19350 12178
rect 19402 12126 19404 12178
rect 19348 12012 19404 12126
rect 19012 11946 19068 11956
rect 19348 11946 19404 11956
rect 18900 11498 18956 11508
rect 19236 11900 19292 11910
rect 18060 11394 18340 11396
rect 18060 11342 18062 11394
rect 18114 11342 18340 11394
rect 19236 11394 19292 11844
rect 18060 11340 18340 11342
rect 18060 11330 18172 11340
rect 16548 10378 16660 10390
rect 17780 10378 17836 10388
rect 16548 9844 16604 10378
rect 16868 10220 17132 10230
rect 16924 10164 16972 10220
rect 17028 10164 17076 10220
rect 16868 10154 17132 10164
rect 16548 9792 16550 9844
rect 16602 9792 16604 9844
rect 18116 9884 18172 11330
rect 18788 11338 18844 11350
rect 18788 11286 18790 11338
rect 18842 11286 18844 11338
rect 19236 11342 19238 11394
rect 19290 11342 19292 11394
rect 19236 11330 19292 11342
rect 18788 11228 18844 11286
rect 18284 11170 18340 11182
rect 18284 11118 18286 11170
rect 18338 11118 18340 11170
rect 18788 11162 18844 11172
rect 18284 11116 18340 11118
rect 18284 11050 18340 11060
rect 19012 11116 19068 11126
rect 19012 10592 19068 11060
rect 18228 10556 18284 10566
rect 18228 10462 18284 10500
rect 19012 10540 19014 10592
rect 19066 10540 19068 10592
rect 18452 10444 18508 10454
rect 18452 9884 18508 10388
rect 18620 10444 18676 10454
rect 18620 10442 18732 10444
rect 18620 10390 18622 10442
rect 18674 10390 18732 10442
rect 18620 10378 18732 10390
rect 18676 9996 18732 10378
rect 19012 10220 19068 10540
rect 19348 10444 19404 10454
rect 19460 10444 19516 12180
rect 19908 11900 19964 12404
rect 20132 12236 20188 12964
rect 21364 12962 21420 13188
rect 21588 13142 21644 13636
rect 21924 13580 21980 13682
rect 22036 13692 22148 13702
rect 22092 13636 22148 13692
rect 22260 13692 22316 13702
rect 22036 13626 22092 13636
rect 22260 13580 22316 13636
rect 21756 13356 21812 13366
rect 21588 13130 21700 13142
rect 21588 13078 21646 13130
rect 21698 13078 21700 13130
rect 21588 13076 21700 13078
rect 21644 13066 21700 13076
rect 20692 12908 20748 12918
rect 21364 12910 21366 12962
rect 21418 12910 21420 12962
rect 21756 13018 21812 13300
rect 21756 12966 21758 13018
rect 21810 12966 21812 13018
rect 21756 12954 21812 12966
rect 21364 12898 21420 12910
rect 20692 12814 20748 12852
rect 20838 12572 21102 12582
rect 20894 12516 20942 12572
rect 20998 12516 21046 12572
rect 20838 12506 21102 12516
rect 20132 12170 20188 12180
rect 20356 12348 20412 12358
rect 21924 12348 21980 13524
rect 22148 13524 22316 13580
rect 22148 13020 22204 13524
rect 22372 13468 22428 14308
rect 22596 14298 22652 14308
rect 22708 14140 22764 14466
rect 22820 14252 22876 15092
rect 22932 14700 22988 15988
rect 23156 15988 23268 16044
rect 23380 16042 23436 16054
rect 23380 15990 23382 16042
rect 23434 15990 23436 16042
rect 23156 15708 23212 15988
rect 23380 15932 23436 15990
rect 23380 15866 23436 15876
rect 23156 15642 23212 15652
rect 23268 15820 23324 15830
rect 23044 15484 23100 15494
rect 23100 15436 23212 15484
rect 23100 15428 23158 15436
rect 23044 15418 23100 15428
rect 23156 15384 23158 15428
rect 23210 15384 23212 15436
rect 23156 15372 23212 15384
rect 23044 15294 23100 15306
rect 23044 15242 23046 15294
rect 23098 15242 23100 15294
rect 23268 15270 23324 15764
rect 23940 15482 23996 16324
rect 24052 16278 24108 16548
rect 24052 16266 24164 16278
rect 24052 16214 24110 16266
rect 24162 16214 24164 16266
rect 24052 16212 24164 16214
rect 24108 16202 24164 16212
rect 24500 16266 24556 16996
rect 24724 16940 24780 16996
rect 24948 16940 25004 16950
rect 24724 16938 25004 16940
rect 24724 16886 24950 16938
rect 25002 16886 25004 16938
rect 24724 16884 25004 16886
rect 24948 16874 25004 16884
rect 24612 16826 24668 16838
rect 24612 16774 24614 16826
rect 24666 16774 24668 16826
rect 24612 16604 24668 16774
rect 24612 16538 24668 16548
rect 24808 16492 25072 16502
rect 24864 16436 24912 16492
rect 24968 16436 25016 16492
rect 24808 16426 25072 16436
rect 25508 16278 25564 18228
rect 25900 18190 25956 18228
rect 26180 18282 26292 18284
rect 26180 18230 26238 18282
rect 26290 18230 26292 18282
rect 26180 18218 26292 18230
rect 26516 18282 26684 18284
rect 26516 18230 26630 18282
rect 26682 18230 26684 18282
rect 26516 18228 26684 18230
rect 26180 17846 26236 18218
rect 26124 17836 26236 17846
rect 26180 17780 26236 17836
rect 26124 17742 26180 17780
rect 26292 16940 26348 16950
rect 26292 16882 26348 16884
rect 26292 16830 26294 16882
rect 26346 16830 26348 16882
rect 26292 16818 26348 16830
rect 25788 16716 25844 16726
rect 25788 16622 25844 16660
rect 25732 16492 25788 16502
rect 24500 16214 24502 16266
rect 24554 16214 24556 16266
rect 24500 16202 24556 16214
rect 25172 16268 25284 16278
rect 25228 16266 25284 16268
rect 25228 16214 25230 16266
rect 25282 16214 25284 16266
rect 25228 16212 25284 16214
rect 25508 16266 25620 16278
rect 25508 16214 25566 16266
rect 25618 16214 25620 16266
rect 25508 16212 25620 16214
rect 25172 16202 25284 16212
rect 25564 16202 25620 16212
rect 23940 15430 23942 15482
rect 23994 15430 23996 15482
rect 23940 15418 23996 15430
rect 24612 16156 24668 16166
rect 24612 15484 24668 16100
rect 25396 16154 25452 16166
rect 25396 16102 25398 16154
rect 25450 16102 25452 16154
rect 24780 16042 24836 16054
rect 24780 15990 24782 16042
rect 24834 15990 24836 16042
rect 24780 15932 24836 15990
rect 24780 15866 24836 15876
rect 25396 15932 25452 16102
rect 24612 15382 24668 15428
rect 25396 15484 25452 15876
rect 25396 15418 25452 15428
rect 25732 15436 25788 16436
rect 26124 16268 26180 16278
rect 26124 16174 26180 16212
rect 25956 16156 26012 16166
rect 25956 16062 26012 16100
rect 26404 16156 26460 16166
rect 26068 16044 26124 16054
rect 26068 15942 26124 15988
rect 26012 15930 26124 15942
rect 26012 15878 26014 15930
rect 26066 15878 26124 15930
rect 26012 15876 26124 15878
rect 26012 15866 26068 15876
rect 26404 15596 26460 16100
rect 26516 16154 26572 18228
rect 26628 18218 26684 18228
rect 26740 17666 26796 18900
rect 27300 18620 27356 19200
rect 28778 18844 29042 18854
rect 28834 18788 28882 18844
rect 28938 18788 28986 18844
rect 28778 18778 29042 18788
rect 27188 18564 27356 18620
rect 29092 18732 29148 18742
rect 27188 18508 27244 18564
rect 27188 18410 27190 18452
rect 27242 18410 27244 18452
rect 28140 18508 28196 18518
rect 27188 18398 27244 18410
rect 27636 18432 27692 18444
rect 27636 18396 27638 18432
rect 27690 18396 27692 18432
rect 28140 18414 28196 18452
rect 27636 18330 27692 18340
rect 28756 18396 28812 18406
rect 26852 18284 26908 18294
rect 27188 18284 27244 18294
rect 26852 18282 27020 18284
rect 26852 18230 26854 18282
rect 26906 18230 27020 18282
rect 26852 18228 27020 18230
rect 26852 18218 26908 18228
rect 26740 17614 26742 17666
rect 26794 17614 26796 17666
rect 26740 17602 26796 17614
rect 26852 16882 26908 16894
rect 26852 16830 26854 16882
rect 26906 16830 26908 16882
rect 26852 16492 26908 16830
rect 26852 16426 26908 16436
rect 26964 16268 27020 18228
rect 27188 17666 27244 18228
rect 27972 18282 28028 18294
rect 27972 18230 27974 18282
rect 28026 18230 28028 18282
rect 27972 17836 28028 18230
rect 27972 17780 28476 17836
rect 27188 17614 27190 17666
rect 27242 17614 27244 17666
rect 27188 17602 27244 17614
rect 28028 17612 28084 17622
rect 28028 17518 28084 17556
rect 28420 16938 28476 17780
rect 28756 17722 28812 18340
rect 28756 17670 28758 17722
rect 28810 17670 28812 17722
rect 28756 17658 28812 17670
rect 29092 17666 29148 18676
rect 29988 18508 30044 19200
rect 29988 18442 30044 18452
rect 30548 18508 30604 18518
rect 30548 18406 30604 18452
rect 30716 18508 30772 18518
rect 30716 18414 30772 18452
rect 30492 18394 30604 18406
rect 30492 18342 30494 18394
rect 30546 18342 30604 18394
rect 30492 18340 30604 18342
rect 32396 18396 32452 18406
rect 32564 18396 32620 19200
rect 32396 18394 32620 18396
rect 32396 18342 32398 18394
rect 32450 18342 32620 18394
rect 32396 18340 32620 18342
rect 30492 18330 30548 18340
rect 32396 18330 32452 18340
rect 29372 18284 29428 18294
rect 29092 17614 29094 17666
rect 29146 17614 29148 17666
rect 29092 17602 29148 17614
rect 29316 18282 29428 18284
rect 29316 18230 29374 18282
rect 29426 18230 29428 18282
rect 29316 18218 29428 18230
rect 29484 18284 29540 18294
rect 28778 17276 29042 17286
rect 28834 17220 28882 17276
rect 28938 17220 28986 17276
rect 28778 17210 29042 17220
rect 28420 16886 28422 16938
rect 28474 16886 28476 16938
rect 28420 16874 28476 16886
rect 26964 16202 27020 16212
rect 27244 16716 27300 16726
rect 27244 16266 27300 16660
rect 27692 16716 27748 16726
rect 27692 16622 27748 16660
rect 27244 16214 27246 16266
rect 27298 16214 27300 16266
rect 27244 16202 27300 16214
rect 28476 16492 28532 16502
rect 28476 16266 28532 16436
rect 28476 16214 28478 16266
rect 28530 16214 28532 16266
rect 28476 16202 28532 16214
rect 26516 16102 26518 16154
rect 26570 16102 26572 16154
rect 26516 16090 26572 16102
rect 26740 16156 26796 16166
rect 28364 16156 28420 16166
rect 26740 15596 26796 16100
rect 28084 16154 28420 16156
rect 28084 16102 28366 16154
rect 28418 16102 28420 16154
rect 28084 16100 28420 16102
rect 28084 16098 28140 16100
rect 28084 16046 28086 16098
rect 28138 16046 28140 16098
rect 28364 16090 28420 16100
rect 28868 16098 28924 16110
rect 28084 16034 28140 16046
rect 28868 16046 28870 16098
rect 28922 16046 28924 16098
rect 26404 15540 26572 15596
rect 25732 15384 25734 15436
rect 25786 15384 25788 15436
rect 24556 15370 24668 15382
rect 24556 15318 24558 15370
rect 24610 15318 24668 15370
rect 24556 15316 24668 15318
rect 25116 15372 25172 15382
rect 25564 15372 25620 15382
rect 25732 15372 25788 15384
rect 25508 15370 25620 15372
rect 24556 15306 24612 15316
rect 23044 15036 23100 15242
rect 23212 15258 23324 15270
rect 23212 15206 23214 15258
rect 23266 15206 23324 15258
rect 23212 15204 23324 15206
rect 24892 15260 24948 15270
rect 23212 15194 23268 15204
rect 23436 15148 23492 15186
rect 24892 15166 24948 15204
rect 23436 15082 23492 15092
rect 24332 15148 24444 15158
rect 24332 15146 24388 15148
rect 24332 15094 24334 15146
rect 24386 15094 24388 15146
rect 24332 15092 24388 15094
rect 24332 15082 24444 15092
rect 23044 14970 23100 14980
rect 23324 15036 23380 15046
rect 25116 15036 25172 15316
rect 25340 15314 25396 15326
rect 25340 15262 25342 15314
rect 25394 15262 25396 15314
rect 25340 15147 25396 15262
rect 25284 15091 25396 15147
rect 25508 15318 25566 15370
rect 25618 15318 25620 15370
rect 25508 15306 25620 15318
rect 25116 14980 25228 15036
rect 22932 14634 22988 14644
rect 23044 14812 23100 14822
rect 22932 14530 22988 14542
rect 22932 14478 22934 14530
rect 22986 14478 22988 14530
rect 22932 14476 22988 14478
rect 22932 14410 22988 14420
rect 23044 14424 23100 14756
rect 23044 14372 23046 14424
rect 23098 14372 23100 14424
rect 23044 14360 23100 14372
rect 23324 14362 23380 14980
rect 24808 14924 25072 14934
rect 24864 14868 24912 14924
rect 24968 14868 25016 14924
rect 24808 14858 25072 14868
rect 24612 14812 24668 14822
rect 25172 14812 25228 14980
rect 23884 14700 23940 14710
rect 23324 14310 23326 14362
rect 23378 14310 23380 14362
rect 22820 14196 23044 14252
rect 22708 14084 22876 14140
rect 22484 13916 22540 13926
rect 22484 13580 22540 13860
rect 22652 13916 22708 13926
rect 22652 13822 22708 13860
rect 22484 13514 22540 13524
rect 22148 12954 22204 12964
rect 22260 13412 22428 13468
rect 22820 13468 22876 14084
rect 22988 13858 23044 14196
rect 23212 14028 23268 14038
rect 23324 14028 23380 14310
rect 23268 13972 23380 14028
rect 23492 14698 23940 14700
rect 23492 14646 23886 14698
rect 23938 14646 23940 14698
rect 23492 14644 23940 14646
rect 23212 13970 23268 13972
rect 23212 13918 23214 13970
rect 23266 13918 23268 13970
rect 23212 13906 23268 13918
rect 22988 13806 22990 13858
rect 23042 13806 23044 13858
rect 22988 13794 23044 13806
rect 22260 12974 22316 13412
rect 22820 13402 22876 13412
rect 23268 13356 23324 13366
rect 23492 13356 23548 14644
rect 23884 14634 23940 14644
rect 24052 14588 24108 14598
rect 23660 14532 23716 14542
rect 23604 14530 23716 14532
rect 23604 14478 23662 14530
rect 23714 14478 23716 14530
rect 23604 14466 23716 14478
rect 24052 14484 24054 14532
rect 24106 14484 24108 14532
rect 24052 14472 24108 14484
rect 24388 14530 24444 14542
rect 24388 14478 24390 14530
rect 24442 14478 24444 14530
rect 23604 13804 23660 14466
rect 23940 14408 23996 14420
rect 23716 14364 23772 14374
rect 23940 14364 23942 14408
rect 23994 14364 23996 14408
rect 23772 14308 23884 14364
rect 23716 14298 23772 14308
rect 23604 13738 23660 13748
rect 23716 14028 23772 14038
rect 23604 13580 23660 13590
rect 23716 13580 23772 13972
rect 23828 13916 23884 14308
rect 23940 14298 23996 14308
rect 24052 14252 24108 14262
rect 23828 13860 23940 13916
rect 23884 13746 23940 13860
rect 23884 13694 23886 13746
rect 23938 13694 23940 13746
rect 24052 13802 24108 14196
rect 24052 13750 24054 13802
rect 24106 13750 24108 13802
rect 24052 13738 24108 13750
rect 23884 13682 23940 13694
rect 23604 13578 23772 13580
rect 23604 13526 23606 13578
rect 23658 13526 23772 13578
rect 23604 13524 23772 13526
rect 24052 13668 24108 13680
rect 24052 13616 24054 13668
rect 24106 13616 24108 13668
rect 23604 13514 23660 13524
rect 23492 13300 23604 13356
rect 22596 13186 22652 13198
rect 22260 12922 22262 12974
rect 22314 12922 22316 12974
rect 22260 12910 22316 12922
rect 22372 13132 22428 13142
rect 22372 12358 22428 13076
rect 22596 13134 22598 13186
rect 22650 13134 22652 13186
rect 22484 12950 22540 12962
rect 22484 12908 22486 12950
rect 22538 12908 22540 12950
rect 22484 12842 22540 12852
rect 22204 12348 22260 12358
rect 21924 12346 22260 12348
rect 21924 12294 22206 12346
rect 22258 12294 22260 12346
rect 21924 12292 22260 12294
rect 20020 12124 20076 12134
rect 20020 12030 20076 12068
rect 20356 11900 20412 12292
rect 22204 12282 22260 12292
rect 22316 12346 22428 12358
rect 22316 12294 22318 12346
rect 22370 12294 22428 12346
rect 22316 12292 22428 12294
rect 22316 12282 22372 12292
rect 20748 12236 20804 12246
rect 22596 12236 22652 13134
rect 22820 13020 22876 13030
rect 22820 12922 22822 12964
rect 22874 12922 22876 12964
rect 22820 12910 22876 12922
rect 23268 12962 23324 13300
rect 22988 12908 23044 12918
rect 23268 12910 23270 12962
rect 23322 12910 23324 12962
rect 23268 12898 23324 12910
rect 22988 12814 23044 12852
rect 23548 12738 23604 13300
rect 23828 13244 23884 13254
rect 23828 13130 23884 13188
rect 24052 13132 24108 13616
rect 24388 13580 24444 14478
rect 24612 14252 24668 14756
rect 25116 14756 25228 14812
rect 24836 14700 24892 14710
rect 25116 14700 25172 14756
rect 24836 14364 24892 14644
rect 24556 14196 24668 14252
rect 24780 14308 24892 14364
rect 25060 14644 25172 14700
rect 25284 14700 25340 15091
rect 25508 14812 25564 15306
rect 26012 15260 26068 15270
rect 26012 15166 26068 15204
rect 26516 15258 26572 15540
rect 26516 15206 26518 15258
rect 26570 15206 26572 15258
rect 26684 15540 26796 15596
rect 28308 15932 28364 15942
rect 26684 15314 26740 15540
rect 26684 15262 26686 15314
rect 26738 15262 26740 15314
rect 26684 15250 26740 15262
rect 27412 15372 27468 15382
rect 28308 15316 28364 15876
rect 28868 15932 28924 16046
rect 28868 15866 28924 15876
rect 29316 15820 29372 18218
rect 29484 18190 29540 18228
rect 30100 18284 30156 18294
rect 31332 18284 31388 18294
rect 30100 18190 30156 18228
rect 30884 18282 31388 18284
rect 30884 18230 31334 18282
rect 31386 18230 31388 18282
rect 30884 18228 31388 18230
rect 29932 17612 29988 17622
rect 29932 17518 29988 17556
rect 30772 17610 30828 17622
rect 30772 17558 30774 17610
rect 30826 17558 30828 17610
rect 30772 17500 30828 17558
rect 30772 17434 30828 17444
rect 30884 17164 30940 18228
rect 31332 18218 31388 18228
rect 31724 18284 31836 18294
rect 31724 18282 31780 18284
rect 31724 18230 31726 18282
rect 31778 18230 31780 18282
rect 31724 18228 31780 18230
rect 31724 18218 31836 18228
rect 32004 18282 32060 18294
rect 32004 18230 32006 18282
rect 32058 18230 32060 18282
rect 32004 17836 32060 18230
rect 32004 17770 32060 17780
rect 32116 18284 32172 18294
rect 31332 17668 31388 17678
rect 31220 17666 31388 17668
rect 31220 17614 31334 17666
rect 31386 17614 31388 17666
rect 32116 17622 32172 18228
rect 32564 17846 32620 18340
rect 32508 17834 32620 17846
rect 32508 17782 32510 17834
rect 32562 17782 32620 17834
rect 32508 17780 32620 17782
rect 32508 17770 32564 17780
rect 31220 17612 31388 17614
rect 31332 17602 31388 17612
rect 32060 17610 32172 17622
rect 31220 17546 31276 17556
rect 32060 17558 32062 17610
rect 32114 17558 32172 17610
rect 32060 17556 32172 17558
rect 32060 17546 32116 17556
rect 30772 17108 30940 17164
rect 30996 17498 31052 17510
rect 30996 17446 30998 17498
rect 31050 17446 31052 17498
rect 29540 16882 29596 16894
rect 29540 16830 29542 16882
rect 29594 16830 29596 16882
rect 29540 16828 29596 16830
rect 29540 16762 29596 16772
rect 30044 16714 30100 16726
rect 30044 16662 30046 16714
rect 30098 16662 30100 16714
rect 30044 16156 30100 16662
rect 30772 16156 30828 17108
rect 30884 16940 30940 16950
rect 30996 16940 31052 17446
rect 31332 17500 31388 17510
rect 31332 17011 31388 17444
rect 31332 16959 31334 17011
rect 31386 16959 31388 17011
rect 31332 16947 31388 16959
rect 30884 16938 31164 16940
rect 30884 16886 30886 16938
rect 30938 16886 31164 16938
rect 30884 16884 31164 16886
rect 30884 16874 30940 16884
rect 30044 16100 30268 16156
rect 29708 16044 29764 16054
rect 29708 16042 30044 16044
rect 29708 15990 29710 16042
rect 29762 15990 30044 16042
rect 29708 15988 30044 15990
rect 29708 15978 29764 15988
rect 29316 15754 29372 15764
rect 28778 15708 29042 15718
rect 28834 15652 28882 15708
rect 28938 15652 28986 15708
rect 28778 15642 29042 15652
rect 27412 15314 27580 15316
rect 27412 15262 27414 15314
rect 27466 15262 27580 15314
rect 27412 15260 27580 15262
rect 27412 15250 27468 15260
rect 26516 15194 26572 15206
rect 25620 15148 25676 15158
rect 26348 15148 26404 15158
rect 26292 15146 26404 15148
rect 25620 14924 25676 15092
rect 25788 15090 25844 15102
rect 25788 15038 25790 15090
rect 25842 15038 25844 15090
rect 25788 15036 25844 15038
rect 26292 15094 26350 15146
rect 26402 15094 26404 15146
rect 26292 15082 26404 15094
rect 26740 15148 26796 15158
rect 26292 15036 26348 15082
rect 25788 14980 25900 15036
rect 25620 14868 25788 14924
rect 25508 14746 25564 14756
rect 24556 14028 24612 14196
rect 24556 13970 24612 13972
rect 24556 13918 24558 13970
rect 24610 13918 24612 13970
rect 24556 13896 24612 13918
rect 24780 14140 24836 14308
rect 24780 13970 24836 14084
rect 24780 13918 24782 13970
rect 24834 13918 24836 13970
rect 24780 13906 24836 13918
rect 25060 13916 25116 14644
rect 25284 14634 25340 14644
rect 25340 14532 25396 14542
rect 25564 14532 25620 14542
rect 25060 13749 25116 13860
rect 25060 13697 25062 13749
rect 25114 13697 25116 13749
rect 25060 13685 25116 13697
rect 25172 14530 25396 14532
rect 25172 14478 25342 14530
rect 25394 14478 25396 14530
rect 25172 14476 25396 14478
rect 24500 13580 24556 13590
rect 24388 13578 24556 13580
rect 24388 13526 24502 13578
rect 24554 13526 24556 13578
rect 24388 13524 24556 13526
rect 24500 13514 24556 13524
rect 24808 13356 25072 13366
rect 24864 13300 24912 13356
rect 24968 13300 25016 13356
rect 24808 13290 25072 13300
rect 25172 13244 25228 14476
rect 25340 14466 25396 14476
rect 25508 14530 25620 14532
rect 25508 14478 25566 14530
rect 25618 14478 25620 14530
rect 25508 14466 25620 14478
rect 25508 14364 25564 14466
rect 25396 14308 25564 14364
rect 25620 14364 25676 14374
rect 25732 14364 25788 14868
rect 25844 14588 25900 14980
rect 25844 14522 25900 14532
rect 25956 14980 26348 15036
rect 25956 14586 26012 14980
rect 26124 14812 26180 14822
rect 26124 14700 26180 14756
rect 25956 14534 25958 14586
rect 26010 14534 26012 14586
rect 25956 14522 26012 14534
rect 26068 14698 26180 14700
rect 26068 14646 26126 14698
rect 26178 14646 26180 14698
rect 26068 14634 26180 14646
rect 26572 14700 26684 14710
rect 26572 14698 26628 14700
rect 26572 14646 26574 14698
rect 26626 14646 26628 14698
rect 26572 14644 26628 14646
rect 26572 14634 26684 14644
rect 25620 14362 25788 14364
rect 25620 14310 25622 14362
rect 25674 14310 25788 14362
rect 25620 14308 25788 14310
rect 25396 13804 25452 14308
rect 25620 14298 25676 14308
rect 25396 13738 25452 13748
rect 25508 13804 25564 13814
rect 25508 13802 25676 13804
rect 25508 13750 25510 13802
rect 25562 13750 25676 13802
rect 25508 13748 25676 13750
rect 25508 13738 25564 13748
rect 25508 13668 25564 13680
rect 25508 13616 25510 13668
rect 25562 13616 25564 13668
rect 25172 13178 25228 13188
rect 25340 13578 25396 13590
rect 25340 13526 25342 13578
rect 25394 13526 25396 13578
rect 24164 13132 24220 13142
rect 23828 13078 23830 13130
rect 23882 13078 23884 13130
rect 23828 13066 23884 13078
rect 23940 13076 24164 13132
rect 23044 12684 23100 12694
rect 22596 12180 22764 12236
rect 20748 12142 20804 12180
rect 22708 12134 22764 12180
rect 23044 12190 23100 12628
rect 23548 12686 23550 12738
rect 23602 12686 23604 12738
rect 23548 12470 23604 12686
rect 23772 12738 23828 12750
rect 23772 12686 23774 12738
rect 23826 12686 23828 12738
rect 23772 12684 23828 12686
rect 23548 12460 23660 12470
rect 23548 12404 23604 12460
rect 23604 12346 23660 12404
rect 23604 12294 23606 12346
rect 23658 12294 23660 12346
rect 23604 12282 23660 12294
rect 23772 12348 23828 12628
rect 23772 12282 23828 12292
rect 23044 12138 23046 12190
rect 23098 12138 23100 12190
rect 20636 12124 20692 12134
rect 22708 12122 22820 12134
rect 23044 12126 23100 12138
rect 23380 12166 23436 12178
rect 22708 12070 22766 12122
rect 22818 12070 22820 12122
rect 22708 12068 22820 12070
rect 20636 12030 20692 12068
rect 22764 12058 22820 12068
rect 23380 12114 23382 12166
rect 23434 12114 23436 12166
rect 21532 12012 21588 12022
rect 21924 12012 21980 12022
rect 19908 11844 20076 11900
rect 19684 11587 19740 11599
rect 19684 11564 19686 11587
rect 19738 11564 19740 11587
rect 19684 11495 19740 11508
rect 19796 10668 19852 10678
rect 19796 10574 19852 10612
rect 20020 10610 20076 11844
rect 20356 11834 20412 11844
rect 21252 12010 21588 12012
rect 21252 11958 21534 12010
rect 21586 11958 21588 12010
rect 21252 11956 21588 11958
rect 21140 11382 21196 11394
rect 21140 11330 21142 11382
rect 21194 11330 21196 11382
rect 21140 11228 21196 11330
rect 21140 11162 21196 11172
rect 20838 11004 21102 11014
rect 20894 10948 20942 11004
rect 20998 10948 21046 11004
rect 20838 10938 21102 10948
rect 21252 10780 21308 11956
rect 21532 11946 21588 11956
rect 21812 12010 21980 12012
rect 21812 11958 21926 12010
rect 21978 11958 21980 12010
rect 21812 11956 21980 11958
rect 20804 10724 21308 10780
rect 21364 11564 21420 11574
rect 20804 10678 20860 10724
rect 20020 10558 20022 10610
rect 20074 10558 20076 10610
rect 20748 10666 20860 10678
rect 20748 10614 20750 10666
rect 20802 10614 20860 10666
rect 20748 10612 20860 10614
rect 21364 10622 21420 11508
rect 21812 11452 21868 11956
rect 21924 11946 21980 11956
rect 21756 11396 21868 11452
rect 23156 11928 23212 11940
rect 23156 11876 23158 11928
rect 23210 11876 23212 11928
rect 21756 11394 21812 11396
rect 21756 11342 21758 11394
rect 21810 11342 21812 11394
rect 21756 11330 21812 11342
rect 20748 10602 20804 10612
rect 21364 10570 21366 10622
rect 21418 10570 21420 10622
rect 21364 10558 21420 10570
rect 21476 11228 21532 11238
rect 20020 10546 20076 10558
rect 19348 10442 19516 10444
rect 19348 10390 19350 10442
rect 19402 10390 19516 10442
rect 19348 10388 19516 10390
rect 19348 10332 19404 10388
rect 19348 10266 19404 10276
rect 19012 10154 19068 10164
rect 18676 9940 19516 9996
rect 18452 9828 19404 9884
rect 16548 9780 16604 9792
rect 17444 9814 17500 9826
rect 16884 9772 16940 9782
rect 16884 9678 16940 9716
rect 17444 9762 17446 9814
rect 17498 9762 17500 9814
rect 15876 9658 16268 9660
rect 15876 9606 15878 9658
rect 15930 9606 16268 9658
rect 15876 9604 16268 9606
rect 15876 9594 15932 9604
rect 16268 9042 16324 9054
rect 15876 9030 15932 9042
rect 15876 8978 15878 9030
rect 15930 8978 15932 9030
rect 16268 8990 16270 9042
rect 16322 8990 16324 9042
rect 16268 8988 16324 8990
rect 15876 8428 15932 8978
rect 15876 8362 15932 8372
rect 16100 8932 16324 8988
rect 16100 7642 16156 8932
rect 16868 8652 17132 8662
rect 16924 8596 16972 8652
rect 17028 8596 17076 8652
rect 16868 8586 17132 8596
rect 16660 8428 16716 8438
rect 16100 7590 16102 7642
rect 16154 7590 16156 7642
rect 16100 7578 16156 7590
rect 16212 8314 16268 8326
rect 16212 8262 16214 8314
rect 16266 8262 16268 8314
rect 16212 7644 16268 8262
rect 16212 7578 16268 7588
rect 12348 6906 12404 6916
rect 12628 6914 12684 6926
rect 11900 6850 11956 6862
rect 12628 6862 12630 6914
rect 12682 6862 12684 6914
rect 11676 6748 11732 6758
rect 11676 6746 11788 6748
rect 11676 6694 11678 6746
rect 11730 6694 11788 6746
rect 11676 6682 11788 6694
rect 11732 6636 11788 6682
rect 11620 6524 11676 6534
rect 11620 6430 11676 6468
rect 11396 5798 11398 5850
rect 11450 5798 11452 5850
rect 11396 5786 11452 5798
rect 11340 4508 11396 4518
rect 11060 4506 11396 4508
rect 11060 4454 11342 4506
rect 11394 4454 11396 4506
rect 11060 4452 11396 4454
rect 11732 4508 11788 6580
rect 12292 6678 12348 6690
rect 12292 6626 12294 6678
rect 12346 6626 12348 6678
rect 12068 6412 12124 6422
rect 12068 6074 12124 6356
rect 12068 6022 12070 6074
rect 12122 6022 12124 6074
rect 12068 6010 12124 6022
rect 12180 6300 12236 6310
rect 12180 5516 12236 6244
rect 12180 4518 12236 5460
rect 12292 5180 12348 6626
rect 12516 6678 12572 6690
rect 12516 6636 12518 6678
rect 12570 6636 12572 6678
rect 12516 6570 12572 6580
rect 12628 6412 12684 6862
rect 13076 6748 13132 6758
rect 13300 6748 13356 7252
rect 13916 7308 13972 7318
rect 13916 7214 13972 7252
rect 13132 6692 13356 6748
rect 14420 6748 14476 7404
rect 15652 7418 15764 7430
rect 15652 7366 15710 7418
rect 15762 7366 15764 7418
rect 15652 7364 15764 7366
rect 15708 7354 15764 7364
rect 14756 7306 14812 7318
rect 14756 7254 14758 7306
rect 14810 7254 14812 7306
rect 12852 6678 12908 6690
rect 12852 6626 12854 6678
rect 12906 6626 12908 6678
rect 13076 6650 13078 6692
rect 13130 6650 13132 6692
rect 13076 6638 13132 6650
rect 13636 6678 13692 6690
rect 14420 6682 14476 6692
rect 14644 7084 14700 7094
rect 12852 6524 12908 6626
rect 12516 6356 12684 6412
rect 12740 6468 12908 6524
rect 13636 6626 13638 6678
rect 13690 6626 13692 6678
rect 12516 5918 12572 6356
rect 12516 5866 12518 5918
rect 12570 5866 12572 5918
rect 12516 5854 12572 5866
rect 12740 5740 12796 6468
rect 12898 6300 13162 6310
rect 12954 6244 13002 6300
rect 13058 6244 13106 6300
rect 12898 6234 13162 6244
rect 12852 6076 12908 6086
rect 12852 5982 12908 6020
rect 13636 6076 13692 6626
rect 14308 6076 14364 6086
rect 13636 6010 13692 6020
rect 13972 6074 14364 6076
rect 13972 6022 14310 6074
rect 14362 6022 14364 6074
rect 13972 6020 14364 6022
rect 13524 5888 13580 5900
rect 13524 5836 13526 5888
rect 13578 5836 13580 5888
rect 12740 5674 12796 5684
rect 13300 5740 13356 5750
rect 12740 5180 12796 5190
rect 12292 5114 12348 5124
rect 12628 5178 12796 5180
rect 12628 5126 12742 5178
rect 12794 5126 12796 5178
rect 12628 5124 12796 5126
rect 12012 4508 12068 4518
rect 11732 4506 12068 4508
rect 11732 4454 12014 4506
rect 12066 4454 12068 4506
rect 11732 4452 12068 4454
rect 10052 4298 10054 4350
rect 10106 4298 10108 4350
rect 10052 4286 10108 4298
rect 10948 4352 11004 4452
rect 11340 4442 11396 4452
rect 12012 4442 12068 4452
rect 12124 4506 12236 4518
rect 12124 4454 12126 4506
rect 12178 4454 12236 4506
rect 12124 4452 12236 4454
rect 12516 4956 12572 4966
rect 12516 4456 12572 4900
rect 12124 4442 12180 4452
rect 12516 4404 12518 4456
rect 12570 4404 12572 4456
rect 12516 4392 12572 4404
rect 10948 4346 11340 4352
rect 10948 4294 10950 4346
rect 11002 4338 11340 4346
rect 11002 4296 11286 4338
rect 11002 4294 11004 4296
rect 10668 4282 10724 4294
rect 10948 4282 11004 4294
rect 11284 4286 11286 4296
rect 11338 4286 11340 4338
rect 12404 4338 12460 4350
rect 10668 4230 10670 4282
rect 10722 4230 10724 4282
rect 11284 4274 11340 4286
rect 11676 4282 11732 4294
rect 10332 4172 10388 4182
rect 9940 3502 9942 3554
rect 9994 3502 9996 3554
rect 9940 3490 9996 3502
rect 10052 4060 10108 4070
rect 10052 3448 10108 4004
rect 10332 3610 10388 4116
rect 10668 4172 10724 4230
rect 11676 4230 11678 4282
rect 11730 4230 11732 4282
rect 10668 4106 10724 4116
rect 10780 4172 10836 4182
rect 11676 4172 11732 4230
rect 10780 4170 10892 4172
rect 10780 4118 10782 4170
rect 10834 4118 10892 4170
rect 10780 4106 10892 4118
rect 11676 4106 11732 4116
rect 12404 4286 12406 4338
rect 12458 4286 12460 4338
rect 10836 3724 10892 4106
rect 12404 3948 12460 4286
rect 12404 3882 12460 3892
rect 10836 3658 10892 3668
rect 11284 3836 11340 3846
rect 10332 3558 10334 3610
rect 10386 3558 10388 3610
rect 10332 3546 10388 3558
rect 10052 3396 10054 3448
rect 10106 3396 10108 3448
rect 10052 3384 10108 3396
rect 10164 3500 10220 3510
rect 9828 2662 9830 2714
rect 9882 2662 9884 2714
rect 9828 2650 9884 2662
rect 9940 2716 9996 2726
rect 9492 2100 9772 2156
rect 9604 1974 9660 1986
rect 9604 1932 9606 1974
rect 9658 1932 9660 1974
rect 9604 1866 9660 1876
rect 8484 1596 8540 1606
rect 8484 1214 8540 1540
rect 8820 1372 8876 1382
rect 8820 1278 8876 1316
rect 9716 1370 9772 2100
rect 9940 1820 9996 2660
rect 10164 2044 10220 3444
rect 10780 3387 10836 3398
rect 10108 1988 10220 2044
rect 10724 3386 10836 3387
rect 10724 3334 10782 3386
rect 10834 3334 10836 3386
rect 10724 3322 10836 3334
rect 11116 3388 11172 3426
rect 11116 3322 11172 3332
rect 10108 1986 10164 1988
rect 10108 1934 10110 1986
rect 10162 1934 10164 1986
rect 10108 1922 10164 1934
rect 9940 1764 10108 1820
rect 9716 1318 9718 1370
rect 9770 1318 9772 1370
rect 9716 1306 9772 1318
rect 8484 1162 8486 1214
rect 8538 1162 8540 1214
rect 8484 1150 8540 1162
rect 10052 1214 10108 1764
rect 10724 1596 10780 3322
rect 10724 1530 10780 1540
rect 10836 1708 10892 1718
rect 10836 1370 10892 1652
rect 11284 1382 11340 3780
rect 12292 3724 12404 3734
rect 12348 3722 12404 3724
rect 12348 3670 12350 3722
rect 12402 3670 12404 3722
rect 12348 3668 12404 3670
rect 12628 3724 12684 5124
rect 12740 5114 12796 5124
rect 12898 4732 13162 4742
rect 12954 4676 13002 4732
rect 13058 4676 13106 4732
rect 12898 4666 13162 4676
rect 12796 4508 12852 4518
rect 12796 4414 12852 4452
rect 13300 4294 13356 5684
rect 13412 4954 13468 4966
rect 13412 4902 13414 4954
rect 13466 4902 13468 4954
rect 13412 4732 13468 4902
rect 13524 4956 13580 5836
rect 13860 5852 13916 5862
rect 13860 5758 13916 5796
rect 13524 4890 13580 4900
rect 13804 4954 13860 4966
rect 13804 4902 13806 4954
rect 13858 4902 13860 4954
rect 13412 4666 13468 4676
rect 13804 4620 13860 4902
rect 13804 4554 13860 4564
rect 13972 4508 14028 6020
rect 14308 6010 14364 6020
rect 14644 5850 14700 7028
rect 14756 6860 14812 7254
rect 14756 6794 14812 6804
rect 14980 7308 15036 7318
rect 14644 5798 14646 5850
rect 14698 5798 14700 5850
rect 14140 5740 14196 5750
rect 14644 5740 14700 5798
rect 14140 5646 14196 5684
rect 14364 5682 14420 5694
rect 14364 5630 14366 5682
rect 14418 5630 14420 5682
rect 14644 5674 14700 5684
rect 14980 5918 15036 7252
rect 16660 6972 16716 8372
rect 17276 8428 17332 8466
rect 17276 8362 17332 8372
rect 17444 8428 17500 9762
rect 18004 9814 18060 9826
rect 18116 9818 18172 9828
rect 18004 9772 18006 9814
rect 18058 9772 18060 9814
rect 18004 9706 18060 9716
rect 19348 9210 19404 9828
rect 19348 9158 19350 9210
rect 19402 9158 19404 9210
rect 19348 9146 19404 9158
rect 19460 9212 19516 9940
rect 20356 9882 20412 9894
rect 20356 9830 20358 9882
rect 20410 9830 20412 9882
rect 19628 9212 19684 9222
rect 19460 9210 19684 9212
rect 19460 9158 19630 9210
rect 19682 9158 19684 9210
rect 19460 9156 19684 9158
rect 19628 9146 19684 9156
rect 20356 9210 20412 9830
rect 21028 9884 21084 9894
rect 21476 9884 21532 11172
rect 21868 11228 21924 11238
rect 21868 10666 21924 11172
rect 23156 10780 23212 11876
rect 23156 10714 23212 10724
rect 21868 10614 21870 10666
rect 21922 10614 21924 10666
rect 21868 10602 21924 10614
rect 21700 10442 21756 10454
rect 21700 10390 21702 10442
rect 21754 10390 21756 10442
rect 21700 10108 21756 10390
rect 23380 10444 23436 12114
rect 23940 12122 23996 13076
rect 24164 13038 24220 13076
rect 24612 13132 24668 13142
rect 24500 13020 24556 13030
rect 24500 12950 24556 12964
rect 24500 12898 24502 12950
rect 24554 12898 24556 12950
rect 24500 12796 24556 12898
rect 23940 12070 23942 12122
rect 23994 12070 23996 12122
rect 23940 12058 23996 12070
rect 24388 12740 24500 12796
rect 24388 11676 24444 12740
rect 24500 12730 24556 12740
rect 24612 12358 24668 13076
rect 25340 13132 25396 13526
rect 25508 13580 25564 13616
rect 25508 13514 25564 13524
rect 25340 13066 25396 13076
rect 25620 12962 25676 13748
rect 26068 13758 26124 14634
rect 26348 14586 26404 14598
rect 26348 14534 26350 14586
rect 26402 14534 26404 14586
rect 26348 14532 26404 14534
rect 26740 14586 26796 15092
rect 27524 14710 27580 15260
rect 27916 15260 27972 15270
rect 27916 15166 27972 15204
rect 28252 15260 28364 15316
rect 28756 15484 28812 15494
rect 28756 15370 28812 15428
rect 28756 15318 28758 15370
rect 28810 15318 28812 15370
rect 29988 15382 30044 15988
rect 29988 15370 30100 15382
rect 28756 15306 28812 15318
rect 29204 15314 29260 15326
rect 29988 15318 30046 15370
rect 30098 15318 30100 15370
rect 29988 15316 30100 15318
rect 29204 15262 29206 15314
rect 29258 15262 29260 15314
rect 26740 14534 26742 14586
rect 26794 14534 26796 14586
rect 27412 14700 27468 14710
rect 27524 14698 27636 14710
rect 27524 14646 27582 14698
rect 27634 14646 27636 14698
rect 27524 14644 27636 14646
rect 27412 14608 27468 14644
rect 27580 14634 27636 14644
rect 27804 14700 27860 14710
rect 27412 14556 27414 14608
rect 27466 14556 27468 14608
rect 27804 14606 27860 14644
rect 27916 14700 27972 14710
rect 28252 14700 28308 15260
rect 27916 14698 28308 14700
rect 27916 14646 27918 14698
rect 27970 14646 28254 14698
rect 28306 14646 28308 14698
rect 27916 14644 28308 14646
rect 27916 14634 27972 14644
rect 28252 14634 28308 14644
rect 28364 15148 28420 15158
rect 28364 14698 28420 15092
rect 29204 15148 29260 15262
rect 29204 15082 29260 15092
rect 30044 15148 30100 15316
rect 30212 15260 30268 16100
rect 30772 16090 30828 16100
rect 31108 16116 31164 16884
rect 31220 16863 31276 16875
rect 31220 16811 31222 16863
rect 31274 16811 31276 16863
rect 31220 16716 31276 16811
rect 31220 16650 31276 16660
rect 31500 16828 31556 16838
rect 31500 16266 31556 16772
rect 31500 16214 31502 16266
rect 31554 16214 31556 16266
rect 31500 16202 31556 16214
rect 31108 16064 31110 16116
rect 31162 16064 31164 16116
rect 30548 16044 30604 16054
rect 30548 15950 30604 15988
rect 30772 15930 30828 15942
rect 30772 15878 30774 15930
rect 30826 15878 30828 15930
rect 30772 15484 30828 15878
rect 30772 15418 30828 15428
rect 30884 15372 30940 15382
rect 31108 15372 31164 16064
rect 31332 16044 31388 16054
rect 31332 15443 31388 15988
rect 31332 15391 31334 15443
rect 31386 15391 31388 15443
rect 31332 15379 31388 15391
rect 31612 15930 31668 15942
rect 31612 15878 31614 15930
rect 31666 15878 31668 15930
rect 30884 15370 31164 15372
rect 30884 15318 30886 15370
rect 30938 15318 31164 15370
rect 30884 15316 31164 15318
rect 31612 15372 31668 15878
rect 30884 15306 30940 15316
rect 30212 15194 30268 15204
rect 31220 15295 31276 15307
rect 31612 15306 31668 15316
rect 31220 15260 31222 15295
rect 31274 15260 31276 15295
rect 31220 15194 31276 15204
rect 32340 15296 32396 15308
rect 32340 15244 32342 15296
rect 32394 15244 32396 15296
rect 30044 15082 30100 15092
rect 30996 15148 31052 15158
rect 28364 14646 28366 14698
rect 28418 14646 28420 14698
rect 28364 14634 28420 14646
rect 30996 14710 31052 15092
rect 31836 15148 31892 15158
rect 31836 15054 31892 15092
rect 32004 15146 32060 15158
rect 32004 15094 32006 15146
rect 32058 15094 32060 15146
rect 32004 14812 32060 15094
rect 32340 14924 32396 15244
rect 32340 14858 32396 14868
rect 31836 14756 32060 14812
rect 30996 14698 31108 14710
rect 30996 14646 31054 14698
rect 31106 14646 31108 14698
rect 30996 14644 31108 14646
rect 31052 14634 31108 14644
rect 31836 14698 31892 14756
rect 31836 14646 31838 14698
rect 31890 14646 31892 14698
rect 31836 14634 31892 14646
rect 27412 14544 27468 14556
rect 31724 14588 31780 14598
rect 26740 14532 26796 14534
rect 26348 14476 26796 14532
rect 26908 14530 26964 14542
rect 26908 14478 26910 14530
rect 26962 14478 26964 14530
rect 26908 14028 26964 14478
rect 27244 14530 27300 14542
rect 27244 14478 27246 14530
rect 27298 14478 27300 14530
rect 27244 14364 27300 14478
rect 29316 14530 29372 14542
rect 29316 14478 29318 14530
rect 29370 14478 29372 14530
rect 31724 14494 31780 14532
rect 27244 14298 27300 14308
rect 27524 14364 27580 14374
rect 26908 13962 26964 13972
rect 27524 13914 27580 14308
rect 28700 14364 28756 14374
rect 28700 14270 28756 14308
rect 28812 14364 28868 14374
rect 29316 14364 29372 14478
rect 29932 14476 29988 14486
rect 30772 14476 30828 14486
rect 29932 14474 30044 14476
rect 29932 14422 29934 14474
rect 29986 14422 30044 14474
rect 29932 14410 30044 14422
rect 30772 14474 31052 14476
rect 30772 14422 30774 14474
rect 30826 14422 31052 14474
rect 30772 14420 31052 14422
rect 30772 14410 30828 14420
rect 28812 14362 29260 14364
rect 28812 14310 28814 14362
rect 28866 14310 29260 14362
rect 28812 14308 29260 14310
rect 28812 14298 28868 14308
rect 28778 14140 29042 14150
rect 28834 14084 28882 14140
rect 28938 14084 28986 14140
rect 28778 14074 29042 14084
rect 27524 13862 27526 13914
rect 27578 13862 27580 13914
rect 27524 13850 27580 13862
rect 27804 13916 27860 13926
rect 27804 13822 27860 13860
rect 26068 13706 26070 13758
rect 26122 13706 26124 13758
rect 24780 12908 24836 12918
rect 24780 12814 24836 12852
rect 25620 12910 25622 12962
rect 25674 12910 25676 12962
rect 25788 13578 25844 13590
rect 25788 13526 25790 13578
rect 25842 13526 25844 13578
rect 25788 13020 25844 13526
rect 26068 13132 26124 13706
rect 26068 13066 26124 13076
rect 26292 13758 26460 13804
rect 26292 13748 26406 13758
rect 25788 12954 25844 12964
rect 25620 12908 25676 12910
rect 26124 12908 26180 12918
rect 25620 12842 25676 12852
rect 26068 12906 26180 12908
rect 26068 12854 26126 12906
rect 26178 12854 26180 12906
rect 26068 12842 26180 12854
rect 24556 12346 24668 12358
rect 24556 12294 24558 12346
rect 24610 12294 24668 12346
rect 24556 12292 24668 12294
rect 25060 12796 25116 12806
rect 24556 12282 24612 12292
rect 25060 12178 25116 12740
rect 24500 12124 24556 12134
rect 25060 12126 25062 12178
rect 25114 12126 25116 12178
rect 25060 12114 25116 12126
rect 24500 12030 24556 12068
rect 24668 12010 24724 12022
rect 24668 11958 24670 12010
rect 24722 11958 24724 12010
rect 24668 11900 24724 11958
rect 24668 11834 24724 11844
rect 25788 12010 25844 12022
rect 25788 11958 25790 12010
rect 25842 11958 25844 12010
rect 24808 11788 25072 11798
rect 24864 11732 24912 11788
rect 24968 11732 25016 11788
rect 24808 11722 25072 11732
rect 25788 11676 25844 11958
rect 24388 11620 24668 11676
rect 24052 11452 24108 11462
rect 23716 11450 24108 11452
rect 23716 11398 24054 11450
rect 24106 11398 24108 11450
rect 23716 11396 24108 11398
rect 23548 10444 23604 10454
rect 23380 10442 23604 10444
rect 23380 10390 23550 10442
rect 23602 10390 23604 10442
rect 23380 10388 23604 10390
rect 23548 10332 23604 10388
rect 23548 10266 23604 10276
rect 21700 10052 21868 10108
rect 21028 9770 21084 9828
rect 21028 9718 21030 9770
rect 21082 9718 21084 9770
rect 21028 9706 21084 9718
rect 21364 9838 21532 9884
rect 21364 9786 21366 9838
rect 21418 9828 21532 9838
rect 21812 9838 21868 10052
rect 21418 9786 21420 9828
rect 21364 9660 21420 9786
rect 21812 9786 21814 9838
rect 21866 9786 21868 9838
rect 21812 9774 21868 9786
rect 23716 9660 23772 11396
rect 24052 11386 24108 11396
rect 24612 11340 24668 11620
rect 25788 11610 25844 11620
rect 26068 11676 26124 12842
rect 26292 12684 26348 13748
rect 26404 13706 26406 13748
rect 26458 13706 26460 13758
rect 29204 13746 29260 14308
rect 29316 14298 29372 14308
rect 29988 13814 30044 14410
rect 30996 13916 31052 14420
rect 31444 14362 31500 14374
rect 31444 14310 31446 14362
rect 31498 14310 31500 14362
rect 31108 13916 31164 13926
rect 30996 13914 31164 13916
rect 30996 13862 31110 13914
rect 31162 13862 31164 13914
rect 30996 13860 31164 13862
rect 31108 13850 31164 13860
rect 29988 13804 30100 13814
rect 29988 13802 30492 13804
rect 29988 13750 30046 13802
rect 30098 13750 30492 13802
rect 29988 13748 30492 13750
rect 26404 13694 26460 13706
rect 26628 13734 26684 13746
rect 26628 13682 26630 13734
rect 26682 13682 26684 13734
rect 29204 13694 29206 13746
rect 29258 13694 29260 13746
rect 30044 13738 30100 13748
rect 29204 13682 29260 13694
rect 26404 13580 26460 13590
rect 26404 13496 26460 13524
rect 26404 13444 26406 13496
rect 26458 13444 26460 13496
rect 26404 13432 26460 13444
rect 26628 13468 26684 13682
rect 27076 13580 27188 13590
rect 27132 13578 27188 13580
rect 27132 13526 27134 13578
rect 27186 13526 27188 13578
rect 27132 13524 27188 13526
rect 27076 13514 27188 13524
rect 27916 13580 27972 13590
rect 28252 13580 28308 13590
rect 27916 13578 28308 13580
rect 27916 13526 27918 13578
rect 27970 13526 28254 13578
rect 28306 13526 28308 13578
rect 27916 13524 28308 13526
rect 27916 13514 27972 13524
rect 26628 13402 26684 13412
rect 27300 13468 27356 13478
rect 27188 13132 27244 13142
rect 27188 12962 27244 13076
rect 26292 12618 26348 12628
rect 26852 12906 26908 12918
rect 26852 12854 26854 12906
rect 26906 12854 26908 12906
rect 26852 12346 26908 12854
rect 27188 12910 27190 12962
rect 27242 12910 27244 12962
rect 27188 12684 27244 12910
rect 27300 12856 27356 13412
rect 28252 13132 28308 13524
rect 28364 13580 28420 13590
rect 28364 13578 28476 13580
rect 28364 13526 28366 13578
rect 28418 13526 28476 13578
rect 28364 13514 28476 13526
rect 28420 13244 28476 13514
rect 28420 13188 28588 13244
rect 28252 13066 28308 13076
rect 28532 12962 28588 13188
rect 27300 12804 27302 12856
rect 27354 12804 27356 12856
rect 28028 12908 28084 12918
rect 28532 12910 28534 12962
rect 28586 12910 28588 12962
rect 28532 12898 28588 12910
rect 29204 13132 29260 13142
rect 28028 12814 28084 12852
rect 27300 12792 27356 12804
rect 27580 12796 27636 12806
rect 27916 12796 27972 12806
rect 27580 12794 27804 12796
rect 27580 12742 27582 12794
rect 27634 12742 27804 12794
rect 27580 12740 27804 12742
rect 27580 12730 27636 12740
rect 27188 12628 27524 12684
rect 26852 12294 26854 12346
rect 26906 12294 26908 12346
rect 26852 12282 26908 12294
rect 27468 12234 27524 12628
rect 27468 12182 27470 12234
rect 27522 12182 27524 12234
rect 27188 12160 27244 12172
rect 27468 12170 27524 12182
rect 26628 12124 26684 12134
rect 26628 12030 26684 12068
rect 27188 12124 27190 12160
rect 27242 12124 27244 12160
rect 26068 11610 26124 11620
rect 25284 11450 25340 11462
rect 25284 11398 25286 11450
rect 25338 11398 25340 11450
rect 24724 11340 24780 11350
rect 24612 11338 24780 11340
rect 24612 11286 24726 11338
rect 24778 11286 24780 11338
rect 24612 11284 24780 11286
rect 24724 11274 24780 11284
rect 25284 10790 25340 11398
rect 26852 11452 26908 11462
rect 26852 11358 26908 11396
rect 26572 11282 26628 11294
rect 26572 11230 26574 11282
rect 26626 11230 26628 11282
rect 23996 10780 24052 10790
rect 23996 10686 24052 10724
rect 24556 10780 24612 10790
rect 24556 10686 24612 10724
rect 25284 10780 25396 10790
rect 25340 10778 25396 10780
rect 25340 10726 25342 10778
rect 25394 10726 25396 10778
rect 25340 10724 25396 10726
rect 26572 10780 26628 11230
rect 26572 10724 26684 10780
rect 25284 10714 25396 10724
rect 25284 10648 25340 10714
rect 24108 10556 24164 10566
rect 24108 10462 24164 10500
rect 24892 10556 24948 10566
rect 24892 10462 24948 10500
rect 25452 10556 25508 10566
rect 25844 10556 25900 10566
rect 25452 10554 25900 10556
rect 25452 10502 25454 10554
rect 25506 10502 25846 10554
rect 25898 10502 25900 10554
rect 25452 10500 25900 10502
rect 25452 10490 25508 10500
rect 25844 10490 25900 10500
rect 26068 10556 26124 10566
rect 24444 10444 24500 10454
rect 24444 10350 24500 10388
rect 25004 10444 25060 10482
rect 25004 10378 25060 10388
rect 25956 10444 26012 10454
rect 24808 10220 25072 10230
rect 24864 10164 24912 10220
rect 24968 10164 25016 10220
rect 24808 10154 25072 10164
rect 24836 9996 24892 10006
rect 24164 9884 24220 9894
rect 21252 9604 21420 9660
rect 23492 9604 23772 9660
rect 24052 9882 24220 9884
rect 24052 9830 24166 9882
rect 24218 9830 24220 9882
rect 24052 9828 24220 9830
rect 20838 9436 21102 9446
rect 20894 9380 20942 9436
rect 20998 9380 21046 9436
rect 20838 9370 21102 9380
rect 20356 9158 20358 9210
rect 20410 9158 20412 9210
rect 20356 9146 20412 9158
rect 20692 9024 20748 9036
rect 19964 8988 20020 8998
rect 18676 8876 18732 8886
rect 19740 8876 19796 8886
rect 18676 8874 18956 8876
rect 18676 8822 18678 8874
rect 18730 8822 18956 8874
rect 18676 8820 18956 8822
rect 18676 8810 18732 8820
rect 17444 8362 17500 8372
rect 18900 8426 18956 8820
rect 19740 8874 19852 8876
rect 19740 8822 19742 8874
rect 19794 8822 19852 8874
rect 19740 8810 19852 8822
rect 18900 8374 18902 8426
rect 18954 8374 18956 8426
rect 18900 8362 18956 8374
rect 19796 8336 19852 8810
rect 17556 8316 17612 8326
rect 17556 8222 17612 8260
rect 17948 8316 18004 8326
rect 18620 8316 18676 8326
rect 19292 8316 19348 8326
rect 17948 8314 18172 8316
rect 17948 8262 17950 8314
rect 18002 8262 18172 8314
rect 17948 8260 18172 8262
rect 17948 8250 18004 8260
rect 16884 8204 16940 8214
rect 16884 8110 16940 8148
rect 17668 7700 18060 7756
rect 17444 7644 17500 7654
rect 17668 7644 17724 7700
rect 16996 7642 17724 7644
rect 16884 7580 16940 7592
rect 16884 7532 16886 7580
rect 16938 7532 16940 7580
rect 16884 7466 16940 7476
rect 16996 7590 17446 7642
rect 17498 7590 17724 7642
rect 16996 7588 17724 7590
rect 16996 7318 17052 7588
rect 17164 7420 17220 7430
rect 17164 7418 17276 7420
rect 17164 7366 17166 7418
rect 17218 7366 17276 7418
rect 17164 7354 17276 7366
rect 16940 7306 17052 7318
rect 16940 7254 16942 7306
rect 16994 7254 17052 7306
rect 16940 7252 17052 7254
rect 16940 7242 16996 7252
rect 16868 7084 17132 7094
rect 16924 7028 16972 7084
rect 17028 7028 17076 7084
rect 16868 7018 17132 7028
rect 16660 6916 16828 6972
rect 16772 6870 16828 6916
rect 15988 6860 16044 6870
rect 16772 6858 16884 6870
rect 16772 6806 16830 6858
rect 16882 6806 16884 6858
rect 16772 6804 16884 6806
rect 15988 6766 16044 6804
rect 16828 6794 16884 6804
rect 17220 6636 17276 7354
rect 17220 6570 17276 6580
rect 14980 5866 14982 5918
rect 15034 5866 15036 5918
rect 16660 6522 16716 6534
rect 16660 6470 16662 6522
rect 16714 6470 16716 6522
rect 14364 5516 14420 5630
rect 14364 5450 14420 5460
rect 14980 5348 15036 5866
rect 15540 5894 15596 5906
rect 15540 5852 15542 5894
rect 15594 5852 15596 5894
rect 15540 5786 15596 5796
rect 16380 5740 16436 5750
rect 14644 5292 15036 5348
rect 15372 5516 15428 5526
rect 15372 5346 15428 5460
rect 15372 5294 15374 5346
rect 15426 5294 15428 5346
rect 14532 5180 14588 5190
rect 14532 5086 14588 5124
rect 14140 4956 14196 4966
rect 14140 4862 14196 4900
rect 13972 4442 14028 4452
rect 14644 4406 14700 5292
rect 15372 5282 15428 5294
rect 15764 5236 16044 5292
rect 14756 5224 14812 5236
rect 14756 5172 14758 5224
rect 14810 5172 14812 5224
rect 14756 4732 14812 5172
rect 14868 5180 14924 5190
rect 14868 4956 14924 5124
rect 15596 5180 15652 5218
rect 15596 5114 15652 5124
rect 14980 5068 15036 5078
rect 15036 5012 15148 5068
rect 14980 5002 15036 5012
rect 14868 4890 14924 4900
rect 14756 4666 14812 4676
rect 14532 4396 14588 4406
rect 14644 4394 14756 4406
rect 14644 4342 14702 4394
rect 14754 4342 14756 4394
rect 14644 4340 14756 4342
rect 14532 4298 14534 4340
rect 14586 4298 14588 4340
rect 13076 4284 13132 4294
rect 12740 3724 12796 3734
rect 12628 3722 12796 3724
rect 12628 3670 12742 3722
rect 12794 3670 12796 3722
rect 12628 3668 12796 3670
rect 11732 3656 11788 3668
rect 12292 3658 12404 3668
rect 12740 3658 12796 3668
rect 11508 3610 11564 3622
rect 11508 3558 11510 3610
rect 11562 3558 11564 3610
rect 11508 3387 11564 3558
rect 11732 3612 11734 3656
rect 11786 3612 11788 3656
rect 11732 3546 11788 3556
rect 13076 3554 13132 4228
rect 13244 4282 13356 4294
rect 13244 4230 13246 4282
rect 13298 4230 13356 4282
rect 13244 4228 13356 4230
rect 13412 4284 13468 4294
rect 13916 4284 13972 4294
rect 14140 4284 14196 4294
rect 13244 4218 13300 4228
rect 13412 4190 13468 4228
rect 13860 4282 13972 4284
rect 13860 4230 13918 4282
rect 13970 4230 13972 4282
rect 13860 4218 13972 4230
rect 14084 4282 14196 4284
rect 14084 4230 14142 4282
rect 14194 4230 14196 4282
rect 14084 4218 14196 4230
rect 13580 4170 13636 4182
rect 13580 4118 13582 4170
rect 13634 4118 13636 4170
rect 13076 3502 13078 3554
rect 13130 3502 13132 3554
rect 13076 3490 13132 3502
rect 13188 3948 13244 3958
rect 10836 1318 10838 1370
rect 10890 1318 10892 1370
rect 10836 1306 10892 1318
rect 11228 1370 11340 1382
rect 11228 1318 11230 1370
rect 11282 1318 11340 1370
rect 11228 1316 11340 1318
rect 11396 3331 11564 3387
rect 13188 3448 13244 3892
rect 13468 3836 13524 3846
rect 13580 3836 13636 4118
rect 13524 3780 13636 3836
rect 13468 3610 13524 3780
rect 13468 3558 13470 3610
rect 13522 3558 13524 3610
rect 13468 3546 13524 3558
rect 13748 3556 13804 3566
rect 13860 3556 13916 4218
rect 14084 3724 14140 4218
rect 14308 4088 14364 4100
rect 14028 3666 14140 3724
rect 14028 3614 14030 3666
rect 14082 3614 14140 3666
rect 14028 3602 14140 3614
rect 13748 3554 13916 3556
rect 13188 3396 13190 3448
rect 13242 3396 13244 3448
rect 13188 3384 13244 3396
rect 13748 3502 13750 3554
rect 13802 3502 13916 3554
rect 13748 3500 13916 3502
rect 13748 3388 13804 3500
rect 11228 1306 11284 1316
rect 10052 1162 10054 1214
rect 10106 1162 10108 1214
rect 10052 1150 10108 1162
rect 10500 1184 10556 1196
rect 10500 1148 10502 1184
rect 10554 1148 10556 1184
rect 10500 1082 10556 1092
rect 11396 1036 11452 3331
rect 13748 3322 13804 3332
rect 12898 3164 13162 3174
rect 12954 3108 13002 3164
rect 13058 3108 13106 3164
rect 12898 3098 13162 3108
rect 13468 2828 13524 2838
rect 12180 2758 12236 2770
rect 12180 2706 12182 2758
rect 12234 2706 12236 2758
rect 12068 2268 12124 2278
rect 11508 2156 11564 2166
rect 11508 1932 11564 2100
rect 12068 2044 12124 2212
rect 11508 1876 11620 1932
rect 11564 1426 11620 1876
rect 11564 1374 11566 1426
rect 11618 1374 11620 1426
rect 11564 1362 11620 1374
rect 8372 980 8540 1036
rect 5796 952 5852 980
rect 5796 900 5798 952
rect 5850 900 5852 952
rect 5796 888 5852 900
rect 8484 800 8540 980
rect 11396 970 11452 980
rect 11956 1146 12012 1158
rect 11956 1094 11958 1146
rect 12010 1094 12012 1146
rect 11956 1036 12012 1094
rect 12068 1102 12124 1988
rect 12180 1372 12236 2706
rect 12740 2758 12796 2770
rect 12740 2706 12742 2758
rect 12794 2706 12796 2758
rect 12404 2044 12460 2054
rect 12404 1950 12460 1988
rect 12740 1932 12796 2706
rect 13244 2604 13300 2614
rect 13468 2604 13524 2772
rect 13244 2602 13524 2604
rect 13244 2550 13246 2602
rect 13298 2550 13470 2602
rect 13522 2550 13524 2602
rect 13244 2548 13524 2550
rect 13244 2538 13356 2548
rect 13468 2538 13524 2548
rect 14084 2770 14140 3602
rect 14084 2718 14086 2770
rect 14138 2718 14140 2770
rect 12740 1866 12796 1876
rect 13076 2268 13132 2278
rect 13076 1930 13132 2212
rect 13076 1878 13078 1930
rect 13130 1878 13132 1930
rect 13076 1866 13132 1878
rect 13300 1974 13356 2538
rect 14084 2156 14140 2718
rect 14084 2090 14140 2100
rect 14196 4060 14252 4070
rect 14196 3610 14252 4004
rect 14196 3558 14198 3610
rect 14250 3558 14252 3610
rect 14196 2882 14252 3558
rect 14308 4036 14310 4088
rect 14362 4036 14364 4088
rect 14308 3612 14364 4036
rect 14532 4060 14588 4298
rect 14700 4284 14756 4340
rect 15092 4326 15148 5012
rect 15652 5010 15708 5022
rect 15652 4958 15654 5010
rect 15706 4958 15708 5010
rect 15652 4956 15708 4958
rect 15764 4956 15820 5236
rect 15988 5180 16044 5236
rect 15988 5124 16100 5180
rect 16044 5122 16100 5124
rect 14700 4218 14756 4228
rect 14868 4284 14924 4294
rect 14532 3994 14588 4004
rect 14588 3836 14644 3846
rect 14588 3722 14644 3780
rect 14588 3670 14590 3722
rect 14642 3670 14644 3722
rect 14588 3658 14644 3670
rect 14308 3546 14364 3556
rect 14196 2830 14198 2882
rect 14250 2830 14252 2882
rect 13300 1932 13302 1974
rect 13354 1932 13356 1974
rect 13300 1866 13356 1876
rect 13860 1974 13916 1986
rect 13860 1922 13862 1974
rect 13914 1922 13916 1974
rect 13860 1708 13916 1922
rect 13860 1642 13916 1652
rect 12898 1596 13162 1606
rect 12954 1540 13002 1596
rect 13058 1540 13106 1596
rect 12898 1530 13162 1540
rect 12180 1306 12236 1316
rect 14084 1372 14140 1382
rect 14196 1372 14252 2830
rect 14868 2828 14924 4228
rect 15092 4274 15094 4326
rect 15146 4274 15148 4326
rect 14868 2762 14924 2772
rect 14980 3542 15036 3554
rect 14980 3490 14982 3542
rect 15034 3490 15036 3542
rect 14868 2604 14924 2614
rect 14980 2604 15036 3490
rect 15092 3500 15148 4274
rect 15316 4900 15820 4956
rect 15876 5110 15932 5122
rect 15876 5058 15878 5110
rect 15930 5058 15932 5110
rect 16044 5070 16046 5122
rect 16098 5070 16100 5122
rect 16044 5058 16100 5070
rect 16380 5122 16436 5684
rect 16660 5516 16716 6470
rect 16660 5450 16716 5460
rect 16868 5516 17132 5526
rect 16924 5460 16972 5516
rect 17028 5460 17076 5516
rect 16868 5450 17132 5460
rect 16604 5180 16660 5190
rect 16380 5070 16382 5122
rect 16434 5070 16436 5122
rect 15316 4350 15372 4900
rect 15876 4508 15932 5058
rect 16380 4732 16436 5070
rect 16380 4666 16436 4676
rect 16548 5178 16660 5180
rect 16548 5126 16606 5178
rect 16658 5126 16660 5178
rect 16548 5114 16660 5126
rect 17332 5180 17388 7588
rect 17444 7578 17500 7588
rect 17780 7532 17836 7542
rect 17780 7434 17782 7476
rect 17834 7434 17836 7476
rect 17780 6748 17836 7434
rect 18004 7420 18060 7700
rect 18116 7654 18172 8260
rect 18620 8314 18732 8316
rect 18620 8262 18622 8314
rect 18674 8262 18732 8314
rect 18620 8250 18732 8262
rect 19292 8314 19516 8316
rect 19292 8262 19294 8314
rect 19346 8262 19516 8314
rect 19292 8260 19516 8262
rect 19292 8250 19348 8260
rect 18228 8092 18284 8102
rect 18228 8090 18396 8092
rect 18228 8038 18230 8090
rect 18282 8038 18396 8090
rect 18228 8036 18396 8038
rect 18228 8026 18284 8036
rect 18116 7642 18228 7654
rect 18116 7590 18174 7642
rect 18226 7590 18228 7642
rect 18116 7588 18228 7590
rect 18172 7578 18228 7588
rect 18116 7474 18172 7486
rect 18116 7422 18118 7474
rect 18170 7422 18172 7474
rect 18116 7420 18172 7422
rect 18004 7364 18172 7420
rect 17780 6682 17836 6692
rect 17892 6972 17948 6982
rect 17892 6708 17948 6916
rect 18340 6860 18396 8036
rect 18508 7644 18564 7654
rect 18508 7550 18564 7588
rect 18676 7084 18732 8250
rect 19460 8092 19516 8260
rect 19740 8314 19852 8336
rect 19740 8262 19742 8314
rect 19794 8262 19852 8314
rect 19740 8250 19852 8262
rect 19964 8314 20020 8932
rect 20356 8988 20412 8998
rect 19964 8262 19966 8314
rect 20018 8262 20020 8314
rect 19964 8250 20020 8262
rect 20132 8316 20188 8326
rect 19796 8204 19852 8250
rect 19628 8092 19684 8102
rect 19460 8090 19684 8092
rect 19460 8038 19630 8090
rect 19682 8038 19684 8090
rect 19460 8036 19684 8038
rect 19628 8026 19684 8036
rect 19572 7644 19628 7654
rect 19796 7644 19852 8148
rect 19572 7642 19852 7644
rect 19572 7590 19574 7642
rect 19626 7590 19852 7642
rect 19572 7588 19852 7590
rect 19572 7578 19628 7588
rect 19236 7456 19292 7468
rect 18844 7420 18900 7430
rect 18844 7326 18900 7364
rect 19236 7420 19238 7456
rect 19290 7420 19292 7456
rect 19236 7354 19292 7364
rect 19852 7308 19908 7318
rect 19796 7306 19908 7308
rect 19796 7254 19854 7306
rect 19906 7254 19908 7306
rect 19796 7242 19908 7254
rect 18676 7028 18956 7084
rect 17892 6656 17894 6708
rect 17946 6656 17948 6708
rect 17892 6644 17948 6656
rect 18004 6804 18396 6860
rect 17892 5852 17948 5862
rect 18004 5852 18060 6804
rect 18676 6748 18732 6758
rect 18676 6656 18678 6692
rect 18730 6656 18732 6692
rect 17892 5850 18060 5852
rect 17892 5798 17894 5850
rect 17946 5798 18060 5850
rect 17892 5796 18060 5798
rect 18228 6636 18284 6646
rect 18676 6644 18732 6656
rect 17892 5786 17948 5796
rect 18228 5190 18284 6580
rect 18564 6188 18620 6198
rect 18564 6074 18620 6132
rect 18564 6022 18566 6074
rect 18618 6022 18620 6074
rect 18564 6010 18620 6022
rect 18788 5852 18844 5862
rect 18564 5796 18788 5852
rect 17332 5122 17388 5124
rect 15876 4452 16044 4508
rect 15316 4298 15318 4350
rect 15370 4298 15372 4350
rect 15092 3434 15148 3444
rect 15204 3778 15260 3790
rect 15204 3726 15206 3778
rect 15258 3726 15260 3778
rect 15204 3052 15260 3726
rect 15316 3566 15372 4298
rect 15652 4326 15708 4338
rect 15652 4274 15654 4326
rect 15706 4274 15708 4326
rect 15316 3514 15318 3566
rect 15370 3514 15372 3566
rect 15316 3502 15372 3514
rect 15428 4088 15484 4100
rect 15428 4036 15430 4088
rect 15482 4036 15484 4088
rect 15204 2996 15372 3052
rect 14868 2602 15036 2604
rect 14868 2550 14870 2602
rect 14922 2550 15036 2602
rect 14868 2548 15036 2550
rect 15204 2826 15260 2838
rect 15204 2774 15206 2826
rect 15258 2774 15260 2826
rect 14868 2538 14924 2548
rect 15204 1932 15260 2774
rect 15204 1866 15260 1876
rect 15316 1596 15372 2996
rect 15428 2716 15484 4036
rect 15652 3724 15708 4274
rect 15876 4326 15932 4338
rect 15876 4284 15878 4326
rect 15930 4284 15932 4326
rect 15876 4218 15932 4228
rect 15988 3948 16044 4452
rect 16548 4396 16604 5114
rect 17332 5070 17334 5122
rect 17386 5070 17388 5122
rect 17724 5180 17780 5190
rect 18172 5180 18284 5190
rect 17724 5178 18284 5180
rect 17724 5126 17726 5178
rect 17778 5126 18174 5178
rect 18226 5126 18284 5178
rect 17724 5124 18284 5126
rect 17724 5114 17780 5124
rect 18172 5114 18284 5124
rect 17332 5048 17388 5070
rect 16660 5010 16716 5022
rect 16660 4958 16662 5010
rect 16714 4958 16716 5010
rect 16660 4956 16716 4958
rect 16660 4890 16716 4900
rect 17444 5004 17500 5016
rect 17444 4952 17446 5004
rect 17498 4952 17500 5004
rect 17444 4844 17500 4952
rect 17444 4778 17500 4788
rect 17892 4956 17948 4966
rect 15652 3658 15708 3668
rect 15932 3892 16044 3948
rect 16436 4326 16492 4338
rect 16548 4330 16604 4340
rect 16436 4274 16438 4326
rect 16490 4274 16492 4326
rect 15932 3836 15988 3892
rect 15932 3666 15988 3780
rect 15932 3614 15934 3666
rect 15986 3614 15988 3666
rect 15932 3602 15988 3614
rect 16156 3612 16212 3622
rect 16156 3554 16212 3556
rect 15540 3542 15596 3554
rect 15540 3500 15542 3542
rect 15594 3500 15596 3542
rect 16156 3502 16158 3554
rect 16210 3502 16212 3554
rect 16156 3490 16212 3502
rect 15540 3434 15596 3444
rect 15428 2660 15596 2716
rect 15316 1530 15372 1540
rect 15428 1820 15484 1830
rect 14812 1372 14868 1382
rect 14084 1370 14868 1372
rect 14084 1318 14086 1370
rect 14138 1318 14814 1370
rect 14866 1318 14868 1370
rect 14084 1316 14868 1318
rect 14084 1306 14140 1316
rect 14812 1306 14868 1316
rect 13356 1260 13412 1270
rect 13356 1166 13412 1204
rect 13748 1260 13804 1270
rect 13748 1146 13804 1204
rect 12068 1090 12180 1102
rect 12068 1046 12126 1090
rect 12124 1038 12126 1046
rect 12178 1038 12180 1090
rect 13748 1094 13750 1146
rect 13802 1094 13804 1146
rect 13748 1082 13804 1094
rect 14476 1148 14532 1158
rect 14476 1054 14532 1092
rect 15204 1148 15260 1158
rect 15204 1054 15260 1092
rect 15428 1100 15484 1764
rect 12124 1026 12180 1038
rect 15428 1048 15430 1100
rect 15482 1048 15484 1100
rect 15540 1148 15596 2660
rect 15876 2604 15932 2614
rect 15876 2510 15932 2548
rect 16212 2042 16268 2054
rect 16212 1990 16214 2042
rect 16266 1990 16268 2042
rect 16212 1372 16268 1990
rect 16212 1306 16268 1316
rect 16436 1370 16492 4274
rect 17220 4284 17276 4294
rect 16868 3948 17132 3958
rect 16924 3892 16972 3948
rect 17028 3892 17076 3948
rect 16868 3882 17132 3892
rect 16548 3724 16604 3734
rect 16548 3630 16604 3668
rect 17220 3568 17276 4228
rect 17332 3568 17388 3578
rect 17220 3566 17388 3568
rect 17220 3514 17334 3566
rect 17386 3514 17388 3566
rect 17220 3512 17388 3514
rect 16868 2380 17132 2390
rect 16924 2324 16972 2380
rect 17028 2324 17076 2380
rect 16868 2314 17132 2324
rect 17220 2166 17276 3512
rect 17332 3502 17388 3512
rect 17892 3566 17948 4900
rect 18228 4956 18284 5114
rect 18452 5180 18508 5190
rect 18452 5078 18454 5124
rect 18506 5078 18508 5124
rect 18452 5066 18508 5078
rect 18228 4890 18284 4900
rect 18340 5004 18396 5016
rect 18340 4952 18342 5004
rect 18394 4952 18396 5004
rect 18340 4396 18396 4952
rect 18340 4330 18396 4340
rect 18564 4172 18620 5796
rect 18788 5758 18844 5796
rect 18788 5180 18844 5190
rect 18788 5122 18844 5124
rect 18788 5070 18790 5122
rect 18842 5070 18844 5122
rect 18788 5058 18844 5070
rect 18900 5016 18956 7028
rect 19236 6972 19292 6982
rect 19236 6870 19292 6916
rect 19796 6972 19852 7242
rect 19796 6906 19852 6916
rect 19236 6858 19348 6870
rect 19236 6806 19294 6858
rect 19346 6806 19348 6858
rect 19236 6794 19348 6806
rect 19012 6522 19068 6534
rect 19012 6470 19014 6522
rect 19066 6470 19068 6522
rect 19012 6412 19068 6470
rect 19012 6346 19068 6356
rect 19236 5862 19292 6794
rect 20132 6748 20188 8260
rect 20356 8102 20412 8932
rect 20692 8972 20694 9024
rect 20746 8972 20748 9024
rect 20524 8428 20580 8438
rect 20692 8428 20748 8972
rect 20524 8426 20748 8428
rect 20524 8374 20526 8426
rect 20578 8374 20748 8426
rect 20524 8372 20748 8374
rect 20972 8428 21028 8438
rect 21252 8428 21308 9604
rect 22260 9212 22316 9222
rect 21588 9148 21644 9160
rect 21588 9100 21590 9148
rect 21642 9100 21644 9148
rect 22260 9118 22316 9156
rect 23492 9210 23548 9604
rect 23492 9158 23494 9210
rect 23546 9158 23548 9210
rect 23492 9146 23548 9158
rect 23156 9100 23212 9110
rect 21588 9034 21644 9044
rect 21700 9034 21756 9046
rect 21420 8988 21476 8998
rect 21420 8894 21476 8932
rect 21700 8982 21702 9034
rect 21754 8982 21756 9034
rect 23156 9002 23158 9044
rect 23210 9002 23212 9044
rect 23156 8990 23212 9002
rect 20972 8426 21308 8428
rect 20972 8374 20974 8426
rect 21026 8374 21308 8426
rect 20972 8372 21308 8374
rect 20524 8362 20580 8372
rect 20972 8362 21028 8372
rect 21252 8316 21308 8372
rect 20804 8258 20860 8270
rect 20804 8206 20806 8258
rect 20858 8206 20860 8258
rect 21252 8250 21308 8260
rect 20804 8204 20860 8206
rect 20804 8138 20860 8148
rect 21700 8204 21756 8982
rect 22652 8876 22708 8886
rect 22652 8874 22764 8876
rect 22652 8822 22654 8874
rect 22706 8822 22764 8874
rect 22652 8810 22764 8822
rect 22036 8370 22092 8382
rect 22036 8318 22038 8370
rect 22090 8318 22092 8370
rect 22036 8316 22092 8318
rect 22036 8250 22092 8260
rect 22372 8258 22428 8270
rect 20356 8090 20468 8102
rect 20356 8038 20414 8090
rect 20466 8038 20468 8090
rect 20356 8036 20468 8038
rect 20244 7644 20300 7654
rect 20412 7644 20468 8036
rect 20838 7868 21102 7878
rect 20894 7812 20942 7868
rect 20998 7812 21046 7868
rect 20838 7802 21102 7812
rect 20300 7588 20468 7644
rect 20244 7550 20300 7588
rect 21700 7474 21756 8148
rect 21924 8204 21980 8214
rect 21924 7592 21980 8148
rect 21924 7540 21926 7592
rect 21978 7540 21980 7592
rect 21924 7528 21980 7540
rect 22372 8206 22374 8258
rect 22426 8206 22428 8258
rect 22372 7542 22428 8206
rect 22708 7654 22764 8810
rect 24052 8426 24108 9828
rect 24164 9818 24220 9828
rect 24836 9770 24892 9940
rect 25956 9826 26012 10388
rect 25228 9772 25284 9782
rect 25452 9772 25508 9782
rect 24836 9718 24838 9770
rect 24890 9718 24892 9770
rect 24836 9706 24892 9718
rect 25172 9770 25508 9772
rect 25172 9718 25230 9770
rect 25282 9718 25454 9770
rect 25506 9718 25508 9770
rect 25956 9774 25958 9826
rect 26010 9774 26012 9826
rect 25956 9762 26012 9774
rect 25172 9716 25508 9718
rect 25172 9706 25284 9716
rect 25452 9706 25508 9716
rect 24052 8374 24054 8426
rect 24106 8374 24108 8426
rect 24052 8362 24108 8374
rect 24164 8986 24220 8998
rect 24164 8934 24166 8986
rect 24218 8934 24220 8986
rect 24164 8876 24220 8934
rect 24164 8427 24220 8820
rect 24808 8652 25072 8662
rect 24864 8596 24912 8652
rect 24968 8596 25016 8652
rect 24808 8586 25072 8596
rect 24164 8371 24332 8427
rect 24276 8326 24332 8371
rect 24276 8314 24388 8326
rect 24276 8262 24334 8314
rect 24386 8262 24388 8314
rect 24276 8260 24388 8262
rect 23716 8246 23772 8258
rect 24332 8250 24388 8260
rect 24500 8316 24556 8326
rect 23716 8204 23718 8246
rect 23770 8204 23772 8246
rect 23716 8138 23772 8148
rect 24500 8152 24556 8260
rect 24500 8100 24502 8152
rect 24554 8100 24556 8152
rect 24500 8088 24556 8100
rect 24612 8250 24668 8262
rect 24612 8198 24614 8250
rect 24666 8198 24668 8250
rect 22708 7644 22876 7654
rect 22708 7642 22820 7644
rect 22708 7590 22766 7642
rect 22818 7590 22820 7642
rect 22708 7588 22820 7590
rect 22764 7578 22876 7588
rect 22372 7530 22484 7542
rect 22372 7478 22430 7530
rect 22482 7478 22484 7530
rect 22372 7476 22484 7478
rect 21700 7422 21702 7474
rect 21754 7422 21756 7474
rect 22428 7466 22484 7476
rect 23380 7456 23436 7468
rect 21700 7410 21756 7422
rect 22092 7420 22148 7430
rect 22092 7418 22204 7420
rect 22092 7366 22094 7418
rect 22146 7366 22204 7418
rect 22092 7354 22204 7366
rect 21700 6860 21756 6870
rect 20132 6702 20300 6748
rect 20132 6692 20246 6702
rect 20244 6650 20246 6692
rect 20298 6650 20300 6702
rect 19684 6636 19740 6646
rect 19684 6542 19740 6580
rect 19796 6412 19852 6422
rect 19180 5850 19292 5862
rect 19180 5798 19182 5850
rect 19234 5798 19292 5850
rect 19180 5796 19292 5798
rect 19684 5852 19740 5862
rect 19180 5786 19236 5796
rect 19684 5758 19740 5796
rect 18900 4964 18902 5016
rect 18954 4964 18956 5016
rect 19796 5068 19852 6356
rect 20244 6076 20300 6650
rect 20860 6690 20916 6702
rect 20860 6638 20862 6690
rect 20914 6638 20916 6690
rect 20860 6636 20916 6638
rect 20860 6580 21308 6636
rect 20838 6300 21102 6310
rect 20894 6244 20942 6300
rect 20998 6244 21046 6300
rect 20838 6234 21102 6244
rect 20244 6020 20468 6076
rect 20356 5962 20468 6020
rect 21252 6074 21308 6580
rect 21252 6022 21254 6074
rect 21306 6022 21308 6074
rect 21252 6010 21308 6022
rect 20356 5910 20414 5962
rect 20466 5910 20468 5962
rect 20356 5898 20468 5910
rect 20020 5852 20076 5862
rect 20020 5738 20076 5796
rect 20020 5686 20022 5738
rect 20074 5686 20076 5738
rect 20020 5674 20076 5686
rect 19964 5292 20020 5302
rect 19964 5234 20020 5236
rect 19964 5182 19966 5234
rect 20018 5182 20020 5234
rect 19964 5170 20020 5182
rect 19796 5012 20076 5068
rect 18900 4952 18956 4964
rect 19180 4956 19236 4966
rect 19180 4862 19236 4900
rect 19516 4954 19572 4966
rect 19516 4902 19518 4954
rect 19570 4902 19572 4954
rect 19516 4732 19572 4902
rect 19516 4666 19572 4676
rect 19628 4954 19684 4966
rect 19628 4902 19630 4954
rect 19682 4902 19684 4954
rect 19628 4508 19684 4902
rect 19628 4442 19684 4452
rect 19740 4844 19796 4854
rect 19740 4506 19796 4788
rect 19740 4454 19742 4506
rect 19794 4454 19796 4506
rect 19740 4442 19796 4454
rect 19460 4396 19516 4406
rect 19236 4394 19516 4396
rect 19236 4342 19462 4394
rect 19514 4342 19516 4394
rect 19236 4340 19516 4342
rect 18564 3568 18620 4116
rect 18788 4172 18844 4182
rect 18788 4078 18844 4116
rect 17892 3514 17894 3566
rect 17946 3514 17948 3566
rect 17892 3502 17948 3514
rect 18340 3512 18620 3568
rect 18172 2770 18228 2782
rect 18172 2718 18174 2770
rect 18226 2718 18228 2770
rect 18172 2716 18228 2718
rect 17556 2660 18228 2716
rect 17220 2156 17332 2166
rect 17220 2100 17276 2156
rect 17276 2024 17332 2100
rect 16436 1318 16438 1370
rect 16490 1318 16492 1370
rect 16436 1306 16492 1318
rect 16604 1820 16660 1830
rect 16604 1258 16660 1764
rect 16884 1820 16940 1830
rect 16884 1726 16940 1764
rect 16604 1206 16606 1258
rect 16658 1206 16660 1258
rect 16604 1194 16660 1206
rect 17220 1596 17276 1606
rect 17220 1214 17276 1540
rect 17556 1370 17612 2660
rect 18340 2604 18396 3512
rect 17948 2548 18396 2604
rect 18676 2828 18732 2838
rect 18676 2758 18732 2772
rect 18676 2706 18678 2758
rect 18730 2706 18732 2758
rect 17948 2042 18004 2548
rect 18564 2156 18620 2166
rect 18676 2156 18732 2706
rect 19236 2716 19292 4340
rect 19460 4330 19516 4340
rect 20020 4346 20076 5012
rect 20188 4898 20244 4910
rect 20188 4846 20190 4898
rect 20242 4846 20244 4898
rect 20188 4348 20244 4846
rect 20356 4620 20412 5898
rect 21588 5888 21644 5900
rect 20580 5852 20636 5862
rect 20580 5516 20636 5796
rect 20356 4554 20412 4564
rect 20468 5460 20636 5516
rect 21588 5836 21590 5888
rect 21642 5836 21644 5888
rect 20020 4294 20022 4346
rect 20074 4294 20076 4346
rect 19852 4170 19908 4182
rect 19852 4118 19854 4170
rect 19906 4118 19908 4170
rect 19852 4060 19908 4118
rect 19460 4004 19908 4060
rect 19460 2726 19516 4004
rect 19796 3836 19852 3846
rect 19796 3500 19852 3780
rect 19628 2828 19684 2838
rect 19628 2734 19684 2772
rect 19236 2650 19292 2660
rect 19404 2714 19516 2726
rect 19404 2662 19406 2714
rect 19458 2662 19516 2714
rect 19404 2660 19516 2662
rect 19404 2650 19460 2660
rect 19012 2604 19068 2614
rect 19012 2510 19068 2548
rect 18620 2100 18732 2156
rect 19124 2156 19180 2166
rect 17948 1990 17950 2042
rect 18002 1990 18004 2042
rect 17948 1978 18004 1990
rect 18340 2044 18396 2054
rect 18340 1986 18396 1988
rect 18340 1934 18342 1986
rect 18394 1934 18396 1986
rect 18564 1998 18620 2100
rect 18564 1946 18566 1998
rect 18618 1946 18620 1998
rect 18564 1934 18620 1946
rect 19012 2044 19068 2054
rect 18340 1922 18396 1934
rect 18284 1820 18340 1830
rect 18284 1818 18844 1820
rect 18284 1766 18286 1818
rect 18338 1766 18844 1818
rect 18284 1764 18844 1766
rect 18284 1754 18340 1764
rect 18452 1596 18508 1606
rect 17556 1318 17558 1370
rect 17610 1318 17612 1370
rect 17556 1306 17612 1318
rect 17780 1372 17836 1382
rect 17780 1278 17836 1316
rect 18116 1372 18172 1382
rect 17220 1162 17222 1214
rect 17274 1162 17276 1214
rect 16044 1148 16100 1158
rect 17220 1150 17276 1162
rect 18116 1214 18172 1316
rect 18452 1370 18508 1540
rect 18452 1318 18454 1370
rect 18506 1318 18508 1370
rect 18452 1306 18508 1318
rect 18116 1162 18118 1214
rect 18170 1162 18172 1214
rect 18116 1150 18172 1162
rect 18788 1214 18844 1764
rect 19012 1372 19068 1988
rect 19124 1998 19180 2100
rect 19124 1946 19126 1998
rect 19178 1946 19180 1998
rect 19124 1934 19180 1946
rect 19124 1372 19180 1382
rect 19012 1370 19180 1372
rect 19012 1318 19126 1370
rect 19178 1318 19180 1370
rect 19012 1316 19180 1318
rect 19796 1372 19852 3444
rect 20020 2828 20076 4294
rect 20132 4292 20244 4348
rect 20132 3836 20188 4292
rect 20356 4172 20412 4182
rect 20356 4078 20412 4116
rect 20132 3770 20188 3780
rect 20244 3612 20300 3622
rect 20020 2762 20076 2772
rect 20132 3610 20300 3612
rect 20132 3558 20246 3610
rect 20298 3558 20300 3610
rect 20132 3556 20300 3558
rect 19908 2716 19964 2726
rect 19908 2614 19964 2660
rect 19908 2602 20020 2614
rect 19908 2550 19966 2602
rect 20018 2550 20020 2602
rect 19908 2548 20020 2550
rect 19964 2538 20020 2548
rect 20020 1372 20076 1382
rect 19796 1370 20076 1372
rect 19796 1318 20022 1370
rect 20074 1318 20076 1370
rect 19796 1316 20076 1318
rect 18788 1162 18790 1214
rect 18842 1162 18844 1214
rect 18788 1150 18844 1162
rect 15540 1146 16100 1148
rect 15540 1094 16046 1146
rect 16098 1094 16100 1146
rect 15540 1092 16100 1094
rect 16044 1082 16100 1092
rect 19124 1148 19180 1316
rect 20020 1306 20076 1316
rect 19124 1082 19180 1092
rect 15428 1036 15484 1048
rect 19516 1036 19572 1046
rect 19740 1036 19796 1046
rect 19516 1034 19740 1036
rect 11956 970 12012 980
rect 19516 982 19518 1034
rect 19570 982 19740 1034
rect 19516 980 19740 982
rect 19516 970 19572 980
rect 19740 942 19796 980
rect 8928 812 9192 822
rect 868 634 924 644
rect 8456 0 8568 800
rect 8984 756 9032 812
rect 9088 756 9136 812
rect 8928 746 9192 756
rect 16868 812 17132 822
rect 16924 756 16972 812
rect 17028 756 17076 812
rect 16868 746 17132 756
rect 20132 586 20188 3556
rect 20244 3546 20300 3556
rect 20300 2940 20356 2950
rect 20468 2940 20524 5460
rect 21588 5404 21644 5836
rect 20580 5348 21644 5404
rect 20580 5290 20636 5348
rect 20580 5238 20582 5290
rect 20634 5238 20636 5290
rect 20580 5226 20636 5238
rect 21196 5234 21252 5246
rect 21196 5182 21198 5234
rect 21250 5182 21252 5234
rect 21196 5180 21252 5182
rect 21364 5180 21420 5190
rect 21700 5180 21756 6804
rect 22036 6748 22092 6758
rect 22036 6076 22092 6692
rect 22148 6636 22204 7354
rect 23380 7404 23382 7456
rect 23434 7404 23436 7456
rect 23044 7308 23100 7318
rect 23044 7306 23212 7308
rect 23044 7254 23046 7306
rect 23098 7254 23212 7306
rect 23044 7252 23212 7254
rect 23044 7242 23100 7252
rect 23156 6858 23212 7252
rect 23380 7196 23436 7404
rect 23380 7130 23436 7140
rect 23940 7420 23996 7430
rect 24612 7420 24668 8198
rect 25172 8204 25228 9706
rect 25732 9660 25788 9670
rect 25732 8986 25788 9604
rect 25732 8934 25734 8986
rect 25786 8934 25788 8986
rect 26068 9042 26124 10500
rect 26628 10444 26684 10724
rect 27188 10612 27244 12068
rect 27300 11676 27356 11686
rect 27300 11413 27356 11620
rect 27300 11361 27302 11413
rect 27354 11361 27356 11413
rect 27300 11349 27356 11361
rect 27412 11452 27468 11462
rect 27412 11288 27468 11396
rect 27412 11236 27414 11288
rect 27466 11236 27468 11288
rect 27412 11224 27468 11236
rect 27748 10612 27804 12740
rect 27916 12702 27972 12740
rect 28778 12572 29042 12582
rect 28834 12516 28882 12572
rect 28938 12516 28986 12572
rect 28778 12506 29042 12516
rect 29204 12178 29260 13076
rect 30436 13030 30492 13748
rect 31444 13728 31500 14310
rect 30772 13690 30828 13702
rect 30772 13638 30774 13690
rect 30826 13638 30828 13690
rect 30212 13020 30268 13030
rect 30436 13018 30548 13030
rect 30436 12966 30494 13018
rect 30546 12966 30548 13018
rect 30436 12964 30548 12966
rect 30212 12926 30268 12964
rect 30492 12954 30548 12964
rect 30772 13020 30828 13638
rect 30772 12954 30828 12964
rect 31444 13676 31446 13728
rect 31498 13676 31500 13728
rect 31444 13020 31500 13676
rect 31444 12954 31500 12964
rect 32004 14028 32060 14038
rect 29372 12908 29428 12918
rect 29372 12906 29484 12908
rect 29372 12854 29374 12906
rect 29426 12854 29484 12906
rect 29372 12842 29484 12854
rect 28644 12160 28700 12172
rect 28308 12124 28364 12134
rect 28308 12030 28364 12068
rect 28644 12124 28646 12160
rect 28698 12124 28700 12160
rect 29204 12126 29206 12178
rect 29258 12126 29260 12178
rect 29204 12114 29260 12126
rect 29428 12124 29484 12842
rect 30772 12833 30828 12845
rect 30772 12781 30774 12833
rect 30826 12781 30828 12833
rect 30772 12234 30828 12781
rect 32004 12346 32060 13972
rect 32004 12294 32006 12346
rect 32058 12294 32060 12346
rect 32004 12282 32060 12294
rect 30772 12182 30774 12234
rect 30826 12182 30828 12234
rect 30772 12170 30828 12182
rect 32340 12160 32396 12172
rect 28644 12058 28700 12068
rect 29428 12058 29484 12068
rect 30044 12124 30100 12134
rect 30044 12030 30100 12068
rect 32340 12108 32342 12160
rect 32394 12108 32396 12160
rect 31836 12012 31892 12022
rect 31836 11918 31892 11956
rect 32340 12012 32396 12108
rect 32340 11946 32396 11956
rect 32116 11900 32172 11910
rect 28778 11004 29042 11014
rect 28834 10948 28882 11004
rect 28938 10948 28986 11004
rect 28778 10938 29042 10948
rect 27188 10556 27356 10612
rect 27748 10556 27916 10612
rect 27300 10554 27356 10556
rect 27300 10502 27302 10554
rect 27354 10502 27356 10554
rect 27300 10490 27356 10502
rect 26628 10378 26684 10388
rect 27132 10444 27188 10464
rect 27748 10444 27804 10454
rect 27132 10386 27188 10388
rect 27132 10334 27134 10386
rect 27186 10334 27188 10386
rect 27132 10108 27188 10334
rect 27524 10442 27804 10444
rect 27524 10390 27750 10442
rect 27802 10390 27804 10442
rect 27524 10388 27804 10390
rect 27132 10052 27244 10108
rect 26572 9772 26628 9782
rect 26572 9678 26628 9716
rect 26964 9772 27020 9782
rect 27188 9772 27244 10052
rect 27300 9772 27356 9782
rect 27188 9770 27356 9772
rect 27188 9718 27302 9770
rect 27354 9718 27356 9770
rect 27188 9716 27356 9718
rect 26068 8990 26070 9042
rect 26122 8990 26124 9042
rect 26068 8978 26124 8990
rect 26740 9548 26796 9558
rect 25732 8922 25788 8934
rect 25452 8818 25508 8830
rect 25452 8766 25454 8818
rect 25506 8766 25508 8818
rect 25452 8540 25508 8766
rect 25396 8484 25564 8540
rect 25284 8316 25340 8326
rect 25284 8222 25340 8260
rect 25172 8138 25228 8148
rect 25396 7980 25452 8484
rect 25508 8316 25564 8484
rect 25508 8250 25564 8260
rect 26572 8316 26628 8326
rect 26572 8222 26628 8260
rect 26740 8314 26796 9492
rect 26964 9110 27020 9716
rect 27300 9548 27356 9716
rect 27300 9482 27356 9492
rect 26908 9098 27020 9110
rect 26908 9046 26910 9098
rect 26962 9046 27020 9098
rect 26908 9044 27020 9046
rect 27524 9100 27580 10388
rect 27748 10378 27804 10388
rect 27860 9996 27916 10556
rect 28084 10592 28140 10604
rect 28084 10540 28086 10592
rect 28138 10540 28140 10592
rect 28084 10444 28140 10540
rect 28084 10378 28140 10388
rect 27860 9930 27916 9940
rect 32004 9996 32060 10006
rect 27804 9772 27860 9782
rect 27804 9678 27860 9716
rect 27692 9660 27748 9670
rect 27692 9566 27748 9604
rect 28778 9436 29042 9446
rect 28834 9380 28882 9436
rect 28938 9380 28986 9436
rect 28778 9370 29042 9380
rect 32004 9210 32060 9940
rect 32004 9158 32006 9210
rect 32058 9158 32060 9210
rect 32004 9146 32060 9158
rect 27636 9100 27692 9110
rect 27524 9098 27692 9100
rect 27524 9046 27638 9098
rect 27690 9046 27692 9098
rect 27524 9044 27692 9046
rect 26908 9034 26964 9044
rect 27636 9034 27692 9044
rect 31836 8876 31892 8886
rect 31836 8782 31892 8820
rect 32116 8427 32172 11844
rect 26740 8262 26742 8314
rect 26794 8262 26796 8314
rect 26740 8250 26796 8262
rect 32004 8371 32172 8427
rect 32228 10332 32284 10342
rect 25116 7924 25452 7980
rect 26068 8204 26124 8214
rect 25116 7644 25172 7924
rect 25116 7586 25172 7588
rect 25116 7534 25118 7586
rect 25170 7534 25172 7586
rect 25116 7512 25172 7534
rect 25788 7586 25844 7598
rect 25788 7534 25790 7586
rect 25842 7534 25844 7586
rect 25788 7532 25844 7534
rect 23940 7418 24668 7420
rect 23940 7366 23942 7418
rect 23994 7366 24668 7418
rect 23940 7364 24668 7366
rect 25396 7476 25844 7532
rect 26068 7542 26124 8148
rect 28778 7868 29042 7878
rect 28834 7812 28882 7868
rect 28938 7812 28986 7868
rect 28778 7802 29042 7812
rect 26068 7532 26180 7542
rect 26068 7530 26460 7532
rect 26068 7478 26126 7530
rect 26178 7478 26460 7530
rect 26068 7476 26460 7478
rect 25396 7418 25452 7476
rect 26124 7466 26180 7476
rect 25396 7366 25398 7418
rect 25450 7366 25452 7418
rect 23156 6806 23158 6858
rect 23210 6806 23212 6858
rect 23156 6794 23212 6806
rect 22820 6748 22876 6758
rect 22148 6570 22204 6580
rect 22596 6636 22652 6646
rect 21196 5124 21308 5180
rect 21252 4956 21308 5124
rect 21364 5086 21420 5124
rect 21588 5124 21756 5180
rect 21812 6074 22092 6076
rect 21812 6022 22038 6074
rect 22090 6022 22092 6074
rect 21812 6020 22092 6022
rect 21588 4956 21644 5124
rect 21812 4966 21868 6020
rect 22036 6010 22092 6020
rect 21252 4900 21644 4956
rect 20838 4732 21102 4742
rect 20894 4676 20942 4732
rect 20998 4676 21046 4732
rect 20838 4666 21102 4676
rect 21196 4620 21252 4630
rect 20580 4508 20636 4518
rect 20580 4172 20636 4452
rect 20692 4396 20748 4406
rect 20692 4298 20694 4340
rect 20746 4298 20748 4340
rect 21196 4396 21252 4564
rect 21588 4506 21644 4900
rect 21756 4954 21868 4966
rect 21756 4902 21758 4954
rect 21810 4902 21868 4954
rect 21756 4900 21868 4902
rect 22092 4954 22148 4966
rect 22092 4902 22094 4954
rect 22146 4902 22148 4954
rect 21756 4890 21812 4900
rect 22092 4844 22148 4902
rect 22092 4778 22148 4788
rect 21588 4454 21590 4506
rect 21642 4454 21644 4506
rect 21588 4442 21644 4454
rect 21196 4394 21308 4396
rect 21196 4342 21198 4394
rect 21250 4342 21308 4394
rect 21196 4330 21308 4342
rect 20692 4286 20748 4298
rect 20580 4116 20748 4172
rect 20300 2938 20524 2940
rect 20300 2886 20302 2938
rect 20354 2886 20524 2938
rect 20300 2884 20524 2886
rect 20300 2874 20356 2884
rect 20580 2828 20636 2838
rect 20580 2726 20582 2772
rect 20634 2726 20636 2772
rect 20580 2714 20636 2726
rect 20412 2604 20468 2614
rect 20412 2602 20524 2604
rect 20412 2550 20414 2602
rect 20466 2550 20524 2602
rect 20412 2538 20524 2550
rect 20356 2380 20412 2390
rect 20356 1146 20412 2324
rect 20468 2044 20524 2538
rect 20692 2380 20748 4116
rect 21252 3566 21308 4330
rect 22260 4172 22316 4182
rect 22260 4078 22316 4116
rect 21252 3514 21254 3566
rect 21306 3514 21308 3566
rect 20916 3500 20972 3510
rect 20916 3406 20972 3444
rect 20838 3164 21102 3174
rect 20894 3108 20942 3164
rect 20998 3108 21046 3164
rect 20838 3098 21102 3108
rect 21252 2782 21308 3514
rect 21756 3554 21812 3566
rect 21756 3502 21758 3554
rect 21810 3502 21812 3554
rect 21756 3500 21812 3502
rect 21756 3444 22204 3500
rect 21252 2730 21254 2782
rect 21306 2730 21308 2782
rect 21252 2604 21308 2730
rect 21812 3276 21868 3286
rect 21812 2782 21868 3220
rect 21812 2730 21814 2782
rect 21866 2730 21868 2782
rect 21812 2718 21868 2730
rect 21252 2538 21308 2548
rect 20692 2314 20748 2324
rect 20468 1988 21420 2044
rect 20838 1596 21102 1606
rect 20894 1540 20942 1596
rect 20998 1540 21046 1596
rect 20838 1530 21102 1540
rect 21364 1214 21420 1988
rect 21476 2042 21532 2054
rect 21476 1990 21478 2042
rect 21530 1990 21532 2042
rect 21476 1708 21532 1990
rect 22148 1930 22204 3444
rect 22596 2044 22652 6580
rect 22708 6524 22764 6534
rect 22708 5850 22764 6468
rect 22708 5798 22710 5850
rect 22762 5798 22764 5850
rect 22708 5786 22764 5798
rect 22820 5238 22876 6692
rect 23828 6636 23884 6646
rect 23828 6522 23884 6580
rect 23828 6470 23830 6522
rect 23882 6470 23884 6522
rect 22820 5186 22822 5238
rect 22874 5186 22876 5238
rect 23436 5292 23492 5302
rect 22820 5174 22876 5186
rect 23044 5180 23100 5190
rect 23044 5086 23100 5124
rect 23436 5010 23492 5236
rect 23828 5292 23884 6470
rect 23940 6300 23996 7364
rect 25396 7354 25452 7366
rect 25396 7196 25452 7206
rect 24808 7084 25072 7094
rect 24864 7028 24912 7084
rect 24968 7028 25016 7084
rect 24808 7018 25072 7028
rect 24332 6860 24388 6870
rect 24332 6766 24388 6804
rect 24108 6748 24164 6758
rect 24108 6654 24164 6692
rect 24556 6690 24612 6702
rect 24556 6638 24558 6690
rect 24610 6638 24612 6690
rect 25284 6690 25340 6702
rect 24556 6636 24612 6638
rect 24556 6570 24612 6580
rect 24724 6670 24780 6682
rect 24724 6618 24726 6670
rect 24778 6618 24780 6670
rect 23940 5852 23996 6244
rect 23940 5786 23996 5796
rect 24052 6522 24108 6534
rect 24052 6470 24054 6522
rect 24106 6470 24108 6522
rect 24052 5628 24108 6470
rect 24724 5740 24780 6618
rect 25284 6638 25286 6690
rect 25338 6638 25340 6690
rect 25284 6412 25340 6638
rect 25396 6584 25452 7140
rect 26292 6682 26348 6694
rect 25396 6532 25398 6584
rect 25450 6532 25452 6584
rect 26180 6636 26236 6646
rect 25396 6520 25452 6532
rect 25676 6522 25732 6534
rect 26012 6524 26068 6534
rect 25284 6346 25340 6356
rect 25676 6470 25678 6522
rect 25730 6470 25732 6522
rect 25676 6300 25732 6470
rect 25956 6522 26068 6524
rect 25956 6470 26014 6522
rect 26066 6470 26068 6522
rect 26180 6532 26182 6580
rect 26234 6532 26236 6580
rect 26180 6520 26236 6532
rect 26292 6630 26294 6682
rect 26346 6630 26348 6682
rect 25956 6458 26068 6470
rect 25956 6300 26012 6458
rect 26292 6412 26348 6630
rect 26292 6346 26348 6356
rect 25732 6244 26012 6300
rect 25676 6234 25732 6244
rect 25060 5894 25116 5906
rect 25060 5852 25062 5894
rect 25114 5852 25116 5894
rect 25060 5786 25116 5796
rect 25508 5894 25564 5906
rect 25508 5842 25510 5894
rect 25562 5842 25564 5894
rect 24052 5562 24108 5572
rect 24612 5684 24780 5740
rect 23828 5226 23884 5236
rect 24612 5180 24668 5684
rect 24808 5516 25072 5526
rect 24864 5460 24912 5516
rect 24968 5460 25016 5516
rect 24808 5450 25072 5460
rect 24724 5180 24780 5190
rect 25508 5180 25564 5842
rect 25844 5852 25900 5862
rect 25844 5758 25900 5796
rect 24612 5178 24780 5180
rect 24612 5126 24726 5178
rect 24778 5126 24780 5178
rect 24612 5124 24780 5126
rect 23436 4958 23438 5010
rect 23490 4958 23492 5010
rect 23436 4946 23492 4958
rect 23772 4954 23828 4966
rect 23772 4902 23774 4954
rect 23826 4902 23828 4954
rect 23772 4732 23828 4902
rect 24388 4956 24444 4966
rect 24388 4862 24444 4900
rect 24612 4956 24668 4966
rect 23772 4666 23828 4676
rect 24612 4350 24668 4900
rect 24724 4508 24780 5124
rect 24724 4442 24780 4452
rect 25172 5124 25564 5180
rect 25956 5190 26012 6244
rect 26068 6300 26124 6310
rect 26068 5404 26124 6244
rect 26404 5974 26460 7476
rect 26964 6678 27020 6690
rect 26964 6636 26966 6678
rect 27018 6636 27020 6678
rect 26964 6570 27020 6580
rect 26628 6524 26684 6534
rect 26628 6430 26684 6468
rect 28778 6300 29042 6310
rect 28834 6244 28882 6300
rect 28938 6244 28986 6300
rect 28778 6234 29042 6244
rect 26404 5962 26516 5974
rect 26404 5910 26462 5962
rect 26514 5910 26516 5962
rect 26404 5908 26516 5910
rect 26460 5898 26516 5908
rect 26236 5740 26292 5750
rect 26236 5738 26348 5740
rect 26236 5686 26238 5738
rect 26290 5686 26348 5738
rect 26236 5674 26348 5686
rect 26292 5404 26348 5674
rect 26068 5348 26236 5404
rect 26292 5348 26460 5404
rect 26180 5190 26236 5348
rect 25956 5178 26068 5190
rect 25956 5126 26014 5178
rect 26066 5126 26068 5178
rect 25956 5124 26068 5126
rect 26180 5178 26292 5190
rect 26180 5126 26238 5178
rect 26290 5126 26292 5178
rect 26180 5124 26292 5126
rect 24612 4298 24614 4350
rect 24666 4298 24668 4350
rect 24612 4286 24668 4298
rect 25172 4326 25228 5124
rect 25620 5110 25676 5122
rect 26012 5114 26068 5124
rect 26236 5114 26292 5124
rect 25620 5058 25622 5110
rect 25674 5058 25676 5110
rect 25284 4956 25340 4966
rect 25284 4862 25340 4900
rect 25620 4844 25676 5058
rect 25620 4778 25676 4788
rect 26180 5004 26236 5016
rect 26180 4952 26182 5004
rect 26234 4952 26236 5004
rect 25172 4274 25174 4326
rect 25226 4274 25228 4326
rect 25172 4060 25228 4274
rect 25508 4508 25564 4518
rect 25396 4172 25452 4182
rect 25396 4078 25452 4116
rect 24808 3948 25072 3958
rect 24864 3892 24912 3948
rect 24968 3892 25016 3948
rect 24808 3882 25072 3892
rect 24052 3612 24108 3622
rect 23492 3610 24108 3612
rect 23492 3558 24054 3610
rect 24106 3558 24108 3610
rect 23492 3556 24108 3558
rect 23268 2268 23324 2278
rect 23268 2166 23324 2212
rect 23212 2154 23324 2166
rect 23212 2102 23214 2154
rect 23266 2102 23324 2154
rect 23212 2100 23324 2102
rect 23212 2090 23268 2100
rect 22764 2044 22820 2054
rect 23100 2044 23156 2054
rect 22596 2042 23100 2044
rect 22372 1986 22428 2008
rect 22372 1934 22374 1986
rect 22426 1934 22428 1986
rect 22372 1932 22428 1934
rect 22148 1878 22150 1930
rect 22202 1878 22204 1930
rect 22148 1866 22204 1878
rect 22260 1876 22372 1932
rect 22596 1990 22766 2042
rect 22818 1990 23100 2042
rect 22596 1988 23100 1990
rect 22260 1708 22316 1876
rect 22372 1866 22428 1876
rect 22484 1868 22540 1880
rect 22484 1816 22486 1868
rect 22538 1816 22540 1868
rect 21476 1642 21532 1652
rect 22036 1652 22316 1708
rect 22372 1708 22428 1718
rect 21756 1484 21812 1494
rect 21756 1370 21812 1428
rect 21756 1318 21758 1370
rect 21810 1318 21812 1370
rect 21756 1306 21812 1318
rect 21924 1308 21980 1320
rect 21364 1162 21366 1214
rect 21418 1162 21420 1214
rect 21924 1260 21926 1308
rect 21978 1260 21980 1308
rect 21924 1194 21980 1204
rect 22036 1194 22092 1652
rect 22372 1370 22428 1652
rect 22372 1318 22374 1370
rect 22426 1318 22428 1370
rect 22372 1306 22428 1318
rect 22484 1372 22540 1816
rect 22596 1484 22652 1988
rect 22764 1978 22820 1988
rect 23100 1912 23156 1988
rect 23380 1978 23436 1990
rect 23380 1932 23382 1978
rect 23434 1932 23436 1978
rect 23380 1866 23436 1876
rect 23268 1708 23324 1718
rect 23268 1484 23324 1652
rect 22596 1418 22652 1428
rect 23156 1428 23324 1484
rect 22484 1306 22540 1316
rect 21364 1150 21420 1162
rect 20356 1094 20358 1146
rect 20410 1094 20412 1146
rect 20356 1082 20412 1094
rect 22036 1148 22038 1194
rect 22090 1148 22092 1194
rect 22708 1260 22764 1270
rect 22708 1162 22710 1204
rect 22762 1162 22764 1204
rect 22708 1150 22764 1162
rect 23156 1214 23212 1428
rect 23492 1370 23548 3556
rect 24052 3546 24108 3556
rect 24724 3388 24780 3398
rect 24724 3294 24780 3332
rect 24836 2940 24892 2950
rect 24836 2846 24892 2884
rect 24164 2604 24220 2614
rect 24164 2510 24220 2548
rect 25060 2604 25116 2642
rect 25060 2538 25116 2548
rect 24332 2492 24388 2502
rect 24332 2154 24388 2436
rect 25172 2492 25228 4004
rect 25508 3747 25564 4452
rect 26180 4396 26236 4952
rect 26404 4732 26460 5348
rect 31836 5068 31892 5078
rect 31836 5066 31948 5068
rect 31836 5014 31838 5066
rect 31890 5014 31948 5066
rect 31836 5002 31948 5014
rect 31892 4956 31948 5002
rect 31892 4890 31948 4900
rect 32004 4954 32060 8371
rect 32004 4902 32006 4954
rect 32058 4902 32060 4954
rect 32004 4890 32060 4902
rect 26404 4666 26460 4676
rect 28778 4732 29042 4742
rect 28834 4676 28882 4732
rect 28938 4676 28986 4732
rect 28778 4666 29042 4676
rect 25844 4340 26236 4396
rect 25844 4294 25900 4340
rect 25788 4282 25900 4294
rect 25788 4230 25790 4282
rect 25842 4230 25900 4282
rect 25788 4228 25900 4230
rect 25788 4218 25844 4228
rect 26012 4170 26068 4182
rect 26012 4118 26014 4170
rect 26066 4118 26068 4170
rect 26012 4060 26068 4118
rect 26012 3994 26068 4004
rect 25508 3695 25510 3747
rect 25562 3695 25564 3747
rect 25508 3683 25564 3695
rect 25844 3554 25900 3566
rect 25620 3498 25676 3510
rect 25620 3446 25622 3498
rect 25674 3446 25676 3498
rect 25620 2940 25676 3446
rect 25844 3502 25846 3554
rect 25898 3502 25900 3554
rect 25844 3388 25900 3502
rect 25844 3322 25900 3332
rect 28778 3164 29042 3174
rect 28834 3108 28882 3164
rect 28938 3108 28986 3164
rect 28778 3098 29042 3108
rect 25620 2874 25676 2884
rect 25172 2426 25228 2436
rect 25396 2752 25452 2764
rect 25396 2700 25398 2752
rect 25450 2700 25452 2752
rect 24808 2380 25072 2390
rect 24864 2324 24912 2380
rect 24968 2324 25016 2380
rect 24808 2314 25072 2324
rect 25396 2268 25452 2700
rect 25676 2604 25732 2614
rect 25900 2604 25956 2614
rect 25676 2602 25956 2604
rect 25676 2550 25678 2602
rect 25730 2550 25902 2602
rect 25954 2550 25956 2602
rect 25676 2548 25956 2550
rect 25676 2492 25732 2548
rect 25900 2538 25956 2548
rect 25676 2426 25732 2436
rect 25396 2202 25452 2212
rect 24332 2102 24334 2154
rect 24386 2102 24388 2154
rect 24332 2090 24388 2102
rect 25620 2156 25676 2166
rect 23772 2044 23828 2054
rect 23772 1950 23828 1988
rect 24052 1978 24108 1990
rect 24052 1932 24054 1978
rect 24106 1932 24108 1978
rect 23940 1868 23996 1880
rect 23940 1816 23942 1868
rect 23994 1816 23996 1868
rect 24052 1866 24108 1876
rect 23940 1708 23996 1816
rect 23940 1642 23996 1652
rect 23492 1318 23494 1370
rect 23546 1318 23548 1370
rect 23492 1306 23548 1318
rect 25620 1370 25676 2100
rect 32004 2156 32060 2166
rect 32228 2156 32284 10276
rect 32340 9024 32396 9036
rect 32340 8972 32342 9024
rect 32394 8972 32396 9024
rect 32340 8876 32396 8972
rect 32340 8427 32396 8820
rect 32340 8371 32508 8427
rect 32452 8316 32508 8371
rect 32452 8250 32508 8260
rect 32340 5110 32396 5122
rect 32340 5058 32342 5110
rect 32394 5058 32396 5110
rect 32340 4956 32396 5058
rect 32340 4890 32396 4900
rect 32004 2154 32284 2156
rect 32004 2102 32006 2154
rect 32058 2102 32284 2154
rect 32004 2100 32284 2102
rect 32004 2090 32060 2100
rect 32340 1974 32396 1986
rect 31836 1930 31892 1942
rect 31836 1878 31838 1930
rect 31890 1878 31892 1930
rect 31836 1708 31892 1878
rect 31836 1642 31892 1652
rect 32340 1922 32342 1974
rect 32394 1922 32396 1974
rect 32340 1708 32396 1922
rect 32340 1642 32396 1652
rect 28778 1596 29042 1606
rect 28834 1540 28882 1596
rect 28938 1540 28986 1596
rect 28778 1530 29042 1540
rect 25620 1318 25622 1370
rect 25674 1318 25676 1370
rect 25620 1306 25676 1318
rect 23156 1162 23158 1214
rect 23210 1162 23212 1214
rect 23156 1150 23212 1162
rect 25956 1184 26012 1196
rect 22036 1082 22092 1092
rect 25956 1132 25958 1184
rect 26010 1132 26012 1184
rect 20132 534 20134 586
rect 20186 534 20188 586
rect 20132 522 20188 534
rect 21028 1034 21084 1046
rect 21028 982 21030 1034
rect 21082 982 21084 1034
rect 21028 586 21084 982
rect 25508 1036 25564 1046
rect 24808 812 25072 822
rect 24864 756 24912 812
rect 24968 756 25016 812
rect 25508 800 25564 980
rect 25956 1036 26012 1132
rect 25956 970 26012 980
rect 26236 1036 26292 1046
rect 26236 942 26292 980
rect 24808 746 25072 756
rect 21028 534 21030 586
rect 21082 534 21084 586
rect 21028 522 21084 534
rect 25480 0 25592 800
<< via2 >>
rect 1204 18452 1260 18508
rect 1428 19012 1484 19068
rect 1876 18618 1932 18620
rect 1876 18566 1878 18618
rect 1878 18566 1930 18618
rect 1930 18566 1932 18618
rect 1876 18564 1932 18566
rect 1540 18462 1596 18508
rect 1540 18452 1542 18462
rect 1542 18452 1594 18462
rect 1594 18452 1596 18462
rect 3388 18506 3444 18508
rect 3388 18454 3390 18506
rect 3390 18454 3442 18506
rect 3442 18454 3444 18506
rect 3388 18452 3444 18454
rect 1428 18340 1484 18396
rect 2940 18394 2996 18396
rect 2940 18342 2942 18394
rect 2942 18342 2994 18394
rect 2994 18342 2996 18394
rect 2940 18340 2996 18342
rect 4958 18842 5014 18844
rect 4958 18790 4960 18842
rect 4960 18790 5012 18842
rect 5012 18790 5014 18842
rect 4958 18788 5014 18790
rect 5062 18842 5118 18844
rect 5062 18790 5064 18842
rect 5064 18790 5116 18842
rect 5116 18790 5118 18842
rect 5062 18788 5118 18790
rect 5166 18842 5222 18844
rect 5166 18790 5168 18842
rect 5168 18790 5220 18842
rect 5220 18790 5222 18842
rect 5166 18788 5222 18790
rect 3892 18340 3948 18396
rect 4508 18394 4564 18396
rect 4508 18342 4510 18394
rect 4510 18342 4562 18394
rect 4562 18342 4564 18394
rect 4508 18340 4564 18342
rect 1652 18228 1708 18284
rect 2716 18282 2772 18284
rect 2716 18230 2718 18282
rect 2718 18230 2770 18282
rect 2770 18230 2772 18282
rect 2716 18228 2772 18230
rect 4340 18282 4396 18284
rect 2548 18116 2604 18172
rect 2100 18004 2156 18060
rect 4340 18230 4342 18282
rect 4342 18230 4394 18282
rect 4394 18230 4396 18282
rect 4340 18228 4396 18230
rect 6300 18282 6356 18284
rect 6300 18230 6302 18282
rect 6302 18230 6354 18282
rect 6354 18230 6356 18282
rect 6300 18228 6356 18230
rect 3164 18004 3220 18060
rect 2660 17780 2716 17836
rect 3724 17780 3780 17836
rect 1540 16894 1596 16940
rect 1540 16884 1542 16894
rect 1542 16884 1594 16894
rect 1594 16884 1596 16894
rect 1876 17498 1932 17500
rect 1876 17446 1878 17498
rect 1878 17446 1930 17498
rect 1930 17446 1932 17498
rect 1876 17444 1932 17446
rect 2548 17610 2604 17612
rect 2548 17558 2550 17610
rect 2550 17558 2602 17610
rect 2602 17558 2604 17610
rect 2548 17556 2604 17558
rect 3724 17610 3780 17612
rect 3724 17558 3726 17610
rect 3726 17558 3778 17610
rect 3778 17558 3780 17610
rect 3724 17556 3780 17558
rect 5852 17834 5908 17836
rect 5852 17782 5854 17834
rect 5854 17782 5906 17834
rect 5906 17782 5908 17834
rect 5852 17780 5908 17782
rect 3388 17498 3444 17500
rect 3388 17446 3390 17498
rect 3390 17446 3442 17498
rect 3442 17446 3444 17498
rect 3388 17444 3444 17446
rect 4958 17274 5014 17276
rect 4958 17222 4960 17274
rect 4960 17222 5012 17274
rect 5012 17222 5014 17274
rect 4958 17220 5014 17222
rect 5062 17274 5118 17276
rect 5062 17222 5064 17274
rect 5064 17222 5116 17274
rect 5116 17222 5118 17274
rect 5062 17220 5118 17222
rect 5166 17274 5222 17276
rect 5166 17222 5168 17274
rect 5168 17222 5220 17274
rect 5220 17222 5222 17274
rect 5166 17220 5222 17222
rect 3500 16996 3556 17052
rect 7140 17780 7196 17836
rect 6804 17722 6860 17724
rect 6804 17670 6806 17722
rect 6806 17670 6858 17722
rect 6858 17670 6860 17722
rect 6804 17668 6860 17670
rect 6412 17610 6468 17612
rect 6412 17558 6414 17610
rect 6414 17558 6466 17610
rect 6466 17558 6468 17610
rect 6412 17556 6468 17558
rect 5964 17498 6020 17500
rect 5964 17446 5966 17498
rect 5966 17446 6018 17498
rect 6018 17446 6020 17498
rect 5964 17444 6020 17446
rect 6300 17220 6356 17276
rect 6692 17444 6748 17500
rect 6356 16996 6412 17052
rect 1428 16660 1484 16716
rect 2044 16714 2100 16716
rect 2044 16662 2046 16714
rect 2046 16662 2098 16714
rect 2098 16662 2100 16714
rect 2044 16660 2100 16662
rect 6916 17220 6972 17276
rect 3164 16714 3220 16716
rect 3164 16662 3166 16714
rect 3166 16662 3218 16714
rect 3218 16662 3220 16714
rect 3164 16660 3220 16662
rect 3724 16660 3780 16716
rect 2548 16117 2604 16156
rect 2548 16100 2550 16117
rect 2550 16100 2602 16117
rect 2602 16100 2604 16117
rect 1540 15540 1596 15596
rect 1204 14308 1260 14364
rect 1204 13412 1260 13468
rect 1596 13636 1652 13692
rect 1316 13076 1372 13132
rect 1316 12180 1372 12236
rect 2268 15764 2324 15820
rect 2884 15370 2940 15372
rect 2884 15318 2886 15370
rect 2886 15318 2938 15370
rect 2938 15318 2940 15370
rect 2884 15316 2940 15318
rect 2100 15092 2156 15148
rect 2884 14868 2940 14924
rect 3220 15316 3276 15372
rect 3108 15204 3164 15260
rect 1876 13748 1932 13804
rect 1764 13188 1820 13244
rect 1708 12906 1764 12908
rect 1708 12854 1710 12906
rect 1710 12854 1762 12906
rect 1762 12854 1764 12906
rect 1708 12852 1764 12854
rect 2324 13524 2380 13580
rect 1876 12404 1932 12460
rect 1596 12234 1652 12236
rect 1596 12182 1598 12234
rect 1598 12182 1650 12234
rect 1650 12182 1652 12234
rect 1596 12180 1652 12182
rect 2436 13018 2492 13020
rect 2436 12966 2438 13018
rect 2438 12966 2490 13018
rect 2490 12966 2492 13018
rect 2436 12964 2492 12966
rect 2660 12852 2716 12908
rect 2324 12234 2380 12236
rect 2324 12182 2326 12234
rect 2326 12182 2378 12234
rect 2378 12182 2380 12234
rect 2324 12180 2380 12182
rect 1876 11956 1932 12012
rect 1372 11844 1428 11900
rect 2212 11620 2268 11676
rect 2660 11620 2716 11676
rect 2324 11508 2380 11564
rect 4900 16660 4956 16716
rect 6636 16266 6692 16268
rect 6636 16214 6638 16266
rect 6638 16214 6690 16266
rect 6690 16214 6692 16266
rect 6636 16212 6692 16214
rect 4958 15706 5014 15708
rect 4958 15654 4960 15706
rect 4960 15654 5012 15706
rect 5012 15654 5014 15706
rect 4958 15652 5014 15654
rect 5062 15706 5118 15708
rect 5062 15654 5064 15706
rect 5064 15654 5116 15706
rect 5116 15654 5118 15706
rect 5062 15652 5118 15654
rect 5166 15706 5222 15708
rect 5166 15654 5168 15706
rect 5168 15654 5220 15706
rect 5220 15654 5222 15706
rect 5166 15652 5222 15654
rect 6468 15482 6524 15484
rect 6468 15430 6470 15482
rect 6470 15430 6522 15482
rect 6522 15430 6524 15482
rect 6468 15428 6524 15430
rect 5516 15370 5572 15372
rect 5516 15318 5518 15370
rect 5518 15318 5570 15370
rect 5570 15318 5572 15370
rect 5516 15316 5572 15318
rect 7252 17556 7308 17612
rect 11172 18676 11228 18732
rect 9996 18564 10052 18620
rect 10164 18506 10220 18508
rect 10164 18454 10166 18506
rect 10166 18454 10218 18506
rect 10218 18454 10220 18506
rect 10164 18452 10220 18454
rect 9044 18228 9100 18284
rect 9268 18228 9324 18284
rect 8928 18058 8984 18060
rect 8928 18006 8930 18058
rect 8930 18006 8982 18058
rect 8982 18006 8984 18058
rect 8928 18004 8984 18006
rect 9032 18058 9088 18060
rect 9032 18006 9034 18058
rect 9034 18006 9086 18058
rect 9086 18006 9088 18058
rect 9032 18004 9088 18006
rect 9136 18058 9192 18060
rect 9136 18006 9138 18058
rect 9138 18006 9190 18058
rect 9190 18006 9192 18058
rect 9136 18004 9192 18006
rect 8708 17780 8764 17836
rect 7924 17668 7980 17724
rect 9492 17685 9548 17724
rect 9492 17668 9494 17685
rect 9494 17668 9546 17685
rect 9546 17668 9548 17685
rect 8092 17108 8148 17164
rect 8372 17556 8428 17612
rect 8932 17610 8988 17612
rect 8932 17558 8934 17610
rect 8934 17558 8986 17610
rect 8986 17558 8988 17610
rect 8932 17556 8988 17558
rect 8596 17220 8652 17276
rect 9436 17108 9492 17164
rect 8928 16490 8984 16492
rect 8928 16438 8930 16490
rect 8930 16438 8982 16490
rect 8982 16438 8984 16490
rect 8928 16436 8984 16438
rect 9032 16490 9088 16492
rect 9032 16438 9034 16490
rect 9034 16438 9086 16490
rect 9086 16438 9088 16490
rect 9032 16436 9088 16438
rect 9136 16490 9192 16492
rect 9136 16438 9138 16490
rect 9138 16438 9190 16490
rect 9190 16438 9192 16490
rect 9136 16436 9192 16438
rect 8876 16154 8932 16156
rect 8876 16102 8878 16154
rect 8878 16102 8930 16154
rect 8930 16102 8932 16154
rect 8876 16100 8932 16102
rect 7364 15652 7420 15708
rect 7140 15540 7196 15596
rect 4060 15258 4116 15260
rect 4060 15206 4062 15258
rect 4062 15206 4114 15258
rect 4114 15206 4116 15258
rect 4060 15204 4116 15206
rect 6132 15244 6134 15260
rect 6134 15244 6186 15260
rect 6186 15244 6188 15260
rect 6916 15316 6972 15372
rect 6132 15204 6188 15244
rect 5404 15146 5460 15148
rect 5404 15094 5406 15146
rect 5406 15094 5458 15146
rect 5458 15094 5460 15146
rect 5404 15092 5460 15094
rect 7532 15258 7588 15260
rect 7532 15206 7534 15258
rect 7534 15206 7586 15258
rect 7586 15206 7588 15258
rect 7532 15204 7588 15206
rect 8876 15876 8932 15932
rect 8708 15428 8764 15484
rect 8596 15316 8652 15372
rect 7924 15204 7980 15260
rect 8092 15092 8148 15148
rect 3500 14308 3556 14364
rect 2996 13636 3052 13692
rect 4004 13524 4060 13580
rect 3164 12740 3220 12796
rect 5012 14308 5068 14364
rect 5516 14196 5572 14252
rect 4958 14138 5014 14140
rect 4958 14086 4960 14138
rect 4960 14086 5012 14138
rect 5012 14086 5014 14138
rect 4958 14084 5014 14086
rect 5062 14138 5118 14140
rect 5062 14086 5064 14138
rect 5064 14086 5116 14138
rect 5116 14086 5118 14138
rect 5062 14084 5118 14086
rect 5166 14138 5222 14140
rect 5166 14086 5168 14138
rect 5168 14086 5220 14138
rect 5220 14086 5222 14138
rect 5166 14084 5222 14086
rect 6244 14196 6300 14252
rect 5852 13690 5908 13692
rect 5852 13638 5854 13690
rect 5854 13638 5906 13690
rect 5906 13638 5908 13690
rect 5852 13636 5908 13638
rect 4620 13412 4676 13468
rect 5404 13578 5460 13580
rect 5404 13526 5406 13578
rect 5406 13526 5458 13578
rect 5458 13526 5460 13578
rect 5404 13524 5460 13526
rect 5964 13578 6020 13580
rect 5964 13526 5966 13578
rect 5966 13526 6018 13578
rect 6018 13526 6020 13578
rect 5964 13524 6020 13526
rect 4564 13018 4620 13020
rect 4564 12966 4566 13018
rect 4566 12966 4618 13018
rect 4618 12966 4620 13018
rect 4564 12964 4620 12966
rect 4116 12740 4172 12796
rect 4228 12234 4284 12236
rect 4228 12182 4230 12234
rect 4230 12182 4282 12234
rect 4282 12182 4284 12234
rect 4228 12180 4284 12182
rect 3276 11562 3332 11564
rect 3276 11510 3278 11562
rect 3278 11510 3330 11562
rect 3330 11510 3332 11562
rect 3276 11508 3332 11510
rect 6356 13860 6412 13916
rect 8260 14308 8316 14364
rect 8596 14868 8652 14924
rect 8036 14084 8092 14140
rect 7476 13972 7532 14028
rect 6916 13758 6972 13804
rect 6916 13748 6918 13758
rect 6918 13748 6970 13758
rect 6970 13748 6972 13758
rect 7252 13682 7254 13692
rect 7254 13682 7306 13692
rect 7306 13682 7308 13692
rect 7252 13636 7308 13682
rect 7140 13524 7196 13580
rect 6860 13188 6916 13244
rect 6636 13130 6692 13132
rect 6636 13078 6638 13130
rect 6638 13078 6690 13130
rect 6690 13078 6692 13130
rect 6636 13076 6692 13078
rect 7028 13076 7084 13132
rect 7588 13130 7644 13132
rect 7588 13078 7590 13130
rect 7590 13078 7642 13130
rect 7642 13078 7644 13130
rect 7588 13076 7644 13078
rect 5404 12740 5460 12796
rect 4958 12570 5014 12572
rect 4958 12518 4960 12570
rect 4960 12518 5012 12570
rect 5012 12518 5014 12570
rect 4958 12516 5014 12518
rect 5062 12570 5118 12572
rect 5062 12518 5064 12570
rect 5064 12518 5116 12570
rect 5116 12518 5118 12570
rect 5062 12516 5118 12518
rect 5166 12570 5222 12572
rect 5166 12518 5168 12570
rect 5168 12518 5220 12570
rect 5220 12518 5222 12570
rect 5166 12516 5222 12518
rect 6468 12404 6524 12460
rect 6244 12292 6300 12348
rect 5852 12234 5908 12236
rect 5852 12182 5854 12234
rect 5854 12182 5906 12234
rect 5906 12182 5908 12234
rect 5852 12180 5908 12182
rect 7196 12346 7252 12348
rect 7196 12294 7198 12346
rect 7198 12294 7250 12346
rect 7250 12294 7252 12346
rect 7196 12292 7252 12294
rect 5516 12010 5572 12012
rect 5516 11958 5518 12010
rect 5518 11958 5570 12010
rect 5570 11958 5572 12010
rect 5516 11956 5572 11958
rect 7084 12010 7140 12012
rect 7084 11958 7086 12010
rect 7086 11958 7138 12010
rect 7138 11958 7140 12010
rect 7084 11956 7140 11958
rect 4676 11620 4732 11676
rect 8148 13914 8204 13916
rect 8148 13862 8150 13914
rect 8150 13862 8202 13914
rect 8202 13862 8204 13914
rect 8148 13860 8204 13862
rect 8428 13748 8484 13804
rect 8204 13690 8260 13692
rect 8204 13638 8206 13690
rect 8206 13638 8258 13690
rect 8258 13638 8260 13690
rect 9436 15146 9492 15148
rect 9436 15094 9438 15146
rect 9438 15094 9490 15146
rect 9490 15094 9492 15146
rect 9436 15092 9492 15094
rect 8928 14922 8984 14924
rect 8928 14870 8930 14922
rect 8930 14870 8982 14922
rect 8982 14870 8984 14922
rect 8928 14868 8984 14870
rect 9032 14922 9088 14924
rect 9032 14870 9034 14922
rect 9034 14870 9086 14922
rect 9086 14870 9088 14922
rect 9032 14868 9088 14870
rect 9136 14922 9192 14924
rect 9136 14870 9138 14922
rect 9138 14870 9190 14922
rect 9190 14870 9192 14922
rect 9136 14868 9192 14870
rect 10164 18228 10220 18284
rect 11340 18564 11396 18620
rect 12898 18842 12954 18844
rect 12898 18790 12900 18842
rect 12900 18790 12952 18842
rect 12952 18790 12954 18842
rect 12898 18788 12954 18790
rect 13002 18842 13058 18844
rect 13002 18790 13004 18842
rect 13004 18790 13056 18842
rect 13056 18790 13058 18842
rect 13002 18788 13058 18790
rect 13106 18842 13162 18844
rect 13106 18790 13108 18842
rect 13108 18790 13160 18842
rect 13160 18790 13162 18842
rect 13106 18788 13162 18790
rect 11732 18380 11734 18396
rect 11734 18380 11786 18396
rect 11786 18380 11788 18396
rect 11732 18340 11788 18380
rect 12516 18340 12572 18396
rect 10052 17834 10108 17836
rect 10052 17782 10054 17834
rect 10054 17782 10106 17834
rect 10106 17782 10108 17834
rect 10052 17780 10108 17782
rect 9828 17332 9884 17388
rect 10388 17602 10390 17612
rect 10390 17602 10442 17612
rect 10442 17602 10444 17612
rect 10388 17556 10444 17602
rect 10612 18228 10668 18284
rect 10780 18282 10836 18284
rect 10780 18230 10782 18282
rect 10782 18230 10834 18282
rect 10834 18230 10836 18282
rect 10780 18228 10836 18230
rect 10948 18116 11004 18172
rect 11172 18116 11228 18172
rect 10612 18004 10668 18060
rect 10612 17556 10668 17612
rect 10780 17610 10836 17612
rect 10780 17558 10782 17610
rect 10782 17558 10834 17610
rect 10834 17558 10836 17610
rect 10780 17556 10836 17558
rect 11060 17444 11116 17500
rect 10108 16436 10164 16492
rect 10724 17108 10780 17164
rect 10612 16884 10668 16940
rect 11788 17834 11844 17836
rect 11788 17782 11790 17834
rect 11790 17782 11842 17834
rect 11842 17782 11844 17834
rect 11788 17780 11844 17782
rect 11508 17556 11564 17612
rect 11284 16884 11340 16940
rect 11396 16772 11452 16828
rect 11004 16266 11060 16268
rect 11004 16214 11006 16266
rect 11006 16214 11058 16266
rect 11058 16214 11060 16266
rect 11004 16212 11060 16214
rect 11172 16212 11228 16268
rect 11620 16996 11676 17052
rect 11956 16826 12012 16828
rect 11956 16774 11958 16826
rect 11958 16774 12010 16826
rect 12010 16774 12012 16826
rect 11956 16772 12012 16774
rect 11620 16660 11676 16716
rect 12404 18116 12460 18172
rect 13300 18340 13356 18396
rect 15988 18900 16044 18956
rect 15652 18676 15708 18732
rect 14196 18340 14252 18396
rect 14028 17780 14084 17836
rect 14420 18116 14476 18172
rect 15316 18340 15372 18396
rect 15092 18282 15148 18284
rect 15092 18230 15094 18282
rect 15094 18230 15146 18282
rect 15146 18230 15148 18282
rect 15092 18228 15148 18230
rect 14868 17780 14924 17836
rect 14980 17685 15036 17724
rect 14980 17668 14982 17685
rect 14982 17668 15034 17685
rect 15034 17668 15036 17685
rect 15428 17834 15484 17836
rect 15428 17782 15430 17834
rect 15430 17782 15482 17834
rect 15482 17782 15484 17834
rect 15428 17780 15484 17782
rect 12292 17050 12348 17052
rect 12292 16998 12294 17050
rect 12294 16998 12346 17050
rect 12346 16998 12348 17050
rect 12292 16996 12348 16998
rect 12404 16548 12460 16604
rect 12124 16266 12180 16268
rect 12124 16214 12126 16266
rect 12126 16214 12178 16266
rect 12178 16214 12180 16266
rect 12124 16212 12180 16214
rect 11620 16100 11676 16156
rect 11788 16154 11844 16156
rect 11788 16102 11790 16154
rect 11790 16102 11842 16154
rect 11842 16102 11844 16154
rect 11788 16100 11844 16102
rect 12572 16212 12628 16268
rect 12628 15652 12684 15708
rect 12516 15438 12572 15484
rect 12516 15428 12518 15438
rect 12518 15428 12570 15438
rect 12570 15428 12572 15438
rect 10612 15243 10614 15260
rect 10614 15243 10666 15260
rect 10666 15243 10668 15260
rect 10612 15204 10668 15243
rect 11060 15204 11116 15260
rect 9604 14756 9660 14812
rect 10052 14644 10108 14700
rect 9380 14362 9436 14364
rect 9380 14310 9382 14362
rect 9382 14310 9434 14362
rect 9434 14310 9436 14362
rect 9380 14308 9436 14310
rect 10052 14084 10108 14140
rect 10164 14420 10220 14476
rect 9828 13972 9884 14028
rect 9492 13914 9548 13916
rect 9492 13862 9494 13914
rect 9494 13862 9546 13914
rect 9546 13862 9548 13914
rect 9492 13860 9548 13862
rect 8204 13636 8260 13638
rect 8596 13636 8652 13692
rect 9940 13636 9996 13692
rect 9044 13524 9100 13580
rect 8260 13300 8316 13356
rect 8928 13354 8984 13356
rect 8928 13302 8930 13354
rect 8930 13302 8982 13354
rect 8982 13302 8984 13354
rect 8928 13300 8984 13302
rect 9032 13354 9088 13356
rect 9032 13302 9034 13354
rect 9034 13302 9086 13354
rect 9086 13302 9088 13354
rect 9032 13300 9088 13302
rect 9136 13354 9192 13356
rect 9136 13302 9138 13354
rect 9138 13302 9190 13354
rect 9190 13302 9192 13354
rect 9136 13300 9192 13302
rect 8652 13188 8708 13244
rect 8876 13130 8932 13132
rect 8876 13078 8878 13130
rect 8878 13078 8930 13130
rect 8930 13078 8932 13130
rect 8876 13076 8932 13078
rect 10108 12906 10164 12908
rect 10108 12854 10110 12906
rect 10110 12854 10162 12906
rect 10162 12854 10164 12906
rect 10108 12852 10164 12854
rect 9884 12794 9940 12796
rect 9884 12742 9886 12794
rect 9886 12742 9938 12794
rect 9938 12742 9940 12794
rect 9884 12740 9940 12742
rect 8260 12292 8316 12348
rect 7924 11956 7980 12012
rect 4564 11508 4620 11564
rect 3108 11396 3164 11452
rect 1540 9940 1596 9996
rect 1316 9268 1372 9324
rect 1540 9268 1596 9324
rect 1876 9268 1932 9324
rect 2996 10554 3052 10556
rect 2996 10502 2998 10554
rect 2998 10502 3050 10554
rect 3050 10502 3052 10554
rect 2996 10500 3052 10502
rect 4452 11413 4508 11452
rect 4452 11396 4454 11413
rect 4454 11396 4506 11413
rect 4506 11396 4508 11413
rect 6244 11396 6300 11452
rect 6804 11396 6860 11452
rect 5796 11284 5852 11340
rect 4958 11002 5014 11004
rect 4958 10950 4960 11002
rect 4960 10950 5012 11002
rect 5012 10950 5014 11002
rect 4958 10948 5014 10950
rect 5062 11002 5118 11004
rect 5062 10950 5064 11002
rect 5064 10950 5116 11002
rect 5116 10950 5118 11002
rect 5062 10948 5118 10950
rect 5166 11002 5222 11004
rect 5166 10950 5168 11002
rect 5168 10950 5220 11002
rect 5220 10950 5222 11002
rect 5166 10948 5222 10950
rect 2548 9940 2604 9996
rect 3556 10612 3612 10668
rect 4228 10666 4284 10668
rect 4228 10614 4230 10666
rect 4230 10614 4282 10666
rect 4282 10614 4284 10666
rect 4228 10612 4284 10614
rect 3444 9098 3500 9100
rect 3444 9046 3446 9098
rect 3446 9046 3498 9098
rect 3498 9046 3500 9098
rect 3444 9044 3500 9046
rect 4788 10500 4844 10556
rect 5460 10388 5516 10444
rect 4060 9994 4116 9996
rect 4060 9942 4062 9994
rect 4062 9942 4114 9994
rect 4114 9942 4116 9994
rect 4060 9940 4116 9942
rect 4564 9604 4620 9660
rect 5460 10164 5516 10220
rect 4900 10052 4956 10108
rect 5908 10052 5964 10108
rect 4788 9716 4844 9772
rect 5068 9770 5124 9772
rect 5068 9718 5070 9770
rect 5070 9718 5122 9770
rect 5122 9718 5124 9770
rect 5068 9716 5124 9718
rect 4958 9434 5014 9436
rect 4958 9382 4960 9434
rect 4960 9382 5012 9434
rect 5012 9382 5014 9434
rect 4958 9380 5014 9382
rect 5062 9434 5118 9436
rect 5062 9382 5064 9434
rect 5064 9382 5116 9434
rect 5116 9382 5118 9434
rect 5062 9380 5118 9382
rect 5166 9434 5222 9436
rect 5166 9382 5168 9434
rect 5168 9382 5220 9434
rect 5220 9382 5222 9434
rect 5166 9380 5222 9382
rect 4564 9044 4620 9100
rect 5908 9882 5964 9884
rect 5908 9830 5910 9882
rect 5910 9830 5962 9882
rect 5962 9830 5964 9882
rect 5908 9828 5964 9830
rect 7140 11620 7196 11676
rect 7252 11396 7308 11452
rect 7028 10612 7084 10668
rect 6468 9940 6524 9996
rect 7252 10052 7308 10108
rect 8036 11172 8092 11228
rect 8820 12108 8822 12124
rect 8822 12108 8874 12124
rect 8874 12108 8876 12124
rect 8820 12068 8876 12108
rect 9492 11956 9548 12012
rect 9268 11844 9324 11900
rect 8928 11786 8984 11788
rect 8928 11734 8930 11786
rect 8930 11734 8982 11786
rect 8982 11734 8984 11786
rect 8928 11732 8984 11734
rect 9032 11786 9088 11788
rect 9032 11734 9034 11786
rect 9034 11734 9086 11786
rect 9086 11734 9088 11786
rect 9032 11732 9088 11734
rect 9136 11786 9192 11788
rect 9136 11734 9138 11786
rect 9138 11734 9190 11786
rect 9190 11734 9192 11786
rect 9136 11732 9192 11734
rect 9324 11620 9380 11676
rect 10052 12068 10108 12124
rect 9716 11508 9772 11564
rect 10500 13748 10556 13804
rect 10948 14644 11004 14700
rect 10780 14420 10836 14476
rect 12068 15250 12070 15260
rect 12070 15250 12122 15260
rect 12122 15250 12124 15260
rect 12068 15204 12124 15250
rect 11396 14980 11452 15036
rect 12236 15092 12292 15148
rect 11732 14980 11788 15036
rect 11508 14868 11564 14924
rect 11172 14644 11228 14700
rect 10444 13018 10500 13020
rect 10444 12966 10446 13018
rect 10446 12966 10498 13018
rect 10498 12966 10500 13018
rect 10444 12964 10500 12966
rect 10276 12180 10332 12236
rect 10612 12068 10668 12124
rect 10500 11956 10556 12012
rect 10052 11508 10108 11564
rect 10276 11396 10332 11452
rect 8708 11284 8764 11340
rect 8148 11060 8204 11116
rect 9436 11284 9492 11340
rect 11340 14420 11396 14476
rect 11844 14756 11900 14812
rect 11732 14420 11788 14476
rect 11284 14084 11340 14140
rect 11508 14084 11564 14140
rect 11508 13748 11564 13804
rect 12628 14980 12684 15036
rect 12180 14780 12236 14812
rect 12180 14756 12182 14780
rect 12182 14756 12234 14780
rect 12234 14756 12236 14780
rect 12180 14466 12182 14476
rect 12182 14466 12234 14476
rect 12234 14466 12236 14476
rect 12180 14420 12236 14466
rect 11396 13524 11452 13580
rect 12404 14644 12460 14700
rect 12516 14420 12572 14476
rect 12124 13578 12180 13580
rect 12124 13526 12126 13578
rect 12126 13526 12178 13578
rect 12178 13526 12180 13578
rect 12124 13524 12180 13526
rect 12012 13412 12068 13468
rect 11508 13300 11564 13356
rect 11396 12964 11452 13020
rect 11956 12852 12012 12908
rect 12068 12740 12124 12796
rect 11732 12404 11788 12460
rect 11620 12068 11676 12124
rect 12292 12740 12348 12796
rect 12180 11956 12236 12012
rect 12068 11844 12124 11900
rect 11508 11620 11564 11676
rect 11844 11732 11900 11788
rect 10948 11562 11004 11564
rect 10948 11510 10950 11562
rect 10950 11510 11002 11562
rect 11002 11510 11004 11562
rect 10948 11508 11004 11510
rect 11396 11508 11452 11564
rect 10836 11396 10892 11452
rect 11060 11396 11116 11452
rect 11620 11508 11676 11564
rect 9660 11172 9716 11228
rect 9940 10948 9996 11004
rect 8260 10554 8316 10556
rect 8260 10502 8262 10554
rect 8262 10502 8314 10554
rect 8314 10502 8316 10554
rect 8260 10500 8316 10502
rect 9100 10442 9156 10444
rect 9100 10390 9102 10442
rect 9102 10390 9154 10442
rect 9154 10390 9156 10442
rect 9100 10388 9156 10390
rect 8928 10218 8984 10220
rect 8928 10166 8930 10218
rect 8930 10166 8982 10218
rect 8982 10166 8984 10218
rect 8928 10164 8984 10166
rect 9032 10218 9088 10220
rect 9032 10166 9034 10218
rect 9034 10166 9086 10218
rect 9086 10166 9088 10218
rect 9032 10164 9088 10166
rect 9136 10218 9192 10220
rect 9136 10166 9138 10218
rect 9138 10166 9190 10218
rect 9190 10166 9192 10218
rect 9136 10164 9192 10166
rect 7476 9940 7532 9996
rect 8092 10052 8148 10108
rect 1316 8036 1372 8092
rect 1204 6916 1260 6972
rect 868 2548 924 2604
rect 1484 7028 1540 7084
rect 2436 7028 2492 7084
rect 1988 6916 2044 6972
rect 2268 6916 2324 6972
rect 1652 6468 1708 6524
rect 4956 8314 5012 8316
rect 4956 8262 4958 8314
rect 4958 8262 5010 8314
rect 5010 8262 5012 8314
rect 4956 8260 5012 8262
rect 7756 9882 7812 9884
rect 7756 9830 7758 9882
rect 7758 9830 7810 9882
rect 7810 9830 7812 9882
rect 8316 9940 8372 9996
rect 7756 9828 7812 9830
rect 6468 8932 6524 8988
rect 6356 8708 6412 8764
rect 6132 8484 6188 8540
rect 5908 8260 5964 8316
rect 4340 8090 4396 8092
rect 4340 8038 4342 8090
rect 4342 8038 4394 8090
rect 4394 8038 4396 8090
rect 4340 8036 4396 8038
rect 4958 7866 5014 7868
rect 4958 7814 4960 7866
rect 4960 7814 5012 7866
rect 5012 7814 5014 7866
rect 4958 7812 5014 7814
rect 5062 7866 5118 7868
rect 5062 7814 5064 7866
rect 5064 7814 5116 7866
rect 5116 7814 5118 7866
rect 5062 7812 5118 7814
rect 5166 7866 5222 7868
rect 5166 7814 5168 7866
rect 5168 7814 5220 7866
rect 5220 7814 5222 7866
rect 5166 7812 5222 7814
rect 4452 7700 4508 7756
rect 2324 6074 2380 6076
rect 2324 6022 2326 6074
rect 2326 6022 2378 6074
rect 2378 6022 2380 6074
rect 2324 6020 2380 6022
rect 1484 5738 1540 5740
rect 1484 5686 1486 5738
rect 1486 5686 1538 5738
rect 1538 5686 1540 5738
rect 1484 5684 1540 5686
rect 1484 5460 1540 5516
rect 1988 5684 2044 5740
rect 2492 5738 2548 5740
rect 2492 5686 2494 5738
rect 2494 5686 2546 5738
rect 2546 5686 2548 5738
rect 2492 5684 2548 5686
rect 1988 5236 2044 5292
rect 2156 5348 2212 5404
rect 2548 5348 2604 5404
rect 1708 4564 1764 4620
rect 2380 4900 2436 4956
rect 2212 4676 2268 4732
rect 2100 4564 2156 4620
rect 2212 4460 2268 4508
rect 2212 4452 2214 4460
rect 2214 4452 2266 4460
rect 2266 4452 2268 4460
rect 1484 4282 1540 4284
rect 1484 4230 1486 4282
rect 1486 4230 1538 4282
rect 1538 4230 1540 4282
rect 1484 4228 1540 4230
rect 2548 4452 2604 4508
rect 1708 4116 1764 4172
rect 1540 4004 1596 4060
rect 1764 3668 1820 3724
rect 2380 3668 2436 3724
rect 2772 6020 2828 6076
rect 3220 7306 3276 7308
rect 3220 7254 3222 7306
rect 3222 7254 3274 7306
rect 3274 7254 3276 7306
rect 3220 7252 3276 7254
rect 3108 7028 3164 7084
rect 4060 7364 4116 7420
rect 4004 6692 4060 6748
rect 3444 6626 3446 6636
rect 3446 6626 3498 6636
rect 3498 6626 3500 6636
rect 3444 6580 3500 6626
rect 3724 6634 3780 6636
rect 3724 6582 3726 6634
rect 3726 6582 3778 6634
rect 3778 6582 3780 6634
rect 3724 6580 3780 6582
rect 2996 5236 3052 5292
rect 2884 5012 2940 5068
rect 3220 5236 3276 5292
rect 3444 5684 3500 5740
rect 2772 4340 2828 4396
rect 2996 4676 3052 4732
rect 3220 4676 3276 4732
rect 3332 4564 3388 4620
rect 4116 6580 4172 6636
rect 4452 6692 4508 6748
rect 4956 7140 5012 7196
rect 5684 7588 5740 7644
rect 8708 9994 8764 9996
rect 8708 9942 8710 9994
rect 8710 9942 8762 9994
rect 8762 9942 8764 9994
rect 8708 9940 8764 9942
rect 8820 9716 8876 9772
rect 8260 9492 8316 9548
rect 8036 9268 8092 9324
rect 7588 9210 7644 9212
rect 7588 9158 7590 9210
rect 7590 9158 7642 9210
rect 7642 9158 7644 9210
rect 7588 9156 7644 9158
rect 7532 8986 7588 8988
rect 7532 8934 7534 8986
rect 7534 8934 7586 8986
rect 7586 8934 7588 8986
rect 7532 8932 7588 8934
rect 7924 8986 7980 8988
rect 7924 8934 7926 8986
rect 7926 8934 7978 8986
rect 7978 8934 7980 8986
rect 7924 8932 7980 8934
rect 7308 8708 7364 8764
rect 7420 8484 7476 8540
rect 7028 8260 7084 8316
rect 6580 7588 6636 7644
rect 6804 7700 6860 7756
rect 6020 7530 6076 7532
rect 6020 7478 6022 7530
rect 6022 7478 6074 7530
rect 6074 7478 6076 7530
rect 6020 7476 6076 7478
rect 6692 7476 6748 7532
rect 5460 7252 5516 7308
rect 6356 7140 6412 7196
rect 6468 7364 6524 7420
rect 5348 6804 5404 6860
rect 5236 6468 5292 6524
rect 4340 6356 4396 6412
rect 4958 6298 5014 6300
rect 4958 6246 4960 6298
rect 4960 6246 5012 6298
rect 5012 6246 5014 6298
rect 4958 6244 5014 6246
rect 5062 6298 5118 6300
rect 5062 6246 5064 6298
rect 5064 6246 5116 6298
rect 5116 6246 5118 6298
rect 5062 6244 5118 6246
rect 5166 6298 5222 6300
rect 5166 6246 5168 6298
rect 5168 6246 5220 6298
rect 5220 6246 5222 6298
rect 5166 6244 5222 6246
rect 6244 6804 6300 6860
rect 5684 6580 5740 6636
rect 6132 6580 6188 6636
rect 6188 6356 6244 6412
rect 4732 6074 4788 6076
rect 4732 6022 4734 6074
rect 4734 6022 4786 6074
rect 4786 6022 4788 6074
rect 4732 6020 4788 6022
rect 3836 5178 3892 5180
rect 3836 5126 3838 5178
rect 3838 5126 3890 5178
rect 3890 5126 3892 5178
rect 3836 5124 3892 5126
rect 3556 4564 3612 4620
rect 3668 4900 3724 4956
rect 2996 3780 3052 3836
rect 1876 3444 1932 3500
rect 2436 3444 2492 3500
rect 3332 4004 3388 4060
rect 3780 4350 3836 4396
rect 3780 4340 3782 4350
rect 3782 4340 3834 4350
rect 3834 4340 3836 4350
rect 4004 4490 4006 4508
rect 4006 4490 4058 4508
rect 4058 4490 4060 4508
rect 4004 4452 4060 4490
rect 3220 2602 3276 2604
rect 3220 2550 3222 2602
rect 3222 2550 3274 2602
rect 3274 2550 3276 2602
rect 3220 2548 3276 2550
rect 2660 2436 2716 2492
rect 3332 2324 3388 2380
rect 7252 7364 7308 7420
rect 6972 7028 7028 7084
rect 6804 6916 6860 6972
rect 8148 9156 8204 9212
rect 10332 10836 10388 10892
rect 10164 10612 10220 10668
rect 10052 10164 10108 10220
rect 9436 9882 9492 9884
rect 9436 9830 9438 9882
rect 9438 9830 9490 9882
rect 9490 9830 9492 9882
rect 9436 9828 9492 9830
rect 10164 9940 10220 9996
rect 10276 10052 10332 10108
rect 10164 9716 10220 9772
rect 9604 9658 9660 9660
rect 9604 9606 9606 9658
rect 9606 9606 9658 9658
rect 9658 9606 9660 9658
rect 9604 9604 9660 9606
rect 8260 8820 8316 8876
rect 8148 8708 8204 8764
rect 8372 8932 8428 8988
rect 8540 8820 8596 8876
rect 9100 8874 9156 8876
rect 9100 8822 9102 8874
rect 9102 8822 9154 8874
rect 9154 8822 9156 8874
rect 9100 8820 9156 8822
rect 8484 8372 8540 8428
rect 8928 8650 8984 8652
rect 8928 8598 8930 8650
rect 8930 8598 8982 8650
rect 8982 8598 8984 8650
rect 8928 8596 8984 8598
rect 9032 8650 9088 8652
rect 9032 8598 9034 8650
rect 9034 8598 9086 8650
rect 9086 8598 9088 8650
rect 9032 8596 9088 8598
rect 9136 8650 9192 8652
rect 9136 8598 9138 8650
rect 9138 8598 9190 8650
rect 9190 8598 9192 8650
rect 9136 8596 9192 8598
rect 9268 8596 9324 8652
rect 9772 8596 9828 8652
rect 11396 11338 11452 11340
rect 11396 11286 11398 11338
rect 11398 11286 11450 11338
rect 11450 11286 11452 11338
rect 11396 11284 11452 11286
rect 11508 11172 11564 11228
rect 11396 10836 11452 10892
rect 10892 10442 10948 10444
rect 10892 10390 10894 10442
rect 10894 10390 10946 10442
rect 10946 10390 10948 10442
rect 10892 10388 10948 10390
rect 10780 10052 10836 10108
rect 11228 10052 11284 10108
rect 12012 11284 12068 11340
rect 12852 17444 12908 17500
rect 12898 17274 12954 17276
rect 12898 17222 12900 17274
rect 12900 17222 12952 17274
rect 12952 17222 12954 17274
rect 12898 17220 12954 17222
rect 13002 17274 13058 17276
rect 13002 17222 13004 17274
rect 13004 17222 13056 17274
rect 13056 17222 13058 17274
rect 13002 17220 13058 17222
rect 13106 17274 13162 17276
rect 13106 17222 13108 17274
rect 13108 17222 13160 17274
rect 13160 17222 13162 17274
rect 13106 17220 13162 17222
rect 13300 16884 13356 16940
rect 12908 16714 12964 16716
rect 12908 16662 12910 16714
rect 12910 16662 12962 16714
rect 12962 16662 12964 16714
rect 12908 16660 12964 16662
rect 13748 16324 13804 16380
rect 14140 16884 14196 16940
rect 15092 17444 15148 17500
rect 15428 16772 15484 16828
rect 14140 16324 14196 16380
rect 14868 16548 14924 16604
rect 12898 15706 12954 15708
rect 12898 15654 12900 15706
rect 12900 15654 12952 15706
rect 12952 15654 12954 15706
rect 12898 15652 12954 15654
rect 13002 15706 13058 15708
rect 13002 15654 13004 15706
rect 13004 15654 13056 15706
rect 13056 15654 13058 15706
rect 13002 15652 13058 15654
rect 13106 15706 13162 15708
rect 13106 15654 13108 15706
rect 13108 15654 13160 15706
rect 13160 15654 13162 15706
rect 13106 15652 13162 15654
rect 13412 15092 13468 15148
rect 13300 14756 13356 14812
rect 13188 14698 13244 14700
rect 13188 14646 13190 14698
rect 13190 14646 13242 14698
rect 13242 14646 13244 14698
rect 13188 14644 13244 14646
rect 12852 14420 12908 14476
rect 13748 15540 13804 15596
rect 14644 15540 14700 15596
rect 14980 16100 15036 16156
rect 14364 15428 14420 15484
rect 14588 15370 14644 15372
rect 14588 15318 14590 15370
rect 14590 15318 14642 15370
rect 14642 15318 14644 15370
rect 14588 15316 14644 15318
rect 13804 15258 13860 15260
rect 13804 15206 13806 15258
rect 13806 15206 13858 15258
rect 13858 15206 13860 15258
rect 13804 15204 13860 15206
rect 15092 15764 15148 15820
rect 13636 15092 13692 15148
rect 14028 14756 14084 14812
rect 14308 14644 14364 14700
rect 13524 14308 13580 14364
rect 12898 14138 12954 14140
rect 12898 14086 12900 14138
rect 12900 14086 12952 14138
rect 12952 14086 12954 14138
rect 12898 14084 12954 14086
rect 13002 14138 13058 14140
rect 13002 14086 13004 14138
rect 13004 14086 13056 14138
rect 13056 14086 13058 14138
rect 13002 14084 13058 14086
rect 13106 14138 13162 14140
rect 13106 14086 13108 14138
rect 13108 14086 13160 14138
rect 13160 14086 13162 14138
rect 13106 14084 13162 14086
rect 13412 13748 13468 13804
rect 13636 13802 13692 13804
rect 13636 13750 13638 13802
rect 13638 13750 13690 13802
rect 13690 13750 13692 13802
rect 13636 13748 13692 13750
rect 14084 14354 14086 14364
rect 14086 14354 14138 14364
rect 14138 14354 14140 14364
rect 14084 14308 14140 14354
rect 13300 13300 13356 13356
rect 13636 13188 13692 13244
rect 13020 12794 13076 12796
rect 13020 12742 13022 12794
rect 13022 12742 13074 12794
rect 13074 12742 13076 12794
rect 13020 12740 13076 12742
rect 13636 12628 13692 12684
rect 12898 12570 12954 12572
rect 12898 12518 12900 12570
rect 12900 12518 12952 12570
rect 12952 12518 12954 12570
rect 12898 12516 12954 12518
rect 13002 12570 13058 12572
rect 13002 12518 13004 12570
rect 13004 12518 13056 12570
rect 13056 12518 13058 12570
rect 13002 12516 13058 12518
rect 13106 12570 13162 12572
rect 13106 12518 13108 12570
rect 13108 12518 13160 12570
rect 13160 12518 13162 12570
rect 13106 12516 13162 12518
rect 12628 12404 12684 12460
rect 12516 12234 12572 12236
rect 12516 12182 12518 12234
rect 12518 12182 12570 12234
rect 12570 12182 12572 12234
rect 12516 12180 12572 12182
rect 12796 11844 12852 11900
rect 12740 11620 12796 11676
rect 12964 11508 13020 11564
rect 12404 11284 12460 11340
rect 13748 12740 13804 12796
rect 14196 13188 14252 13244
rect 14196 12964 14252 13020
rect 14532 14420 14588 14476
rect 14532 13524 14588 13580
rect 15820 18452 15876 18508
rect 16548 18676 16604 18732
rect 18004 18564 18060 18620
rect 19236 18564 19292 18620
rect 16436 18394 16492 18396
rect 16436 18342 16438 18394
rect 16438 18342 16490 18394
rect 16490 18342 16492 18394
rect 16436 18340 16492 18342
rect 16604 18394 16660 18396
rect 16604 18342 16606 18394
rect 16606 18342 16658 18394
rect 16658 18342 16660 18394
rect 16604 18340 16660 18342
rect 15876 17668 15932 17724
rect 16212 18228 16268 18284
rect 16100 17722 16156 17724
rect 16100 17670 16102 17722
rect 16102 17670 16154 17722
rect 16154 17670 16156 17722
rect 16100 17668 16156 17670
rect 16436 18116 16492 18172
rect 16212 17444 16268 17500
rect 16324 18004 16380 18060
rect 16868 18058 16924 18060
rect 16868 18006 16870 18058
rect 16870 18006 16922 18058
rect 16922 18006 16924 18058
rect 16868 18004 16924 18006
rect 16972 18058 17028 18060
rect 16972 18006 16974 18058
rect 16974 18006 17026 18058
rect 17026 18006 17028 18058
rect 16972 18004 17028 18006
rect 17076 18058 17132 18060
rect 17076 18006 17078 18058
rect 17078 18006 17130 18058
rect 17130 18006 17132 18058
rect 17076 18004 17132 18006
rect 18228 18340 18284 18396
rect 18620 18394 18676 18396
rect 18620 18342 18622 18394
rect 18622 18342 18674 18394
rect 18674 18342 18676 18394
rect 18620 18340 18676 18342
rect 21868 18900 21924 18956
rect 20838 18842 20894 18844
rect 20838 18790 20840 18842
rect 20840 18790 20892 18842
rect 20892 18790 20894 18842
rect 20838 18788 20894 18790
rect 20942 18842 20998 18844
rect 20942 18790 20944 18842
rect 20944 18790 20996 18842
rect 20996 18790 20998 18842
rect 20942 18788 20998 18790
rect 21046 18842 21102 18844
rect 21046 18790 21048 18842
rect 21048 18790 21100 18842
rect 21100 18790 21102 18842
rect 21046 18788 21102 18790
rect 19460 18452 19516 18508
rect 21140 18462 21196 18508
rect 21140 18452 21142 18462
rect 21142 18452 21194 18462
rect 21194 18452 21196 18462
rect 18004 18116 18060 18172
rect 16772 16996 16828 17052
rect 15820 16266 15876 16268
rect 15820 16214 15822 16266
rect 15822 16214 15874 16266
rect 15874 16214 15876 16266
rect 15820 16212 15876 16214
rect 15932 16100 15988 16156
rect 17220 16894 17276 16940
rect 17220 16884 17222 16894
rect 17222 16884 17274 16894
rect 17274 16884 17276 16894
rect 16772 16714 16828 16716
rect 16772 16662 16774 16714
rect 16774 16662 16826 16714
rect 16826 16662 16828 16714
rect 16772 16660 16828 16662
rect 18396 17722 18452 17724
rect 18396 17670 18398 17722
rect 18398 17670 18450 17722
rect 18450 17670 18452 17722
rect 18396 17668 18452 17670
rect 18788 17610 18844 17612
rect 18788 17558 18790 17610
rect 18790 17558 18842 17610
rect 18842 17558 18844 17610
rect 18788 17556 18844 17558
rect 17780 17444 17836 17500
rect 17836 17220 17892 17276
rect 18004 16938 18060 16940
rect 18004 16886 18006 16938
rect 18006 16886 18058 16938
rect 18058 16886 18060 16938
rect 18004 16884 18060 16886
rect 23100 18618 23156 18620
rect 23100 18566 23102 18618
rect 23102 18566 23154 18618
rect 23154 18566 23156 18618
rect 23100 18564 23156 18566
rect 22596 18462 22652 18508
rect 22596 18452 22598 18462
rect 22598 18452 22650 18462
rect 22650 18452 22652 18462
rect 23996 18506 24052 18508
rect 23996 18454 23998 18506
rect 23998 18454 24050 18506
rect 24050 18454 24052 18506
rect 23996 18452 24052 18454
rect 26740 18900 26796 18956
rect 25788 18676 25844 18732
rect 23772 18394 23828 18396
rect 19516 17834 19572 17836
rect 19516 17782 19518 17834
rect 19518 17782 19570 17834
rect 19570 17782 19572 17834
rect 19516 17780 19572 17782
rect 20020 18228 20076 18284
rect 19740 17780 19796 17836
rect 19908 18116 19964 18172
rect 19236 17444 19292 17500
rect 17556 16714 17612 16716
rect 17556 16662 17558 16714
rect 17558 16662 17610 16714
rect 17610 16662 17612 16714
rect 17556 16660 17612 16662
rect 16868 16490 16924 16492
rect 16868 16438 16870 16490
rect 16870 16438 16922 16490
rect 16922 16438 16924 16490
rect 16868 16436 16924 16438
rect 16972 16490 17028 16492
rect 16972 16438 16974 16490
rect 16974 16438 17026 16490
rect 17026 16438 17028 16490
rect 16972 16436 17028 16438
rect 17076 16490 17132 16492
rect 17076 16438 17078 16490
rect 17078 16438 17130 16490
rect 17130 16438 17132 16490
rect 17076 16436 17132 16438
rect 15428 15764 15484 15820
rect 15316 15316 15372 15372
rect 15652 15540 15708 15596
rect 16212 15764 16268 15820
rect 16212 15540 16268 15596
rect 16100 15428 16156 15484
rect 16324 15428 16380 15484
rect 15652 15204 15708 15260
rect 15204 15092 15260 15148
rect 15092 13972 15148 14028
rect 15204 14420 15260 14476
rect 15316 14308 15372 14364
rect 15540 14868 15596 14924
rect 16324 14980 16380 15036
rect 15204 13748 15260 13804
rect 15428 13688 15430 13692
rect 15430 13688 15482 13692
rect 15482 13688 15484 13692
rect 15428 13636 15484 13688
rect 14756 13524 14812 13580
rect 15036 13578 15092 13580
rect 15036 13526 15038 13578
rect 15038 13526 15090 13578
rect 15090 13526 15092 13578
rect 15036 13524 15092 13526
rect 16100 13972 16156 14028
rect 15652 13412 15708 13468
rect 14756 13300 14812 13356
rect 14308 12852 14364 12908
rect 14644 13188 14700 13244
rect 14532 12740 14588 12796
rect 14084 12516 14140 12572
rect 14420 12068 14476 12124
rect 13524 11508 13580 11564
rect 13300 11396 13356 11452
rect 14308 11508 14364 11564
rect 11732 10164 11788 10220
rect 11620 10052 11676 10108
rect 11900 10052 11956 10108
rect 11060 9940 11116 9996
rect 11508 9716 11564 9772
rect 11732 9828 11788 9884
rect 11172 9492 11228 9548
rect 11900 9604 11956 9660
rect 11900 9268 11956 9324
rect 11620 8982 11622 8988
rect 11622 8982 11674 8988
rect 11674 8982 11676 8988
rect 11620 8932 11676 8982
rect 12292 9828 12348 9884
rect 12180 9492 12236 9548
rect 12572 11226 12628 11228
rect 12572 11174 12574 11226
rect 12574 11174 12626 11226
rect 12626 11174 12628 11226
rect 12572 11172 12628 11174
rect 13300 11172 13356 11228
rect 12898 11002 12954 11004
rect 12898 10950 12900 11002
rect 12900 10950 12952 11002
rect 12952 10950 12954 11002
rect 12898 10948 12954 10950
rect 13002 11002 13058 11004
rect 13002 10950 13004 11002
rect 13004 10950 13056 11002
rect 13056 10950 13058 11002
rect 13002 10948 13058 10950
rect 13106 11002 13162 11004
rect 13106 10950 13108 11002
rect 13108 10950 13160 11002
rect 13160 10950 13162 11002
rect 13106 10948 13162 10950
rect 13300 10948 13356 11004
rect 13412 10836 13468 10892
rect 13580 11060 13636 11116
rect 12852 10724 12908 10780
rect 15316 12852 15372 12908
rect 15540 13076 15596 13132
rect 15540 12852 15596 12908
rect 15540 12628 15596 12684
rect 15092 11620 15148 11676
rect 14476 11226 14532 11228
rect 14476 11174 14478 11226
rect 14478 11174 14530 11226
rect 14530 11174 14532 11226
rect 14476 11172 14532 11174
rect 14140 10724 14196 10780
rect 14308 10724 14364 10780
rect 12572 10554 12628 10556
rect 12572 10502 12574 10554
rect 12574 10502 12626 10554
rect 12626 10502 12628 10554
rect 12572 10500 12628 10502
rect 15988 13748 16044 13804
rect 16100 13412 16156 13468
rect 16772 16042 16828 16044
rect 16772 15990 16774 16042
rect 16774 15990 16826 16042
rect 16826 15990 16828 16042
rect 16772 15988 16828 15990
rect 16772 15764 16828 15820
rect 16996 15540 17052 15596
rect 23772 18342 23774 18394
rect 23774 18342 23826 18394
rect 23826 18342 23828 18394
rect 23772 18340 23828 18342
rect 26628 18340 26684 18396
rect 21364 17780 21420 17836
rect 20916 17602 20918 17612
rect 20918 17602 20970 17612
rect 20970 17602 20972 17612
rect 20916 17556 20972 17602
rect 20838 17274 20894 17276
rect 20838 17222 20840 17274
rect 20840 17222 20892 17274
rect 20892 17222 20894 17274
rect 20838 17220 20894 17222
rect 20942 17274 20998 17276
rect 20942 17222 20944 17274
rect 20944 17222 20996 17274
rect 20996 17222 20998 17274
rect 20942 17220 20998 17222
rect 21046 17274 21102 17276
rect 21046 17222 21048 17274
rect 21048 17222 21100 17274
rect 21100 17222 21102 17274
rect 21046 17220 21102 17222
rect 20020 16772 20076 16828
rect 18564 16660 18620 16716
rect 19292 16548 19348 16604
rect 19460 16436 19516 16492
rect 17780 16324 17836 16380
rect 17612 16154 17668 16156
rect 17612 16102 17614 16154
rect 17614 16102 17666 16154
rect 17666 16102 17668 16154
rect 17612 16100 17668 16102
rect 17388 15764 17444 15820
rect 17556 15764 17612 15820
rect 18620 16324 18676 16380
rect 17892 16100 17948 16156
rect 18004 15988 18060 16044
rect 18340 16100 18396 16156
rect 19292 16324 19348 16380
rect 18788 16212 18844 16268
rect 16604 14980 16660 15036
rect 18620 15540 18676 15596
rect 18732 15764 18788 15820
rect 18116 15370 18172 15372
rect 18116 15318 18118 15370
rect 18118 15318 18170 15370
rect 18170 15318 18172 15370
rect 18116 15316 18172 15318
rect 18564 15248 18566 15260
rect 18566 15248 18618 15260
rect 18618 15248 18620 15260
rect 17220 15092 17276 15148
rect 17612 15146 17668 15148
rect 16868 14922 16924 14924
rect 16868 14870 16870 14922
rect 16870 14870 16922 14922
rect 16922 14870 16924 14922
rect 16868 14868 16924 14870
rect 16972 14922 17028 14924
rect 16972 14870 16974 14922
rect 16974 14870 17026 14922
rect 17026 14870 17028 14922
rect 16972 14868 17028 14870
rect 17076 14922 17132 14924
rect 17076 14870 17078 14922
rect 17078 14870 17130 14922
rect 17130 14870 17132 14922
rect 17076 14868 17132 14870
rect 16548 13972 16604 14028
rect 16324 13524 16380 13580
rect 16436 13412 16492 13468
rect 17612 15094 17614 15146
rect 17614 15094 17666 15146
rect 17666 15094 17668 15146
rect 17612 15092 17668 15094
rect 18564 15204 18620 15248
rect 17388 14644 17444 14700
rect 17556 14756 17612 14812
rect 17388 14474 17444 14476
rect 17388 14422 17390 14474
rect 17390 14422 17442 14474
rect 17442 14422 17444 14474
rect 17388 14420 17444 14422
rect 17388 13860 17444 13916
rect 17108 13578 17164 13580
rect 17108 13526 17110 13578
rect 17110 13526 17162 13578
rect 17162 13526 17164 13578
rect 17108 13524 17164 13526
rect 16868 13354 16924 13356
rect 16868 13302 16870 13354
rect 16870 13302 16922 13354
rect 16922 13302 16924 13354
rect 16868 13300 16924 13302
rect 16972 13354 17028 13356
rect 16972 13302 16974 13354
rect 16974 13302 17026 13354
rect 17026 13302 17028 13354
rect 16972 13300 17028 13302
rect 17076 13354 17132 13356
rect 17076 13302 17078 13354
rect 17078 13302 17130 13354
rect 17130 13302 17132 13354
rect 17076 13300 17132 13302
rect 16380 12852 16436 12908
rect 16212 12628 16268 12684
rect 16996 12852 17052 12908
rect 15652 12114 15654 12124
rect 15654 12114 15706 12124
rect 15706 12114 15708 12124
rect 15652 12068 15708 12114
rect 15316 11284 15372 11340
rect 13804 10554 13860 10556
rect 12796 10442 12852 10444
rect 12796 10390 12798 10442
rect 12798 10390 12850 10442
rect 12850 10390 12852 10442
rect 12796 10388 12852 10390
rect 12852 10164 12908 10220
rect 12852 9994 12908 9996
rect 12852 9942 12854 9994
rect 12854 9942 12906 9994
rect 12906 9942 12908 9994
rect 12852 9940 12908 9942
rect 12516 9882 12572 9884
rect 12516 9830 12518 9882
rect 12518 9830 12570 9882
rect 12570 9830 12572 9882
rect 12516 9828 12572 9830
rect 13804 10502 13806 10554
rect 13806 10502 13858 10554
rect 13858 10502 13860 10554
rect 13804 10500 13860 10502
rect 13692 10276 13748 10332
rect 13412 9828 13468 9884
rect 12292 9604 12348 9660
rect 12292 9044 12348 9100
rect 10276 8484 10332 8540
rect 8708 8194 8710 8204
rect 8710 8194 8762 8204
rect 8762 8194 8764 8204
rect 8708 8148 8764 8194
rect 8932 7642 8988 7644
rect 8932 7590 8934 7642
rect 8934 7590 8986 7642
rect 8986 7590 8988 7642
rect 8932 7588 8988 7590
rect 7028 6804 7084 6860
rect 7644 7306 7700 7308
rect 7644 7254 7646 7306
rect 7646 7254 7698 7306
rect 7698 7254 7700 7306
rect 7644 7252 7700 7254
rect 7420 6804 7476 6860
rect 8204 7306 8260 7308
rect 8204 7254 8206 7306
rect 8206 7254 8258 7306
rect 8258 7254 8260 7306
rect 8204 7252 8260 7254
rect 9156 7306 9212 7308
rect 9156 7254 9158 7306
rect 9158 7254 9210 7306
rect 9210 7254 9212 7306
rect 9156 7252 9212 7254
rect 8928 7082 8984 7084
rect 8928 7030 8930 7082
rect 8930 7030 8982 7082
rect 8982 7030 8984 7082
rect 8928 7028 8984 7030
rect 9032 7082 9088 7084
rect 9032 7030 9034 7082
rect 9034 7030 9086 7082
rect 9086 7030 9088 7082
rect 9032 7028 9088 7030
rect 9136 7082 9192 7084
rect 9136 7030 9138 7082
rect 9138 7030 9190 7082
rect 9190 7030 9192 7082
rect 9136 7028 9192 7030
rect 7924 6804 7980 6860
rect 7700 6580 7756 6636
rect 6804 6468 6860 6524
rect 8148 6692 8204 6748
rect 7700 6244 7756 6300
rect 8036 6468 8092 6524
rect 7420 5962 7476 5964
rect 4508 5178 4564 5180
rect 4508 5126 4510 5178
rect 4510 5126 4562 5178
rect 4562 5126 4564 5178
rect 4508 5124 4564 5126
rect 4676 5460 4732 5516
rect 5404 5348 5460 5404
rect 4676 5124 4732 5180
rect 4788 5236 4844 5292
rect 4452 4676 4508 4732
rect 5908 5460 5964 5516
rect 7420 5910 7422 5962
rect 7422 5910 7474 5962
rect 7474 5910 7476 5962
rect 7420 5908 7476 5910
rect 6188 5236 6244 5292
rect 6916 5290 6972 5292
rect 6916 5238 6918 5290
rect 6918 5238 6970 5290
rect 6970 5238 6972 5290
rect 6916 5236 6972 5238
rect 5516 5124 5572 5180
rect 7140 5738 7196 5740
rect 7140 5686 7142 5738
rect 7142 5686 7194 5738
rect 7194 5686 7196 5738
rect 7140 5684 7196 5686
rect 7308 5178 7364 5180
rect 7308 5126 7310 5178
rect 7310 5126 7362 5178
rect 7362 5126 7364 5178
rect 7308 5124 7364 5126
rect 4900 5012 4956 5068
rect 5068 4954 5124 4956
rect 5068 4902 5070 4954
rect 5070 4902 5122 4954
rect 5122 4902 5124 4954
rect 5068 4900 5124 4902
rect 4788 4676 4844 4732
rect 4958 4730 5014 4732
rect 4958 4678 4960 4730
rect 4960 4678 5012 4730
rect 5012 4678 5014 4730
rect 4958 4676 5014 4678
rect 5062 4730 5118 4732
rect 5062 4678 5064 4730
rect 5064 4678 5116 4730
rect 5116 4678 5118 4730
rect 5062 4676 5118 4678
rect 5166 4730 5222 4732
rect 5166 4678 5168 4730
rect 5168 4678 5220 4730
rect 5220 4678 5222 4730
rect 5166 4676 5222 4678
rect 4116 3780 4172 3836
rect 4340 3780 4396 3836
rect 4116 3444 4172 3500
rect 5908 4952 5910 4956
rect 5910 4952 5962 4956
rect 5962 4952 5964 4956
rect 5908 4900 5964 4952
rect 6076 4788 6132 4844
rect 5348 4564 5404 4620
rect 6748 4954 6804 4956
rect 6748 4902 6750 4954
rect 6750 4902 6802 4954
rect 6802 4902 6804 4954
rect 6748 4900 6804 4902
rect 6524 4564 6580 4620
rect 4788 3722 4844 3724
rect 4788 3670 4790 3722
rect 4790 3670 4842 3722
rect 4842 3670 4844 3722
rect 4788 3668 4844 3670
rect 4900 3556 4956 3612
rect 6244 4456 6300 4508
rect 6244 4452 6246 4456
rect 6246 4452 6298 4456
rect 6298 4452 6300 4456
rect 6244 4004 6300 4060
rect 5796 3892 5852 3948
rect 4004 2324 4060 2380
rect 6412 3780 6468 3836
rect 2436 1930 2492 1932
rect 2436 1878 2438 1930
rect 2438 1878 2490 1930
rect 2490 1878 2492 1930
rect 2436 1876 2492 1878
rect 2548 1540 2604 1596
rect 4340 2772 4396 2828
rect 5348 3220 5404 3276
rect 4958 3162 5014 3164
rect 4958 3110 4960 3162
rect 4960 3110 5012 3162
rect 5012 3110 5014 3162
rect 4958 3108 5014 3110
rect 5062 3162 5118 3164
rect 5062 3110 5064 3162
rect 5064 3110 5116 3162
rect 5116 3110 5118 3162
rect 5062 3108 5118 3110
rect 5166 3162 5222 3164
rect 5166 3110 5168 3162
rect 5168 3110 5220 3162
rect 5220 3110 5222 3162
rect 5166 3108 5222 3110
rect 6076 3610 6132 3612
rect 6076 3558 6078 3610
rect 6078 3558 6130 3610
rect 6130 3558 6132 3610
rect 6076 3556 6132 3558
rect 6300 3498 6356 3500
rect 6300 3446 6302 3498
rect 6302 3446 6354 3498
rect 6354 3446 6356 3498
rect 6300 3444 6356 3446
rect 6860 4452 6916 4508
rect 8596 6580 8652 6636
rect 8484 6522 8540 6524
rect 8484 6470 8486 6522
rect 8486 6470 8538 6522
rect 8538 6470 8540 6522
rect 8484 6468 8540 6470
rect 8148 6356 8204 6412
rect 7812 5124 7868 5180
rect 8372 5908 8428 5964
rect 8036 5012 8092 5068
rect 7700 4788 7756 4844
rect 7924 4788 7980 4844
rect 7252 4564 7308 4620
rect 7084 4394 7140 4396
rect 7084 4342 7086 4394
rect 7086 4342 7138 4394
rect 7138 4342 7140 4394
rect 7084 4340 7140 4342
rect 7364 4340 7420 4396
rect 6804 4170 6860 4172
rect 6804 4118 6806 4170
rect 6806 4118 6858 4170
rect 6858 4118 6860 4170
rect 6804 4116 6860 4118
rect 7252 3892 7308 3948
rect 6916 3780 6972 3836
rect 6692 3668 6748 3724
rect 5796 3220 5852 3276
rect 6356 3220 6412 3276
rect 5348 2772 5404 2828
rect 4564 2548 4620 2604
rect 4788 2660 4844 2716
rect 5796 2772 5852 2828
rect 4788 2154 4844 2156
rect 4788 2102 4790 2154
rect 4790 2102 4842 2154
rect 4842 2102 4844 2154
rect 4788 2100 4844 2102
rect 5460 2100 5516 2156
rect 5572 2324 5628 2380
rect 4452 1764 4508 1820
rect 4958 1594 5014 1596
rect 4958 1542 4960 1594
rect 4960 1542 5012 1594
rect 5012 1542 5014 1594
rect 4958 1540 5014 1542
rect 5062 1594 5118 1596
rect 5062 1542 5064 1594
rect 5064 1542 5116 1594
rect 5116 1542 5118 1594
rect 5062 1540 5118 1542
rect 5166 1594 5222 1596
rect 5166 1542 5168 1594
rect 5168 1542 5220 1594
rect 5220 1542 5222 1594
rect 5166 1540 5222 1542
rect 4676 1132 4678 1148
rect 4678 1132 4730 1148
rect 4730 1132 4732 1148
rect 4676 1092 4732 1132
rect 5796 1876 5852 1932
rect 6356 2212 6412 2268
rect 6132 1876 6188 1932
rect 7028 3498 7084 3500
rect 7028 3446 7030 3498
rect 7030 3446 7082 3498
rect 7082 3446 7084 3498
rect 7028 3444 7084 3446
rect 6916 2772 6972 2828
rect 7140 3108 7196 3164
rect 7588 4340 7644 4396
rect 8148 4788 8204 4844
rect 8260 5460 8316 5516
rect 9940 7588 9996 7644
rect 9380 6580 9436 6636
rect 8820 6132 8876 6188
rect 8820 5908 8876 5964
rect 9044 6468 9100 6524
rect 10388 7140 10444 7196
rect 9828 6580 9884 6636
rect 9604 6522 9660 6524
rect 9604 6470 9606 6522
rect 9606 6470 9658 6522
rect 9658 6470 9660 6522
rect 9604 6468 9660 6470
rect 8484 5290 8540 5292
rect 8484 5238 8486 5290
rect 8486 5238 8538 5290
rect 8538 5238 8540 5290
rect 8484 5236 8540 5238
rect 7588 4116 7644 4172
rect 8372 3892 8428 3948
rect 7476 3556 7532 3612
rect 7588 3332 7644 3388
rect 6804 2660 6860 2716
rect 6804 1988 6860 2044
rect 7028 2660 7084 2716
rect 7812 3108 7868 3164
rect 8260 3332 8316 3388
rect 7196 2436 7252 2492
rect 7252 2212 7308 2268
rect 6972 1764 7028 1820
rect 7700 2548 7756 2604
rect 8928 5514 8984 5516
rect 8928 5462 8930 5514
rect 8930 5462 8982 5514
rect 8982 5462 8984 5514
rect 8928 5460 8984 5462
rect 9032 5514 9088 5516
rect 9032 5462 9034 5514
rect 9034 5462 9086 5514
rect 9086 5462 9088 5514
rect 9032 5460 9088 5462
rect 9136 5514 9192 5516
rect 9136 5462 9138 5514
rect 9138 5462 9190 5514
rect 9190 5462 9192 5514
rect 9136 5460 9192 5462
rect 8708 5236 8764 5292
rect 10332 6634 10388 6636
rect 10332 6582 10334 6634
rect 10334 6582 10386 6634
rect 10386 6582 10388 6634
rect 10332 6580 10388 6582
rect 9940 6468 9996 6524
rect 12516 9492 12572 9548
rect 13468 9492 13524 9548
rect 12898 9434 12954 9436
rect 12898 9382 12900 9434
rect 12900 9382 12952 9434
rect 12952 9382 12954 9434
rect 12898 9380 12954 9382
rect 13002 9434 13058 9436
rect 13002 9382 13004 9434
rect 13004 9382 13056 9434
rect 13056 9382 13058 9434
rect 13002 9380 13058 9382
rect 13106 9434 13162 9436
rect 13106 9382 13108 9434
rect 13108 9382 13160 9434
rect 13160 9382 13162 9434
rect 13106 9380 13162 9382
rect 14084 9940 14140 9996
rect 13916 9658 13972 9660
rect 13916 9606 13918 9658
rect 13918 9606 13970 9658
rect 13970 9606 13972 9658
rect 13916 9604 13972 9606
rect 14756 10724 14812 10780
rect 14756 10500 14812 10556
rect 14868 10388 14924 10444
rect 15148 10276 15204 10332
rect 14924 10052 14980 10108
rect 14420 9492 14476 9548
rect 14532 9754 14534 9772
rect 14534 9754 14586 9772
rect 14586 9754 14588 9772
rect 14532 9716 14588 9754
rect 13580 9268 13636 9324
rect 12628 9210 12684 9212
rect 12628 9158 12630 9210
rect 12630 9158 12682 9210
rect 12682 9158 12684 9210
rect 12628 9156 12684 9158
rect 13188 9156 13244 9212
rect 12404 8932 12460 8988
rect 12292 8314 12348 8316
rect 12292 8262 12294 8314
rect 12294 8262 12346 8314
rect 12346 8262 12348 8314
rect 12292 8260 12348 8262
rect 12180 8148 12236 8204
rect 11620 7700 11676 7756
rect 12796 8986 12852 8988
rect 12796 8934 12798 8986
rect 12798 8934 12850 8986
rect 12850 8934 12852 8986
rect 12796 8932 12852 8934
rect 12964 8596 13020 8652
rect 13972 9098 14028 9100
rect 13972 9046 13974 9098
rect 13974 9046 14026 9098
rect 14026 9046 14028 9098
rect 13972 9044 14028 9046
rect 14420 9054 14476 9100
rect 14420 9044 14422 9054
rect 14422 9044 14474 9054
rect 14474 9044 14476 9054
rect 13356 8986 13412 8988
rect 13356 8934 13358 8986
rect 13358 8934 13410 8986
rect 13410 8934 13412 8986
rect 13356 8932 13412 8934
rect 12898 7866 12954 7868
rect 12898 7814 12900 7866
rect 12900 7814 12952 7866
rect 12952 7814 12954 7866
rect 12898 7812 12954 7814
rect 13002 7866 13058 7868
rect 13002 7814 13004 7866
rect 13004 7814 13056 7866
rect 13056 7814 13058 7866
rect 13002 7812 13058 7814
rect 13106 7866 13162 7868
rect 13106 7814 13108 7866
rect 13108 7814 13160 7866
rect 13160 7814 13162 7866
rect 13106 7812 13162 7814
rect 10836 7252 10892 7308
rect 10668 7028 10724 7084
rect 10836 6916 10892 6972
rect 10500 6356 10556 6412
rect 10668 6020 10724 6076
rect 10948 5572 11004 5628
rect 10052 4564 10108 4620
rect 9940 4452 9996 4508
rect 9380 4004 9436 4060
rect 8928 3946 8984 3948
rect 8928 3894 8930 3946
rect 8930 3894 8982 3946
rect 8982 3894 8984 3946
rect 8928 3892 8984 3894
rect 9032 3946 9088 3948
rect 9032 3894 9034 3946
rect 9034 3894 9086 3946
rect 9086 3894 9088 3946
rect 9032 3892 9088 3894
rect 9136 3946 9192 3948
rect 9136 3894 9138 3946
rect 9138 3894 9190 3946
rect 9190 3894 9192 3946
rect 9136 3892 9192 3894
rect 9492 3780 9548 3836
rect 9268 3556 9324 3612
rect 7700 1876 7756 1932
rect 7924 1988 7980 2044
rect 8148 1764 8204 1820
rect 9492 3332 9548 3388
rect 9660 3610 9716 3612
rect 9660 3558 9662 3610
rect 9662 3558 9714 3610
rect 9714 3558 9716 3610
rect 9660 3556 9716 3558
rect 8092 1146 8148 1148
rect 8092 1094 8094 1146
rect 8094 1094 8146 1146
rect 8146 1094 8148 1146
rect 8092 1092 8148 1094
rect 8652 2826 8708 2828
rect 8652 2774 8654 2826
rect 8654 2774 8706 2826
rect 8706 2774 8708 2826
rect 8652 2772 8708 2774
rect 9156 2826 9212 2828
rect 9156 2774 9158 2826
rect 9158 2774 9210 2826
rect 9210 2774 9212 2826
rect 9156 2772 9212 2774
rect 8876 2714 8932 2716
rect 8876 2662 8878 2714
rect 8878 2662 8930 2714
rect 8930 2662 8932 2714
rect 8876 2660 8932 2662
rect 8928 2378 8984 2380
rect 8928 2326 8930 2378
rect 8930 2326 8982 2378
rect 8982 2326 8984 2378
rect 8928 2324 8984 2326
rect 9032 2378 9088 2380
rect 9032 2326 9034 2378
rect 9034 2326 9086 2378
rect 9086 2326 9088 2378
rect 9032 2324 9088 2326
rect 9136 2378 9192 2380
rect 9136 2326 9138 2378
rect 9138 2326 9190 2378
rect 9190 2326 9192 2378
rect 9136 2324 9192 2326
rect 9604 2772 9660 2828
rect 10948 4452 11004 4508
rect 11956 7404 11958 7420
rect 11958 7404 12010 7420
rect 12010 7404 12012 7420
rect 12796 7418 12852 7420
rect 11956 7364 12012 7404
rect 11284 7140 11340 7196
rect 11900 7028 11956 7084
rect 12796 7366 12798 7418
rect 12798 7366 12850 7418
rect 12850 7366 12852 7418
rect 12796 7364 12852 7366
rect 12516 7252 12572 7308
rect 14644 9658 14700 9660
rect 14644 9606 14646 9658
rect 14646 9606 14698 9658
rect 14698 9606 14700 9658
rect 14644 9604 14700 9606
rect 14756 9492 14812 9548
rect 14644 9054 14700 9100
rect 14644 9044 14646 9054
rect 14646 9044 14698 9054
rect 14698 9044 14700 9054
rect 14980 9828 15036 9884
rect 15876 11508 15932 11564
rect 15988 12068 16044 12124
rect 15540 10724 15596 10780
rect 15484 10500 15540 10556
rect 15484 10164 15540 10220
rect 15316 9716 15372 9772
rect 15428 9492 15484 9548
rect 15316 9044 15372 9100
rect 14868 8596 14924 8652
rect 14532 8148 14588 8204
rect 15428 7642 15484 7644
rect 15428 7590 15430 7642
rect 15430 7590 15482 7642
rect 15482 7590 15484 7642
rect 15428 7588 15484 7590
rect 15092 7486 15148 7532
rect 15092 7476 15094 7486
rect 15094 7476 15146 7486
rect 15146 7476 15148 7486
rect 16436 12114 16438 12124
rect 16438 12114 16490 12124
rect 16490 12114 16492 12124
rect 16436 12068 16492 12114
rect 17668 14644 17724 14700
rect 18956 15540 19012 15596
rect 18116 14644 18172 14700
rect 18620 14474 18676 14476
rect 18620 14422 18622 14474
rect 18622 14422 18674 14474
rect 18674 14422 18676 14474
rect 18620 14420 18676 14422
rect 17780 13860 17836 13916
rect 17668 13636 17724 13692
rect 17892 13748 17948 13804
rect 18396 14362 18452 14364
rect 18396 14310 18398 14362
rect 18398 14310 18450 14362
rect 18450 14310 18452 14362
rect 18396 14308 18452 14310
rect 17556 13412 17612 13468
rect 17332 12516 17388 12572
rect 17444 13188 17500 13244
rect 17892 13300 17948 13356
rect 19572 15540 19628 15596
rect 22036 18004 22092 18060
rect 22988 18282 23044 18284
rect 22988 18230 22990 18282
rect 22990 18230 23042 18282
rect 23042 18230 23044 18282
rect 22988 18228 23044 18230
rect 22260 18116 22316 18172
rect 23212 17834 23268 17836
rect 23212 17782 23214 17834
rect 23214 17782 23266 17834
rect 23266 17782 23268 17834
rect 23212 17780 23268 17782
rect 21980 16996 22036 17052
rect 19908 16212 19964 16268
rect 20524 16660 20580 16716
rect 20412 16548 20468 16604
rect 20636 16324 20692 16380
rect 19796 15652 19852 15708
rect 21308 16714 21364 16716
rect 21308 16662 21310 16714
rect 21310 16662 21362 16714
rect 21362 16662 21364 16714
rect 21308 16660 21364 16662
rect 22260 16812 22262 16828
rect 22262 16812 22314 16828
rect 22314 16812 22316 16828
rect 24808 18058 24864 18060
rect 24808 18006 24810 18058
rect 24810 18006 24862 18058
rect 24862 18006 24864 18058
rect 24808 18004 24864 18006
rect 24912 18058 24968 18060
rect 24912 18006 24914 18058
rect 24914 18006 24966 18058
rect 24966 18006 24968 18058
rect 24912 18004 24968 18006
rect 25016 18058 25072 18060
rect 25016 18006 25018 18058
rect 25018 18006 25070 18058
rect 25070 18006 25072 18058
rect 25016 18004 25072 18006
rect 23604 16884 23660 16940
rect 22260 16772 22316 16812
rect 22596 16548 22652 16604
rect 21756 16436 21812 16492
rect 21028 16212 21084 16268
rect 20838 15706 20894 15708
rect 20838 15654 20840 15706
rect 20840 15654 20892 15706
rect 20892 15654 20894 15706
rect 20838 15652 20894 15654
rect 20942 15706 20998 15708
rect 20942 15654 20944 15706
rect 20944 15654 20996 15706
rect 20996 15654 20998 15706
rect 20942 15652 20998 15654
rect 21046 15706 21102 15708
rect 21046 15654 21048 15706
rect 21048 15654 21100 15706
rect 21100 15654 21102 15706
rect 21046 15652 21102 15654
rect 22652 16324 22708 16380
rect 23884 16714 23940 16716
rect 23884 16662 23886 16714
rect 23886 16662 23938 16714
rect 23938 16662 23940 16714
rect 23884 16660 23940 16662
rect 24724 17560 24780 17612
rect 24724 17556 24726 17560
rect 24726 17556 24778 17560
rect 24778 17556 24780 17560
rect 25284 17610 25340 17612
rect 25284 17558 25286 17610
rect 25286 17558 25338 17610
rect 25338 17558 25340 17610
rect 25284 17556 25340 17558
rect 24388 16660 24444 16716
rect 24052 16548 24108 16604
rect 21812 16212 21868 16268
rect 20580 15540 20636 15596
rect 21196 15540 21252 15596
rect 21532 16154 21588 16156
rect 21532 16102 21534 16154
rect 21534 16102 21586 16154
rect 21586 16102 21588 16154
rect 21532 16100 21588 16102
rect 22260 16212 22316 16268
rect 22820 16212 22876 16268
rect 23380 16212 23436 16268
rect 23772 16154 23828 16156
rect 23772 16102 23774 16154
rect 23774 16102 23826 16154
rect 23826 16102 23828 16154
rect 23772 16100 23828 16102
rect 21532 15540 21588 15596
rect 22372 15540 22428 15596
rect 21700 15428 21756 15484
rect 21364 15316 21420 15372
rect 19572 15092 19628 15148
rect 19292 14698 19348 14700
rect 19292 14646 19294 14698
rect 19294 14646 19346 14698
rect 19346 14646 19348 14698
rect 19292 14644 19348 14646
rect 19852 14868 19908 14924
rect 20244 14756 20300 14812
rect 18900 14196 18956 14252
rect 18172 13300 18228 13356
rect 18452 13300 18508 13356
rect 18340 13188 18396 13244
rect 18564 13188 18620 13244
rect 18116 13076 18172 13132
rect 17780 12906 17836 12908
rect 17780 12854 17782 12906
rect 17782 12854 17834 12906
rect 17834 12854 17836 12906
rect 17780 12852 17836 12854
rect 17556 12740 17612 12796
rect 18004 12628 18060 12684
rect 18228 12852 18284 12908
rect 18340 12740 18396 12796
rect 16212 11956 16268 12012
rect 16884 11956 16940 12012
rect 17892 12180 17948 12236
rect 19012 14084 19068 14140
rect 19124 14308 19180 14364
rect 18788 13758 18844 13804
rect 18788 13748 18790 13758
rect 18790 13748 18842 13758
rect 18842 13748 18844 13758
rect 20692 14980 20748 15036
rect 20580 14644 20636 14700
rect 20244 14196 20300 14252
rect 20468 14466 20470 14476
rect 20470 14466 20522 14476
rect 20522 14466 20524 14476
rect 20468 14420 20524 14466
rect 20468 14196 20524 14252
rect 21084 14980 21140 15036
rect 21252 14980 21308 15036
rect 21532 15146 21588 15148
rect 21532 15094 21534 15146
rect 21534 15094 21586 15146
rect 21586 15094 21588 15146
rect 21532 15092 21588 15094
rect 22036 15204 22092 15260
rect 21252 14308 21308 14364
rect 21644 14698 21700 14700
rect 21644 14646 21646 14698
rect 21646 14646 21698 14698
rect 21698 14646 21700 14698
rect 21644 14644 21700 14646
rect 21980 14756 22036 14812
rect 22204 14644 22260 14700
rect 21700 14420 21756 14476
rect 20838 14138 20894 14140
rect 20838 14086 20840 14138
rect 20840 14086 20892 14138
rect 20892 14086 20894 14138
rect 20838 14084 20894 14086
rect 20942 14138 20998 14140
rect 20942 14086 20944 14138
rect 20944 14086 20996 14138
rect 20996 14086 20998 14138
rect 20942 14084 20998 14086
rect 21046 14138 21102 14140
rect 21046 14086 21048 14138
rect 21048 14086 21100 14138
rect 21100 14086 21102 14138
rect 21046 14084 21102 14086
rect 21700 14084 21756 14140
rect 20524 13690 20580 13692
rect 20524 13638 20526 13690
rect 20526 13638 20578 13690
rect 20578 13638 20580 13690
rect 22428 14586 22484 14588
rect 22428 14534 22430 14586
rect 22430 14534 22482 14586
rect 22482 14534 22484 14586
rect 22428 14532 22484 14534
rect 22764 15370 22820 15372
rect 22764 15318 22766 15370
rect 22766 15318 22818 15370
rect 22818 15318 22820 15370
rect 22764 15316 22820 15318
rect 22036 14196 22092 14252
rect 20524 13636 20580 13638
rect 18900 13188 18956 13244
rect 19348 13188 19404 13244
rect 19180 13018 19236 13020
rect 19180 12966 19182 13018
rect 19182 12966 19234 13018
rect 19234 12966 19236 13018
rect 19180 12964 19236 12966
rect 19740 13018 19796 13020
rect 19740 12966 19742 13018
rect 19742 12966 19794 13018
rect 19794 12966 19796 13018
rect 19740 12964 19796 12966
rect 20748 13578 20804 13580
rect 20748 13526 20750 13578
rect 20750 13526 20802 13578
rect 20802 13526 20804 13578
rect 20748 13524 20804 13526
rect 21364 13412 21420 13468
rect 20468 13188 20524 13244
rect 21364 13188 21420 13244
rect 21028 13130 21084 13132
rect 21028 13078 21030 13130
rect 21030 13078 21082 13130
rect 21082 13078 21084 13130
rect 21028 13076 21084 13078
rect 18676 12292 18732 12348
rect 18508 12122 18564 12124
rect 18508 12070 18510 12122
rect 18510 12070 18562 12122
rect 18562 12070 18564 12122
rect 18508 12068 18564 12070
rect 16868 11786 16924 11788
rect 16868 11734 16870 11786
rect 16870 11734 16922 11786
rect 16922 11734 16924 11786
rect 16868 11732 16924 11734
rect 16972 11786 17028 11788
rect 16972 11734 16974 11786
rect 16974 11734 17026 11786
rect 17026 11734 17028 11786
rect 16972 11732 17028 11734
rect 17076 11786 17132 11788
rect 17076 11734 17078 11786
rect 17078 11734 17130 11786
rect 17130 11734 17132 11786
rect 17076 11732 17132 11734
rect 16436 11284 16492 11340
rect 16940 11284 16996 11340
rect 17668 12010 17724 12012
rect 17668 11958 17670 12010
rect 17670 11958 17722 12010
rect 17722 11958 17724 12010
rect 17668 11956 17724 11958
rect 17388 11620 17444 11676
rect 17500 11562 17556 11564
rect 17500 11510 17502 11562
rect 17502 11510 17554 11562
rect 17554 11510 17556 11562
rect 17500 11508 17556 11510
rect 18284 11956 18340 12012
rect 18004 11620 18060 11676
rect 15988 9828 16044 9884
rect 15764 9716 15820 9772
rect 17332 10554 17388 10556
rect 17332 10502 17334 10554
rect 17334 10502 17386 10554
rect 17386 10502 17388 10554
rect 17332 10500 17388 10502
rect 19124 12292 19180 12348
rect 19908 12404 19964 12460
rect 19012 12180 19068 12236
rect 19348 11956 19404 12012
rect 19460 12180 19516 12236
rect 18900 11508 18956 11564
rect 19236 11844 19292 11900
rect 17780 10388 17836 10444
rect 16868 10218 16924 10220
rect 16868 10166 16870 10218
rect 16870 10166 16922 10218
rect 16922 10166 16924 10218
rect 16868 10164 16924 10166
rect 16972 10218 17028 10220
rect 16972 10166 16974 10218
rect 16974 10166 17026 10218
rect 17026 10166 17028 10218
rect 16972 10164 17028 10166
rect 17076 10218 17132 10220
rect 17076 10166 17078 10218
rect 17078 10166 17130 10218
rect 17130 10166 17132 10218
rect 17076 10164 17132 10166
rect 18788 11172 18844 11228
rect 18284 11060 18340 11116
rect 19012 11060 19068 11116
rect 18228 10554 18284 10556
rect 18228 10502 18230 10554
rect 18230 10502 18282 10554
rect 18282 10502 18284 10554
rect 18228 10500 18284 10502
rect 18116 9828 18172 9884
rect 18452 10388 18508 10444
rect 22036 13636 22092 13692
rect 22260 13690 22316 13692
rect 22260 13638 22262 13690
rect 22262 13638 22314 13690
rect 22314 13638 22316 13690
rect 22260 13636 22316 13638
rect 21924 13524 21980 13580
rect 21756 13300 21812 13356
rect 20692 12906 20748 12908
rect 20692 12854 20694 12906
rect 20694 12854 20746 12906
rect 20746 12854 20748 12906
rect 20692 12852 20748 12854
rect 20838 12570 20894 12572
rect 20838 12518 20840 12570
rect 20840 12518 20892 12570
rect 20892 12518 20894 12570
rect 20838 12516 20894 12518
rect 20942 12570 20998 12572
rect 20942 12518 20944 12570
rect 20944 12518 20996 12570
rect 20996 12518 20998 12570
rect 20942 12516 20998 12518
rect 21046 12570 21102 12572
rect 21046 12518 21048 12570
rect 21048 12518 21100 12570
rect 21100 12518 21102 12570
rect 21046 12516 21102 12518
rect 20132 12180 20188 12236
rect 20356 12346 20412 12348
rect 20356 12294 20358 12346
rect 20358 12294 20410 12346
rect 20410 12294 20412 12346
rect 20356 12292 20412 12294
rect 23380 15876 23436 15932
rect 23156 15652 23212 15708
rect 23268 15764 23324 15820
rect 23044 15428 23100 15484
rect 24612 16548 24668 16604
rect 24808 16490 24864 16492
rect 24808 16438 24810 16490
rect 24810 16438 24862 16490
rect 24862 16438 24864 16490
rect 24808 16436 24864 16438
rect 24912 16490 24968 16492
rect 24912 16438 24914 16490
rect 24914 16438 24966 16490
rect 24966 16438 24968 16490
rect 24912 16436 24968 16438
rect 25016 16490 25072 16492
rect 25016 16438 25018 16490
rect 25018 16438 25070 16490
rect 25070 16438 25072 16490
rect 25016 16436 25072 16438
rect 25900 18282 25956 18284
rect 25900 18230 25902 18282
rect 25902 18230 25954 18282
rect 25954 18230 25956 18282
rect 25900 18228 25956 18230
rect 26124 17834 26180 17836
rect 26124 17782 26126 17834
rect 26126 17782 26178 17834
rect 26178 17782 26180 17834
rect 26124 17780 26180 17782
rect 26292 16884 26348 16940
rect 25788 16714 25844 16716
rect 25788 16662 25790 16714
rect 25790 16662 25842 16714
rect 25842 16662 25844 16714
rect 25788 16660 25844 16662
rect 25732 16436 25788 16492
rect 25172 16212 25228 16268
rect 24612 16100 24668 16156
rect 24780 15876 24836 15932
rect 25396 15876 25452 15932
rect 24612 15428 24668 15484
rect 25396 15428 25452 15484
rect 26124 16266 26180 16268
rect 26124 16214 26126 16266
rect 26126 16214 26178 16266
rect 26178 16214 26180 16266
rect 26124 16212 26180 16214
rect 25956 16154 26012 16156
rect 25956 16102 25958 16154
rect 25958 16102 26010 16154
rect 26010 16102 26012 16154
rect 25956 16100 26012 16102
rect 26404 16100 26460 16156
rect 26068 15988 26124 16044
rect 28778 18842 28834 18844
rect 28778 18790 28780 18842
rect 28780 18790 28832 18842
rect 28832 18790 28834 18842
rect 28778 18788 28834 18790
rect 28882 18842 28938 18844
rect 28882 18790 28884 18842
rect 28884 18790 28936 18842
rect 28936 18790 28938 18842
rect 28882 18788 28938 18790
rect 28986 18842 29042 18844
rect 28986 18790 28988 18842
rect 28988 18790 29040 18842
rect 29040 18790 29042 18842
rect 28986 18788 29042 18790
rect 29092 18676 29148 18732
rect 27188 18462 27244 18508
rect 27188 18452 27190 18462
rect 27190 18452 27242 18462
rect 27242 18452 27244 18462
rect 28140 18506 28196 18508
rect 28140 18454 28142 18506
rect 28142 18454 28194 18506
rect 28194 18454 28196 18506
rect 28140 18452 28196 18454
rect 27636 18380 27638 18396
rect 27638 18380 27690 18396
rect 27690 18380 27692 18396
rect 27636 18340 27692 18380
rect 28756 18340 28812 18396
rect 26852 16436 26908 16492
rect 27188 18228 27244 18284
rect 28028 17610 28084 17612
rect 28028 17558 28030 17610
rect 28030 17558 28082 17610
rect 28082 17558 28084 17610
rect 28028 17556 28084 17558
rect 29988 18452 30044 18508
rect 30548 18452 30604 18508
rect 30716 18506 30772 18508
rect 30716 18454 30718 18506
rect 30718 18454 30770 18506
rect 30770 18454 30772 18506
rect 30716 18452 30772 18454
rect 29484 18282 29540 18284
rect 29484 18230 29486 18282
rect 29486 18230 29538 18282
rect 29538 18230 29540 18282
rect 29484 18228 29540 18230
rect 28778 17274 28834 17276
rect 28778 17222 28780 17274
rect 28780 17222 28832 17274
rect 28832 17222 28834 17274
rect 28778 17220 28834 17222
rect 28882 17274 28938 17276
rect 28882 17222 28884 17274
rect 28884 17222 28936 17274
rect 28936 17222 28938 17274
rect 28882 17220 28938 17222
rect 28986 17274 29042 17276
rect 28986 17222 28988 17274
rect 28988 17222 29040 17274
rect 29040 17222 29042 17274
rect 28986 17220 29042 17222
rect 26964 16212 27020 16268
rect 27244 16660 27300 16716
rect 27692 16714 27748 16716
rect 27692 16662 27694 16714
rect 27694 16662 27746 16714
rect 27746 16662 27748 16714
rect 27692 16660 27748 16662
rect 28476 16436 28532 16492
rect 26740 16100 26796 16156
rect 25116 15370 25172 15372
rect 25116 15318 25118 15370
rect 25118 15318 25170 15370
rect 25170 15318 25172 15370
rect 25116 15316 25172 15318
rect 24892 15258 24948 15260
rect 24892 15206 24894 15258
rect 24894 15206 24946 15258
rect 24946 15206 24948 15258
rect 24892 15204 24948 15206
rect 23436 15146 23492 15148
rect 23436 15094 23438 15146
rect 23438 15094 23490 15146
rect 23490 15094 23492 15146
rect 23436 15092 23492 15094
rect 24388 15092 24444 15148
rect 23044 14980 23100 15036
rect 23324 14980 23380 15036
rect 22932 14644 22988 14700
rect 23044 14756 23100 14812
rect 22932 14420 22988 14476
rect 24808 14922 24864 14924
rect 24808 14870 24810 14922
rect 24810 14870 24862 14922
rect 24862 14870 24864 14922
rect 24808 14868 24864 14870
rect 24912 14922 24968 14924
rect 24912 14870 24914 14922
rect 24914 14870 24966 14922
rect 24966 14870 24968 14922
rect 24912 14868 24968 14870
rect 25016 14922 25072 14924
rect 25016 14870 25018 14922
rect 25018 14870 25070 14922
rect 25070 14870 25072 14922
rect 25016 14868 25072 14870
rect 24612 14756 24668 14812
rect 22484 13860 22540 13916
rect 22652 13914 22708 13916
rect 22652 13862 22654 13914
rect 22654 13862 22706 13914
rect 22706 13862 22708 13914
rect 22652 13860 22708 13862
rect 22484 13524 22540 13580
rect 22148 12964 22204 13020
rect 23212 13972 23268 14028
rect 22820 13412 22876 13468
rect 23268 13300 23324 13356
rect 24052 14536 24108 14588
rect 24052 14532 24054 14536
rect 24054 14532 24106 14536
rect 24106 14532 24108 14536
rect 23716 14308 23772 14364
rect 23604 13748 23660 13804
rect 23716 13972 23772 14028
rect 23940 14356 23942 14364
rect 23942 14356 23994 14364
rect 23994 14356 23996 14364
rect 23940 14308 23996 14356
rect 24052 14196 24108 14252
rect 22372 13076 22428 13132
rect 22484 12898 22486 12908
rect 22486 12898 22538 12908
rect 22538 12898 22540 12908
rect 22484 12852 22540 12898
rect 20020 12122 20076 12124
rect 20020 12070 20022 12122
rect 20022 12070 20074 12122
rect 20074 12070 20076 12122
rect 20020 12068 20076 12070
rect 20748 12234 20804 12236
rect 20748 12182 20750 12234
rect 20750 12182 20802 12234
rect 20802 12182 20804 12234
rect 20748 12180 20804 12182
rect 22820 12974 22876 13020
rect 22820 12964 22822 12974
rect 22822 12964 22874 12974
rect 22874 12964 22876 12974
rect 22988 12906 23044 12908
rect 22988 12854 22990 12906
rect 22990 12854 23042 12906
rect 23042 12854 23044 12906
rect 22988 12852 23044 12854
rect 23828 13188 23884 13244
rect 24836 14644 24892 14700
rect 26012 15258 26068 15260
rect 26012 15206 26014 15258
rect 26014 15206 26066 15258
rect 26066 15206 26068 15258
rect 26012 15204 26068 15206
rect 28308 15876 28364 15932
rect 27412 15316 27468 15372
rect 28868 15876 28924 15932
rect 30100 18282 30156 18284
rect 30100 18230 30102 18282
rect 30102 18230 30154 18282
rect 30154 18230 30156 18282
rect 30100 18228 30156 18230
rect 29932 17610 29988 17612
rect 29932 17558 29934 17610
rect 29934 17558 29986 17610
rect 29986 17558 29988 17610
rect 29932 17556 29988 17558
rect 30772 17444 30828 17500
rect 31780 18228 31836 18284
rect 32004 17780 32060 17836
rect 32116 18228 32172 18284
rect 31220 17556 31276 17612
rect 29540 16772 29596 16828
rect 31332 17444 31388 17500
rect 29316 15764 29372 15820
rect 28778 15706 28834 15708
rect 28778 15654 28780 15706
rect 28780 15654 28832 15706
rect 28832 15654 28834 15706
rect 28778 15652 28834 15654
rect 28882 15706 28938 15708
rect 28882 15654 28884 15706
rect 28884 15654 28936 15706
rect 28936 15654 28938 15706
rect 28882 15652 28938 15654
rect 28986 15706 29042 15708
rect 28986 15654 28988 15706
rect 28988 15654 29040 15706
rect 29040 15654 29042 15706
rect 28986 15652 29042 15654
rect 25620 15092 25676 15148
rect 26740 15092 26796 15148
rect 25508 14756 25564 14812
rect 25284 14644 25340 14700
rect 24556 13972 24612 14028
rect 24780 14084 24836 14140
rect 25060 13860 25116 13916
rect 24808 13354 24864 13356
rect 24808 13302 24810 13354
rect 24810 13302 24862 13354
rect 24862 13302 24864 13354
rect 24808 13300 24864 13302
rect 24912 13354 24968 13356
rect 24912 13302 24914 13354
rect 24914 13302 24966 13354
rect 24966 13302 24968 13354
rect 24912 13300 24968 13302
rect 25016 13354 25072 13356
rect 25016 13302 25018 13354
rect 25018 13302 25070 13354
rect 25070 13302 25072 13354
rect 25016 13300 25072 13302
rect 25844 14532 25900 14588
rect 26124 14756 26180 14812
rect 26628 14644 26684 14700
rect 25396 13748 25452 13804
rect 25172 13188 25228 13244
rect 24164 13130 24220 13132
rect 24164 13078 24166 13130
rect 24166 13078 24218 13130
rect 24218 13078 24220 13130
rect 24164 13076 24220 13078
rect 23044 12628 23100 12684
rect 23772 12628 23828 12684
rect 23604 12404 23660 12460
rect 23772 12292 23828 12348
rect 20636 12122 20692 12124
rect 20636 12070 20638 12122
rect 20638 12070 20690 12122
rect 20690 12070 20692 12122
rect 20636 12068 20692 12070
rect 19684 11535 19686 11564
rect 19686 11535 19738 11564
rect 19738 11535 19740 11564
rect 19684 11508 19740 11535
rect 19796 10666 19852 10668
rect 19796 10614 19798 10666
rect 19798 10614 19850 10666
rect 19850 10614 19852 10666
rect 19796 10612 19852 10614
rect 20356 11844 20412 11900
rect 21140 11172 21196 11228
rect 20838 11002 20894 11004
rect 20838 10950 20840 11002
rect 20840 10950 20892 11002
rect 20892 10950 20894 11002
rect 20838 10948 20894 10950
rect 20942 11002 20998 11004
rect 20942 10950 20944 11002
rect 20944 10950 20996 11002
rect 20996 10950 20998 11002
rect 20942 10948 20998 10950
rect 21046 11002 21102 11004
rect 21046 10950 21048 11002
rect 21048 10950 21100 11002
rect 21100 10950 21102 11002
rect 21046 10948 21102 10950
rect 21364 11508 21420 11564
rect 21476 11172 21532 11228
rect 19348 10276 19404 10332
rect 19012 10164 19068 10220
rect 16884 9770 16940 9772
rect 16884 9718 16886 9770
rect 16886 9718 16938 9770
rect 16938 9718 16940 9770
rect 16884 9716 16940 9718
rect 15876 8372 15932 8428
rect 16868 8650 16924 8652
rect 16868 8598 16870 8650
rect 16870 8598 16922 8650
rect 16922 8598 16924 8650
rect 16868 8596 16924 8598
rect 16972 8650 17028 8652
rect 16972 8598 16974 8650
rect 16974 8598 17026 8650
rect 17026 8598 17028 8650
rect 16972 8596 17028 8598
rect 17076 8650 17132 8652
rect 17076 8598 17078 8650
rect 17078 8598 17130 8650
rect 17130 8598 17132 8650
rect 17076 8596 17132 8598
rect 16660 8372 16716 8428
rect 16212 7588 16268 7644
rect 13300 7252 13356 7308
rect 12348 6916 12404 6972
rect 11732 6580 11788 6636
rect 11620 6522 11676 6524
rect 11620 6470 11622 6522
rect 11622 6470 11674 6522
rect 11674 6470 11676 6522
rect 11620 6468 11676 6470
rect 12068 6356 12124 6412
rect 12180 6244 12236 6300
rect 12180 5460 12236 5516
rect 12516 6626 12518 6636
rect 12518 6626 12570 6636
rect 12570 6626 12572 6636
rect 12516 6580 12572 6626
rect 13916 7306 13972 7308
rect 13916 7254 13918 7306
rect 13918 7254 13970 7306
rect 13970 7254 13972 7306
rect 13916 7252 13972 7254
rect 13076 6702 13132 6748
rect 13076 6692 13078 6702
rect 13078 6692 13130 6702
rect 13130 6692 13132 6702
rect 14420 6692 14476 6748
rect 14644 7028 14700 7084
rect 12898 6298 12954 6300
rect 12898 6246 12900 6298
rect 12900 6246 12952 6298
rect 12952 6246 12954 6298
rect 12898 6244 12954 6246
rect 13002 6298 13058 6300
rect 13002 6246 13004 6298
rect 13004 6246 13056 6298
rect 13056 6246 13058 6298
rect 13002 6244 13058 6246
rect 13106 6298 13162 6300
rect 13106 6246 13108 6298
rect 13108 6246 13160 6298
rect 13160 6246 13162 6298
rect 13106 6244 13162 6246
rect 12852 6074 12908 6076
rect 12852 6022 12854 6074
rect 12854 6022 12906 6074
rect 12906 6022 12908 6074
rect 12852 6020 12908 6022
rect 13636 6020 13692 6076
rect 12740 5684 12796 5740
rect 13300 5684 13356 5740
rect 12292 5124 12348 5180
rect 12516 4900 12572 4956
rect 10332 4116 10388 4172
rect 10052 4004 10108 4060
rect 10668 4116 10724 4172
rect 11676 4116 11732 4172
rect 12404 3892 12460 3948
rect 10836 3668 10892 3724
rect 11284 3780 11340 3836
rect 10164 3444 10220 3500
rect 9940 2660 9996 2716
rect 9604 1922 9606 1932
rect 9606 1922 9658 1932
rect 9658 1922 9660 1932
rect 9604 1876 9660 1922
rect 8484 1540 8540 1596
rect 8820 1370 8876 1372
rect 8820 1318 8822 1370
rect 8822 1318 8874 1370
rect 8874 1318 8876 1370
rect 8820 1316 8876 1318
rect 11116 3386 11172 3388
rect 11116 3334 11118 3386
rect 11118 3334 11170 3386
rect 11170 3334 11172 3386
rect 11116 3332 11172 3334
rect 10724 1540 10780 1596
rect 10836 1652 10892 1708
rect 12292 3668 12348 3724
rect 12898 4730 12954 4732
rect 12898 4678 12900 4730
rect 12900 4678 12952 4730
rect 12952 4678 12954 4730
rect 12898 4676 12954 4678
rect 13002 4730 13058 4732
rect 13002 4678 13004 4730
rect 13004 4678 13056 4730
rect 13056 4678 13058 4730
rect 13002 4676 13058 4678
rect 13106 4730 13162 4732
rect 13106 4678 13108 4730
rect 13108 4678 13160 4730
rect 13160 4678 13162 4730
rect 13106 4676 13162 4678
rect 12796 4506 12852 4508
rect 12796 4454 12798 4506
rect 12798 4454 12850 4506
rect 12850 4454 12852 4506
rect 12796 4452 12852 4454
rect 13860 5850 13916 5852
rect 13860 5798 13862 5850
rect 13862 5798 13914 5850
rect 13914 5798 13916 5850
rect 13860 5796 13916 5798
rect 13524 4900 13580 4956
rect 13412 4676 13468 4732
rect 13804 4564 13860 4620
rect 14756 6804 14812 6860
rect 14980 7252 15036 7308
rect 14140 5738 14196 5740
rect 14140 5686 14142 5738
rect 14142 5686 14194 5738
rect 14194 5686 14196 5738
rect 14140 5684 14196 5686
rect 14644 5684 14700 5740
rect 17276 8426 17332 8428
rect 17276 8374 17278 8426
rect 17278 8374 17330 8426
rect 17330 8374 17332 8426
rect 17276 8372 17332 8374
rect 18004 9762 18006 9772
rect 18006 9762 18058 9772
rect 18058 9762 18060 9772
rect 18004 9716 18060 9762
rect 21868 11172 21924 11228
rect 23156 10724 23212 10780
rect 24612 13076 24668 13132
rect 24500 12964 24556 13020
rect 24500 12740 24556 12796
rect 25508 13524 25564 13580
rect 25340 13076 25396 13132
rect 27916 15258 27972 15260
rect 27916 15206 27918 15258
rect 27918 15206 27970 15258
rect 27970 15206 27972 15258
rect 27916 15204 27972 15206
rect 28756 15428 28812 15484
rect 27412 14644 27468 14700
rect 27804 14698 27860 14700
rect 27804 14646 27806 14698
rect 27806 14646 27858 14698
rect 27858 14646 27860 14698
rect 27804 14644 27860 14646
rect 28364 15092 28420 15148
rect 29204 15092 29260 15148
rect 30772 16100 30828 16156
rect 31220 16660 31276 16716
rect 31500 16772 31556 16828
rect 30548 16042 30604 16044
rect 30548 15990 30550 16042
rect 30550 15990 30602 16042
rect 30602 15990 30604 16042
rect 30548 15988 30604 15990
rect 30772 15428 30828 15484
rect 31332 15988 31388 16044
rect 31612 15316 31668 15372
rect 30212 15204 30268 15260
rect 31220 15243 31222 15260
rect 31222 15243 31274 15260
rect 31274 15243 31276 15260
rect 31220 15204 31276 15243
rect 30044 15092 30100 15148
rect 30996 15092 31052 15148
rect 31836 15146 31892 15148
rect 31836 15094 31838 15146
rect 31838 15094 31890 15146
rect 31890 15094 31892 15146
rect 31836 15092 31892 15094
rect 32340 14868 32396 14924
rect 31724 14586 31780 14588
rect 31724 14534 31726 14586
rect 31726 14534 31778 14586
rect 31778 14534 31780 14586
rect 31724 14532 31780 14534
rect 27244 14308 27300 14364
rect 27524 14308 27580 14364
rect 26908 13972 26964 14028
rect 28700 14362 28756 14364
rect 28700 14310 28702 14362
rect 28702 14310 28754 14362
rect 28754 14310 28756 14362
rect 28700 14308 28756 14310
rect 28778 14138 28834 14140
rect 28778 14086 28780 14138
rect 28780 14086 28832 14138
rect 28832 14086 28834 14138
rect 28778 14084 28834 14086
rect 28882 14138 28938 14140
rect 28882 14086 28884 14138
rect 28884 14086 28936 14138
rect 28936 14086 28938 14138
rect 28882 14084 28938 14086
rect 28986 14138 29042 14140
rect 28986 14086 28988 14138
rect 28988 14086 29040 14138
rect 29040 14086 29042 14138
rect 28986 14084 29042 14086
rect 27804 13914 27860 13916
rect 27804 13862 27806 13914
rect 27806 13862 27858 13914
rect 27858 13862 27860 13914
rect 27804 13860 27860 13862
rect 24780 12906 24836 12908
rect 24780 12854 24782 12906
rect 24782 12854 24834 12906
rect 24834 12854 24836 12906
rect 24780 12852 24836 12854
rect 26068 13076 26124 13132
rect 25788 12964 25844 13020
rect 25620 12852 25676 12908
rect 25060 12740 25116 12796
rect 24500 12122 24556 12124
rect 24500 12070 24502 12122
rect 24502 12070 24554 12122
rect 24554 12070 24556 12122
rect 24500 12068 24556 12070
rect 24668 11844 24724 11900
rect 24808 11786 24864 11788
rect 24808 11734 24810 11786
rect 24810 11734 24862 11786
rect 24862 11734 24864 11786
rect 24808 11732 24864 11734
rect 24912 11786 24968 11788
rect 24912 11734 24914 11786
rect 24914 11734 24966 11786
rect 24966 11734 24968 11786
rect 24912 11732 24968 11734
rect 25016 11786 25072 11788
rect 25016 11734 25018 11786
rect 25018 11734 25070 11786
rect 25070 11734 25072 11786
rect 25016 11732 25072 11734
rect 23548 10276 23604 10332
rect 21028 9828 21084 9884
rect 25788 11620 25844 11676
rect 29316 14308 29372 14364
rect 26404 13524 26460 13580
rect 27076 13524 27132 13580
rect 26628 13412 26684 13468
rect 27300 13412 27356 13468
rect 27188 13076 27244 13132
rect 26292 12628 26348 12684
rect 28252 13076 28308 13132
rect 28028 12906 28084 12908
rect 28028 12854 28030 12906
rect 28030 12854 28082 12906
rect 28082 12854 28084 12906
rect 29204 13076 29260 13132
rect 28028 12852 28084 12854
rect 26628 12122 26684 12124
rect 26628 12070 26630 12122
rect 26630 12070 26682 12122
rect 26682 12070 26684 12122
rect 26628 12068 26684 12070
rect 27188 12108 27190 12124
rect 27190 12108 27242 12124
rect 27242 12108 27244 12124
rect 27188 12068 27244 12108
rect 26068 11620 26124 11676
rect 26852 11450 26908 11452
rect 26852 11398 26854 11450
rect 26854 11398 26906 11450
rect 26906 11398 26908 11450
rect 26852 11396 26908 11398
rect 23996 10778 24052 10780
rect 23996 10726 23998 10778
rect 23998 10726 24050 10778
rect 24050 10726 24052 10778
rect 23996 10724 24052 10726
rect 24556 10778 24612 10780
rect 24556 10726 24558 10778
rect 24558 10726 24610 10778
rect 24610 10726 24612 10778
rect 24556 10724 24612 10726
rect 25284 10724 25340 10780
rect 24108 10554 24164 10556
rect 24108 10502 24110 10554
rect 24110 10502 24162 10554
rect 24162 10502 24164 10554
rect 24108 10500 24164 10502
rect 24892 10554 24948 10556
rect 24892 10502 24894 10554
rect 24894 10502 24946 10554
rect 24946 10502 24948 10554
rect 24892 10500 24948 10502
rect 26068 10500 26124 10556
rect 24444 10442 24500 10444
rect 24444 10390 24446 10442
rect 24446 10390 24498 10442
rect 24498 10390 24500 10442
rect 24444 10388 24500 10390
rect 25004 10442 25060 10444
rect 25004 10390 25006 10442
rect 25006 10390 25058 10442
rect 25058 10390 25060 10442
rect 25004 10388 25060 10390
rect 25956 10388 26012 10444
rect 24808 10218 24864 10220
rect 24808 10166 24810 10218
rect 24810 10166 24862 10218
rect 24862 10166 24864 10218
rect 24808 10164 24864 10166
rect 24912 10218 24968 10220
rect 24912 10166 24914 10218
rect 24914 10166 24966 10218
rect 24966 10166 24968 10218
rect 24912 10164 24968 10166
rect 25016 10218 25072 10220
rect 25016 10166 25018 10218
rect 25018 10166 25070 10218
rect 25070 10166 25072 10218
rect 25016 10164 25072 10166
rect 24836 9940 24892 9996
rect 20838 9434 20894 9436
rect 20838 9382 20840 9434
rect 20840 9382 20892 9434
rect 20892 9382 20894 9434
rect 20838 9380 20894 9382
rect 20942 9434 20998 9436
rect 20942 9382 20944 9434
rect 20944 9382 20996 9434
rect 20996 9382 20998 9434
rect 20942 9380 20998 9382
rect 21046 9434 21102 9436
rect 21046 9382 21048 9434
rect 21048 9382 21100 9434
rect 21100 9382 21102 9434
rect 21046 9380 21102 9382
rect 19964 8986 20020 8988
rect 19964 8934 19966 8986
rect 19966 8934 20018 8986
rect 20018 8934 20020 8986
rect 19964 8932 20020 8934
rect 17444 8372 17500 8428
rect 17556 8314 17612 8316
rect 17556 8262 17558 8314
rect 17558 8262 17610 8314
rect 17610 8262 17612 8314
rect 17556 8260 17612 8262
rect 16884 8202 16940 8204
rect 16884 8150 16886 8202
rect 16886 8150 16938 8202
rect 16938 8150 16940 8202
rect 16884 8148 16940 8150
rect 16884 7528 16886 7532
rect 16886 7528 16938 7532
rect 16938 7528 16940 7532
rect 16884 7476 16940 7528
rect 16868 7082 16924 7084
rect 16868 7030 16870 7082
rect 16870 7030 16922 7082
rect 16922 7030 16924 7082
rect 16868 7028 16924 7030
rect 16972 7082 17028 7084
rect 16972 7030 16974 7082
rect 16974 7030 17026 7082
rect 17026 7030 17028 7082
rect 16972 7028 17028 7030
rect 17076 7082 17132 7084
rect 17076 7030 17078 7082
rect 17078 7030 17130 7082
rect 17130 7030 17132 7082
rect 17076 7028 17132 7030
rect 15988 6858 16044 6860
rect 15988 6806 15990 6858
rect 15990 6806 16042 6858
rect 16042 6806 16044 6858
rect 15988 6804 16044 6806
rect 17220 6580 17276 6636
rect 14364 5460 14420 5516
rect 15540 5842 15542 5852
rect 15542 5842 15594 5852
rect 15594 5842 15596 5852
rect 15540 5796 15596 5842
rect 16380 5684 16436 5740
rect 15372 5460 15428 5516
rect 14532 5178 14588 5180
rect 14532 5126 14534 5178
rect 14534 5126 14586 5178
rect 14586 5126 14588 5178
rect 14532 5124 14588 5126
rect 14140 4954 14196 4956
rect 14140 4902 14142 4954
rect 14142 4902 14194 4954
rect 14194 4902 14196 4954
rect 14140 4900 14196 4902
rect 13972 4452 14028 4508
rect 14868 5124 14924 5180
rect 15596 5178 15652 5180
rect 15596 5126 15598 5178
rect 15598 5126 15650 5178
rect 15650 5126 15652 5178
rect 15596 5124 15652 5126
rect 14980 5012 15036 5068
rect 14868 4900 14924 4956
rect 14756 4676 14812 4732
rect 14532 4350 14588 4396
rect 14532 4340 14534 4350
rect 14534 4340 14586 4350
rect 14586 4340 14588 4350
rect 13076 4228 13132 4284
rect 11732 3604 11734 3612
rect 11734 3604 11786 3612
rect 11786 3604 11788 3612
rect 11732 3556 11788 3604
rect 13412 4282 13468 4284
rect 13412 4230 13414 4282
rect 13414 4230 13466 4282
rect 13466 4230 13468 4282
rect 13412 4228 13468 4230
rect 13188 3892 13244 3948
rect 13468 3780 13524 3836
rect 13748 3332 13804 3388
rect 10500 1132 10502 1148
rect 10502 1132 10554 1148
rect 10554 1132 10556 1148
rect 10500 1092 10556 1132
rect 12898 3162 12954 3164
rect 12898 3110 12900 3162
rect 12900 3110 12952 3162
rect 12952 3110 12954 3162
rect 12898 3108 12954 3110
rect 13002 3162 13058 3164
rect 13002 3110 13004 3162
rect 13004 3110 13056 3162
rect 13056 3110 13058 3162
rect 13002 3108 13058 3110
rect 13106 3162 13162 3164
rect 13106 3110 13108 3162
rect 13108 3110 13160 3162
rect 13160 3110 13162 3162
rect 13106 3108 13162 3110
rect 13468 2772 13524 2828
rect 12068 2212 12124 2268
rect 11508 2100 11564 2156
rect 12068 1988 12124 2044
rect 11396 980 11452 1036
rect 12404 2042 12460 2044
rect 12404 1990 12406 2042
rect 12406 1990 12458 2042
rect 12458 1990 12460 2042
rect 12404 1988 12460 1990
rect 12740 1876 12796 1932
rect 13076 2212 13132 2268
rect 14084 2100 14140 2156
rect 14196 4004 14252 4060
rect 14700 4228 14756 4284
rect 14868 4228 14924 4284
rect 14532 4004 14588 4060
rect 14588 3780 14644 3836
rect 14308 3556 14364 3612
rect 13300 1922 13302 1932
rect 13302 1922 13354 1932
rect 13354 1922 13356 1932
rect 13300 1876 13356 1922
rect 13860 1652 13916 1708
rect 12898 1594 12954 1596
rect 12898 1542 12900 1594
rect 12900 1542 12952 1594
rect 12952 1542 12954 1594
rect 12898 1540 12954 1542
rect 13002 1594 13058 1596
rect 13002 1542 13004 1594
rect 13004 1542 13056 1594
rect 13056 1542 13058 1594
rect 13002 1540 13058 1542
rect 13106 1594 13162 1596
rect 13106 1542 13108 1594
rect 13108 1542 13160 1594
rect 13160 1542 13162 1594
rect 13106 1540 13162 1542
rect 12180 1316 12236 1372
rect 14868 2772 14924 2828
rect 16660 5460 16716 5516
rect 16868 5514 16924 5516
rect 16868 5462 16870 5514
rect 16870 5462 16922 5514
rect 16922 5462 16924 5514
rect 16868 5460 16924 5462
rect 16972 5514 17028 5516
rect 16972 5462 16974 5514
rect 16974 5462 17026 5514
rect 17026 5462 17028 5514
rect 16972 5460 17028 5462
rect 17076 5514 17132 5516
rect 17076 5462 17078 5514
rect 17078 5462 17130 5514
rect 17130 5462 17132 5514
rect 17076 5460 17132 5462
rect 16380 4676 16436 4732
rect 17780 7486 17836 7532
rect 17780 7476 17782 7486
rect 17782 7476 17834 7486
rect 17834 7476 17836 7486
rect 17780 6692 17836 6748
rect 17892 6916 17948 6972
rect 18508 7642 18564 7644
rect 18508 7590 18510 7642
rect 18510 7590 18562 7642
rect 18562 7590 18564 7642
rect 18508 7588 18564 7590
rect 20356 8932 20412 8988
rect 20132 8260 20188 8316
rect 19796 8148 19852 8204
rect 18844 7418 18900 7420
rect 18844 7366 18846 7418
rect 18846 7366 18898 7418
rect 18898 7366 18900 7418
rect 18844 7364 18900 7366
rect 19236 7404 19238 7420
rect 19238 7404 19290 7420
rect 19290 7404 19292 7420
rect 19236 7364 19292 7404
rect 18676 6708 18732 6748
rect 18676 6692 18678 6708
rect 18678 6692 18730 6708
rect 18730 6692 18732 6708
rect 18228 6634 18284 6636
rect 18228 6582 18230 6634
rect 18230 6582 18282 6634
rect 18282 6582 18284 6634
rect 18228 6580 18284 6582
rect 18564 6132 18620 6188
rect 18788 5850 18844 5852
rect 18788 5798 18790 5850
rect 18790 5798 18842 5850
rect 18842 5798 18844 5850
rect 18788 5796 18844 5798
rect 17332 5124 17388 5180
rect 15092 3444 15148 3500
rect 15204 1876 15260 1932
rect 15876 4274 15878 4284
rect 15878 4274 15930 4284
rect 15930 4274 15932 4284
rect 15876 4228 15932 4274
rect 16660 4900 16716 4956
rect 17444 4788 17500 4844
rect 17892 4900 17948 4956
rect 16548 4340 16604 4396
rect 15652 3668 15708 3724
rect 15932 3780 15988 3836
rect 16156 3556 16212 3612
rect 15540 3490 15542 3500
rect 15542 3490 15594 3500
rect 15594 3490 15596 3500
rect 15540 3444 15596 3490
rect 15316 1540 15372 1596
rect 15428 1764 15484 1820
rect 13356 1258 13412 1260
rect 13356 1206 13358 1258
rect 13358 1206 13410 1258
rect 13410 1206 13412 1258
rect 13356 1204 13412 1206
rect 13748 1204 13804 1260
rect 11956 980 12012 1036
rect 14476 1146 14532 1148
rect 14476 1094 14478 1146
rect 14478 1094 14530 1146
rect 14530 1094 14532 1146
rect 14476 1092 14532 1094
rect 15204 1146 15260 1148
rect 15204 1094 15206 1146
rect 15206 1094 15258 1146
rect 15258 1094 15260 1146
rect 15204 1092 15260 1094
rect 15876 2602 15932 2604
rect 15876 2550 15878 2602
rect 15878 2550 15930 2602
rect 15930 2550 15932 2602
rect 15876 2548 15932 2550
rect 16212 1316 16268 1372
rect 17220 4228 17276 4284
rect 16868 3946 16924 3948
rect 16868 3894 16870 3946
rect 16870 3894 16922 3946
rect 16922 3894 16924 3946
rect 16868 3892 16924 3894
rect 16972 3946 17028 3948
rect 16972 3894 16974 3946
rect 16974 3894 17026 3946
rect 17026 3894 17028 3946
rect 16972 3892 17028 3894
rect 17076 3946 17132 3948
rect 17076 3894 17078 3946
rect 17078 3894 17130 3946
rect 17130 3894 17132 3946
rect 17076 3892 17132 3894
rect 16548 3722 16604 3724
rect 16548 3670 16550 3722
rect 16550 3670 16602 3722
rect 16602 3670 16604 3722
rect 16548 3668 16604 3670
rect 16868 2378 16924 2380
rect 16868 2326 16870 2378
rect 16870 2326 16922 2378
rect 16922 2326 16924 2378
rect 16868 2324 16924 2326
rect 16972 2378 17028 2380
rect 16972 2326 16974 2378
rect 16974 2326 17026 2378
rect 17026 2326 17028 2378
rect 16972 2324 17028 2326
rect 17076 2378 17132 2380
rect 17076 2326 17078 2378
rect 17078 2326 17130 2378
rect 17130 2326 17132 2378
rect 17076 2324 17132 2326
rect 18452 5130 18508 5180
rect 18452 5124 18454 5130
rect 18454 5124 18506 5130
rect 18506 5124 18508 5130
rect 18228 4900 18284 4956
rect 18340 4340 18396 4396
rect 18788 5124 18844 5180
rect 19236 6916 19292 6972
rect 19796 6916 19852 6972
rect 19012 6356 19068 6412
rect 22260 9210 22316 9212
rect 22260 9158 22262 9210
rect 22262 9158 22314 9210
rect 22314 9158 22316 9210
rect 22260 9156 22316 9158
rect 21588 9096 21590 9100
rect 21590 9096 21642 9100
rect 21642 9096 21644 9100
rect 21588 9044 21644 9096
rect 23156 9054 23212 9100
rect 21420 8986 21476 8988
rect 21420 8934 21422 8986
rect 21422 8934 21474 8986
rect 21474 8934 21476 8986
rect 21420 8932 21476 8934
rect 23156 9044 23158 9054
rect 23158 9044 23210 9054
rect 23210 9044 23212 9054
rect 21252 8260 21308 8316
rect 20804 8148 20860 8204
rect 22036 8260 22092 8316
rect 21700 8148 21756 8204
rect 20838 7866 20894 7868
rect 20838 7814 20840 7866
rect 20840 7814 20892 7866
rect 20892 7814 20894 7866
rect 20838 7812 20894 7814
rect 20942 7866 20998 7868
rect 20942 7814 20944 7866
rect 20944 7814 20996 7866
rect 20996 7814 20998 7866
rect 20942 7812 20998 7814
rect 21046 7866 21102 7868
rect 21046 7814 21048 7866
rect 21048 7814 21100 7866
rect 21100 7814 21102 7866
rect 21046 7812 21102 7814
rect 20244 7642 20300 7644
rect 20244 7590 20246 7642
rect 20246 7590 20298 7642
rect 20298 7590 20300 7642
rect 20244 7588 20300 7590
rect 21924 8148 21980 8204
rect 24164 8820 24220 8876
rect 24808 8650 24864 8652
rect 24808 8598 24810 8650
rect 24810 8598 24862 8650
rect 24862 8598 24864 8650
rect 24808 8596 24864 8598
rect 24912 8650 24968 8652
rect 24912 8598 24914 8650
rect 24914 8598 24966 8650
rect 24966 8598 24968 8650
rect 24912 8596 24968 8598
rect 25016 8650 25072 8652
rect 25016 8598 25018 8650
rect 25018 8598 25070 8650
rect 25070 8598 25072 8650
rect 25016 8596 25072 8598
rect 24500 8260 24556 8316
rect 23716 8194 23718 8204
rect 23718 8194 23770 8204
rect 23770 8194 23772 8204
rect 23716 8148 23772 8194
rect 22820 7588 22876 7644
rect 21700 6804 21756 6860
rect 19684 6634 19740 6636
rect 19684 6582 19686 6634
rect 19686 6582 19738 6634
rect 19738 6582 19740 6634
rect 19684 6580 19740 6582
rect 19796 6356 19852 6412
rect 19684 5850 19740 5852
rect 19684 5798 19686 5850
rect 19686 5798 19738 5850
rect 19738 5798 19740 5850
rect 19684 5796 19740 5798
rect 20838 6298 20894 6300
rect 20838 6246 20840 6298
rect 20840 6246 20892 6298
rect 20892 6246 20894 6298
rect 20838 6244 20894 6246
rect 20942 6298 20998 6300
rect 20942 6246 20944 6298
rect 20944 6246 20996 6298
rect 20996 6246 20998 6298
rect 20942 6244 20998 6246
rect 21046 6298 21102 6300
rect 21046 6246 21048 6298
rect 21048 6246 21100 6298
rect 21100 6246 21102 6298
rect 21046 6244 21102 6246
rect 20020 5796 20076 5852
rect 19964 5236 20020 5292
rect 19180 4954 19236 4956
rect 19180 4902 19182 4954
rect 19182 4902 19234 4954
rect 19234 4902 19236 4954
rect 19180 4900 19236 4902
rect 19516 4676 19572 4732
rect 19628 4452 19684 4508
rect 19740 4788 19796 4844
rect 18564 4116 18620 4172
rect 18788 4170 18844 4172
rect 18788 4118 18790 4170
rect 18790 4118 18842 4170
rect 18842 4118 18844 4170
rect 18788 4116 18844 4118
rect 17276 2154 17332 2156
rect 17276 2102 17278 2154
rect 17278 2102 17330 2154
rect 17330 2102 17332 2154
rect 17276 2100 17332 2102
rect 16604 1764 16660 1820
rect 16884 1818 16940 1820
rect 16884 1766 16886 1818
rect 16886 1766 16938 1818
rect 16938 1766 16940 1818
rect 16884 1764 16940 1766
rect 17220 1540 17276 1596
rect 18676 2772 18732 2828
rect 20580 5796 20636 5852
rect 20356 4564 20412 4620
rect 19796 3780 19852 3836
rect 19796 3444 19852 3500
rect 19628 2826 19684 2828
rect 19628 2774 19630 2826
rect 19630 2774 19682 2826
rect 19682 2774 19684 2826
rect 19628 2772 19684 2774
rect 19236 2660 19292 2716
rect 19012 2602 19068 2604
rect 19012 2550 19014 2602
rect 19014 2550 19066 2602
rect 19066 2550 19068 2602
rect 19012 2548 19068 2550
rect 18564 2100 18620 2156
rect 19124 2100 19180 2156
rect 18340 1988 18396 2044
rect 19012 1988 19068 2044
rect 18452 1540 18508 1596
rect 17780 1370 17836 1372
rect 17780 1318 17782 1370
rect 17782 1318 17834 1370
rect 17834 1318 17836 1370
rect 17780 1316 17836 1318
rect 18116 1316 18172 1372
rect 20356 4170 20412 4172
rect 20356 4118 20358 4170
rect 20358 4118 20410 4170
rect 20410 4118 20412 4170
rect 20356 4116 20412 4118
rect 20132 3780 20188 3836
rect 20020 2772 20076 2828
rect 19908 2660 19964 2716
rect 19124 1092 19180 1148
rect 19740 1034 19796 1036
rect 19740 982 19742 1034
rect 19742 982 19794 1034
rect 19794 982 19796 1034
rect 19740 980 19796 982
rect 8928 810 8984 812
rect 868 644 924 700
rect 8928 758 8930 810
rect 8930 758 8982 810
rect 8982 758 8984 810
rect 8928 756 8984 758
rect 9032 810 9088 812
rect 9032 758 9034 810
rect 9034 758 9086 810
rect 9086 758 9088 810
rect 9032 756 9088 758
rect 9136 810 9192 812
rect 9136 758 9138 810
rect 9138 758 9190 810
rect 9190 758 9192 810
rect 9136 756 9192 758
rect 16868 810 16924 812
rect 16868 758 16870 810
rect 16870 758 16922 810
rect 16922 758 16924 810
rect 16868 756 16924 758
rect 16972 810 17028 812
rect 16972 758 16974 810
rect 16974 758 17026 810
rect 17026 758 17028 810
rect 16972 756 17028 758
rect 17076 810 17132 812
rect 17076 758 17078 810
rect 17078 758 17130 810
rect 17130 758 17132 810
rect 17076 756 17132 758
rect 22036 6692 22092 6748
rect 23380 7140 23436 7196
rect 25732 9604 25788 9660
rect 27300 11620 27356 11676
rect 27412 11396 27468 11452
rect 27916 12794 27972 12796
rect 27916 12742 27918 12794
rect 27918 12742 27970 12794
rect 27970 12742 27972 12794
rect 27916 12740 27972 12742
rect 28778 12570 28834 12572
rect 28778 12518 28780 12570
rect 28780 12518 28832 12570
rect 28832 12518 28834 12570
rect 28778 12516 28834 12518
rect 28882 12570 28938 12572
rect 28882 12518 28884 12570
rect 28884 12518 28936 12570
rect 28936 12518 28938 12570
rect 28882 12516 28938 12518
rect 28986 12570 29042 12572
rect 28986 12518 28988 12570
rect 28988 12518 29040 12570
rect 29040 12518 29042 12570
rect 28986 12516 29042 12518
rect 30212 13018 30268 13020
rect 30212 12966 30214 13018
rect 30214 12966 30266 13018
rect 30266 12966 30268 13018
rect 30212 12964 30268 12966
rect 30772 12964 30828 13020
rect 31444 12964 31500 13020
rect 32004 13972 32060 14028
rect 28308 12122 28364 12124
rect 28308 12070 28310 12122
rect 28310 12070 28362 12122
rect 28362 12070 28364 12122
rect 28308 12068 28364 12070
rect 28644 12108 28646 12124
rect 28646 12108 28698 12124
rect 28698 12108 28700 12124
rect 28644 12068 28700 12108
rect 29428 12068 29484 12124
rect 30044 12122 30100 12124
rect 30044 12070 30046 12122
rect 30046 12070 30098 12122
rect 30098 12070 30100 12122
rect 30044 12068 30100 12070
rect 31836 12010 31892 12012
rect 31836 11958 31838 12010
rect 31838 11958 31890 12010
rect 31890 11958 31892 12010
rect 31836 11956 31892 11958
rect 32340 11956 32396 12012
rect 32116 11844 32172 11900
rect 28778 11002 28834 11004
rect 28778 10950 28780 11002
rect 28780 10950 28832 11002
rect 28832 10950 28834 11002
rect 28778 10948 28834 10950
rect 28882 11002 28938 11004
rect 28882 10950 28884 11002
rect 28884 10950 28936 11002
rect 28936 10950 28938 11002
rect 28882 10948 28938 10950
rect 28986 11002 29042 11004
rect 28986 10950 28988 11002
rect 28988 10950 29040 11002
rect 29040 10950 29042 11002
rect 28986 10948 29042 10950
rect 26628 10388 26684 10444
rect 27132 10388 27188 10444
rect 26572 9770 26628 9772
rect 26572 9718 26574 9770
rect 26574 9718 26626 9770
rect 26626 9718 26628 9770
rect 26572 9716 26628 9718
rect 26964 9716 27020 9772
rect 26740 9492 26796 9548
rect 25284 8314 25340 8316
rect 25284 8262 25286 8314
rect 25286 8262 25338 8314
rect 25338 8262 25340 8314
rect 25284 8260 25340 8262
rect 25172 8148 25228 8204
rect 25508 8260 25564 8316
rect 26572 8314 26628 8316
rect 26572 8262 26574 8314
rect 26574 8262 26626 8314
rect 26626 8262 26628 8314
rect 26572 8260 26628 8262
rect 27300 9492 27356 9548
rect 28084 10388 28140 10444
rect 27860 9940 27916 9996
rect 32004 9940 32060 9996
rect 27804 9770 27860 9772
rect 27804 9718 27806 9770
rect 27806 9718 27858 9770
rect 27858 9718 27860 9770
rect 27804 9716 27860 9718
rect 27692 9658 27748 9660
rect 27692 9606 27694 9658
rect 27694 9606 27746 9658
rect 27746 9606 27748 9658
rect 27692 9604 27748 9606
rect 28778 9434 28834 9436
rect 28778 9382 28780 9434
rect 28780 9382 28832 9434
rect 28832 9382 28834 9434
rect 28778 9380 28834 9382
rect 28882 9434 28938 9436
rect 28882 9382 28884 9434
rect 28884 9382 28936 9434
rect 28936 9382 28938 9434
rect 28882 9380 28938 9382
rect 28986 9434 29042 9436
rect 28986 9382 28988 9434
rect 28988 9382 29040 9434
rect 29040 9382 29042 9434
rect 28986 9380 29042 9382
rect 31836 8874 31892 8876
rect 31836 8822 31838 8874
rect 31838 8822 31890 8874
rect 31890 8822 31892 8874
rect 31836 8820 31892 8822
rect 32228 10276 32284 10332
rect 26068 8148 26124 8204
rect 25116 7588 25172 7644
rect 28778 7866 28834 7868
rect 28778 7814 28780 7866
rect 28780 7814 28832 7866
rect 28832 7814 28834 7866
rect 28778 7812 28834 7814
rect 28882 7866 28938 7868
rect 28882 7814 28884 7866
rect 28884 7814 28936 7866
rect 28936 7814 28938 7866
rect 28882 7812 28938 7814
rect 28986 7866 29042 7868
rect 28986 7814 28988 7866
rect 28988 7814 29040 7866
rect 29040 7814 29042 7866
rect 28986 7812 29042 7814
rect 22820 6692 22876 6748
rect 22148 6580 22204 6636
rect 22596 6580 22652 6636
rect 21364 5178 21420 5180
rect 21364 5126 21366 5178
rect 21366 5126 21418 5178
rect 21418 5126 21420 5178
rect 21364 5124 21420 5126
rect 20838 4730 20894 4732
rect 20838 4678 20840 4730
rect 20840 4678 20892 4730
rect 20892 4678 20894 4730
rect 20838 4676 20894 4678
rect 20942 4730 20998 4732
rect 20942 4678 20944 4730
rect 20944 4678 20996 4730
rect 20996 4678 20998 4730
rect 20942 4676 20998 4678
rect 21046 4730 21102 4732
rect 21046 4678 21048 4730
rect 21048 4678 21100 4730
rect 21100 4678 21102 4730
rect 21046 4676 21102 4678
rect 21196 4564 21252 4620
rect 20580 4452 20636 4508
rect 20692 4350 20748 4396
rect 20692 4340 20694 4350
rect 20694 4340 20746 4350
rect 20746 4340 20748 4350
rect 22092 4788 22148 4844
rect 20580 2778 20636 2828
rect 20580 2772 20582 2778
rect 20582 2772 20634 2778
rect 20634 2772 20636 2778
rect 20356 2324 20412 2380
rect 22260 4170 22316 4172
rect 22260 4118 22262 4170
rect 22262 4118 22314 4170
rect 22314 4118 22316 4170
rect 22260 4116 22316 4118
rect 20916 3498 20972 3500
rect 20916 3446 20918 3498
rect 20918 3446 20970 3498
rect 20970 3446 20972 3498
rect 20916 3444 20972 3446
rect 20838 3162 20894 3164
rect 20838 3110 20840 3162
rect 20840 3110 20892 3162
rect 20892 3110 20894 3162
rect 20838 3108 20894 3110
rect 20942 3162 20998 3164
rect 20942 3110 20944 3162
rect 20944 3110 20996 3162
rect 20996 3110 20998 3162
rect 20942 3108 20998 3110
rect 21046 3162 21102 3164
rect 21046 3110 21048 3162
rect 21048 3110 21100 3162
rect 21100 3110 21102 3162
rect 21046 3108 21102 3110
rect 21812 3220 21868 3276
rect 21252 2548 21308 2604
rect 20692 2324 20748 2380
rect 20838 1594 20894 1596
rect 20838 1542 20840 1594
rect 20840 1542 20892 1594
rect 20892 1542 20894 1594
rect 20838 1540 20894 1542
rect 20942 1594 20998 1596
rect 20942 1542 20944 1594
rect 20944 1542 20996 1594
rect 20996 1542 20998 1594
rect 20942 1540 20998 1542
rect 21046 1594 21102 1596
rect 21046 1542 21048 1594
rect 21048 1542 21100 1594
rect 21100 1542 21102 1594
rect 21046 1540 21102 1542
rect 22708 6468 22764 6524
rect 23828 6580 23884 6636
rect 23436 5236 23492 5292
rect 23044 5178 23100 5180
rect 23044 5126 23046 5178
rect 23046 5126 23098 5178
rect 23098 5126 23100 5178
rect 23044 5124 23100 5126
rect 25396 7140 25452 7196
rect 24808 7082 24864 7084
rect 24808 7030 24810 7082
rect 24810 7030 24862 7082
rect 24862 7030 24864 7082
rect 24808 7028 24864 7030
rect 24912 7082 24968 7084
rect 24912 7030 24914 7082
rect 24914 7030 24966 7082
rect 24966 7030 24968 7082
rect 24912 7028 24968 7030
rect 25016 7082 25072 7084
rect 25016 7030 25018 7082
rect 25018 7030 25070 7082
rect 25070 7030 25072 7082
rect 25016 7028 25072 7030
rect 24332 6858 24388 6860
rect 24332 6806 24334 6858
rect 24334 6806 24386 6858
rect 24386 6806 24388 6858
rect 24332 6804 24388 6806
rect 24108 6746 24164 6748
rect 24108 6694 24110 6746
rect 24110 6694 24162 6746
rect 24162 6694 24164 6746
rect 24108 6692 24164 6694
rect 24556 6580 24612 6636
rect 23940 6244 23996 6300
rect 23940 5796 23996 5852
rect 26180 6584 26236 6636
rect 26180 6580 26182 6584
rect 26182 6580 26234 6584
rect 26234 6580 26236 6584
rect 25284 6356 25340 6412
rect 26292 6356 26348 6412
rect 25676 6244 25732 6300
rect 25060 5842 25062 5852
rect 25062 5842 25114 5852
rect 25114 5842 25116 5852
rect 25060 5796 25116 5842
rect 24052 5572 24108 5628
rect 23828 5236 23884 5292
rect 24808 5514 24864 5516
rect 24808 5462 24810 5514
rect 24810 5462 24862 5514
rect 24862 5462 24864 5514
rect 24808 5460 24864 5462
rect 24912 5514 24968 5516
rect 24912 5462 24914 5514
rect 24914 5462 24966 5514
rect 24966 5462 24968 5514
rect 24912 5460 24968 5462
rect 25016 5514 25072 5516
rect 25016 5462 25018 5514
rect 25018 5462 25070 5514
rect 25070 5462 25072 5514
rect 25016 5460 25072 5462
rect 25844 5850 25900 5852
rect 25844 5798 25846 5850
rect 25846 5798 25898 5850
rect 25898 5798 25900 5850
rect 25844 5796 25900 5798
rect 24388 4954 24444 4956
rect 24388 4902 24390 4954
rect 24390 4902 24442 4954
rect 24442 4902 24444 4954
rect 24388 4900 24444 4902
rect 24612 4900 24668 4956
rect 23772 4676 23828 4732
rect 24724 4452 24780 4508
rect 26068 6244 26124 6300
rect 26964 6626 26966 6636
rect 26966 6626 27018 6636
rect 27018 6626 27020 6636
rect 26964 6580 27020 6626
rect 26628 6522 26684 6524
rect 26628 6470 26630 6522
rect 26630 6470 26682 6522
rect 26682 6470 26684 6522
rect 26628 6468 26684 6470
rect 28778 6298 28834 6300
rect 28778 6246 28780 6298
rect 28780 6246 28832 6298
rect 28832 6246 28834 6298
rect 28778 6244 28834 6246
rect 28882 6298 28938 6300
rect 28882 6246 28884 6298
rect 28884 6246 28936 6298
rect 28936 6246 28938 6298
rect 28882 6244 28938 6246
rect 28986 6298 29042 6300
rect 28986 6246 28988 6298
rect 28988 6246 29040 6298
rect 29040 6246 29042 6298
rect 28986 6244 29042 6246
rect 25284 4954 25340 4956
rect 25284 4902 25286 4954
rect 25286 4902 25338 4954
rect 25338 4902 25340 4954
rect 25284 4900 25340 4902
rect 25620 4788 25676 4844
rect 25508 4452 25564 4508
rect 25396 4170 25452 4172
rect 25396 4118 25398 4170
rect 25398 4118 25450 4170
rect 25450 4118 25452 4170
rect 25396 4116 25452 4118
rect 25172 4004 25228 4060
rect 24808 3946 24864 3948
rect 24808 3894 24810 3946
rect 24810 3894 24862 3946
rect 24862 3894 24864 3946
rect 24808 3892 24864 3894
rect 24912 3946 24968 3948
rect 24912 3894 24914 3946
rect 24914 3894 24966 3946
rect 24966 3894 24968 3946
rect 24912 3892 24968 3894
rect 25016 3946 25072 3948
rect 25016 3894 25018 3946
rect 25018 3894 25070 3946
rect 25070 3894 25072 3946
rect 25016 3892 25072 3894
rect 23268 2212 23324 2268
rect 23100 2042 23156 2044
rect 22372 1876 22428 1932
rect 23100 1990 23102 2042
rect 23102 1990 23154 2042
rect 23154 1990 23156 2042
rect 23100 1988 23156 1990
rect 21476 1652 21532 1708
rect 22372 1652 22428 1708
rect 21756 1428 21812 1484
rect 21924 1256 21926 1260
rect 21926 1256 21978 1260
rect 21978 1256 21980 1260
rect 21924 1204 21980 1256
rect 23380 1926 23382 1932
rect 23382 1926 23434 1932
rect 23434 1926 23436 1932
rect 23380 1876 23436 1926
rect 23268 1652 23324 1708
rect 22596 1428 22652 1484
rect 22484 1316 22540 1372
rect 22708 1214 22764 1260
rect 22708 1204 22710 1214
rect 22710 1204 22762 1214
rect 22762 1204 22764 1214
rect 24724 3386 24780 3388
rect 24724 3334 24726 3386
rect 24726 3334 24778 3386
rect 24778 3334 24780 3386
rect 24724 3332 24780 3334
rect 24836 2938 24892 2940
rect 24836 2886 24838 2938
rect 24838 2886 24890 2938
rect 24890 2886 24892 2938
rect 24836 2884 24892 2886
rect 24164 2602 24220 2604
rect 24164 2550 24166 2602
rect 24166 2550 24218 2602
rect 24218 2550 24220 2602
rect 24164 2548 24220 2550
rect 25060 2602 25116 2604
rect 25060 2550 25062 2602
rect 25062 2550 25114 2602
rect 25114 2550 25116 2602
rect 25060 2548 25116 2550
rect 24332 2436 24388 2492
rect 31892 4900 31948 4956
rect 26404 4676 26460 4732
rect 28778 4730 28834 4732
rect 28778 4678 28780 4730
rect 28780 4678 28832 4730
rect 28832 4678 28834 4730
rect 28778 4676 28834 4678
rect 28882 4730 28938 4732
rect 28882 4678 28884 4730
rect 28884 4678 28936 4730
rect 28936 4678 28938 4730
rect 28882 4676 28938 4678
rect 28986 4730 29042 4732
rect 28986 4678 28988 4730
rect 28988 4678 29040 4730
rect 29040 4678 29042 4730
rect 28986 4676 29042 4678
rect 26012 4004 26068 4060
rect 25844 3332 25900 3388
rect 28778 3162 28834 3164
rect 28778 3110 28780 3162
rect 28780 3110 28832 3162
rect 28832 3110 28834 3162
rect 28778 3108 28834 3110
rect 28882 3162 28938 3164
rect 28882 3110 28884 3162
rect 28884 3110 28936 3162
rect 28936 3110 28938 3162
rect 28882 3108 28938 3110
rect 28986 3162 29042 3164
rect 28986 3110 28988 3162
rect 28988 3110 29040 3162
rect 29040 3110 29042 3162
rect 28986 3108 29042 3110
rect 25620 2884 25676 2940
rect 25172 2436 25228 2492
rect 24808 2378 24864 2380
rect 24808 2326 24810 2378
rect 24810 2326 24862 2378
rect 24862 2326 24864 2378
rect 24808 2324 24864 2326
rect 24912 2378 24968 2380
rect 24912 2326 24914 2378
rect 24914 2326 24966 2378
rect 24966 2326 24968 2378
rect 24912 2324 24968 2326
rect 25016 2378 25072 2380
rect 25016 2326 25018 2378
rect 25018 2326 25070 2378
rect 25070 2326 25072 2378
rect 25016 2324 25072 2326
rect 25676 2436 25732 2492
rect 25396 2212 25452 2268
rect 25620 2100 25676 2156
rect 23772 2042 23828 2044
rect 23772 1990 23774 2042
rect 23774 1990 23826 2042
rect 23826 1990 23828 2042
rect 23772 1988 23828 1990
rect 24052 1926 24054 1932
rect 24054 1926 24106 1932
rect 24106 1926 24108 1932
rect 24052 1876 24108 1926
rect 23940 1652 23996 1708
rect 32340 8820 32396 8876
rect 32452 8260 32508 8316
rect 32340 4900 32396 4956
rect 31836 1652 31892 1708
rect 32340 1652 32396 1708
rect 28778 1594 28834 1596
rect 28778 1542 28780 1594
rect 28780 1542 28832 1594
rect 28832 1542 28834 1594
rect 28778 1540 28834 1542
rect 28882 1594 28938 1596
rect 28882 1542 28884 1594
rect 28884 1542 28936 1594
rect 28936 1542 28938 1594
rect 28882 1540 28938 1542
rect 28986 1594 29042 1596
rect 28986 1542 28988 1594
rect 28988 1542 29040 1594
rect 29040 1542 29042 1594
rect 28986 1540 29042 1542
rect 22036 1142 22038 1148
rect 22038 1142 22090 1148
rect 22090 1142 22092 1148
rect 22036 1092 22092 1142
rect 25508 980 25564 1036
rect 24808 810 24864 812
rect 24808 758 24810 810
rect 24810 758 24862 810
rect 24862 758 24864 810
rect 24808 756 24864 758
rect 24912 810 24968 812
rect 24912 758 24914 810
rect 24914 758 24966 810
rect 24966 758 24968 810
rect 24912 756 24968 758
rect 25016 810 25072 812
rect 25016 758 25018 810
rect 25018 758 25070 810
rect 25070 758 25072 810
rect 25956 980 26012 1036
rect 26236 1034 26292 1036
rect 26236 982 26238 1034
rect 26238 982 26290 1034
rect 26290 982 26292 1034
rect 26236 980 26292 982
rect 25016 756 25072 758
<< metal3 >>
rect 0 19292 800 19320
rect 0 19236 1484 19292
rect 0 19208 800 19236
rect 1428 19068 1484 19236
rect 1418 19012 1428 19068
rect 1484 19012 1494 19068
rect 15978 18900 15988 18956
rect 16044 18900 21868 18956
rect 21924 18900 26740 18956
rect 26796 18900 26806 18956
rect 4948 18788 4958 18844
rect 5014 18788 5062 18844
rect 5118 18788 5166 18844
rect 5222 18788 5232 18844
rect 12888 18788 12898 18844
rect 12954 18788 13002 18844
rect 13058 18788 13106 18844
rect 13162 18788 13172 18844
rect 20828 18788 20838 18844
rect 20894 18788 20942 18844
rect 20998 18788 21046 18844
rect 21102 18788 21112 18844
rect 28768 18788 28778 18844
rect 28834 18788 28882 18844
rect 28938 18788 28986 18844
rect 29042 18788 29052 18844
rect 11162 18676 11172 18732
rect 11228 18676 15652 18732
rect 15708 18676 15718 18732
rect 16538 18676 16548 18732
rect 16604 18676 25788 18732
rect 25844 18676 29092 18732
rect 29148 18676 29158 18732
rect 1866 18564 1876 18620
rect 1932 18564 9996 18620
rect 10052 18564 10062 18620
rect 11330 18564 11340 18620
rect 11396 18564 18004 18620
rect 18060 18564 18070 18620
rect 19226 18564 19236 18620
rect 19292 18564 23100 18620
rect 23156 18564 23166 18620
rect 1194 18452 1204 18508
rect 1260 18452 1540 18508
rect 1596 18452 3388 18508
rect 3444 18452 3454 18508
rect 10154 18452 10164 18508
rect 10220 18452 15820 18508
rect 15876 18452 15886 18508
rect 19450 18452 19460 18508
rect 19516 18452 21140 18508
rect 21196 18452 21206 18508
rect 22586 18452 22596 18508
rect 22652 18452 23996 18508
rect 24052 18452 24062 18508
rect 27178 18452 27188 18508
rect 27244 18452 28140 18508
rect 28196 18452 28206 18508
rect 29978 18452 29988 18508
rect 30044 18452 30548 18508
rect 30604 18452 30716 18508
rect 30772 18452 30782 18508
rect 21140 18396 21196 18452
rect 1418 18340 1428 18396
rect 1484 18340 2940 18396
rect 2996 18340 3006 18396
rect 3882 18340 3892 18396
rect 3948 18340 4508 18396
rect 4564 18340 4574 18396
rect 11722 18340 11732 18396
rect 11788 18340 12516 18396
rect 12572 18340 12582 18396
rect 13262 18340 13300 18396
rect 13356 18340 13366 18396
rect 14186 18340 14196 18396
rect 14252 18340 15316 18396
rect 15372 18340 15382 18396
rect 16426 18340 16436 18396
rect 16492 18340 16502 18396
rect 16594 18340 16604 18396
rect 16660 18340 18228 18396
rect 18284 18340 18294 18396
rect 18442 18340 18452 18396
rect 18508 18340 18620 18396
rect 18676 18340 18686 18396
rect 21140 18340 23772 18396
rect 23828 18340 23838 18396
rect 26618 18340 26628 18396
rect 26684 18340 27636 18396
rect 27692 18340 28756 18396
rect 28812 18340 28822 18396
rect 16436 18284 16492 18340
rect 33200 18284 34000 18312
rect 1642 18228 1652 18284
rect 1708 18228 2716 18284
rect 2772 18228 2782 18284
rect 4302 18228 4340 18284
rect 4396 18228 4406 18284
rect 6290 18228 6300 18284
rect 6356 18228 9044 18284
rect 9100 18228 9268 18284
rect 9324 18228 9334 18284
rect 10154 18228 10164 18284
rect 10220 18228 10612 18284
rect 10668 18228 10678 18284
rect 10770 18228 10780 18284
rect 10836 18228 15092 18284
rect 15148 18228 15158 18284
rect 16202 18228 16212 18284
rect 16268 18228 18284 18284
rect 20010 18228 20020 18284
rect 20076 18228 22988 18284
rect 23044 18228 23054 18284
rect 25890 18228 25900 18284
rect 25956 18228 27188 18284
rect 27244 18228 27254 18284
rect 29474 18228 29484 18284
rect 29540 18228 30100 18284
rect 30156 18228 30166 18284
rect 31770 18228 31780 18284
rect 31836 18228 32116 18284
rect 32172 18228 34000 18284
rect 2510 18116 2548 18172
rect 2604 18116 2614 18172
rect 4106 18116 4116 18172
rect 4172 18116 10948 18172
rect 11004 18116 11014 18172
rect 11162 18116 11172 18172
rect 11228 18116 12404 18172
rect 12460 18116 14420 18172
rect 14476 18116 16436 18172
rect 16492 18116 16502 18172
rect 16660 18116 18004 18172
rect 18060 18116 18070 18172
rect 0 18060 800 18088
rect 16660 18060 16716 18116
rect 18228 18060 18284 18228
rect 33200 18200 34000 18228
rect 19898 18116 19908 18172
rect 19964 18116 22260 18172
rect 22316 18116 22326 18172
rect 0 18004 2100 18060
rect 2156 18004 3164 18060
rect 3220 18004 3230 18060
rect 8918 18004 8928 18060
rect 8984 18004 9032 18060
rect 9088 18004 9136 18060
rect 9192 18004 9202 18060
rect 10602 18004 10612 18060
rect 10668 18004 16324 18060
rect 16380 18004 16716 18060
rect 16858 18004 16868 18060
rect 16924 18004 16972 18060
rect 17028 18004 17076 18060
rect 17132 18004 17142 18060
rect 18228 18004 22036 18060
rect 22092 18004 22102 18060
rect 24798 18004 24808 18060
rect 24864 18004 24912 18060
rect 24968 18004 25016 18060
rect 25072 18004 25082 18060
rect 0 17976 800 18004
rect 2650 17780 2660 17836
rect 2716 17780 3724 17836
rect 3780 17780 3790 17836
rect 5842 17780 5852 17836
rect 5908 17780 7140 17836
rect 7196 17780 7206 17836
rect 8698 17780 8708 17836
rect 8764 17780 10052 17836
rect 10108 17780 10118 17836
rect 11778 17780 11788 17836
rect 11844 17780 14028 17836
rect 14084 17724 14140 17836
rect 14858 17780 14868 17836
rect 14924 17780 15428 17836
rect 15484 17780 15494 17836
rect 19506 17780 19516 17836
rect 19572 17780 19740 17836
rect 19796 17780 21364 17836
rect 21420 17780 21430 17836
rect 23202 17780 23212 17836
rect 23268 17780 26124 17836
rect 26180 17780 26190 17836
rect 31891 17780 32004 17836
rect 32060 17780 32070 17836
rect 31891 17724 31947 17780
rect 2548 17668 6804 17724
rect 6860 17668 6870 17724
rect 7914 17668 7924 17724
rect 7980 17668 9492 17724
rect 9548 17668 9558 17724
rect 14084 17668 14980 17724
rect 15036 17668 15046 17724
rect 15866 17668 15876 17724
rect 15932 17668 16100 17724
rect 16156 17668 16166 17724
rect 18386 17668 18396 17724
rect 18452 17668 31947 17724
rect 2548 17612 2604 17668
rect 2538 17556 2548 17612
rect 2604 17556 2614 17612
rect 3714 17556 3724 17612
rect 3836 17556 3846 17612
rect 6402 17556 6412 17612
rect 6468 17556 7252 17612
rect 7308 17556 7318 17612
rect 8362 17556 8372 17612
rect 8428 17556 8932 17612
rect 8988 17556 10388 17612
rect 10444 17556 10454 17612
rect 10602 17556 10612 17612
rect 10668 17556 10678 17612
rect 10770 17556 10780 17612
rect 10836 17556 11508 17612
rect 11564 17556 11574 17612
rect 18778 17556 18788 17612
rect 18844 17556 20916 17612
rect 20972 17556 20982 17612
rect 24714 17556 24724 17612
rect 24780 17556 25284 17612
rect 25340 17556 25350 17612
rect 28018 17556 28028 17612
rect 28084 17556 29932 17612
rect 29988 17556 31220 17612
rect 31276 17556 31286 17612
rect 1866 17444 1876 17500
rect 1932 17444 3388 17500
rect 3444 17444 3454 17500
rect 5954 17444 5964 17500
rect 6020 17444 6692 17500
rect 6748 17444 6758 17500
rect 9828 17388 9884 17556
rect 10612 17388 10668 17556
rect 11050 17444 11060 17500
rect 11116 17444 12852 17500
rect 12908 17444 12918 17500
rect 15082 17444 15092 17500
rect 15148 17444 16212 17500
rect 16268 17444 16278 17500
rect 17770 17444 17780 17500
rect 17836 17444 19236 17500
rect 19292 17444 19302 17500
rect 30762 17444 30772 17500
rect 30828 17444 31332 17500
rect 31388 17444 31398 17500
rect 9818 17332 9828 17388
rect 9884 17332 9894 17388
rect 10612 17332 15147 17388
rect 15091 17276 15147 17332
rect 4948 17220 4958 17276
rect 5014 17220 5062 17276
rect 5118 17220 5166 17276
rect 5222 17220 5232 17276
rect 6290 17220 6300 17276
rect 6356 17220 6916 17276
rect 6972 17220 8596 17276
rect 8652 17220 8662 17276
rect 12888 17220 12898 17276
rect 12954 17220 13002 17276
rect 13058 17220 13106 17276
rect 13162 17220 13172 17276
rect 15091 17220 17836 17276
rect 17892 17220 17902 17276
rect 20828 17220 20838 17276
rect 20894 17220 20942 17276
rect 20998 17220 21046 17276
rect 21102 17220 21112 17276
rect 28768 17220 28778 17276
rect 28834 17220 28882 17276
rect 28938 17220 28986 17276
rect 29042 17220 29052 17276
rect 8082 17108 8092 17164
rect 8148 17108 9436 17164
rect 9492 17108 10724 17164
rect 10780 17108 10790 17164
rect 3490 16996 3500 17052
rect 3556 16996 4788 17052
rect 4844 16996 4854 17052
rect 6318 16996 6356 17052
rect 6412 16996 6422 17052
rect 11610 16996 11620 17052
rect 11676 16996 12292 17052
rect 12348 16996 12358 17052
rect 16762 16996 16772 17052
rect 16828 16996 21980 17052
rect 22036 16996 22046 17052
rect 1530 16884 1540 16940
rect 1596 16884 1606 16940
rect 10602 16884 10612 16940
rect 10668 16884 11284 16940
rect 11340 16884 13300 16940
rect 13356 16884 13366 16940
rect 14130 16884 14140 16940
rect 14196 16884 17220 16940
rect 17276 16884 17286 16940
rect 17994 16884 18004 16940
rect 18060 16884 18116 16940
rect 18172 16884 18182 16940
rect 23594 16884 23604 16940
rect 23660 16884 26292 16940
rect 26348 16884 26358 16940
rect 0 16828 800 16856
rect 1540 16828 1596 16884
rect 0 16772 1596 16828
rect 11386 16772 11396 16828
rect 11452 16772 11956 16828
rect 12012 16772 12022 16828
rect 14980 16772 15428 16828
rect 15484 16772 15494 16828
rect 20010 16772 20020 16828
rect 20076 16772 21308 16828
rect 0 16744 800 16772
rect 14980 16716 15036 16772
rect 1418 16660 1428 16716
rect 1484 16660 2044 16716
rect 2100 16660 2110 16716
rect 3154 16660 3164 16716
rect 3220 16660 3724 16716
rect 3780 16660 4900 16716
rect 4956 16660 4966 16716
rect 11610 16660 11620 16716
rect 11676 16660 12740 16716
rect 12796 16660 12806 16716
rect 12898 16660 12908 16716
rect 12964 16660 15036 16716
rect 16538 16660 16548 16716
rect 16604 16660 16772 16716
rect 16828 16660 16838 16716
rect 17546 16660 17556 16716
rect 17612 16660 18564 16716
rect 18620 16660 18630 16716
rect 19124 16660 20524 16716
rect 20580 16660 20590 16716
rect 21252 16660 21308 16772
rect 21476 16772 22260 16828
rect 22316 16772 22326 16828
rect 29530 16772 29540 16828
rect 29596 16772 31500 16828
rect 31556 16772 31566 16828
rect 21364 16660 21374 16716
rect 19124 16604 19180 16660
rect 21476 16604 21532 16772
rect 23874 16660 23884 16716
rect 23940 16660 24388 16716
rect 24444 16660 25788 16716
rect 25844 16660 25854 16716
rect 27234 16660 27244 16716
rect 27300 16660 27692 16716
rect 27748 16660 31220 16716
rect 31276 16660 31286 16716
rect 12394 16548 12404 16604
rect 12460 16548 14868 16604
rect 14924 16548 14934 16604
rect 16660 16548 19180 16604
rect 19282 16548 19292 16604
rect 19348 16548 20412 16604
rect 20468 16548 21532 16604
rect 22586 16548 22596 16604
rect 22652 16548 24052 16604
rect 24108 16548 24612 16604
rect 24668 16548 24678 16604
rect 16660 16492 16716 16548
rect 8918 16436 8928 16492
rect 8984 16436 9032 16492
rect 9088 16436 9136 16492
rect 9192 16436 9202 16492
rect 10098 16436 10108 16492
rect 10164 16436 13300 16492
rect 13356 16436 13366 16492
rect 15091 16436 16716 16492
rect 16858 16436 16868 16492
rect 16924 16436 16972 16492
rect 17028 16436 17076 16492
rect 17132 16436 17142 16492
rect 19450 16436 19460 16492
rect 19516 16436 21756 16492
rect 21812 16436 21822 16492
rect 24798 16436 24808 16492
rect 24864 16436 24912 16492
rect 24968 16436 25016 16492
rect 25072 16436 25082 16492
rect 25722 16436 25732 16492
rect 25788 16436 26852 16492
rect 26908 16436 28476 16492
rect 28532 16436 28542 16492
rect 15091 16380 15147 16436
rect 8474 16324 8484 16380
rect 8540 16324 13748 16380
rect 13804 16324 14140 16380
rect 14196 16324 14206 16380
rect 14308 16324 15147 16380
rect 15204 16324 17780 16380
rect 17836 16324 17846 16380
rect 18610 16324 18620 16380
rect 18676 16324 19292 16380
rect 19348 16324 19358 16380
rect 20626 16324 20636 16380
rect 20692 16324 22260 16380
rect 22316 16324 22652 16380
rect 22708 16324 22718 16380
rect 14308 16268 14364 16324
rect 15204 16268 15260 16324
rect 17780 16268 17836 16324
rect 6626 16212 6636 16268
rect 6692 16212 8764 16268
rect 10042 16212 10052 16268
rect 10108 16212 11004 16268
rect 11060 16212 11070 16268
rect 11162 16212 11172 16268
rect 11228 16212 11266 16268
rect 12114 16212 12124 16268
rect 12180 16212 12572 16268
rect 12628 16212 12638 16268
rect 12730 16212 12740 16268
rect 12796 16212 14364 16268
rect 14746 16212 14756 16268
rect 14812 16212 15260 16268
rect 15418 16212 15428 16268
rect 15484 16212 15820 16268
rect 15876 16212 15886 16268
rect 17780 16212 18620 16268
rect 18778 16212 18788 16268
rect 18844 16212 19908 16268
rect 19964 16212 21028 16268
rect 21084 16212 21094 16268
rect 21802 16212 21812 16268
rect 21868 16212 22260 16268
rect 22316 16212 22326 16268
rect 22782 16212 22820 16268
rect 22876 16212 22886 16268
rect 23370 16212 23380 16268
rect 23436 16212 25172 16268
rect 25228 16212 25238 16268
rect 26114 16212 26124 16268
rect 26180 16212 26964 16268
rect 27020 16212 27030 16268
rect 2538 16100 2548 16156
rect 2604 16100 8484 16156
rect 8540 16100 8550 16156
rect 8708 16044 8764 16212
rect 11172 16156 11228 16212
rect 14756 16156 14812 16212
rect 18564 16156 18620 16212
rect 8866 16100 8876 16156
rect 8932 16100 11228 16156
rect 11582 16100 11620 16156
rect 11676 16100 11686 16156
rect 11778 16100 11788 16156
rect 11844 16100 14812 16156
rect 14970 16100 14980 16156
rect 15036 16100 15932 16156
rect 15988 16100 15998 16156
rect 16772 16100 17612 16156
rect 17668 16100 17892 16156
rect 17948 16100 17958 16156
rect 18302 16100 18340 16156
rect 18396 16100 18406 16156
rect 18564 16100 21532 16156
rect 21588 16100 21598 16156
rect 23706 16100 23716 16156
rect 23828 16100 24612 16156
rect 24668 16100 25956 16156
rect 26012 16100 26404 16156
rect 26460 16100 26470 16156
rect 26730 16100 26740 16156
rect 26796 16100 30772 16156
rect 30828 16100 30838 16156
rect 16772 16044 16828 16100
rect 8708 15988 9100 16044
rect 11386 15988 11396 16044
rect 11452 15988 16548 16044
rect 16604 15988 16614 16044
rect 16762 15988 16772 16044
rect 16828 15988 16838 16044
rect 17994 15988 18004 16044
rect 18060 15988 26068 16044
rect 26124 15988 26134 16044
rect 30538 15988 30548 16044
rect 30604 15988 31332 16044
rect 31388 15988 31398 16044
rect 9044 15932 9100 15988
rect 7578 15876 7588 15932
rect 7644 15876 8876 15932
rect 8932 15876 8942 15932
rect 9044 15876 23380 15932
rect 23436 15876 23446 15932
rect 24602 15876 24612 15932
rect 24668 15876 24780 15932
rect 24836 15876 25396 15932
rect 25452 15876 25462 15932
rect 28298 15876 28308 15932
rect 28364 15876 28868 15932
rect 28924 15876 28934 15932
rect 2258 15764 2268 15820
rect 2324 15764 14140 15820
rect 15082 15764 15092 15820
rect 15148 15764 15428 15820
rect 15484 15764 16212 15820
rect 16268 15764 16278 15820
rect 16762 15764 16772 15820
rect 16828 15764 17388 15820
rect 17444 15764 17454 15820
rect 17546 15764 17556 15820
rect 17612 15764 17650 15820
rect 18722 15764 18732 15820
rect 18788 15764 22820 15820
rect 22876 15764 22886 15820
rect 23258 15764 23268 15820
rect 23324 15764 29316 15820
rect 29372 15764 29382 15820
rect 14084 15708 14140 15764
rect 4948 15652 4958 15708
rect 5014 15652 5062 15708
rect 5118 15652 5166 15708
rect 5222 15652 5232 15708
rect 7354 15652 7364 15708
rect 7420 15652 12628 15708
rect 12684 15652 12694 15708
rect 12888 15652 12898 15708
rect 12954 15652 13002 15708
rect 13058 15652 13106 15708
rect 13162 15652 13172 15708
rect 14084 15652 19796 15708
rect 19852 15652 19862 15708
rect 20828 15652 20838 15708
rect 20894 15652 20942 15708
rect 20998 15652 21046 15708
rect 21102 15652 21112 15708
rect 21252 15652 22484 15708
rect 22540 15652 22550 15708
rect 23146 15652 23156 15708
rect 23212 15652 23222 15708
rect 28768 15652 28778 15708
rect 28834 15652 28882 15708
rect 28938 15652 28986 15708
rect 29042 15652 29052 15708
rect 0 15596 800 15624
rect 0 15540 1540 15596
rect 1596 15540 1606 15596
rect 7130 15540 7140 15596
rect 7196 15540 13748 15596
rect 13804 15540 13814 15596
rect 14634 15540 14644 15596
rect 14700 15540 15652 15596
rect 15708 15540 15718 15596
rect 16202 15540 16212 15596
rect 16268 15540 16996 15596
rect 17052 15540 17062 15596
rect 18554 15540 18564 15596
rect 18676 15540 18686 15596
rect 18946 15540 18956 15596
rect 19012 15540 19572 15596
rect 19628 15540 19638 15596
rect 20570 15540 20580 15596
rect 20636 15540 21196 15596
rect 21252 15540 21308 15652
rect 23156 15596 23212 15652
rect 21466 15540 21476 15596
rect 21588 15540 21598 15596
rect 22362 15540 22372 15596
rect 22428 15540 23212 15596
rect 0 15512 800 15540
rect 6458 15428 6468 15484
rect 6524 15428 8708 15484
rect 8764 15428 8774 15484
rect 12478 15428 12516 15484
rect 12572 15428 12582 15484
rect 14354 15428 14364 15484
rect 14420 15428 14924 15484
rect 16062 15428 16100 15484
rect 16156 15428 16166 15484
rect 16314 15428 16324 15484
rect 16380 15428 21700 15484
rect 21756 15428 21766 15484
rect 23006 15428 23044 15484
rect 23100 15428 23110 15484
rect 24490 15428 24500 15484
rect 24556 15428 24612 15484
rect 24668 15428 24678 15484
rect 25386 15428 25396 15484
rect 25452 15428 26796 15484
rect 28746 15428 28756 15484
rect 28812 15428 30772 15484
rect 30828 15428 30838 15484
rect 14868 15372 14924 15428
rect 2874 15316 2884 15372
rect 2940 15316 3220 15372
rect 3276 15316 5516 15372
rect 5572 15316 5582 15372
rect 6906 15316 6916 15372
rect 6972 15316 8596 15372
rect 8652 15316 8662 15372
rect 14578 15316 14588 15372
rect 14700 15316 14710 15372
rect 14868 15316 15204 15372
rect 15260 15316 15316 15372
rect 15372 15316 15382 15372
rect 18106 15316 18116 15372
rect 18172 15316 21364 15372
rect 21420 15316 21430 15372
rect 22754 15316 22764 15372
rect 22820 15316 25116 15372
rect 25172 15316 25182 15372
rect 3098 15204 3108 15260
rect 3164 15204 4060 15260
rect 4116 15204 6132 15260
rect 6188 15204 6198 15260
rect 7522 15204 7532 15260
rect 7588 15204 7924 15260
rect 7980 15204 10612 15260
rect 10668 15204 10678 15260
rect 11050 15204 11060 15260
rect 11116 15204 12068 15260
rect 12124 15204 12134 15260
rect 13794 15204 13804 15260
rect 13860 15204 15428 15260
rect 15484 15204 15494 15260
rect 15642 15204 15652 15260
rect 15708 15204 17836 15260
rect 18554 15204 18564 15260
rect 18620 15204 18676 15260
rect 18732 15204 18742 15260
rect 21242 15204 21252 15260
rect 21308 15204 22036 15260
rect 22092 15204 22102 15260
rect 23491 15204 24892 15260
rect 24948 15204 26012 15260
rect 26068 15204 26180 15260
rect 17780 15148 17836 15204
rect 23491 15148 23547 15204
rect 2090 15092 2100 15148
rect 2156 15092 5404 15148
rect 5460 15092 5470 15148
rect 8082 15092 8092 15148
rect 8148 15092 9436 15148
rect 9492 15092 9502 15148
rect 12226 15092 12236 15148
rect 12292 15092 13412 15148
rect 13468 15092 13478 15148
rect 13626 15092 13636 15148
rect 13692 15092 15204 15148
rect 15260 15092 15270 15148
rect 16090 15092 16100 15148
rect 16156 15092 17220 15148
rect 17276 15092 17612 15148
rect 17668 15092 17678 15148
rect 17780 15092 19572 15148
rect 19628 15092 19638 15148
rect 19786 15092 19796 15148
rect 19852 15092 21532 15148
rect 21588 15092 23436 15148
rect 23492 15092 23547 15148
rect 24378 15092 24388 15148
rect 24444 15092 25620 15148
rect 25676 15092 25686 15148
rect 16324 15036 16380 15092
rect 10938 14980 10948 15036
rect 11004 14980 11396 15036
rect 11452 14980 11462 15036
rect 11722 14980 11732 15036
rect 11788 14980 12628 15036
rect 12684 14980 14532 15036
rect 14588 14980 14598 15036
rect 16314 14980 16324 15036
rect 16380 14980 16390 15036
rect 16594 14980 16604 15036
rect 16660 14980 20692 15036
rect 20748 14980 21084 15036
rect 21140 14980 21150 15036
rect 21242 14980 21252 15036
rect 21308 14980 21346 15036
rect 23034 14980 23044 15036
rect 23100 14980 23324 15036
rect 23380 14980 23390 15036
rect 2874 14868 2884 14924
rect 2940 14868 8596 14924
rect 8652 14868 8662 14924
rect 8918 14868 8928 14924
rect 8984 14868 9032 14924
rect 9088 14868 9136 14924
rect 9192 14868 9202 14924
rect 11470 14868 11508 14924
rect 11564 14868 11574 14924
rect 13300 14868 15540 14924
rect 15596 14868 15606 14924
rect 16858 14868 16868 14924
rect 16924 14868 16972 14924
rect 17028 14868 17076 14924
rect 17132 14868 17142 14924
rect 18554 14868 18564 14924
rect 18620 14868 19852 14924
rect 19964 14868 19974 14924
rect 21476 14868 24668 14924
rect 24798 14868 24808 14924
rect 24864 14868 24912 14924
rect 24968 14868 25016 14924
rect 25072 14868 25082 14924
rect 13300 14812 13356 14868
rect 21476 14812 21532 14868
rect 24612 14812 24668 14868
rect 26124 14812 26180 15204
rect 26740 15148 26796 15428
rect 27402 15316 27412 15372
rect 27468 15316 31612 15372
rect 31668 15316 31678 15372
rect 27906 15204 27916 15260
rect 27972 15204 30212 15260
rect 30268 15204 31220 15260
rect 31276 15204 31286 15260
rect 26730 15092 26740 15148
rect 26796 15092 26806 15148
rect 28354 15092 28364 15148
rect 28420 15092 29204 15148
rect 29260 15092 29270 15148
rect 30034 15092 30044 15148
rect 30100 15092 30996 15148
rect 31052 15092 31062 15148
rect 31826 15092 31836 15148
rect 31892 15092 31947 15148
rect 31891 14924 31947 15092
rect 33200 14924 34000 14952
rect 31891 14868 32340 14924
rect 32396 14868 34000 14924
rect 33200 14840 34000 14868
rect 9594 14756 9604 14812
rect 9660 14756 11844 14812
rect 11900 14756 11910 14812
rect 12142 14756 12180 14812
rect 12236 14756 12246 14812
rect 12404 14756 13300 14812
rect 13356 14756 13366 14812
rect 14018 14756 14028 14812
rect 14084 14756 17556 14812
rect 17612 14756 17622 14812
rect 20234 14756 20244 14812
rect 20300 14756 21532 14812
rect 21970 14756 21980 14812
rect 22036 14756 23044 14812
rect 23100 14756 23110 14812
rect 24602 14756 24612 14812
rect 24668 14756 25508 14812
rect 25564 14756 25574 14812
rect 26114 14756 26124 14812
rect 26180 14756 26190 14812
rect 12404 14700 12460 14756
rect 10042 14644 10052 14700
rect 10108 14644 10948 14700
rect 11004 14644 11014 14700
rect 11162 14644 11172 14700
rect 11228 14644 12404 14700
rect 12460 14644 12470 14700
rect 12730 14644 12740 14700
rect 12796 14644 13188 14700
rect 13244 14644 13254 14700
rect 14298 14644 14308 14700
rect 14364 14644 17388 14700
rect 17444 14644 17668 14700
rect 17724 14644 18116 14700
rect 18172 14644 18182 14700
rect 18442 14644 18452 14700
rect 18508 14644 19292 14700
rect 19348 14644 19796 14700
rect 19852 14644 19862 14700
rect 20570 14644 20580 14700
rect 20636 14644 21476 14700
rect 21532 14644 21542 14700
rect 21634 14644 21644 14700
rect 21700 14644 22204 14700
rect 22260 14644 22270 14700
rect 22922 14644 22932 14700
rect 22988 14644 22998 14700
rect 24826 14644 24836 14700
rect 24892 14644 25284 14700
rect 25340 14644 25350 14700
rect 26618 14644 26628 14700
rect 26684 14644 27412 14700
rect 27468 14644 27478 14700
rect 27626 14644 27636 14700
rect 27692 14644 27804 14700
rect 27860 14644 27870 14700
rect 22932 14588 22988 14644
rect 11340 14532 21756 14588
rect 22418 14532 22428 14588
rect 22484 14532 24052 14588
rect 24108 14532 24118 14588
rect 25834 14532 25844 14588
rect 25900 14532 31724 14588
rect 31780 14532 31790 14588
rect 11340 14476 11396 14532
rect 21700 14476 21756 14532
rect 10154 14420 10164 14476
rect 10220 14420 10780 14476
rect 10836 14420 11340 14476
rect 11396 14420 11406 14476
rect 11722 14420 11732 14476
rect 11788 14420 12180 14476
rect 12236 14420 12246 14476
rect 12506 14420 12516 14476
rect 12572 14420 12852 14476
rect 12908 14420 12918 14476
rect 14522 14420 14532 14476
rect 14588 14420 15204 14476
rect 15260 14420 15270 14476
rect 17378 14420 17388 14476
rect 17444 14420 18452 14476
rect 18508 14420 18518 14476
rect 18610 14420 18620 14476
rect 18676 14420 20468 14476
rect 20524 14420 20534 14476
rect 21690 14420 21700 14476
rect 21756 14420 22932 14476
rect 22988 14420 22998 14476
rect 0 14364 800 14392
rect 0 14308 1204 14364
rect 1260 14308 1270 14364
rect 3490 14308 3500 14364
rect 3556 14308 5012 14364
rect 5068 14308 5078 14364
rect 8250 14308 8260 14364
rect 8316 14308 9380 14364
rect 9436 14308 9446 14364
rect 13514 14308 13524 14364
rect 13580 14308 14084 14364
rect 14140 14308 14150 14364
rect 14522 14308 14532 14364
rect 14588 14308 15147 14364
rect 15306 14308 15316 14364
rect 15372 14308 18396 14364
rect 18452 14308 18462 14364
rect 19114 14308 19124 14364
rect 19180 14308 21252 14364
rect 21308 14308 21318 14364
rect 21466 14308 21476 14364
rect 21532 14308 23716 14364
rect 23772 14308 23782 14364
rect 23930 14308 23940 14364
rect 23996 14308 27244 14364
rect 27300 14308 27310 14364
rect 27514 14308 27524 14364
rect 27580 14308 28700 14364
rect 28756 14308 29316 14364
rect 29372 14308 29382 14364
rect 0 14280 800 14308
rect 15091 14252 15147 14308
rect 5506 14196 5516 14252
rect 5572 14196 6244 14252
rect 6300 14196 14252 14252
rect 15091 14196 18564 14252
rect 18620 14196 18630 14252
rect 18890 14196 18900 14252
rect 18956 14196 20244 14252
rect 20300 14196 20310 14252
rect 20458 14196 20468 14252
rect 20524 14196 21756 14252
rect 22026 14196 22036 14252
rect 22092 14196 24052 14252
rect 24108 14196 24118 14252
rect 14196 14140 14252 14196
rect 21700 14140 21756 14196
rect 4948 14084 4958 14140
rect 5014 14084 5062 14140
rect 5118 14084 5166 14140
rect 5222 14084 5232 14140
rect 8026 14084 8036 14140
rect 8092 14084 10052 14140
rect 10108 14084 11284 14140
rect 11340 14084 11508 14140
rect 11564 14084 11574 14140
rect 12888 14084 12898 14140
rect 12954 14084 13002 14140
rect 13058 14084 13106 14140
rect 13162 14084 13172 14140
rect 14196 14084 19012 14140
rect 19068 14084 19078 14140
rect 20828 14084 20838 14140
rect 20894 14084 20942 14140
rect 20998 14084 21046 14140
rect 21102 14084 21112 14140
rect 21690 14084 21700 14140
rect 21756 14084 24780 14140
rect 24836 14084 24846 14140
rect 28768 14084 28778 14140
rect 28834 14084 28882 14140
rect 28938 14084 28986 14140
rect 29042 14084 29052 14140
rect 7466 13972 7476 14028
rect 7532 13972 9828 14028
rect 9884 13972 15092 14028
rect 15148 13972 16100 14028
rect 16156 13972 16166 14028
rect 16538 13972 16548 14028
rect 16604 13972 23212 14028
rect 23268 13972 23278 14028
rect 23706 13972 23716 14028
rect 23772 13972 24556 14028
rect 24612 13972 24622 14028
rect 26898 13972 26908 14028
rect 26964 13972 32004 14028
rect 32060 13972 32070 14028
rect 6346 13860 6356 13916
rect 6412 13860 8148 13916
rect 8204 13860 8214 13916
rect 9482 13860 9492 13916
rect 9548 13860 17388 13916
rect 17444 13860 17454 13916
rect 17770 13860 17780 13916
rect 17836 13860 22484 13916
rect 22540 13860 22550 13916
rect 22642 13860 22652 13916
rect 22708 13860 25060 13916
rect 25116 13860 25126 13916
rect 26842 13860 26852 13916
rect 26908 13860 27804 13916
rect 27860 13860 27870 13916
rect 1866 13748 1876 13804
rect 1932 13748 6916 13804
rect 6972 13748 6982 13804
rect 8418 13748 8428 13804
rect 8484 13748 10500 13804
rect 10556 13748 10566 13804
rect 11498 13748 11508 13804
rect 11564 13748 13412 13804
rect 13468 13748 13478 13804
rect 13626 13748 13636 13804
rect 13692 13748 13702 13804
rect 15194 13748 15204 13804
rect 15260 13748 15988 13804
rect 16044 13748 16054 13804
rect 17882 13748 17892 13804
rect 17948 13748 18788 13804
rect 18844 13748 18854 13804
rect 20131 13748 23604 13804
rect 23660 13748 23670 13804
rect 25386 13748 25396 13804
rect 25452 13748 25462 13804
rect 13412 13692 13468 13748
rect 13636 13692 13692 13748
rect 20131 13692 20187 13748
rect 1586 13636 1596 13692
rect 1652 13636 2996 13692
rect 3052 13636 5852 13692
rect 5908 13636 5918 13692
rect 7242 13636 7252 13692
rect 7308 13636 8148 13692
rect 8260 13636 8270 13692
rect 8586 13636 8596 13692
rect 8652 13636 9940 13692
rect 9996 13636 10006 13692
rect 13412 13636 13580 13692
rect 13636 13636 15428 13692
rect 15484 13636 17668 13692
rect 17724 13636 20187 13692
rect 20458 13636 20468 13692
rect 20580 13636 22036 13692
rect 22092 13636 22102 13692
rect 22250 13636 22260 13692
rect 22316 13636 22354 13692
rect 13524 13580 13580 13636
rect 25396 13580 25452 13748
rect 2314 13524 2324 13580
rect 2380 13524 3668 13580
rect 3724 13524 3734 13580
rect 3994 13524 4004 13580
rect 4060 13524 5404 13580
rect 5460 13524 5470 13580
rect 5954 13524 5964 13580
rect 6020 13524 7140 13580
rect 7196 13524 7206 13580
rect 9034 13524 9044 13580
rect 9100 13524 9110 13580
rect 10938 13524 10948 13580
rect 11004 13524 11396 13580
rect 11452 13524 11462 13580
rect 12114 13524 12124 13580
rect 12180 13524 13300 13580
rect 13356 13524 13366 13580
rect 13524 13524 14532 13580
rect 14588 13524 14598 13580
rect 14746 13524 14756 13580
rect 14812 13524 15036 13580
rect 15092 13524 16324 13580
rect 16380 13524 17108 13580
rect 17164 13524 17174 13580
rect 20738 13524 20748 13580
rect 20804 13524 21924 13580
rect 21980 13524 21990 13580
rect 22474 13524 22484 13580
rect 22540 13524 25508 13580
rect 25564 13524 25574 13580
rect 26394 13524 26404 13580
rect 26460 13524 27076 13580
rect 27132 13524 27142 13580
rect 9044 13468 9100 13524
rect 1194 13412 1204 13468
rect 1260 13412 4620 13468
rect 4676 13412 4686 13468
rect 8260 13412 9100 13468
rect 12002 13412 12012 13468
rect 12068 13412 15652 13468
rect 15708 13412 15718 13468
rect 16090 13412 16100 13468
rect 16156 13412 16436 13468
rect 16492 13412 16502 13468
rect 17546 13412 17556 13468
rect 17612 13412 21364 13468
rect 21420 13412 22820 13468
rect 22876 13412 22886 13468
rect 26618 13412 26628 13468
rect 26684 13412 27300 13468
rect 27356 13412 27366 13468
rect 8260 13356 8316 13412
rect 8250 13300 8260 13356
rect 8316 13300 8326 13356
rect 8918 13300 8928 13356
rect 8984 13300 9032 13356
rect 9088 13300 9136 13356
rect 9192 13300 9202 13356
rect 11498 13300 11508 13356
rect 11564 13300 11620 13356
rect 11676 13300 11686 13356
rect 13290 13300 13300 13356
rect 13356 13300 14420 13356
rect 14718 13300 14756 13356
rect 14812 13300 14822 13356
rect 16858 13300 16868 13356
rect 16924 13300 16972 13356
rect 17028 13300 17076 13356
rect 17132 13300 17142 13356
rect 17882 13300 17892 13356
rect 17948 13300 18172 13356
rect 18228 13300 18238 13356
rect 18442 13300 18452 13356
rect 18508 13300 21756 13356
rect 21812 13300 23268 13356
rect 23324 13300 23334 13356
rect 24798 13300 24808 13356
rect 24864 13300 24912 13356
rect 24968 13300 25016 13356
rect 25072 13300 25082 13356
rect 14364 13244 14420 13300
rect 1754 13188 1764 13244
rect 1820 13188 6860 13244
rect 6916 13188 6926 13244
rect 8642 13188 8652 13244
rect 8708 13188 13636 13244
rect 13692 13188 14196 13244
rect 14252 13188 14262 13244
rect 14364 13188 14644 13244
rect 14700 13188 17444 13244
rect 17500 13188 18340 13244
rect 18396 13188 18406 13244
rect 18554 13188 18564 13244
rect 18620 13188 18900 13244
rect 18956 13188 18966 13244
rect 19338 13188 19348 13244
rect 19404 13188 20468 13244
rect 20524 13188 21364 13244
rect 21420 13188 21430 13244
rect 23818 13188 23828 13244
rect 23884 13188 25172 13244
rect 25228 13188 25238 13244
rect 0 13132 800 13160
rect 0 13076 1316 13132
rect 1372 13076 1382 13132
rect 6626 13076 6636 13132
rect 6692 13076 7028 13132
rect 7084 13076 7588 13132
rect 7644 13076 7654 13132
rect 8866 13076 8876 13132
rect 8932 13076 15540 13132
rect 15596 13076 15606 13132
rect 18106 13076 18116 13132
rect 18172 13076 21028 13132
rect 21084 13076 21094 13132
rect 22362 13076 22372 13132
rect 22428 13076 22932 13132
rect 22988 13076 24164 13132
rect 24220 13076 24230 13132
rect 24602 13076 24612 13132
rect 24668 13076 25340 13132
rect 25396 13076 25406 13132
rect 26058 13076 26068 13132
rect 26124 13076 27188 13132
rect 27244 13076 27254 13132
rect 28242 13076 28252 13132
rect 28308 13076 29204 13132
rect 29260 13076 29270 13132
rect 0 13048 800 13076
rect 2426 12964 2436 13020
rect 2492 12964 4564 13020
rect 4620 12964 4630 13020
rect 10434 12964 10444 13020
rect 10500 12964 11396 13020
rect 11452 12964 12236 13020
rect 14186 12964 14196 13020
rect 14252 12964 19180 13020
rect 19236 12964 19246 13020
rect 19730 12964 19740 13020
rect 19796 12964 22148 13020
rect 22204 12964 22820 13020
rect 22876 12964 22886 13020
rect 24490 12964 24500 13020
rect 24556 12964 25788 13020
rect 25844 12964 25854 13020
rect 30202 12964 30212 13020
rect 30268 12964 30772 13020
rect 30828 12964 31444 13020
rect 31500 12964 31510 13020
rect 12180 12908 12236 12964
rect 1698 12852 1708 12908
rect 1764 12852 2660 12908
rect 2716 12852 2726 12908
rect 10098 12852 10108 12908
rect 10164 12852 11956 12908
rect 12012 12852 12022 12908
rect 12180 12852 14308 12908
rect 14364 12852 14374 12908
rect 14522 12852 14532 12908
rect 14588 12852 15316 12908
rect 15372 12852 15382 12908
rect 15530 12852 15540 12908
rect 15596 12852 16380 12908
rect 16436 12852 16996 12908
rect 17052 12852 17780 12908
rect 17836 12852 18228 12908
rect 18284 12852 18294 12908
rect 18564 12852 20692 12908
rect 20748 12852 20758 12908
rect 22408 12852 22484 12908
rect 22540 12852 22988 12908
rect 23044 12852 23054 12908
rect 24490 12852 24500 12908
rect 24556 12852 24780 12908
rect 24836 12852 24846 12908
rect 25610 12852 25620 12908
rect 25676 12852 28028 12908
rect 28084 12852 28094 12908
rect 3154 12740 3164 12796
rect 3220 12740 4116 12796
rect 4172 12740 5404 12796
rect 5460 12740 5470 12796
rect 9874 12740 9884 12796
rect 9940 12740 12068 12796
rect 12124 12740 12134 12796
rect 12282 12740 12292 12796
rect 12348 12740 13020 12796
rect 13076 12740 13748 12796
rect 13804 12740 14532 12796
rect 14588 12740 14598 12796
rect 17546 12740 17556 12796
rect 17612 12740 18340 12796
rect 18396 12740 18406 12796
rect 13626 12628 13636 12684
rect 13692 12628 15540 12684
rect 15596 12628 16212 12684
rect 16268 12628 18004 12684
rect 18060 12628 18070 12684
rect 18564 12572 18620 12852
rect 18778 12740 18788 12796
rect 18844 12740 24500 12796
rect 24556 12740 24566 12796
rect 25050 12740 25060 12796
rect 25116 12740 27916 12796
rect 27972 12740 27982 12796
rect 19898 12628 19908 12684
rect 19964 12628 23044 12684
rect 23100 12628 23110 12684
rect 23762 12628 23772 12684
rect 23828 12628 26292 12684
rect 26348 12628 26358 12684
rect 4948 12516 4958 12572
rect 5014 12516 5062 12572
rect 5118 12516 5166 12572
rect 5222 12516 5232 12572
rect 12888 12516 12898 12572
rect 12954 12516 13002 12572
rect 13058 12516 13106 12572
rect 13162 12516 13172 12572
rect 13626 12516 13636 12572
rect 13692 12516 14084 12572
rect 14140 12516 16380 12572
rect 17322 12516 17332 12572
rect 17388 12516 18620 12572
rect 20828 12516 20838 12572
rect 20894 12516 20942 12572
rect 20998 12516 21046 12572
rect 21102 12516 21112 12572
rect 28768 12516 28778 12572
rect 28834 12516 28882 12572
rect 28938 12516 28986 12572
rect 29042 12516 29052 12572
rect 1866 12404 1876 12460
rect 1932 12404 6468 12460
rect 6524 12404 6534 12460
rect 11498 12404 11508 12460
rect 11564 12404 11732 12460
rect 11788 12404 12628 12460
rect 12684 12404 13412 12460
rect 13468 12404 14532 12460
rect 14588 12404 14598 12460
rect 16324 12348 16380 12516
rect 17770 12404 17780 12460
rect 17836 12404 18676 12460
rect 18732 12404 18742 12460
rect 18890 12404 18900 12460
rect 18956 12404 19908 12460
rect 19964 12404 23604 12460
rect 23660 12404 23670 12460
rect 6234 12292 6244 12348
rect 6300 12292 7196 12348
rect 7252 12292 8260 12348
rect 8316 12292 8326 12348
rect 16324 12292 18676 12348
rect 18732 12292 19124 12348
rect 19180 12292 19190 12348
rect 20346 12292 20356 12348
rect 20412 12292 23772 12348
rect 23828 12292 23838 12348
rect 1306 12180 1316 12236
rect 1372 12180 1596 12236
rect 1652 12180 1662 12236
rect 2314 12180 2324 12236
rect 2380 12180 4228 12236
rect 4284 12180 4294 12236
rect 5842 12180 5852 12236
rect 5908 12180 10276 12236
rect 10332 12180 10342 12236
rect 12506 12180 12516 12236
rect 12572 12180 16492 12236
rect 17882 12180 17892 12236
rect 17948 12180 19012 12236
rect 19068 12180 19078 12236
rect 19450 12180 19460 12236
rect 19516 12180 20132 12236
rect 20188 12180 20748 12236
rect 20804 12180 20814 12236
rect 16436 12124 16492 12180
rect 8810 12068 8820 12124
rect 8876 12068 10052 12124
rect 10108 12068 10118 12124
rect 10602 12068 10612 12124
rect 10668 12068 11620 12124
rect 11676 12068 11686 12124
rect 14410 12068 14420 12124
rect 14476 12068 15652 12124
rect 15708 12068 15988 12124
rect 16044 12068 16054 12124
rect 16426 12068 16436 12124
rect 16492 12068 17780 12124
rect 17836 12068 17846 12124
rect 18498 12068 18508 12124
rect 18564 12068 20020 12124
rect 20076 12068 20636 12124
rect 20692 12068 20702 12124
rect 24462 12068 24500 12124
rect 24556 12068 24566 12124
rect 26618 12068 26628 12124
rect 26684 12068 27188 12124
rect 27244 12068 28308 12124
rect 28364 12068 28374 12124
rect 28634 12068 28644 12124
rect 28700 12068 29428 12124
rect 29484 12068 30044 12124
rect 30100 12068 30110 12124
rect 1866 11956 1876 12012
rect 1932 11956 5516 12012
rect 5572 11956 5582 12012
rect 7074 11956 7084 12012
rect 7140 11956 7924 12012
rect 7980 11956 9492 12012
rect 9548 11956 10500 12012
rect 10556 11956 12180 12012
rect 12236 11956 12246 12012
rect 16202 11956 16212 12012
rect 16268 11956 16884 12012
rect 16940 11956 16950 12012
rect 17658 11956 17668 12012
rect 17724 11956 18284 12012
rect 18340 11956 19348 12012
rect 19404 11956 19414 12012
rect 31826 11956 31836 12012
rect 31892 11956 32340 12012
rect 32396 11956 32620 12012
rect 0 11900 800 11928
rect 16884 11900 16940 11956
rect 0 11844 1372 11900
rect 1428 11844 1438 11900
rect 9258 11844 9268 11900
rect 9324 11844 9940 11900
rect 9996 11844 11900 11900
rect 12058 11844 12068 11900
rect 12124 11844 12796 11900
rect 12852 11844 15204 11900
rect 15260 11844 16660 11900
rect 16716 11844 16726 11900
rect 16884 11844 19236 11900
rect 19292 11844 20356 11900
rect 20412 11844 20422 11900
rect 24658 11844 24668 11900
rect 24724 11844 32116 11900
rect 32172 11844 32182 11900
rect 0 11816 800 11844
rect 11844 11788 11900 11844
rect 8918 11732 8928 11788
rect 8984 11732 9032 11788
rect 9088 11732 9136 11788
rect 9192 11732 9202 11788
rect 11834 11732 11844 11788
rect 11900 11732 14644 11788
rect 14700 11732 14710 11788
rect 16858 11732 16868 11788
rect 16924 11732 16972 11788
rect 17028 11732 17076 11788
rect 17132 11732 17142 11788
rect 24798 11732 24808 11788
rect 24864 11732 24912 11788
rect 24968 11732 25016 11788
rect 25072 11732 25082 11788
rect 32564 11676 32620 11956
rect 33200 11676 34000 11704
rect 2202 11620 2212 11676
rect 2268 11620 2660 11676
rect 2716 11620 4676 11676
rect 4732 11620 4742 11676
rect 7130 11620 7140 11676
rect 7196 11620 9324 11676
rect 9380 11620 11508 11676
rect 11564 11620 11574 11676
rect 12730 11620 12740 11676
rect 12796 11620 15092 11676
rect 15148 11620 15158 11676
rect 17210 11620 17220 11676
rect 17276 11620 17388 11676
rect 17444 11620 17454 11676
rect 17966 11620 18004 11676
rect 18060 11620 18070 11676
rect 25778 11620 25788 11676
rect 25844 11620 26068 11676
rect 26124 11620 27300 11676
rect 27356 11620 27366 11676
rect 32564 11620 34000 11676
rect 33200 11592 34000 11620
rect 2314 11508 2324 11564
rect 2380 11508 3276 11564
rect 3332 11508 4564 11564
rect 4620 11508 4630 11564
rect 9706 11508 9716 11564
rect 9772 11508 10052 11564
rect 10108 11508 10118 11564
rect 10910 11508 10948 11564
rect 11004 11508 11014 11564
rect 11386 11508 11396 11564
rect 11452 11508 11620 11564
rect 11676 11508 11686 11564
rect 12954 11508 12964 11564
rect 13020 11508 13524 11564
rect 13580 11508 13590 11564
rect 14298 11508 14308 11564
rect 14364 11508 15876 11564
rect 15932 11508 15942 11564
rect 17490 11508 17500 11564
rect 17556 11508 18900 11564
rect 18956 11508 18966 11564
rect 19674 11508 19684 11564
rect 19740 11508 21364 11564
rect 21420 11508 21430 11564
rect 3098 11396 3108 11452
rect 3164 11396 4452 11452
rect 4508 11396 4518 11452
rect 6234 11396 6244 11452
rect 6300 11396 6804 11452
rect 6860 11396 7252 11452
rect 7308 11396 7318 11452
rect 10266 11396 10276 11452
rect 10332 11396 10836 11452
rect 10892 11396 10902 11452
rect 11050 11396 11060 11452
rect 11116 11396 13300 11452
rect 13356 11396 13366 11452
rect 26842 11396 26852 11452
rect 26908 11396 27412 11452
rect 27468 11396 27478 11452
rect 5786 11284 5796 11340
rect 5852 11284 8708 11340
rect 8764 11284 8774 11340
rect 9426 11284 9436 11340
rect 9492 11284 11396 11340
rect 11452 11284 11462 11340
rect 12002 11284 12012 11340
rect 12068 11284 12404 11340
rect 12460 11284 12470 11340
rect 13636 11284 15316 11340
rect 15372 11284 15382 11340
rect 16426 11284 16436 11340
rect 16492 11284 16940 11340
rect 16996 11284 17006 11340
rect 7578 11172 7588 11228
rect 7644 11172 8036 11228
rect 8092 11172 9660 11228
rect 9716 11172 11508 11228
rect 11564 11172 12572 11228
rect 12628 11172 13300 11228
rect 13356 11172 13366 11228
rect 8138 11060 8148 11116
rect 8204 11060 13580 11116
rect 13636 11060 13692 11284
rect 14466 11172 14476 11228
rect 14532 11172 18788 11228
rect 18844 11172 18854 11228
rect 21130 11172 21140 11228
rect 21196 11172 21476 11228
rect 21532 11172 21868 11228
rect 21924 11172 21934 11228
rect 18274 11060 18284 11116
rect 18340 11060 19012 11116
rect 19068 11060 19078 11116
rect 4948 10948 4958 11004
rect 5014 10948 5062 11004
rect 5118 10948 5166 11004
rect 5222 10948 5232 11004
rect 9902 10948 9940 11004
rect 9996 10948 10006 11004
rect 12888 10948 12898 11004
rect 12954 10948 13002 11004
rect 13058 10948 13106 11004
rect 13162 10948 13172 11004
rect 13290 10948 13300 11004
rect 13356 10948 14140 11004
rect 20828 10948 20838 11004
rect 20894 10948 20942 11004
rect 20998 10948 21046 11004
rect 21102 10948 21112 11004
rect 28768 10948 28778 11004
rect 28834 10948 28882 11004
rect 28938 10948 28986 11004
rect 29042 10948 29052 11004
rect 14084 10892 14140 10948
rect 10322 10836 10332 10892
rect 10388 10836 11396 10892
rect 11452 10836 13412 10892
rect 13468 10836 13478 10892
rect 14084 10836 14364 10892
rect 14308 10780 14364 10836
rect 12842 10724 12852 10780
rect 12908 10724 14140 10780
rect 14196 10724 14206 10780
rect 14298 10724 14308 10780
rect 14364 10724 14374 10780
rect 14746 10724 14756 10780
rect 14812 10724 15540 10780
rect 15596 10724 15606 10780
rect 23146 10724 23156 10780
rect 23212 10724 23996 10780
rect 24052 10724 24062 10780
rect 24546 10724 24556 10780
rect 24612 10724 25284 10780
rect 25340 10724 25350 10780
rect 0 10668 800 10696
rect 0 10612 3556 10668
rect 3612 10612 3622 10668
rect 4218 10612 4228 10668
rect 4284 10612 7028 10668
rect 7084 10612 7094 10668
rect 10154 10612 10164 10668
rect 10220 10612 19796 10668
rect 19852 10612 19862 10668
rect 0 10584 800 10612
rect 2986 10500 2996 10556
rect 3052 10500 4788 10556
rect 4844 10500 4854 10556
rect 8222 10500 8260 10556
rect 8316 10500 8326 10556
rect 12562 10500 12572 10556
rect 12628 10500 13636 10556
rect 13692 10500 13702 10556
rect 13794 10500 13804 10556
rect 13860 10500 14756 10556
rect 14812 10500 14822 10556
rect 15474 10500 15484 10556
rect 15540 10500 17332 10556
rect 17388 10500 17398 10556
rect 18190 10500 18228 10556
rect 18284 10500 18294 10556
rect 24098 10500 24108 10556
rect 24164 10500 24892 10556
rect 24948 10500 26068 10556
rect 26124 10500 26134 10556
rect 5450 10388 5460 10444
rect 5516 10388 9100 10444
rect 9156 10388 9166 10444
rect 10882 10388 10892 10444
rect 10948 10388 12796 10444
rect 12852 10388 13692 10444
rect 14858 10388 14868 10444
rect 14924 10388 17780 10444
rect 17836 10388 18452 10444
rect 18508 10388 18518 10444
rect 23482 10388 23492 10444
rect 23548 10388 24444 10444
rect 24500 10388 24510 10444
rect 24994 10388 25004 10444
rect 25060 10388 25956 10444
rect 26012 10388 26022 10444
rect 26618 10388 26628 10444
rect 26684 10388 27132 10444
rect 27188 10388 28084 10444
rect 28140 10388 28150 10444
rect 13636 10276 13692 10388
rect 13748 10276 13758 10332
rect 15138 10276 15148 10332
rect 15204 10276 19348 10332
rect 19404 10276 19414 10332
rect 23538 10276 23548 10332
rect 23604 10276 32228 10332
rect 32284 10276 32294 10332
rect 5422 10164 5460 10220
rect 5516 10164 5526 10220
rect 8918 10164 8928 10220
rect 8984 10164 9032 10220
rect 9088 10164 9136 10220
rect 9192 10164 9202 10220
rect 10042 10164 10052 10220
rect 10108 10164 11732 10220
rect 11788 10164 11798 10220
rect 12842 10164 12852 10220
rect 12908 10164 15484 10220
rect 15540 10164 15550 10220
rect 16858 10164 16868 10220
rect 16924 10164 16972 10220
rect 17028 10164 17076 10220
rect 17132 10164 17142 10220
rect 19002 10164 19012 10220
rect 19068 10164 20187 10220
rect 24798 10164 24808 10220
rect 24864 10164 24912 10220
rect 24968 10164 25016 10220
rect 25072 10164 25082 10220
rect 4890 10052 4900 10108
rect 4956 10052 5908 10108
rect 5964 10052 5974 10108
rect 7242 10052 7252 10108
rect 7308 10052 8092 10108
rect 8148 10052 8158 10108
rect 10266 10052 10276 10108
rect 10332 10052 10780 10108
rect 10836 10052 10846 10108
rect 11218 10052 11228 10108
rect 11284 10052 11620 10108
rect 11676 10052 11686 10108
rect 11890 10052 11900 10108
rect 11956 10052 14924 10108
rect 14980 10052 14990 10108
rect 11284 9996 11340 10052
rect 20131 9996 20187 10164
rect 1530 9940 1540 9996
rect 1596 9940 2548 9996
rect 2604 9940 4060 9996
rect 4172 9940 4182 9996
rect 6458 9940 6468 9996
rect 6524 9940 7476 9996
rect 7532 9940 8316 9996
rect 8372 9940 8382 9996
rect 8698 9940 8708 9996
rect 8764 9940 10164 9996
rect 10220 9940 11060 9996
rect 11116 9940 11126 9996
rect 11284 9940 12852 9996
rect 12908 9940 12918 9996
rect 13402 9940 13412 9996
rect 13468 9940 14084 9996
rect 14140 9940 14150 9996
rect 20131 9940 24836 9996
rect 24892 9940 24902 9996
rect 27850 9940 27860 9996
rect 27916 9940 32004 9996
rect 32060 9940 32070 9996
rect 11284 9884 11340 9940
rect 5898 9828 5908 9884
rect 5964 9828 7588 9884
rect 7644 9828 7654 9884
rect 7746 9828 7756 9884
rect 7812 9828 9436 9884
rect 9492 9828 9502 9884
rect 9940 9828 11340 9884
rect 11722 9828 11732 9884
rect 11788 9828 12292 9884
rect 12348 9828 12516 9884
rect 12572 9828 12582 9884
rect 13402 9828 13412 9884
rect 13468 9828 14980 9884
rect 15036 9828 15988 9884
rect 16044 9828 16054 9884
rect 18106 9828 18116 9884
rect 18172 9828 21028 9884
rect 21084 9828 21094 9884
rect 9940 9772 9996 9828
rect 4778 9716 4788 9772
rect 4844 9716 5068 9772
rect 5124 9716 5348 9772
rect 5404 9716 5414 9772
rect 8810 9716 8820 9772
rect 8876 9716 9996 9772
rect 10154 9716 10164 9772
rect 10220 9716 11508 9772
rect 11564 9716 14532 9772
rect 14588 9716 14598 9772
rect 15306 9716 15316 9772
rect 15372 9716 15764 9772
rect 15820 9716 15830 9772
rect 16874 9716 16884 9772
rect 16940 9716 18004 9772
rect 18060 9716 18070 9772
rect 26562 9716 26572 9772
rect 26628 9716 26964 9772
rect 27020 9716 27804 9772
rect 27860 9716 27870 9772
rect 4554 9604 4564 9660
rect 4620 9604 9604 9660
rect 9660 9604 9670 9660
rect 11890 9604 11900 9660
rect 11956 9604 12292 9660
rect 12348 9604 12358 9660
rect 13906 9604 13916 9660
rect 13972 9604 14644 9660
rect 14700 9604 14710 9660
rect 25722 9604 25732 9660
rect 25788 9604 27692 9660
rect 27748 9604 27758 9660
rect 8250 9492 8260 9548
rect 8316 9492 11172 9548
rect 11228 9492 12180 9548
rect 12236 9492 12516 9548
rect 12572 9492 12582 9548
rect 13458 9492 13468 9548
rect 13524 9492 14420 9548
rect 14476 9492 14486 9548
rect 14746 9492 14756 9548
rect 14812 9492 15428 9548
rect 15484 9492 15494 9548
rect 26730 9492 26740 9548
rect 26796 9492 27300 9548
rect 27356 9492 27366 9548
rect 4948 9380 4958 9436
rect 5014 9380 5062 9436
rect 5118 9380 5166 9436
rect 5222 9380 5232 9436
rect 12888 9380 12898 9436
rect 12954 9380 13002 9436
rect 13058 9380 13106 9436
rect 13162 9380 13172 9436
rect 20828 9380 20838 9436
rect 20894 9380 20942 9436
rect 20998 9380 21046 9436
rect 21102 9380 21112 9436
rect 28768 9380 28778 9436
rect 28834 9380 28882 9436
rect 28938 9380 28986 9436
rect 29042 9380 29052 9436
rect 0 9324 800 9352
rect 0 9268 1316 9324
rect 1372 9268 1540 9324
rect 1596 9268 1606 9324
rect 1866 9268 1876 9324
rect 1932 9268 8036 9324
rect 8092 9268 8102 9324
rect 11890 9268 11900 9324
rect 11956 9268 13580 9324
rect 13636 9268 13646 9324
rect 0 9240 800 9268
rect 7578 9156 7588 9212
rect 7644 9156 8148 9212
rect 8204 9156 8214 9212
rect 12618 9156 12628 9212
rect 12684 9156 13188 9212
rect 13244 9156 13254 9212
rect 22222 9156 22260 9212
rect 22316 9156 22326 9212
rect 3434 9044 3444 9100
rect 3500 9044 4564 9100
rect 4620 9044 4630 9100
rect 12282 9044 12292 9100
rect 12348 9044 13972 9100
rect 14028 9044 14420 9100
rect 14476 9044 14486 9100
rect 14634 9044 14644 9100
rect 14700 9044 15316 9100
rect 15372 9044 15382 9100
rect 21578 9044 21588 9100
rect 21644 9044 23156 9100
rect 23212 9044 23222 9100
rect 6458 8932 6468 8988
rect 6524 8932 7532 8988
rect 7588 8932 7598 8988
rect 7914 8932 7924 8988
rect 7980 8932 8372 8988
rect 8428 8932 8438 8988
rect 11610 8932 11620 8988
rect 11676 8932 12404 8988
rect 12460 8932 12796 8988
rect 12852 8932 13356 8988
rect 13412 8932 13422 8988
rect 19954 8932 19964 8988
rect 20020 8932 20356 8988
rect 20412 8932 21420 8988
rect 21476 8932 21486 8988
rect 7532 8876 7588 8932
rect 7532 8820 8260 8876
rect 8316 8820 8326 8876
rect 8530 8820 8540 8876
rect 8596 8820 9100 8876
rect 9156 8820 9166 8876
rect 18106 8820 18116 8876
rect 18172 8820 24164 8876
rect 24220 8820 24230 8876
rect 31826 8820 31836 8876
rect 31892 8820 32340 8876
rect 32396 8820 32406 8876
rect 6346 8708 6356 8764
rect 6412 8708 7308 8764
rect 7364 8708 8148 8764
rect 8204 8708 8214 8764
rect 8918 8596 8928 8652
rect 8984 8596 9032 8652
rect 9088 8596 9136 8652
rect 9192 8596 9202 8652
rect 9258 8596 9268 8652
rect 9324 8596 9772 8652
rect 9828 8596 12964 8652
rect 13020 8596 14868 8652
rect 14924 8596 14934 8652
rect 16858 8596 16868 8652
rect 16924 8596 16972 8652
rect 17028 8596 17076 8652
rect 17132 8596 17142 8652
rect 24798 8596 24808 8652
rect 24864 8596 24912 8652
rect 24968 8596 25016 8652
rect 25072 8596 25082 8652
rect 6122 8484 6132 8540
rect 6188 8484 7420 8540
rect 7476 8484 10276 8540
rect 10332 8484 10342 8540
rect 7028 8372 8484 8428
rect 8540 8372 8550 8428
rect 15866 8372 15876 8428
rect 15932 8372 16660 8428
rect 16716 8372 17276 8428
rect 17332 8372 17444 8428
rect 17500 8372 20188 8428
rect 7028 8316 7084 8372
rect 20132 8316 20188 8372
rect 33200 8316 34000 8344
rect 4946 8260 4956 8316
rect 5012 8260 5460 8316
rect 5516 8260 5526 8316
rect 5898 8260 5908 8316
rect 5964 8260 7028 8316
rect 7084 8260 7094 8316
rect 12282 8260 12292 8316
rect 12348 8260 17556 8316
rect 17612 8260 17622 8316
rect 20122 8260 20132 8316
rect 20188 8260 21252 8316
rect 21308 8260 22036 8316
rect 22092 8260 24332 8316
rect 24490 8260 24500 8316
rect 24556 8260 25284 8316
rect 25340 8260 25350 8316
rect 25498 8260 25508 8316
rect 25564 8260 26572 8316
rect 26628 8260 26638 8316
rect 32442 8260 32452 8316
rect 32508 8260 34000 8316
rect 24276 8204 24332 8260
rect 33200 8232 34000 8260
rect 8698 8148 8708 8204
rect 8764 8148 12180 8204
rect 12236 8148 12246 8204
rect 14522 8148 14532 8204
rect 14588 8148 16884 8204
rect 16940 8148 16950 8204
rect 19786 8148 19796 8204
rect 19852 8148 20804 8204
rect 20860 8148 21700 8204
rect 21756 8148 21766 8204
rect 21914 8148 21924 8204
rect 21980 8148 23716 8204
rect 23772 8148 23782 8204
rect 24276 8148 25172 8204
rect 25228 8148 26068 8204
rect 26124 8148 26134 8204
rect 0 8092 800 8120
rect 0 8036 1316 8092
rect 1372 8036 1382 8092
rect 4302 8036 4340 8092
rect 4396 8036 4406 8092
rect 0 8008 800 8036
rect 4948 7812 4958 7868
rect 5014 7812 5062 7868
rect 5118 7812 5166 7868
rect 5222 7812 5232 7868
rect 12888 7812 12898 7868
rect 12954 7812 13002 7868
rect 13058 7812 13106 7868
rect 13162 7812 13172 7868
rect 20828 7812 20838 7868
rect 20894 7812 20942 7868
rect 20998 7812 21046 7868
rect 21102 7812 21112 7868
rect 28768 7812 28778 7868
rect 28834 7812 28882 7868
rect 28938 7812 28986 7868
rect 29042 7812 29052 7868
rect 4442 7700 4452 7756
rect 4508 7700 6804 7756
rect 6860 7700 6870 7756
rect 8138 7700 8148 7756
rect 8204 7700 9940 7756
rect 9996 7700 11620 7756
rect 11676 7700 11686 7756
rect 1306 7588 1316 7644
rect 1372 7588 5684 7644
rect 5740 7588 6580 7644
rect 6636 7588 6646 7644
rect 8922 7588 8932 7644
rect 8988 7588 9940 7644
rect 9996 7588 10006 7644
rect 15418 7588 15428 7644
rect 15484 7588 16212 7644
rect 16268 7588 16278 7644
rect 18498 7588 18508 7644
rect 18564 7588 20244 7644
rect 20300 7588 20310 7644
rect 22810 7588 22820 7644
rect 22876 7588 25116 7644
rect 25172 7588 25182 7644
rect 1754 7476 1764 7532
rect 1820 7476 6020 7532
rect 6076 7476 6086 7532
rect 6682 7476 6692 7532
rect 6748 7476 7588 7532
rect 15082 7476 15092 7532
rect 15148 7476 16884 7532
rect 16940 7476 16950 7532
rect 17742 7476 17780 7532
rect 17836 7476 17846 7532
rect 4050 7364 4060 7420
rect 4116 7364 6468 7420
rect 6524 7364 7252 7420
rect 7308 7364 7318 7420
rect 7532 7308 7588 7476
rect 10938 7364 10948 7420
rect 11004 7364 11956 7420
rect 12012 7364 12796 7420
rect 12852 7364 18844 7420
rect 18900 7364 19236 7420
rect 19292 7364 19684 7420
rect 19740 7364 19750 7420
rect 3210 7252 3220 7308
rect 3276 7252 5460 7308
rect 5516 7252 5526 7308
rect 7532 7252 7644 7308
rect 7756 7252 7766 7308
rect 8194 7252 8204 7308
rect 8260 7252 9156 7308
rect 9212 7252 9222 7308
rect 10826 7252 10836 7308
rect 10892 7252 12516 7308
rect 12572 7252 12582 7308
rect 13290 7252 13300 7308
rect 13356 7252 13916 7308
rect 13972 7252 14980 7308
rect 15036 7252 15046 7308
rect 1418 7140 1428 7196
rect 1484 7140 4956 7196
rect 5012 7140 6356 7196
rect 6412 7140 6422 7196
rect 10378 7140 10388 7196
rect 10444 7140 11284 7196
rect 11340 7140 11350 7196
rect 23370 7140 23380 7196
rect 23436 7140 25396 7196
rect 25452 7140 25462 7196
rect 1474 7028 1484 7084
rect 1540 7028 2268 7084
rect 2426 7028 2436 7084
rect 2492 7028 3108 7084
rect 3164 7028 6972 7084
rect 7028 7028 7038 7084
rect 8918 7028 8928 7084
rect 8984 7028 9032 7084
rect 9088 7028 9136 7084
rect 9192 7028 9202 7084
rect 10658 7028 10668 7084
rect 10724 7028 11900 7084
rect 11956 7028 14644 7084
rect 14700 7028 14710 7084
rect 16858 7028 16868 7084
rect 16924 7028 16972 7084
rect 17028 7028 17076 7084
rect 17132 7028 17142 7084
rect 24798 7028 24808 7084
rect 24864 7028 24912 7084
rect 24968 7028 25016 7084
rect 25072 7028 25082 7084
rect 1194 6916 1204 6972
rect 1260 6916 1988 6972
rect 2044 6916 2054 6972
rect 2212 6916 2268 7028
rect 2324 6916 6804 6972
rect 6860 6916 6870 6972
rect 10826 6916 10836 6972
rect 10892 6916 12348 6972
rect 12404 6916 12414 6972
rect 12516 6916 17892 6972
rect 17948 6916 19236 6972
rect 19292 6916 19796 6972
rect 19852 6916 19862 6972
rect 0 6860 800 6888
rect 12516 6860 12572 6916
rect 0 6804 1596 6860
rect 3434 6804 3444 6860
rect 3500 6804 5348 6860
rect 5404 6804 5414 6860
rect 6234 6804 6244 6860
rect 6300 6804 6860 6860
rect 6990 6804 7028 6860
rect 7084 6804 7420 6860
rect 7476 6804 7486 6860
rect 7914 6804 7924 6860
rect 7980 6804 12572 6860
rect 14746 6804 14756 6860
rect 14812 6804 15988 6860
rect 16044 6804 16054 6860
rect 21690 6804 21700 6860
rect 21756 6804 24332 6860
rect 24388 6804 24398 6860
rect 0 6776 800 6804
rect 1540 6636 1596 6804
rect 6804 6748 6860 6804
rect 3994 6692 4004 6748
rect 4060 6692 4452 6748
rect 4508 6692 4518 6748
rect 6804 6692 8148 6748
rect 8204 6692 8214 6748
rect 11508 6692 13076 6748
rect 13132 6692 13142 6748
rect 14382 6692 14420 6748
rect 14476 6692 14486 6748
rect 17770 6692 17780 6748
rect 17836 6692 18676 6748
rect 18732 6692 18742 6748
rect 22026 6692 22036 6748
rect 22092 6692 22820 6748
rect 22876 6692 24108 6748
rect 24164 6692 24174 6748
rect 11508 6636 11564 6692
rect 1540 6580 3444 6636
rect 3500 6580 3724 6636
rect 3780 6580 3790 6636
rect 4106 6580 4116 6636
rect 4172 6580 5684 6636
rect 5740 6580 5750 6636
rect 6122 6580 6132 6636
rect 6188 6580 7700 6636
rect 7756 6580 7766 6636
rect 8586 6580 8596 6636
rect 8652 6580 9380 6636
rect 9436 6580 9828 6636
rect 9884 6580 10332 6636
rect 10388 6580 11564 6636
rect 11722 6580 11732 6636
rect 11788 6580 12516 6636
rect 12572 6580 12582 6636
rect 17210 6580 17220 6636
rect 17276 6580 18228 6636
rect 18284 6580 18294 6636
rect 19674 6580 19684 6636
rect 19740 6580 22148 6636
rect 22204 6580 22596 6636
rect 22652 6580 22662 6636
rect 23818 6580 23828 6636
rect 23884 6580 24556 6636
rect 24612 6580 24622 6636
rect 26170 6580 26180 6636
rect 26236 6580 26964 6636
rect 27020 6580 27030 6636
rect 1642 6468 1652 6524
rect 1708 6468 5236 6524
rect 5292 6468 5302 6524
rect 6794 6468 6804 6524
rect 6860 6468 6916 6524
rect 6972 6468 6982 6524
rect 8026 6468 8036 6524
rect 8092 6468 8484 6524
rect 8540 6468 8550 6524
rect 9034 6468 9044 6524
rect 9100 6468 9604 6524
rect 9660 6468 9670 6524
rect 9930 6468 9940 6524
rect 9996 6468 11620 6524
rect 11676 6468 11686 6524
rect 22698 6468 22708 6524
rect 22764 6468 26628 6524
rect 26684 6468 26694 6524
rect 4330 6356 4340 6412
rect 4396 6356 6188 6412
rect 6244 6356 6254 6412
rect 8138 6356 8148 6412
rect 8204 6356 10500 6412
rect 10556 6356 12068 6412
rect 12124 6356 12134 6412
rect 19002 6356 19012 6412
rect 19068 6356 19796 6412
rect 19852 6356 25284 6412
rect 25340 6356 26292 6412
rect 26348 6356 26358 6412
rect 26068 6300 26124 6356
rect 4948 6244 4958 6300
rect 5014 6244 5062 6300
rect 5118 6244 5166 6300
rect 5222 6244 5232 6300
rect 7690 6244 7700 6300
rect 7756 6244 12180 6300
rect 12236 6244 12246 6300
rect 12888 6244 12898 6300
rect 12954 6244 13002 6300
rect 13058 6244 13106 6300
rect 13162 6244 13172 6300
rect 20828 6244 20838 6300
rect 20894 6244 20942 6300
rect 20998 6244 21046 6300
rect 21102 6244 21112 6300
rect 23930 6244 23940 6300
rect 23996 6244 25676 6300
rect 25732 6244 25742 6300
rect 26058 6244 26068 6300
rect 26124 6244 26134 6300
rect 28768 6244 28778 6300
rect 28834 6244 28882 6300
rect 28938 6244 28986 6300
rect 29042 6244 29052 6300
rect 8810 6132 8820 6188
rect 8876 6132 18564 6188
rect 18620 6132 18630 6188
rect 2314 6020 2324 6076
rect 2380 6020 2772 6076
rect 2828 6020 2838 6076
rect 4722 6020 4732 6076
rect 4788 6020 10668 6076
rect 10724 6020 10734 6076
rect 12842 6020 12852 6076
rect 12908 6020 13636 6076
rect 13692 6020 13702 6076
rect 7410 5908 7420 5964
rect 7476 5908 8372 5964
rect 8428 5908 8438 5964
rect 8810 5908 8820 5964
rect 8876 5908 8886 5964
rect 8820 5740 8876 5908
rect 13850 5796 13860 5852
rect 13916 5796 15540 5852
rect 15596 5796 15606 5852
rect 18778 5796 18788 5852
rect 18844 5796 19684 5852
rect 19740 5796 19750 5852
rect 20010 5796 20020 5852
rect 20076 5796 20580 5852
rect 20636 5796 23940 5852
rect 23996 5796 24006 5852
rect 25050 5796 25060 5852
rect 25116 5796 25844 5852
rect 25900 5796 25910 5852
rect 1474 5684 1484 5740
rect 1540 5684 1988 5740
rect 2044 5684 2054 5740
rect 2212 5684 2492 5740
rect 2548 5684 3444 5740
rect 3500 5684 7140 5740
rect 7196 5684 7206 5740
rect 8260 5684 8876 5740
rect 12730 5684 12740 5740
rect 12796 5684 13300 5740
rect 13356 5684 14140 5740
rect 14196 5684 14206 5740
rect 14634 5684 14644 5740
rect 14700 5684 16380 5740
rect 16436 5684 16446 5740
rect 0 5628 800 5656
rect 0 5572 1204 5628
rect 1260 5572 1270 5628
rect 0 5544 800 5572
rect 2212 5516 2268 5684
rect 8260 5516 8316 5684
rect 10938 5572 10948 5628
rect 11004 5572 24052 5628
rect 24108 5572 24118 5628
rect 1474 5460 1484 5516
rect 1540 5460 2268 5516
rect 2324 5460 4676 5516
rect 4732 5460 4742 5516
rect 5898 5460 5908 5516
rect 5964 5460 8260 5516
rect 8316 5460 8326 5516
rect 8918 5460 8928 5516
rect 8984 5460 9032 5516
rect 9088 5460 9136 5516
rect 9192 5460 9202 5516
rect 12170 5460 12180 5516
rect 12236 5460 14364 5516
rect 14420 5460 15372 5516
rect 15428 5460 16660 5516
rect 16716 5460 16726 5516
rect 16858 5460 16868 5516
rect 16924 5460 16972 5516
rect 17028 5460 17076 5516
rect 17132 5460 17142 5516
rect 24798 5460 24808 5516
rect 24864 5460 24912 5516
rect 24968 5460 25016 5516
rect 25072 5460 25082 5516
rect 2324 5404 2380 5460
rect 2146 5348 2156 5404
rect 2212 5348 2380 5404
rect 2538 5348 2548 5404
rect 2604 5348 5404 5404
rect 5460 5348 5470 5404
rect 1978 5236 1988 5292
rect 2044 5236 2996 5292
rect 3052 5236 3220 5292
rect 3276 5236 3286 5292
rect 3892 5236 4788 5292
rect 4844 5236 4854 5292
rect 6178 5236 6188 5292
rect 6244 5236 6916 5292
rect 6972 5236 6982 5292
rect 8474 5236 8484 5292
rect 8540 5236 8708 5292
rect 8764 5236 8774 5292
rect 19954 5236 19964 5292
rect 20020 5236 23436 5292
rect 23492 5236 23828 5292
rect 23884 5236 23894 5292
rect 3892 5180 3948 5236
rect 3826 5124 3836 5180
rect 3948 5124 3958 5180
rect 4442 5124 4452 5180
rect 4564 5124 4574 5180
rect 4666 5124 4676 5180
rect 4732 5124 5516 5180
rect 5572 5124 5582 5180
rect 7298 5124 7308 5180
rect 7364 5124 7812 5180
rect 7868 5124 7878 5180
rect 12282 5124 12292 5180
rect 12348 5124 14532 5180
rect 14588 5124 14598 5180
rect 14858 5124 14868 5180
rect 14924 5124 15596 5180
rect 15652 5124 15662 5180
rect 17322 5124 17332 5180
rect 17388 5124 18452 5180
rect 18508 5124 18788 5180
rect 18844 5124 18854 5180
rect 21326 5124 21364 5180
rect 21420 5124 23044 5180
rect 23100 5124 23110 5180
rect 14532 5068 14588 5124
rect 2874 5012 2884 5068
rect 2940 5012 4900 5068
rect 4956 5012 4966 5068
rect 8026 5012 8036 5068
rect 8092 5012 13300 5068
rect 13356 5012 14140 5068
rect 14532 5012 14980 5068
rect 15036 5012 15046 5068
rect 2370 4900 2380 4956
rect 2436 4900 3387 4956
rect 3658 4900 3668 4956
rect 3724 4900 5068 4956
rect 5124 4900 5134 4956
rect 5898 4900 5908 4956
rect 5964 4900 6748 4956
rect 6804 4900 6814 4956
rect 12506 4900 12516 4956
rect 12572 4900 13524 4956
rect 13580 4900 13590 4956
rect 14084 4900 14140 5012
rect 23044 4956 23100 5124
rect 33200 4956 34000 4984
rect 14196 4900 14868 4956
rect 14924 4900 14934 4956
rect 16650 4900 16660 4956
rect 16716 4900 17892 4956
rect 17948 4900 17958 4956
rect 18218 4900 18228 4956
rect 18284 4900 19180 4956
rect 19236 4900 19740 4956
rect 23044 4900 24388 4956
rect 24444 4900 24454 4956
rect 24602 4900 24612 4956
rect 24668 4900 25284 4956
rect 25340 4900 25350 4956
rect 31882 4900 31892 4956
rect 31948 4900 32340 4956
rect 32396 4900 34000 4956
rect 3331 4844 3387 4900
rect 3331 4788 4844 4844
rect 6066 4788 6076 4844
rect 6132 4788 7700 4844
rect 7756 4788 7924 4844
rect 7980 4788 8148 4844
rect 8204 4788 13468 4844
rect 14410 4788 14420 4844
rect 14476 4788 17444 4844
rect 17500 4788 17510 4844
rect 19684 4788 19740 4900
rect 33200 4872 34000 4900
rect 19796 4788 19806 4844
rect 22082 4788 22092 4844
rect 22148 4788 25620 4844
rect 25676 4788 25686 4844
rect 4788 4732 4844 4788
rect 13412 4732 13468 4788
rect 2202 4676 2212 4732
rect 2268 4676 2996 4732
rect 3052 4676 3062 4732
rect 3210 4676 3220 4732
rect 3276 4676 4452 4732
rect 4508 4676 4518 4732
rect 4778 4676 4788 4732
rect 4844 4676 4854 4732
rect 4948 4676 4958 4732
rect 5014 4676 5062 4732
rect 5118 4676 5166 4732
rect 5222 4676 5232 4732
rect 12888 4676 12898 4732
rect 12954 4676 13002 4732
rect 13058 4676 13106 4732
rect 13162 4676 13172 4732
rect 13402 4676 13412 4732
rect 13468 4676 14756 4732
rect 14812 4676 14822 4732
rect 16370 4676 16380 4732
rect 16436 4676 19516 4732
rect 19572 4676 19582 4732
rect 20828 4676 20838 4732
rect 20894 4676 20942 4732
rect 20998 4676 21046 4732
rect 21102 4676 21112 4732
rect 23762 4676 23772 4732
rect 23828 4676 26404 4732
rect 26460 4676 26470 4732
rect 28768 4676 28778 4732
rect 28834 4676 28882 4732
rect 28938 4676 28986 4732
rect 29042 4676 29052 4732
rect 1698 4564 1708 4620
rect 1764 4564 2100 4620
rect 2156 4564 3332 4620
rect 3388 4564 3464 4620
rect 3546 4564 3556 4620
rect 3612 4564 5348 4620
rect 5404 4564 5414 4620
rect 6514 4564 6524 4620
rect 6580 4564 7252 4620
rect 7308 4564 7318 4620
rect 10042 4564 10052 4620
rect 10108 4564 13804 4620
rect 13860 4564 13870 4620
rect 20346 4564 20356 4620
rect 20412 4564 21196 4620
rect 21252 4564 21262 4620
rect 2202 4452 2212 4508
rect 2268 4452 2548 4508
rect 2604 4452 4004 4508
rect 4060 4452 4070 4508
rect 6234 4452 6244 4508
rect 6300 4452 6860 4508
rect 6916 4452 6926 4508
rect 9864 4452 9940 4508
rect 9996 4452 10948 4508
rect 11004 4452 11014 4508
rect 12786 4452 12796 4508
rect 12852 4452 13972 4508
rect 14028 4452 14038 4508
rect 19618 4452 19628 4508
rect 19684 4452 20580 4508
rect 20636 4452 24724 4508
rect 24780 4452 25508 4508
rect 25564 4452 25574 4508
rect 0 4396 800 4424
rect 0 4340 1428 4396
rect 1484 4340 1494 4396
rect 2762 4340 2772 4396
rect 2828 4340 3444 4396
rect 3500 4340 3780 4396
rect 3836 4340 3846 4396
rect 7074 4340 7084 4396
rect 7140 4340 7364 4396
rect 7420 4340 7588 4396
rect 7644 4340 7654 4396
rect 14522 4340 14532 4396
rect 14588 4340 16548 4396
rect 16604 4340 16614 4396
rect 18330 4340 18340 4396
rect 18396 4340 20692 4396
rect 20748 4340 20758 4396
rect 0 4312 800 4340
rect 1474 4228 1484 4284
rect 1596 4228 1606 4284
rect 3322 4228 3332 4284
rect 3388 4228 7644 4284
rect 13066 4228 13076 4284
rect 13132 4228 13300 4284
rect 13356 4228 13412 4284
rect 13468 4228 13478 4284
rect 14690 4228 14700 4284
rect 14756 4228 14868 4284
rect 14924 4228 15876 4284
rect 15932 4228 17220 4284
rect 17276 4228 17286 4284
rect 7588 4172 7644 4228
rect 1698 4116 1708 4172
rect 1764 4116 6804 4172
rect 6860 4116 6870 4172
rect 7578 4116 7588 4172
rect 7644 4116 7654 4172
rect 10322 4116 10332 4172
rect 10388 4116 10668 4172
rect 10724 4116 11676 4172
rect 11732 4116 18564 4172
rect 18620 4116 18630 4172
rect 18778 4116 18788 4172
rect 18844 4116 20356 4172
rect 20412 4116 20422 4172
rect 22250 4116 22260 4172
rect 22316 4116 25396 4172
rect 25452 4116 25462 4172
rect 1530 4004 1540 4060
rect 1596 4004 3332 4060
rect 3388 4004 3398 4060
rect 6234 4004 6244 4060
rect 6300 4004 8764 4060
rect 9370 4004 9380 4060
rect 9436 4004 10052 4060
rect 10108 4004 10118 4060
rect 14186 4004 14196 4060
rect 14252 4004 14532 4060
rect 14588 4004 14598 4060
rect 25162 4004 25172 4060
rect 25228 4004 26012 4060
rect 26068 4004 26078 4060
rect 5786 3892 5796 3948
rect 5852 3892 7252 3948
rect 7308 3892 7318 3948
rect 8334 3892 8372 3948
rect 8428 3892 8438 3948
rect 8708 3836 8764 4004
rect 8918 3892 8928 3948
rect 8984 3892 9032 3948
rect 9088 3892 9136 3948
rect 9192 3892 9202 3948
rect 12394 3892 12404 3948
rect 12460 3892 13188 3948
rect 13244 3892 13254 3948
rect 16858 3892 16868 3948
rect 16924 3892 16972 3948
rect 17028 3892 17076 3948
rect 17132 3892 17142 3948
rect 24798 3892 24808 3948
rect 24864 3892 24912 3948
rect 24968 3892 25016 3948
rect 25072 3892 25082 3948
rect 2986 3780 2996 3836
rect 3052 3780 4116 3836
rect 4172 3780 4182 3836
rect 4330 3780 4340 3836
rect 4396 3780 4452 3836
rect 4508 3780 5180 3836
rect 6402 3780 6412 3836
rect 6468 3780 6916 3836
rect 6972 3780 6982 3836
rect 8708 3780 9492 3836
rect 9548 3780 9558 3836
rect 10612 3780 11284 3836
rect 11340 3780 11350 3836
rect 13458 3780 13468 3836
rect 13524 3780 14588 3836
rect 14644 3780 15932 3836
rect 15988 3780 15998 3836
rect 19786 3780 19796 3836
rect 19852 3780 20132 3836
rect 20188 3780 20198 3836
rect 1726 3668 1764 3724
rect 1820 3668 1830 3724
rect 2370 3668 2380 3724
rect 2436 3668 4788 3724
rect 4844 3668 4854 3724
rect 5124 3612 5180 3780
rect 10612 3724 10668 3780
rect 6682 3668 6692 3724
rect 6748 3668 10668 3724
rect 10826 3668 10836 3724
rect 10892 3668 12292 3724
rect 12348 3668 12358 3724
rect 15642 3668 15652 3724
rect 15708 3668 16548 3724
rect 16604 3668 16614 3724
rect 4778 3556 4788 3612
rect 4844 3556 4900 3612
rect 4956 3556 4966 3612
rect 5124 3556 6076 3612
rect 6132 3556 6692 3612
rect 6748 3556 6758 3612
rect 7466 3556 7476 3612
rect 7532 3556 9268 3612
rect 9324 3556 9334 3612
rect 9650 3556 9660 3612
rect 9716 3556 11732 3612
rect 11788 3556 11798 3612
rect 14298 3556 14308 3612
rect 14364 3556 16156 3612
rect 16212 3556 16222 3612
rect 1866 3444 1876 3500
rect 1932 3444 2436 3500
rect 2492 3444 2502 3500
rect 3882 3444 3892 3500
rect 3948 3444 4116 3500
rect 4172 3444 6300 3500
rect 6356 3444 6804 3500
rect 6860 3444 6870 3500
rect 7018 3444 7028 3500
rect 7084 3444 10164 3500
rect 10220 3444 10230 3500
rect 15082 3444 15092 3500
rect 15148 3444 15540 3500
rect 15596 3444 19796 3500
rect 19852 3444 19862 3500
rect 20458 3444 20468 3500
rect 20524 3444 20916 3500
rect 20972 3444 20982 3500
rect 4778 3332 4788 3388
rect 4844 3332 4956 3388
rect 7578 3332 7588 3388
rect 7644 3332 8260 3388
rect 8316 3332 8326 3388
rect 9482 3332 9492 3388
rect 9548 3332 11116 3388
rect 11172 3332 13748 3388
rect 13804 3332 13814 3388
rect 21812 3332 24724 3388
rect 24780 3332 25844 3388
rect 25900 3332 25910 3388
rect 4900 3276 4956 3332
rect 21812 3276 21868 3332
rect 4900 3220 5348 3276
rect 5404 3220 5414 3276
rect 5786 3220 5796 3276
rect 5852 3220 6356 3276
rect 6412 3220 6422 3276
rect 21802 3220 21812 3276
rect 21868 3220 21878 3276
rect 0 3164 800 3192
rect 0 3108 1316 3164
rect 1372 3108 1382 3164
rect 4948 3108 4958 3164
rect 5014 3108 5062 3164
rect 5118 3108 5166 3164
rect 5222 3108 5232 3164
rect 7130 3108 7140 3164
rect 7196 3108 7812 3164
rect 7868 3108 7878 3164
rect 12888 3108 12898 3164
rect 12954 3108 13002 3164
rect 13058 3108 13106 3164
rect 13162 3108 13172 3164
rect 20828 3108 20838 3164
rect 20894 3108 20942 3164
rect 20998 3108 21046 3164
rect 21102 3108 21112 3164
rect 28768 3108 28778 3164
rect 28834 3108 28882 3164
rect 28938 3108 28986 3164
rect 29042 3108 29052 3164
rect 0 3080 800 3108
rect 24826 2884 24836 2940
rect 24892 2884 25620 2940
rect 25676 2884 25686 2940
rect 4302 2772 4340 2828
rect 4396 2772 4406 2828
rect 5338 2772 5348 2828
rect 5404 2772 5796 2828
rect 5852 2772 5862 2828
rect 6906 2772 6916 2828
rect 6972 2772 8652 2828
rect 8708 2772 9156 2828
rect 9212 2772 9604 2828
rect 9660 2772 9670 2828
rect 13458 2772 13468 2828
rect 13524 2772 14868 2828
rect 14924 2772 14934 2828
rect 18666 2772 18676 2828
rect 18732 2772 19628 2828
rect 19684 2716 19740 2828
rect 20010 2772 20020 2828
rect 20076 2772 20580 2828
rect 20636 2772 20646 2828
rect 4778 2660 4788 2716
rect 4844 2660 6804 2716
rect 6860 2660 6870 2716
rect 7018 2660 7028 2716
rect 7084 2660 8876 2716
rect 8932 2660 9940 2716
rect 9996 2660 19236 2716
rect 19292 2660 19302 2716
rect 19684 2660 19908 2716
rect 19964 2660 20187 2716
rect 20131 2604 20187 2660
rect 858 2548 868 2604
rect 924 2548 3220 2604
rect 3276 2548 3286 2604
rect 4554 2548 4564 2604
rect 4620 2548 7700 2604
rect 7756 2548 7766 2604
rect 15866 2548 15876 2604
rect 15932 2548 19012 2604
rect 19068 2548 19078 2604
rect 20131 2548 21252 2604
rect 21308 2548 21318 2604
rect 24154 2548 24164 2604
rect 24220 2548 25060 2604
rect 25116 2548 25126 2604
rect 21252 2492 21308 2548
rect 2650 2436 2660 2492
rect 2716 2436 6916 2492
rect 6972 2436 7196 2492
rect 7252 2436 7262 2492
rect 21252 2436 24332 2492
rect 24388 2436 25172 2492
rect 25228 2436 25676 2492
rect 25732 2436 25742 2492
rect 3322 2324 3332 2380
rect 3388 2324 4004 2380
rect 4060 2324 5572 2380
rect 5628 2324 5638 2380
rect 8918 2324 8928 2380
rect 8984 2324 9032 2380
rect 9088 2324 9136 2380
rect 9192 2324 9202 2380
rect 16858 2324 16868 2380
rect 16924 2324 16972 2380
rect 17028 2324 17076 2380
rect 17132 2324 17142 2380
rect 20346 2324 20356 2380
rect 20412 2324 20692 2380
rect 20748 2324 20758 2380
rect 24798 2324 24808 2380
rect 24864 2324 24912 2380
rect 24968 2324 25016 2380
rect 25072 2324 25082 2380
rect 6346 2212 6356 2268
rect 6412 2212 7252 2268
rect 7308 2212 7318 2268
rect 12058 2212 12068 2268
rect 12124 2212 13076 2268
rect 13132 2212 13142 2268
rect 23258 2212 23268 2268
rect 23324 2212 25396 2268
rect 25452 2212 25462 2268
rect 4778 2100 4788 2156
rect 4844 2100 5460 2156
rect 5516 2100 11508 2156
rect 11564 2100 14084 2156
rect 14140 2100 14150 2156
rect 17266 2100 17276 2156
rect 17332 2100 18564 2156
rect 18620 2100 18630 2156
rect 19114 2100 19124 2156
rect 19180 2100 25620 2156
rect 25676 2100 25686 2156
rect 6794 1988 6804 2044
rect 6860 1988 7924 2044
rect 7980 1988 12068 2044
rect 12124 1988 12134 2044
rect 12394 1988 12404 2044
rect 12460 1988 18172 2044
rect 18330 1988 18340 2044
rect 18396 1988 19012 2044
rect 19068 1988 19078 2044
rect 23090 1988 23100 2044
rect 23156 1988 23772 2044
rect 23828 1988 23838 2044
rect 0 1932 800 1960
rect 0 1876 1596 1932
rect 2426 1876 2436 1932
rect 2492 1876 5796 1932
rect 5852 1876 6132 1932
rect 6188 1876 7700 1932
rect 7756 1876 7766 1932
rect 9594 1876 9604 1932
rect 9660 1876 12740 1932
rect 12796 1876 13300 1932
rect 13356 1876 13366 1932
rect 15091 1876 15204 1932
rect 15260 1876 15270 1932
rect 0 1848 800 1876
rect 1540 1596 1596 1876
rect 15091 1820 15147 1876
rect 4442 1764 4452 1820
rect 4508 1764 6972 1820
rect 7028 1764 8148 1820
rect 8204 1764 15147 1820
rect 15390 1764 15428 1820
rect 15484 1764 16604 1820
rect 16660 1764 16884 1820
rect 16940 1764 16950 1820
rect 18116 1708 18172 1988
rect 22362 1876 22372 1932
rect 22428 1876 23380 1932
rect 23436 1876 24052 1932
rect 24108 1876 24118 1932
rect 33200 1708 34000 1736
rect 10826 1652 10836 1708
rect 10892 1652 13860 1708
rect 13916 1652 13926 1708
rect 18116 1652 18508 1708
rect 21466 1652 21476 1708
rect 21532 1652 22372 1708
rect 22428 1652 22438 1708
rect 23258 1652 23268 1708
rect 23324 1652 23940 1708
rect 23996 1652 24006 1708
rect 31826 1652 31836 1708
rect 31892 1652 32340 1708
rect 32396 1652 34000 1708
rect 18452 1596 18508 1652
rect 33200 1624 34000 1652
rect 1540 1540 2548 1596
rect 2604 1540 2614 1596
rect 4948 1540 4958 1596
rect 5014 1540 5062 1596
rect 5118 1540 5166 1596
rect 5222 1540 5232 1596
rect 8474 1540 8484 1596
rect 8540 1540 10724 1596
rect 10780 1540 10790 1596
rect 12888 1540 12898 1596
rect 12954 1540 13002 1596
rect 13058 1540 13106 1596
rect 13162 1540 13172 1596
rect 15306 1540 15316 1596
rect 15372 1540 17220 1596
rect 17276 1540 17286 1596
rect 18442 1540 18452 1596
rect 18508 1540 18518 1596
rect 20828 1540 20838 1596
rect 20894 1540 20942 1596
rect 20998 1540 21046 1596
rect 21102 1540 21112 1596
rect 28768 1540 28778 1596
rect 28834 1540 28882 1596
rect 28938 1540 28986 1596
rect 29042 1540 29052 1596
rect 21746 1428 21756 1484
rect 21812 1428 22596 1484
rect 22652 1428 22662 1484
rect 8810 1316 8820 1372
rect 8876 1316 12180 1372
rect 12236 1316 12246 1372
rect 16202 1316 16212 1372
rect 16268 1316 17780 1372
rect 17836 1316 17846 1372
rect 18106 1316 18116 1372
rect 18172 1316 22484 1372
rect 22540 1316 22550 1372
rect 1194 1204 1204 1260
rect 1260 1204 3387 1260
rect 12730 1204 12740 1260
rect 12796 1204 13356 1260
rect 13412 1204 13748 1260
rect 13804 1204 13814 1260
rect 21914 1204 21924 1260
rect 21980 1204 22708 1260
rect 22764 1204 22774 1260
rect 3331 1148 3387 1204
rect 3331 1092 4676 1148
rect 4732 1092 8092 1148
rect 8148 1092 8158 1148
rect 10490 1092 10500 1148
rect 10556 1092 14476 1148
rect 14532 1092 14542 1148
rect 15166 1092 15204 1148
rect 15260 1092 15270 1148
rect 19114 1092 19124 1148
rect 19180 1092 22036 1148
rect 22092 1092 22102 1148
rect 15204 1036 15260 1092
rect 11386 980 11396 1036
rect 11452 980 11956 1036
rect 12012 980 15260 1036
rect 19674 980 19684 1036
rect 19796 980 19806 1036
rect 25498 980 25508 1036
rect 25564 980 25956 1036
rect 26012 980 26236 1036
rect 26292 980 26302 1036
rect 8918 756 8928 812
rect 8984 756 9032 812
rect 9088 756 9136 812
rect 9192 756 9202 812
rect 16858 756 16868 812
rect 16924 756 16972 812
rect 17028 756 17076 812
rect 17132 756 17142 812
rect 24798 756 24808 812
rect 24864 756 24912 812
rect 24968 756 25016 812
rect 25072 756 25082 812
rect 0 700 800 728
rect 0 644 868 700
rect 924 644 934 700
rect 0 616 800 644
<< via3 >>
rect 4958 18788 5014 18844
rect 5062 18788 5118 18844
rect 5166 18788 5222 18844
rect 12898 18788 12954 18844
rect 13002 18788 13058 18844
rect 13106 18788 13162 18844
rect 20838 18788 20894 18844
rect 20942 18788 20998 18844
rect 21046 18788 21102 18844
rect 28778 18788 28834 18844
rect 28882 18788 28938 18844
rect 28986 18788 29042 18844
rect 13300 18340 13356 18396
rect 18452 18340 18508 18396
rect 4340 18228 4396 18284
rect 2548 18116 2604 18172
rect 4116 18116 4172 18172
rect 8928 18004 8984 18060
rect 9032 18004 9088 18060
rect 9136 18004 9192 18060
rect 16868 18004 16924 18060
rect 16972 18004 17028 18060
rect 17076 18004 17132 18060
rect 24808 18004 24864 18060
rect 24912 18004 24968 18060
rect 25016 18004 25072 18060
rect 3780 17556 3836 17612
rect 4958 17220 5014 17276
rect 5062 17220 5118 17276
rect 5166 17220 5222 17276
rect 12898 17220 12954 17276
rect 13002 17220 13058 17276
rect 13106 17220 13162 17276
rect 20838 17220 20894 17276
rect 20942 17220 20998 17276
rect 21046 17220 21102 17276
rect 28778 17220 28834 17276
rect 28882 17220 28938 17276
rect 28986 17220 29042 17276
rect 4788 16996 4844 17052
rect 6356 16996 6412 17052
rect 18116 16884 18172 16940
rect 12740 16660 12796 16716
rect 16548 16660 16604 16716
rect 8928 16436 8984 16492
rect 9032 16436 9088 16492
rect 9136 16436 9192 16492
rect 13300 16436 13356 16492
rect 16868 16436 16924 16492
rect 16972 16436 17028 16492
rect 17076 16436 17132 16492
rect 24808 16436 24864 16492
rect 24912 16436 24968 16492
rect 25016 16436 25072 16492
rect 8484 16324 8540 16380
rect 22260 16324 22316 16380
rect 10052 16212 10108 16268
rect 11172 16212 11228 16268
rect 12740 16212 12796 16268
rect 14756 16212 14812 16268
rect 15428 16212 15484 16268
rect 22820 16212 22876 16268
rect 8484 16100 8540 16156
rect 11620 16100 11676 16156
rect 18340 16100 18396 16156
rect 23716 16100 23772 16156
rect 11396 15988 11452 16044
rect 16548 15988 16604 16044
rect 7588 15876 7644 15932
rect 24612 15876 24668 15932
rect 17556 15764 17612 15820
rect 22820 15764 22876 15820
rect 4958 15652 5014 15708
rect 5062 15652 5118 15708
rect 5166 15652 5222 15708
rect 12898 15652 12954 15708
rect 13002 15652 13058 15708
rect 13106 15652 13162 15708
rect 20838 15652 20894 15708
rect 20942 15652 20998 15708
rect 21046 15652 21102 15708
rect 22484 15652 22540 15708
rect 28778 15652 28834 15708
rect 28882 15652 28938 15708
rect 28986 15652 29042 15708
rect 18564 15540 18620 15596
rect 21476 15540 21532 15596
rect 12516 15428 12572 15484
rect 16100 15428 16156 15484
rect 23044 15428 23100 15484
rect 24500 15428 24556 15484
rect 14644 15316 14700 15372
rect 15204 15316 15260 15372
rect 15428 15204 15484 15260
rect 18676 15204 18732 15260
rect 21252 15204 21308 15260
rect 16100 15092 16156 15148
rect 19796 15092 19852 15148
rect 10948 14980 11004 15036
rect 11396 14980 11452 15036
rect 14532 14980 14588 15036
rect 21252 14980 21308 15036
rect 8928 14868 8984 14924
rect 9032 14868 9088 14924
rect 9136 14868 9192 14924
rect 11508 14868 11564 14924
rect 16868 14868 16924 14924
rect 16972 14868 17028 14924
rect 17076 14868 17132 14924
rect 18564 14868 18620 14924
rect 19908 14868 19964 14924
rect 24808 14868 24864 14924
rect 24912 14868 24968 14924
rect 25016 14868 25072 14924
rect 12180 14756 12236 14812
rect 12740 14644 12796 14700
rect 18452 14644 18508 14700
rect 19796 14644 19852 14700
rect 21476 14644 21532 14700
rect 27636 14644 27692 14700
rect 18452 14420 18508 14476
rect 14084 14308 14140 14364
rect 14532 14308 14588 14364
rect 21476 14308 21532 14364
rect 18564 14196 18620 14252
rect 4958 14084 5014 14140
rect 5062 14084 5118 14140
rect 5166 14084 5222 14140
rect 12898 14084 12954 14140
rect 13002 14084 13058 14140
rect 13106 14084 13162 14140
rect 20838 14084 20894 14140
rect 20942 14084 20998 14140
rect 21046 14084 21102 14140
rect 28778 14084 28834 14140
rect 28882 14084 28938 14140
rect 28986 14084 29042 14140
rect 26852 13860 26908 13916
rect 8148 13636 8204 13692
rect 20468 13636 20524 13692
rect 22260 13636 22316 13692
rect 3668 13524 3724 13580
rect 10948 13524 11004 13580
rect 13300 13524 13356 13580
rect 8928 13300 8984 13356
rect 9032 13300 9088 13356
rect 9136 13300 9192 13356
rect 11620 13300 11676 13356
rect 14756 13300 14812 13356
rect 16868 13300 16924 13356
rect 16972 13300 17028 13356
rect 17076 13300 17132 13356
rect 24808 13300 24864 13356
rect 24912 13300 24968 13356
rect 25016 13300 25072 13356
rect 7588 13076 7644 13132
rect 22932 13076 22988 13132
rect 14532 12852 14588 12908
rect 22484 12852 22540 12908
rect 24500 12852 24556 12908
rect 18788 12740 18844 12796
rect 19908 12628 19964 12684
rect 4958 12516 5014 12572
rect 5062 12516 5118 12572
rect 5166 12516 5222 12572
rect 12898 12516 12954 12572
rect 13002 12516 13058 12572
rect 13106 12516 13162 12572
rect 13636 12516 13692 12572
rect 20838 12516 20894 12572
rect 20942 12516 20998 12572
rect 21046 12516 21102 12572
rect 28778 12516 28834 12572
rect 28882 12516 28938 12572
rect 28986 12516 29042 12572
rect 11508 12404 11564 12460
rect 13412 12404 13468 12460
rect 14532 12404 14588 12460
rect 17780 12404 17836 12460
rect 18676 12404 18732 12460
rect 18900 12404 18956 12460
rect 11620 12068 11676 12124
rect 17780 12068 17836 12124
rect 24500 12068 24556 12124
rect 9940 11844 9996 11900
rect 15204 11844 15260 11900
rect 16660 11844 16716 11900
rect 8928 11732 8984 11788
rect 9032 11732 9088 11788
rect 9136 11732 9192 11788
rect 14644 11732 14700 11788
rect 16868 11732 16924 11788
rect 16972 11732 17028 11788
rect 17076 11732 17132 11788
rect 24808 11732 24864 11788
rect 24912 11732 24968 11788
rect 25016 11732 25072 11788
rect 17220 11620 17276 11676
rect 18004 11620 18060 11676
rect 10948 11508 11004 11564
rect 7588 11172 7644 11228
rect 4958 10948 5014 11004
rect 5062 10948 5118 11004
rect 5166 10948 5222 11004
rect 9940 10948 9996 11004
rect 12898 10948 12954 11004
rect 13002 10948 13058 11004
rect 13106 10948 13162 11004
rect 20838 10948 20894 11004
rect 20942 10948 20998 11004
rect 21046 10948 21102 11004
rect 28778 10948 28834 11004
rect 28882 10948 28938 11004
rect 28986 10948 29042 11004
rect 8260 10500 8316 10556
rect 13636 10500 13692 10556
rect 18228 10500 18284 10556
rect 23492 10388 23548 10444
rect 5460 10164 5516 10220
rect 8928 10164 8984 10220
rect 9032 10164 9088 10220
rect 9136 10164 9192 10220
rect 16868 10164 16924 10220
rect 16972 10164 17028 10220
rect 17076 10164 17132 10220
rect 24808 10164 24864 10220
rect 24912 10164 24968 10220
rect 25016 10164 25072 10220
rect 4116 9940 4172 9996
rect 13412 9940 13468 9996
rect 7588 9828 7644 9884
rect 5348 9716 5404 9772
rect 4958 9380 5014 9436
rect 5062 9380 5118 9436
rect 5166 9380 5222 9436
rect 12898 9380 12954 9436
rect 13002 9380 13058 9436
rect 13106 9380 13162 9436
rect 20838 9380 20894 9436
rect 20942 9380 20998 9436
rect 21046 9380 21102 9436
rect 28778 9380 28834 9436
rect 28882 9380 28938 9436
rect 28986 9380 29042 9436
rect 22260 9156 22316 9212
rect 18116 8820 18172 8876
rect 8928 8596 8984 8652
rect 9032 8596 9088 8652
rect 9136 8596 9192 8652
rect 16868 8596 16924 8652
rect 16972 8596 17028 8652
rect 17076 8596 17132 8652
rect 24808 8596 24864 8652
rect 24912 8596 24968 8652
rect 25016 8596 25072 8652
rect 5460 8260 5516 8316
rect 4340 8036 4396 8092
rect 4958 7812 5014 7868
rect 5062 7812 5118 7868
rect 5166 7812 5222 7868
rect 12898 7812 12954 7868
rect 13002 7812 13058 7868
rect 13106 7812 13162 7868
rect 20838 7812 20894 7868
rect 20942 7812 20998 7868
rect 21046 7812 21102 7868
rect 28778 7812 28834 7868
rect 28882 7812 28938 7868
rect 28986 7812 29042 7868
rect 8148 7700 8204 7756
rect 9940 7700 9996 7756
rect 1316 7588 1372 7644
rect 1764 7476 1820 7532
rect 17780 7476 17836 7532
rect 10948 7364 11004 7420
rect 19684 7364 19740 7420
rect 7700 7252 7756 7308
rect 1428 7140 1484 7196
rect 8928 7028 8984 7084
rect 9032 7028 9088 7084
rect 9136 7028 9192 7084
rect 16868 7028 16924 7084
rect 16972 7028 17028 7084
rect 17076 7028 17132 7084
rect 24808 7028 24864 7084
rect 24912 7028 24968 7084
rect 25016 7028 25072 7084
rect 3444 6804 3500 6860
rect 7028 6804 7084 6860
rect 14420 6692 14476 6748
rect 6916 6468 6972 6524
rect 4958 6244 5014 6300
rect 5062 6244 5118 6300
rect 5166 6244 5222 6300
rect 12898 6244 12954 6300
rect 13002 6244 13058 6300
rect 13106 6244 13162 6300
rect 20838 6244 20894 6300
rect 20942 6244 20998 6300
rect 21046 6244 21102 6300
rect 28778 6244 28834 6300
rect 28882 6244 28938 6300
rect 28986 6244 29042 6300
rect 1204 5572 1260 5628
rect 8928 5460 8984 5516
rect 9032 5460 9088 5516
rect 9136 5460 9192 5516
rect 16868 5460 16924 5516
rect 16972 5460 17028 5516
rect 17076 5460 17132 5516
rect 24808 5460 24864 5516
rect 24912 5460 24968 5516
rect 25016 5460 25072 5516
rect 3892 5124 3948 5180
rect 4452 5124 4508 5180
rect 21364 5124 21420 5180
rect 13300 5012 13356 5068
rect 14420 4788 14476 4844
rect 4958 4676 5014 4732
rect 5062 4676 5118 4732
rect 5166 4676 5222 4732
rect 12898 4676 12954 4732
rect 13002 4676 13058 4732
rect 13106 4676 13162 4732
rect 20838 4676 20894 4732
rect 20942 4676 20998 4732
rect 21046 4676 21102 4732
rect 28778 4676 28834 4732
rect 28882 4676 28938 4732
rect 28986 4676 29042 4732
rect 3332 4564 3388 4620
rect 9940 4452 9996 4508
rect 1428 4340 1484 4396
rect 3444 4340 3500 4396
rect 1540 4228 1596 4284
rect 3332 4228 3388 4284
rect 13300 4228 13356 4284
rect 8372 3892 8428 3948
rect 8928 3892 8984 3948
rect 9032 3892 9088 3948
rect 9136 3892 9192 3948
rect 16868 3892 16924 3948
rect 16972 3892 17028 3948
rect 17076 3892 17132 3948
rect 24808 3892 24864 3948
rect 24912 3892 24968 3948
rect 25016 3892 25072 3948
rect 4452 3780 4508 3836
rect 1764 3668 1820 3724
rect 4788 3556 4844 3612
rect 6692 3556 6748 3612
rect 3892 3444 3948 3500
rect 6804 3444 6860 3500
rect 20468 3444 20524 3500
rect 4788 3332 4844 3388
rect 1316 3108 1372 3164
rect 4958 3108 5014 3164
rect 5062 3108 5118 3164
rect 5166 3108 5222 3164
rect 12898 3108 12954 3164
rect 13002 3108 13058 3164
rect 13106 3108 13162 3164
rect 20838 3108 20894 3164
rect 20942 3108 20998 3164
rect 21046 3108 21102 3164
rect 28778 3108 28834 3164
rect 28882 3108 28938 3164
rect 28986 3108 29042 3164
rect 4340 2772 4396 2828
rect 6916 2436 6972 2492
rect 8928 2324 8984 2380
rect 9032 2324 9088 2380
rect 9136 2324 9192 2380
rect 16868 2324 16924 2380
rect 16972 2324 17028 2380
rect 17076 2324 17132 2380
rect 24808 2324 24864 2380
rect 24912 2324 24968 2380
rect 25016 2324 25072 2380
rect 15428 1764 15484 1820
rect 4958 1540 5014 1596
rect 5062 1540 5118 1596
rect 5166 1540 5222 1596
rect 12898 1540 12954 1596
rect 13002 1540 13058 1596
rect 13106 1540 13162 1596
rect 20838 1540 20894 1596
rect 20942 1540 20998 1596
rect 21046 1540 21102 1596
rect 28778 1540 28834 1596
rect 28882 1540 28938 1596
rect 28986 1540 29042 1596
rect 1204 1204 1260 1260
rect 12740 1204 12796 1260
rect 15204 1092 15260 1148
rect 19684 980 19740 1036
rect 8928 756 8984 812
rect 9032 756 9088 812
rect 9136 756 9192 812
rect 16868 756 16924 812
rect 16972 756 17028 812
rect 17076 756 17132 812
rect 24808 756 24864 812
rect 24912 756 24968 812
rect 25016 756 25072 812
<< metal4 >>
rect 4930 18844 5250 18876
rect 4930 18788 4958 18844
rect 5014 18788 5062 18844
rect 5118 18788 5166 18844
rect 5222 18788 5250 18844
rect 4340 18388 4396 18398
rect 4340 18284 4396 18332
rect 4340 18218 4396 18228
rect 2548 18172 2604 18182
rect 2548 16408 2604 18116
rect 4116 18172 4172 18182
rect 2548 16342 2604 16352
rect 3780 17612 3836 17622
rect 3780 15148 3836 17556
rect 3668 15092 3780 15147
rect 3668 15091 3836 15092
rect 3668 13580 3724 15091
rect 3780 15082 3836 15091
rect 3668 13514 3724 13524
rect 4116 9996 4172 18116
rect 4930 17276 5250 18788
rect 8900 18060 9220 18876
rect 8900 18004 8928 18060
rect 8984 18004 9032 18060
rect 9088 18004 9136 18060
rect 9192 18004 9220 18060
rect 4930 17220 4958 17276
rect 5014 17220 5062 17276
rect 5118 17220 5166 17276
rect 5222 17220 5250 17276
rect 4788 17052 4844 17062
rect 4788 16228 4844 16996
rect 4788 16162 4844 16172
rect 4930 17044 5250 17220
rect 4930 16988 4958 17044
rect 5014 16988 5062 17044
rect 5118 16988 5166 17044
rect 5222 16988 5250 17044
rect 4930 16940 5250 16988
rect 6356 17308 6412 17318
rect 6356 17052 6412 17252
rect 6356 16986 6412 16996
rect 4930 16884 4958 16940
rect 5014 16884 5062 16940
rect 5118 16884 5166 16940
rect 5222 16884 5250 16940
rect 4930 16836 5250 16884
rect 4930 16780 4958 16836
rect 5014 16780 5062 16836
rect 5118 16780 5166 16836
rect 5222 16780 5250 16836
rect 4116 9930 4172 9940
rect 4930 15708 5250 16780
rect 8900 16492 9220 18004
rect 12870 18844 13190 18876
rect 12870 18788 12898 18844
rect 12954 18788 13002 18844
rect 13058 18788 13106 18844
rect 13162 18788 13190 18844
rect 12870 17276 13190 18788
rect 12870 17220 12898 17276
rect 12954 17220 13002 17276
rect 13058 17220 13106 17276
rect 13162 17220 13190 17276
rect 12870 17044 13190 17220
rect 12870 16988 12898 17044
rect 12954 16988 13002 17044
rect 13058 16988 13106 17044
rect 13162 16988 13190 17044
rect 12870 16940 13190 16988
rect 12870 16884 12898 16940
rect 12954 16884 13002 16940
rect 13058 16884 13106 16940
rect 13162 16884 13190 16940
rect 12870 16836 13190 16884
rect 12870 16780 12898 16836
rect 12954 16780 13002 16836
rect 13058 16780 13106 16836
rect 13162 16780 13190 16836
rect 8900 16436 8928 16492
rect 8984 16436 9032 16492
rect 9088 16436 9136 16492
rect 9192 16436 9220 16492
rect 8484 16380 8540 16390
rect 8484 16156 8540 16324
rect 8484 16090 8540 16100
rect 4930 15652 4958 15708
rect 5014 15652 5062 15708
rect 5118 15652 5166 15708
rect 5222 15652 5250 15708
rect 4930 14140 5250 15652
rect 4930 14084 4958 14140
rect 5014 14084 5062 14140
rect 5118 14084 5166 14140
rect 5222 14084 5250 14140
rect 4930 12572 5250 14084
rect 7588 15932 7644 15942
rect 7588 13132 7644 15876
rect 8900 14924 9220 16436
rect 12740 16716 12796 16726
rect 10052 16408 10108 16418
rect 10052 16268 10108 16352
rect 10052 16202 10108 16212
rect 11172 16268 11228 16278
rect 11172 16048 11228 16212
rect 12740 16268 12796 16660
rect 12740 16202 12796 16212
rect 11620 16156 11676 16166
rect 11172 15982 11228 15992
rect 11396 16044 11452 16054
rect 8900 14868 8928 14924
rect 8984 14868 9032 14924
rect 9088 14868 9136 14924
rect 9192 14868 9220 14924
rect 8900 14740 9220 14868
rect 8900 14684 8928 14740
rect 8984 14684 9032 14740
rect 9088 14684 9136 14740
rect 9192 14684 9220 14740
rect 8900 14636 9220 14684
rect 8900 14580 8928 14636
rect 8984 14580 9032 14636
rect 9088 14580 9136 14636
rect 9192 14580 9220 14636
rect 8900 14532 9220 14580
rect 8900 14476 8928 14532
rect 8984 14476 9032 14532
rect 9088 14476 9136 14532
rect 9192 14476 9220 14532
rect 7588 13066 7644 13076
rect 8148 13692 8204 13702
rect 4930 12516 4958 12572
rect 5014 12516 5062 12572
rect 5118 12516 5166 12572
rect 5222 12516 5250 12572
rect 4930 12436 5250 12516
rect 4930 12380 4958 12436
rect 5014 12380 5062 12436
rect 5118 12380 5166 12436
rect 5222 12380 5250 12436
rect 4930 12332 5250 12380
rect 4930 12276 4958 12332
rect 5014 12276 5062 12332
rect 5118 12276 5166 12332
rect 5222 12276 5250 12332
rect 4930 12228 5250 12276
rect 4930 12172 4958 12228
rect 5014 12172 5062 12228
rect 5118 12172 5166 12228
rect 5222 12172 5250 12228
rect 4930 11004 5250 12172
rect 4930 10948 4958 11004
rect 5014 10948 5062 11004
rect 5118 10948 5166 11004
rect 5222 10948 5250 11004
rect 4930 9436 5250 10948
rect 7588 11228 7644 11238
rect 5460 10220 5516 10230
rect 5348 9772 5404 9782
rect 5348 9568 5404 9716
rect 5348 9502 5404 9512
rect 4930 9380 4958 9436
rect 5014 9380 5062 9436
rect 5118 9380 5166 9436
rect 5222 9380 5250 9436
rect 4340 8092 4396 8102
rect 1316 7644 1372 7654
rect 1204 5628 1260 5638
rect 1204 1260 1260 5572
rect 1316 3164 1372 7588
rect 1764 7532 1820 7542
rect 1428 7196 1484 7206
rect 1428 4396 1484 7140
rect 1428 4330 1484 4340
rect 1540 4284 1596 4294
rect 1540 3988 1596 4228
rect 1540 3922 1596 3932
rect 1764 3724 1820 7476
rect 3444 6860 3500 6870
rect 3332 4620 3388 4630
rect 3332 4284 3388 4564
rect 3444 4396 3500 6804
rect 3444 4330 3500 4340
rect 3892 5180 3948 5190
rect 3332 4218 3388 4228
rect 1764 3658 1820 3668
rect 3892 3500 3948 5124
rect 3892 3434 3948 3444
rect 1316 3098 1372 3108
rect 4340 2828 4396 8036
rect 4930 7868 5250 9380
rect 5460 8316 5516 10164
rect 7588 9884 7644 11172
rect 7588 9818 7644 9828
rect 5460 8250 5516 8260
rect 4930 7772 4958 7868
rect 5014 7772 5062 7868
rect 5118 7772 5166 7868
rect 5222 7772 5250 7868
rect 4930 7724 5250 7772
rect 4930 7668 4958 7724
rect 5014 7668 5062 7724
rect 5118 7668 5166 7724
rect 5222 7668 5250 7724
rect 8148 7756 8204 13636
rect 8900 13356 9220 14476
rect 8900 13300 8928 13356
rect 8984 13300 9032 13356
rect 9088 13300 9136 13356
rect 9192 13300 9220 13356
rect 8900 11788 9220 13300
rect 10948 15036 11004 15046
rect 10948 13580 11004 14980
rect 11396 15036 11452 15988
rect 11396 14970 11452 14980
rect 8900 11732 8928 11788
rect 8984 11732 9032 11788
rect 9088 11732 9136 11788
rect 9192 11732 9220 11788
rect 8260 10648 8316 10658
rect 8260 10556 8316 10592
rect 8260 10490 8316 10500
rect 8148 7690 8204 7700
rect 8900 10220 9220 11732
rect 9940 11900 9996 11910
rect 9940 11004 9996 11844
rect 9940 10938 9996 10948
rect 10948 11564 11004 13524
rect 11508 14924 11564 14934
rect 11508 12460 11564 14868
rect 11620 13356 11676 16100
rect 12870 15708 13190 16780
rect 13300 18396 13356 18406
rect 13300 16588 13356 18340
rect 16840 18060 17160 18876
rect 20810 18844 21130 18876
rect 20810 18788 20838 18844
rect 20894 18788 20942 18844
rect 20998 18788 21046 18844
rect 21102 18788 21130 18844
rect 18452 18396 18508 18406
rect 18452 18302 18508 18332
rect 16840 18004 16868 18060
rect 16924 18004 16972 18060
rect 17028 18004 17076 18060
rect 17132 18004 17160 18060
rect 13300 16492 13356 16532
rect 13300 16426 13356 16436
rect 16548 16716 16604 16726
rect 12870 15652 12898 15708
rect 12954 15652 13002 15708
rect 13058 15652 13106 15708
rect 13162 15652 13190 15708
rect 12516 15508 12572 15522
rect 12516 15418 12572 15428
rect 12740 15148 12796 15158
rect 12180 14968 12236 14978
rect 12180 14812 12236 14912
rect 12180 14746 12236 14756
rect 12740 14700 12796 15092
rect 12740 14634 12796 14644
rect 11620 13290 11676 13300
rect 12870 14140 13190 15652
rect 14756 16268 14812 16278
rect 14644 15372 14700 15382
rect 14532 15036 14588 15046
rect 12870 14084 12898 14140
rect 12954 14084 13002 14140
rect 13058 14084 13106 14140
rect 13162 14084 13190 14140
rect 11508 12394 11564 12404
rect 12870 12572 13190 14084
rect 14084 14364 14140 14374
rect 12870 12516 12898 12572
rect 12954 12516 13002 12572
rect 13058 12516 13106 12572
rect 13162 12516 13190 12572
rect 12870 12436 13190 12516
rect 12870 12380 12898 12436
rect 12954 12380 13002 12436
rect 13058 12380 13106 12436
rect 13162 12380 13190 12436
rect 12870 12332 13190 12380
rect 12870 12276 12898 12332
rect 12954 12276 13002 12332
rect 13058 12276 13106 12332
rect 13162 12276 13190 12332
rect 12870 12228 13190 12276
rect 12870 12172 12898 12228
rect 12954 12172 13002 12228
rect 13058 12172 13106 12228
rect 13162 12172 13190 12228
rect 8900 10164 8928 10220
rect 8984 10164 9032 10220
rect 9088 10164 9136 10220
rect 9192 10164 9220 10220
rect 8900 10132 9220 10164
rect 8900 10076 8928 10132
rect 8984 10076 9032 10132
rect 9088 10076 9136 10132
rect 9192 10076 9220 10132
rect 8900 10028 9220 10076
rect 8900 9972 8928 10028
rect 8984 9972 9032 10028
rect 9088 9972 9136 10028
rect 9192 9972 9220 10028
rect 8900 9924 9220 9972
rect 8900 9868 8928 9924
rect 8984 9868 9032 9924
rect 9088 9868 9136 9924
rect 9192 9868 9220 9924
rect 8900 8652 9220 9868
rect 8900 8596 8928 8652
rect 8984 8596 9032 8652
rect 9088 8596 9136 8652
rect 9192 8596 9220 8652
rect 4930 7620 5250 7668
rect 4930 7564 4958 7620
rect 5014 7564 5062 7620
rect 5118 7564 5166 7620
rect 5222 7564 5250 7620
rect 4930 6300 5250 7564
rect 7700 7308 7756 7318
rect 7028 6860 7084 6870
rect 4930 6244 4958 6300
rect 5014 6244 5062 6300
rect 5118 6244 5166 6300
rect 5222 6244 5250 6300
rect 4452 5180 4508 5190
rect 4452 3836 4508 5124
rect 4452 3770 4508 3780
rect 4930 4732 5250 6244
rect 4930 4676 4958 4732
rect 5014 4676 5062 4732
rect 5118 4676 5166 4732
rect 5222 4676 5250 4732
rect 4788 3612 4844 3622
rect 4788 3388 4844 3556
rect 4788 3322 4844 3332
rect 4340 2762 4396 2772
rect 4930 3220 5250 4676
rect 6916 6524 6972 6534
rect 6692 4168 6748 4178
rect 6692 3612 6748 4112
rect 6692 3546 6748 3556
rect 6804 3500 6860 3510
rect 6804 3382 6860 3392
rect 4930 3060 4958 3220
rect 5014 3060 5062 3220
rect 5118 3060 5166 3220
rect 5222 3060 5250 3220
rect 4930 3012 5250 3060
rect 4930 2956 4958 3012
rect 5014 2956 5062 3012
rect 5118 2956 5166 3012
rect 5222 2956 5250 3012
rect 1204 1194 1260 1204
rect 4930 1596 5250 2956
rect 6916 2492 6972 6468
rect 7028 4168 7084 6804
rect 7028 4102 7084 4112
rect 7700 3448 7756 7252
rect 8900 7084 9220 8596
rect 8900 7028 8928 7084
rect 8984 7028 9032 7084
rect 9088 7028 9136 7084
rect 9192 7028 9220 7084
rect 8900 5524 9220 7028
rect 8900 5460 8928 5524
rect 8984 5460 9032 5524
rect 9088 5460 9136 5524
rect 9192 5460 9220 5524
rect 8900 5420 9220 5460
rect 8900 5364 8928 5420
rect 8984 5364 9032 5420
rect 9088 5364 9136 5420
rect 9192 5364 9220 5420
rect 8900 5316 9220 5364
rect 8900 5260 8928 5316
rect 8984 5260 9032 5316
rect 9088 5260 9136 5316
rect 9192 5260 9220 5316
rect 8372 3988 8428 3998
rect 8372 3882 8428 3892
rect 8900 3948 9220 5260
rect 9940 7756 9996 7766
rect 9940 4508 9996 7700
rect 10948 7420 11004 11508
rect 11620 12124 11676 12134
rect 11620 11548 11676 12068
rect 11620 11482 11676 11492
rect 10948 7354 11004 7364
rect 12870 11004 13190 12172
rect 12870 10948 12898 11004
rect 12954 10948 13002 11004
rect 13058 10948 13106 11004
rect 13162 10948 13190 11004
rect 12870 9436 13190 10948
rect 13300 13580 13356 13590
rect 13300 10468 13356 13524
rect 13636 12572 13692 12582
rect 13300 10402 13356 10412
rect 13412 12460 13468 12470
rect 13412 9996 13468 12404
rect 13636 10556 13692 12516
rect 14084 11728 14140 14308
rect 14532 14364 14588 14980
rect 14532 14298 14588 14308
rect 14644 14068 14700 15316
rect 14532 12908 14588 12918
rect 14532 12460 14588 12852
rect 14532 12394 14588 12404
rect 14644 11788 14700 14012
rect 14756 13356 14812 16212
rect 15428 16268 15484 16278
rect 14756 13290 14812 13300
rect 15204 15372 15260 15382
rect 15204 11900 15260 15316
rect 15428 15260 15484 16212
rect 16548 16044 16604 16660
rect 16548 15978 16604 15988
rect 16840 16492 17160 18004
rect 16840 16436 16868 16492
rect 16924 16436 16972 16492
rect 17028 16436 17076 16492
rect 17132 16436 17160 16492
rect 15428 15148 15484 15204
rect 15428 15082 15484 15092
rect 16100 15484 16156 15494
rect 16100 15148 16156 15428
rect 16100 15082 16156 15092
rect 16840 14924 17160 16436
rect 17556 17308 17612 17318
rect 17556 15820 17612 17252
rect 20810 17276 21130 18788
rect 20810 17220 20838 17276
rect 20894 17220 20942 17276
rect 20998 17220 21046 17276
rect 21102 17220 21130 17276
rect 20810 17044 21130 17220
rect 20810 16988 20838 17044
rect 20894 16988 20942 17044
rect 20998 16988 21046 17044
rect 21102 16988 21130 17044
rect 17556 15754 17612 15764
rect 18116 16940 18172 16950
rect 16840 14868 16868 14924
rect 16924 14868 16972 14924
rect 17028 14868 17076 14924
rect 17132 14868 17160 14924
rect 16840 14740 17160 14868
rect 16840 14684 16868 14740
rect 16924 14684 16972 14740
rect 17028 14684 17076 14740
rect 17132 14684 17160 14740
rect 16840 14636 17160 14684
rect 16840 14580 16868 14636
rect 16924 14580 16972 14636
rect 17028 14580 17076 14636
rect 17132 14580 17160 14636
rect 16840 14532 17160 14580
rect 16840 14476 16868 14532
rect 16924 14476 16972 14532
rect 17028 14476 17076 14532
rect 17132 14476 17160 14532
rect 16840 13356 17160 14476
rect 16840 13300 16868 13356
rect 16924 13300 16972 13356
rect 17028 13300 17076 13356
rect 17132 13300 17160 13356
rect 15204 11834 15260 11844
rect 16660 12808 16716 12818
rect 16660 11900 16716 12752
rect 16660 11834 16716 11844
rect 14644 11722 14700 11732
rect 16840 11788 17160 13300
rect 16840 11732 16868 11788
rect 16924 11732 16972 11788
rect 17028 11732 17076 11788
rect 17132 11732 17160 11788
rect 17780 12460 17836 12470
rect 17780 12124 17836 12404
rect 14084 11662 14140 11672
rect 13636 10490 13692 10500
rect 13412 9930 13468 9940
rect 16840 10220 17160 11732
rect 17220 11728 17276 11738
rect 17220 11610 17276 11620
rect 16840 10164 16868 10220
rect 16924 10164 16972 10220
rect 17028 10164 17076 10220
rect 17132 10164 17160 10220
rect 16840 10132 17160 10164
rect 16840 10076 16868 10132
rect 16924 10076 16972 10132
rect 17028 10076 17076 10132
rect 17132 10076 17160 10132
rect 16840 10028 17160 10076
rect 16840 9972 16868 10028
rect 16924 9972 16972 10028
rect 17028 9972 17076 10028
rect 17132 9972 17160 10028
rect 12870 9380 12898 9436
rect 12954 9380 13002 9436
rect 13058 9380 13106 9436
rect 13162 9380 13190 9436
rect 12870 7868 13190 9380
rect 12870 7772 12898 7868
rect 12954 7772 13002 7868
rect 13058 7772 13106 7868
rect 13162 7772 13190 7868
rect 12870 7724 13190 7772
rect 12870 7668 12898 7724
rect 12954 7668 13002 7724
rect 13058 7668 13106 7724
rect 13162 7668 13190 7724
rect 12870 7620 13190 7668
rect 12870 7564 12898 7620
rect 12954 7564 13002 7620
rect 13058 7564 13106 7620
rect 13162 7564 13190 7620
rect 9940 4442 9996 4452
rect 12870 6300 13190 7564
rect 16840 9924 17160 9972
rect 16840 9868 16868 9924
rect 16924 9868 16972 9924
rect 17028 9868 17076 9924
rect 17132 9868 17160 9924
rect 16840 8652 17160 9868
rect 16840 8596 16868 8652
rect 16924 8596 16972 8652
rect 17028 8596 17076 8652
rect 17132 8596 17160 8652
rect 16840 7084 17160 8596
rect 17780 7532 17836 12068
rect 18004 11676 18060 11686
rect 18004 11548 18060 11620
rect 18004 11482 18060 11492
rect 18116 8876 18172 16884
rect 20810 16940 21130 16988
rect 20810 16884 20838 16940
rect 20894 16884 20942 16940
rect 20998 16884 21046 16940
rect 21102 16884 21130 16940
rect 20810 16836 21130 16884
rect 20810 16780 20838 16836
rect 20894 16780 20942 16836
rect 20998 16780 21046 16836
rect 21102 16780 21130 16836
rect 18340 16228 18396 16238
rect 18340 16156 18396 16172
rect 18340 16090 18396 16100
rect 20810 15708 21130 16780
rect 24780 18060 25100 18876
rect 24780 18004 24808 18060
rect 24864 18004 24912 18060
rect 24968 18004 25016 18060
rect 25072 18004 25100 18060
rect 23044 16588 23100 16598
rect 20810 15652 20838 15708
rect 20894 15652 20942 15708
rect 20998 15652 21046 15708
rect 21102 15652 21130 15708
rect 18564 15596 18620 15606
rect 18564 15328 18620 15540
rect 18564 15262 18620 15272
rect 18676 15260 18732 15270
rect 18564 14924 18620 14934
rect 18452 14700 18508 14710
rect 18452 14476 18508 14644
rect 18452 14410 18508 14420
rect 18564 14252 18620 14868
rect 18564 14186 18620 14196
rect 18676 12460 18732 15204
rect 18900 15148 18956 15158
rect 18788 12808 18844 12834
rect 18788 12730 18844 12740
rect 18676 12394 18732 12404
rect 18900 12460 18956 15092
rect 19796 15148 19852 15158
rect 19796 14700 19852 15092
rect 19796 14634 19852 14644
rect 19908 14924 19964 14934
rect 19908 12684 19964 14868
rect 20810 14140 21130 15652
rect 22260 16380 22316 16390
rect 21476 15596 21532 15606
rect 21252 15260 21308 15270
rect 21252 15036 21308 15204
rect 21252 14970 21308 14980
rect 21476 14700 21532 15540
rect 21476 14364 21532 14644
rect 21476 14298 21532 14308
rect 20810 14084 20838 14140
rect 20894 14084 20942 14140
rect 20998 14084 21046 14140
rect 21102 14084 21130 14140
rect 20468 14068 20524 14078
rect 20468 13692 20524 14012
rect 20468 13626 20524 13636
rect 19908 12618 19964 12628
rect 18900 12394 18956 12404
rect 20810 12572 21130 14084
rect 22260 13692 22316 16324
rect 22820 16268 22876 16278
rect 22820 15820 22876 16212
rect 22260 13626 22316 13636
rect 22484 15708 22540 15718
rect 22484 12908 22540 15652
rect 22820 15147 22876 15764
rect 23044 15484 23100 16532
rect 24780 16492 25100 18004
rect 24780 16436 24808 16492
rect 24864 16436 24912 16492
rect 24968 16436 25016 16492
rect 25072 16436 25100 16492
rect 23716 16156 23772 16166
rect 23716 16048 23772 16100
rect 23716 15982 23772 15992
rect 24612 15932 24668 15942
rect 23044 15418 23100 15428
rect 24500 15484 24556 15494
rect 22820 15091 22988 15147
rect 22932 13132 22988 15091
rect 22932 13066 22988 13076
rect 22484 12842 22540 12852
rect 24500 12908 24556 15428
rect 24612 15328 24668 15876
rect 24612 15262 24668 15272
rect 20810 12516 20838 12572
rect 20894 12516 20942 12572
rect 20998 12516 21046 12572
rect 21102 12516 21130 12572
rect 20810 12436 21130 12516
rect 20810 12380 20838 12436
rect 20894 12380 20942 12436
rect 20998 12380 21046 12436
rect 21102 12380 21130 12436
rect 20810 12332 21130 12380
rect 20810 12276 20838 12332
rect 20894 12276 20942 12332
rect 20998 12276 21046 12332
rect 21102 12276 21130 12332
rect 20810 12228 21130 12276
rect 20810 12172 20838 12228
rect 20894 12172 20942 12228
rect 20998 12172 21046 12228
rect 21102 12172 21130 12228
rect 20810 11004 21130 12172
rect 24500 12124 24556 12852
rect 24500 12058 24556 12068
rect 24780 14924 25100 16436
rect 28750 18844 29070 18876
rect 28750 18788 28778 18844
rect 28834 18788 28882 18844
rect 28938 18788 28986 18844
rect 29042 18788 29070 18844
rect 28750 17276 29070 18788
rect 28750 17220 28778 17276
rect 28834 17220 28882 17276
rect 28938 17220 28986 17276
rect 29042 17220 29070 17276
rect 28750 17044 29070 17220
rect 28750 16988 28778 17044
rect 28834 16988 28882 17044
rect 28938 16988 28986 17044
rect 29042 16988 29070 17044
rect 28750 16940 29070 16988
rect 28750 16884 28778 16940
rect 28834 16884 28882 16940
rect 28938 16884 28986 16940
rect 29042 16884 29070 16940
rect 28750 16836 29070 16884
rect 28750 16780 28778 16836
rect 28834 16780 28882 16836
rect 28938 16780 28986 16836
rect 29042 16780 29070 16836
rect 28750 15708 29070 16780
rect 28750 15652 28778 15708
rect 28834 15652 28882 15708
rect 28938 15652 28986 15708
rect 29042 15652 29070 15708
rect 27636 15508 27692 15518
rect 24780 14868 24808 14924
rect 24864 14868 24912 14924
rect 24968 14868 25016 14924
rect 25072 14868 25100 14924
rect 24780 14740 25100 14868
rect 24780 14684 24808 14740
rect 24864 14684 24912 14740
rect 24968 14684 25016 14740
rect 25072 14684 25100 14740
rect 24780 14636 25100 14684
rect 24780 14580 24808 14636
rect 24864 14580 24912 14636
rect 24968 14580 25016 14636
rect 25072 14580 25100 14636
rect 24780 14532 25100 14580
rect 24780 14476 24808 14532
rect 24864 14476 24912 14532
rect 24968 14476 25016 14532
rect 25072 14476 25100 14532
rect 24780 13356 25100 14476
rect 26852 14968 26908 14978
rect 26852 13916 26908 14912
rect 27636 14700 27692 15452
rect 27636 14634 27692 14644
rect 26852 13850 26908 13860
rect 28750 14140 29070 15652
rect 28750 14084 28778 14140
rect 28834 14084 28882 14140
rect 28938 14084 28986 14140
rect 29042 14084 29070 14140
rect 24780 13300 24808 13356
rect 24864 13300 24912 13356
rect 24968 13300 25016 13356
rect 25072 13300 25100 13356
rect 20810 10948 20838 11004
rect 20894 10948 20942 11004
rect 20998 10948 21046 11004
rect 21102 10948 21130 11004
rect 18228 10648 18284 10658
rect 18228 10556 18284 10592
rect 18228 10490 18284 10500
rect 18116 8810 18172 8820
rect 20810 9436 21130 10948
rect 24780 11788 25100 13300
rect 24780 11732 24808 11788
rect 24864 11732 24912 11788
rect 24968 11732 25016 11788
rect 25072 11732 25100 11788
rect 23492 10468 23548 10482
rect 23492 10378 23548 10388
rect 24780 10220 25100 11732
rect 24780 10164 24808 10220
rect 24864 10164 24912 10220
rect 24968 10164 25016 10220
rect 25072 10164 25100 10220
rect 24780 10132 25100 10164
rect 24780 10076 24808 10132
rect 24864 10076 24912 10132
rect 24968 10076 25016 10132
rect 25072 10076 25100 10132
rect 24780 10028 25100 10076
rect 24780 9972 24808 10028
rect 24864 9972 24912 10028
rect 24968 9972 25016 10028
rect 25072 9972 25100 10028
rect 24780 9924 25100 9972
rect 24780 9868 24808 9924
rect 24864 9868 24912 9924
rect 24968 9868 25016 9924
rect 25072 9868 25100 9924
rect 20810 9380 20838 9436
rect 20894 9380 20942 9436
rect 20998 9380 21046 9436
rect 21102 9380 21130 9436
rect 17780 7466 17836 7476
rect 20810 7868 21130 9380
rect 22260 9568 22316 9578
rect 22260 9212 22316 9512
rect 22260 9146 22316 9156
rect 20810 7772 20838 7868
rect 20894 7772 20942 7868
rect 20998 7772 21046 7868
rect 21102 7772 21130 7868
rect 20810 7724 21130 7772
rect 20810 7668 20838 7724
rect 20894 7668 20942 7724
rect 20998 7668 21046 7724
rect 21102 7668 21130 7724
rect 20810 7620 21130 7668
rect 20810 7564 20838 7620
rect 20894 7564 20942 7620
rect 20998 7564 21046 7620
rect 21102 7564 21130 7620
rect 16840 7028 16868 7084
rect 16924 7028 16972 7084
rect 17028 7028 17076 7084
rect 17132 7028 17160 7084
rect 12870 6244 12898 6300
rect 12954 6244 13002 6300
rect 13058 6244 13106 6300
rect 13162 6244 13190 6300
rect 12870 4732 13190 6244
rect 14420 6748 14476 6758
rect 12870 4676 12898 4732
rect 12954 4676 13002 4732
rect 13058 4676 13106 4732
rect 13162 4676 13190 4732
rect 8900 3892 8928 3948
rect 8984 3892 9032 3948
rect 9088 3892 9136 3948
rect 9192 3892 9220 3948
rect 7700 3382 7756 3392
rect 6916 2426 6972 2436
rect 4930 1540 4958 1596
rect 5014 1540 5062 1596
rect 5118 1540 5166 1596
rect 5222 1540 5250 1596
rect 4930 724 5250 1540
rect 8900 2380 9220 3892
rect 8900 2324 8928 2380
rect 8984 2324 9032 2380
rect 9088 2324 9136 2380
rect 9192 2324 9220 2380
rect 8900 812 9220 2324
rect 12740 3448 12796 3458
rect 12740 1260 12796 3392
rect 12740 1194 12796 1204
rect 12870 3220 13190 4676
rect 13300 5068 13356 5078
rect 13300 4284 13356 5012
rect 14420 4844 14476 6692
rect 16840 5524 17160 7028
rect 16840 5460 16868 5524
rect 16924 5460 16972 5524
rect 17028 5460 17076 5524
rect 17132 5460 17160 5524
rect 16840 5420 17160 5460
rect 16840 5364 16868 5420
rect 16924 5364 16972 5420
rect 17028 5364 17076 5420
rect 17132 5364 17160 5420
rect 16840 5316 17160 5364
rect 16840 5260 16868 5316
rect 16924 5260 16972 5316
rect 17028 5260 17076 5316
rect 17132 5260 17160 5316
rect 14420 4778 14476 4788
rect 15204 4888 15260 4898
rect 13300 4218 13356 4228
rect 12870 3060 12898 3220
rect 12954 3060 13002 3220
rect 13058 3060 13106 3220
rect 13162 3060 13190 3220
rect 12870 3012 13190 3060
rect 12870 2956 12898 3012
rect 12954 2956 13002 3012
rect 13058 2956 13106 3012
rect 13162 2956 13190 3012
rect 12870 1596 13190 2956
rect 12870 1540 12898 1596
rect 12954 1540 13002 1596
rect 13058 1540 13106 1596
rect 13162 1540 13190 1596
rect 8900 756 8928 812
rect 8984 756 9032 812
rect 9088 756 9136 812
rect 9192 756 9220 812
rect 8900 724 9220 756
rect 12870 724 13190 1540
rect 15204 1148 15260 4832
rect 15428 4168 15484 4178
rect 15428 1820 15484 4112
rect 15428 1754 15484 1764
rect 16840 3948 17160 5260
rect 16840 3892 16868 3948
rect 16924 3892 16972 3948
rect 17028 3892 17076 3948
rect 17132 3892 17160 3948
rect 16840 2380 17160 3892
rect 16840 2324 16868 2380
rect 16924 2324 16972 2380
rect 17028 2324 17076 2380
rect 17132 2324 17160 2380
rect 15204 1082 15260 1092
rect 16840 812 17160 2324
rect 19684 7420 19740 7430
rect 19684 1036 19740 7364
rect 20810 6300 21130 7564
rect 20810 6244 20838 6300
rect 20894 6244 20942 6300
rect 20998 6244 21046 6300
rect 21102 6244 21130 6300
rect 20810 4732 21130 6244
rect 24780 8652 25100 9868
rect 24780 8596 24808 8652
rect 24864 8596 24912 8652
rect 24968 8596 25016 8652
rect 25072 8596 25100 8652
rect 24780 7084 25100 8596
rect 24780 7028 24808 7084
rect 24864 7028 24912 7084
rect 24968 7028 25016 7084
rect 25072 7028 25100 7084
rect 24780 5524 25100 7028
rect 24780 5460 24808 5524
rect 24864 5460 24912 5524
rect 24968 5460 25016 5524
rect 25072 5460 25100 5524
rect 24780 5420 25100 5460
rect 24780 5364 24808 5420
rect 24864 5364 24912 5420
rect 24968 5364 25016 5420
rect 25072 5364 25100 5420
rect 24780 5316 25100 5364
rect 24780 5260 24808 5316
rect 24864 5260 24912 5316
rect 24968 5260 25016 5316
rect 25072 5260 25100 5316
rect 21364 5180 21420 5190
rect 21364 4888 21420 5124
rect 21364 4822 21420 4832
rect 20810 4676 20838 4732
rect 20894 4676 20942 4732
rect 20998 4676 21046 4732
rect 21102 4676 21130 4732
rect 20468 3500 20524 3510
rect 20468 3382 20524 3392
rect 19684 970 19740 980
rect 20810 3220 21130 4676
rect 20810 3060 20838 3220
rect 20894 3060 20942 3220
rect 20998 3060 21046 3220
rect 21102 3060 21130 3220
rect 20810 3012 21130 3060
rect 20810 2956 20838 3012
rect 20894 2956 20942 3012
rect 20998 2956 21046 3012
rect 21102 2956 21130 3012
rect 20810 1596 21130 2956
rect 20810 1540 20838 1596
rect 20894 1540 20942 1596
rect 20998 1540 21046 1596
rect 21102 1540 21130 1596
rect 16840 756 16868 812
rect 16924 756 16972 812
rect 17028 756 17076 812
rect 17132 756 17160 812
rect 16840 724 17160 756
rect 20810 724 21130 1540
rect 24780 3948 25100 5260
rect 24780 3892 24808 3948
rect 24864 3892 24912 3948
rect 24968 3892 25016 3948
rect 25072 3892 25100 3948
rect 24780 2380 25100 3892
rect 24780 2324 24808 2380
rect 24864 2324 24912 2380
rect 24968 2324 25016 2380
rect 25072 2324 25100 2380
rect 24780 812 25100 2324
rect 24780 756 24808 812
rect 24864 756 24912 812
rect 24968 756 25016 812
rect 25072 756 25100 812
rect 24780 724 25100 756
rect 28750 12572 29070 14084
rect 28750 12516 28778 12572
rect 28834 12516 28882 12572
rect 28938 12516 28986 12572
rect 29042 12516 29070 12572
rect 28750 12436 29070 12516
rect 28750 12380 28778 12436
rect 28834 12380 28882 12436
rect 28938 12380 28986 12436
rect 29042 12380 29070 12436
rect 28750 12332 29070 12380
rect 28750 12276 28778 12332
rect 28834 12276 28882 12332
rect 28938 12276 28986 12332
rect 29042 12276 29070 12332
rect 28750 12228 29070 12276
rect 28750 12172 28778 12228
rect 28834 12172 28882 12228
rect 28938 12172 28986 12228
rect 29042 12172 29070 12228
rect 28750 11004 29070 12172
rect 28750 10948 28778 11004
rect 28834 10948 28882 11004
rect 28938 10948 28986 11004
rect 29042 10948 29070 11004
rect 28750 9436 29070 10948
rect 28750 9380 28778 9436
rect 28834 9380 28882 9436
rect 28938 9380 28986 9436
rect 29042 9380 29070 9436
rect 28750 7868 29070 9380
rect 28750 7772 28778 7868
rect 28834 7772 28882 7868
rect 28938 7772 28986 7868
rect 29042 7772 29070 7868
rect 28750 7724 29070 7772
rect 28750 7668 28778 7724
rect 28834 7668 28882 7724
rect 28938 7668 28986 7724
rect 29042 7668 29070 7724
rect 28750 7620 29070 7668
rect 28750 7564 28778 7620
rect 28834 7564 28882 7620
rect 28938 7564 28986 7620
rect 29042 7564 29070 7620
rect 28750 6300 29070 7564
rect 28750 6244 28778 6300
rect 28834 6244 28882 6300
rect 28938 6244 28986 6300
rect 29042 6244 29070 6300
rect 28750 4732 29070 6244
rect 28750 4676 28778 4732
rect 28834 4676 28882 4732
rect 28938 4676 28986 4732
rect 29042 4676 29070 4732
rect 28750 3220 29070 4676
rect 28750 3060 28778 3220
rect 28834 3060 28882 3220
rect 28938 3060 28986 3220
rect 29042 3060 29070 3220
rect 28750 3012 29070 3060
rect 28750 2956 28778 3012
rect 28834 2956 28882 3012
rect 28938 2956 28986 3012
rect 29042 2956 29070 3012
rect 28750 1596 29070 2956
rect 28750 1540 28778 1596
rect 28834 1540 28882 1596
rect 28938 1540 28986 1596
rect 29042 1540 29070 1596
rect 28750 724 29070 1540
<< via4 >>
rect 4340 18332 4396 18388
rect 2548 16352 2604 16408
rect 3780 15092 3836 15148
rect 4788 16172 4844 16228
rect 4958 16988 5014 17044
rect 5062 16988 5118 17044
rect 5166 16988 5222 17044
rect 6356 17252 6412 17308
rect 4958 16884 5014 16940
rect 5062 16884 5118 16940
rect 5166 16884 5222 16940
rect 4958 16780 5014 16836
rect 5062 16780 5118 16836
rect 5166 16780 5222 16836
rect 12898 16988 12954 17044
rect 13002 16988 13058 17044
rect 13106 16988 13162 17044
rect 12898 16884 12954 16940
rect 13002 16884 13058 16940
rect 13106 16884 13162 16940
rect 12898 16780 12954 16836
rect 13002 16780 13058 16836
rect 13106 16780 13162 16836
rect 10052 16352 10108 16408
rect 11172 15992 11228 16048
rect 8928 14684 8984 14740
rect 9032 14684 9088 14740
rect 9136 14684 9192 14740
rect 8928 14580 8984 14636
rect 9032 14580 9088 14636
rect 9136 14580 9192 14636
rect 8928 14476 8984 14532
rect 9032 14476 9088 14532
rect 9136 14476 9192 14532
rect 4958 12380 5014 12436
rect 5062 12380 5118 12436
rect 5166 12380 5222 12436
rect 4958 12276 5014 12332
rect 5062 12276 5118 12332
rect 5166 12276 5222 12332
rect 4958 12172 5014 12228
rect 5062 12172 5118 12228
rect 5166 12172 5222 12228
rect 5348 9512 5404 9568
rect 1540 3932 1596 3988
rect 4958 7812 5014 7828
rect 4958 7772 5014 7812
rect 5062 7812 5118 7828
rect 5062 7772 5118 7812
rect 5166 7812 5222 7828
rect 5166 7772 5222 7812
rect 4958 7668 5014 7724
rect 5062 7668 5118 7724
rect 5166 7668 5222 7724
rect 8260 10592 8316 10648
rect 18452 18340 18508 18388
rect 18452 18332 18508 18340
rect 13300 16532 13356 16588
rect 12516 15484 12572 15508
rect 12516 15452 12572 15484
rect 12740 15092 12796 15148
rect 12180 14912 12236 14968
rect 12898 12380 12954 12436
rect 13002 12380 13058 12436
rect 13106 12380 13162 12436
rect 12898 12276 12954 12332
rect 13002 12276 13058 12332
rect 13106 12276 13162 12332
rect 12898 12172 12954 12228
rect 13002 12172 13058 12228
rect 13106 12172 13162 12228
rect 8928 10076 8984 10132
rect 9032 10076 9088 10132
rect 9136 10076 9192 10132
rect 8928 9972 8984 10028
rect 9032 9972 9088 10028
rect 9136 9972 9192 10028
rect 8928 9868 8984 9924
rect 9032 9868 9088 9924
rect 9136 9868 9192 9924
rect 4958 7564 5014 7620
rect 5062 7564 5118 7620
rect 5166 7564 5222 7620
rect 6692 4112 6748 4168
rect 6804 3444 6860 3448
rect 6804 3392 6860 3444
rect 4958 3164 5014 3220
rect 4958 3108 5014 3116
rect 4958 3060 5014 3108
rect 5062 3164 5118 3220
rect 5062 3108 5118 3116
rect 5062 3060 5118 3108
rect 5166 3164 5222 3220
rect 5166 3108 5222 3116
rect 5166 3060 5222 3108
rect 4958 2956 5014 3012
rect 5062 2956 5118 3012
rect 5166 2956 5222 3012
rect 7028 4112 7084 4168
rect 8928 5516 8984 5524
rect 8928 5468 8984 5516
rect 9032 5516 9088 5524
rect 9032 5468 9088 5516
rect 9136 5516 9192 5524
rect 9136 5468 9192 5516
rect 8928 5364 8984 5420
rect 9032 5364 9088 5420
rect 9136 5364 9192 5420
rect 8928 5260 8984 5316
rect 9032 5260 9088 5316
rect 9136 5260 9192 5316
rect 8372 3948 8428 3988
rect 8372 3932 8428 3948
rect 11620 11492 11676 11548
rect 13300 10412 13356 10468
rect 14644 14012 14700 14068
rect 14084 11672 14140 11728
rect 15428 15092 15484 15148
rect 17556 17252 17612 17308
rect 20838 16988 20894 17044
rect 20942 16988 20998 17044
rect 21046 16988 21102 17044
rect 16868 14684 16924 14740
rect 16972 14684 17028 14740
rect 17076 14684 17132 14740
rect 16868 14580 16924 14636
rect 16972 14580 17028 14636
rect 17076 14580 17132 14636
rect 16868 14476 16924 14532
rect 16972 14476 17028 14532
rect 17076 14476 17132 14532
rect 16660 12752 16716 12808
rect 17220 11676 17276 11728
rect 17220 11672 17276 11676
rect 16868 10076 16924 10132
rect 16972 10076 17028 10132
rect 17076 10076 17132 10132
rect 16868 9972 16924 10028
rect 16972 9972 17028 10028
rect 17076 9972 17132 10028
rect 12898 7812 12954 7828
rect 12898 7772 12954 7812
rect 13002 7812 13058 7828
rect 13002 7772 13058 7812
rect 13106 7812 13162 7828
rect 13106 7772 13162 7812
rect 12898 7668 12954 7724
rect 13002 7668 13058 7724
rect 13106 7668 13162 7724
rect 12898 7564 12954 7620
rect 13002 7564 13058 7620
rect 13106 7564 13162 7620
rect 16868 9868 16924 9924
rect 16972 9868 17028 9924
rect 17076 9868 17132 9924
rect 18004 11492 18060 11548
rect 20838 16884 20894 16940
rect 20942 16884 20998 16940
rect 21046 16884 21102 16940
rect 20838 16780 20894 16836
rect 20942 16780 20998 16836
rect 21046 16780 21102 16836
rect 18340 16172 18396 16228
rect 23044 16532 23100 16588
rect 18564 15272 18620 15328
rect 18900 15092 18956 15148
rect 18788 12796 18844 12808
rect 18788 12752 18844 12796
rect 20468 14012 20524 14068
rect 23716 15992 23772 16048
rect 24612 15272 24668 15328
rect 20838 12380 20894 12436
rect 20942 12380 20998 12436
rect 21046 12380 21102 12436
rect 20838 12276 20894 12332
rect 20942 12276 20998 12332
rect 21046 12276 21102 12332
rect 20838 12172 20894 12228
rect 20942 12172 20998 12228
rect 21046 12172 21102 12228
rect 28778 16988 28834 17044
rect 28882 16988 28938 17044
rect 28986 16988 29042 17044
rect 28778 16884 28834 16940
rect 28882 16884 28938 16940
rect 28986 16884 29042 16940
rect 28778 16780 28834 16836
rect 28882 16780 28938 16836
rect 28986 16780 29042 16836
rect 27636 15452 27692 15508
rect 24808 14684 24864 14740
rect 24912 14684 24968 14740
rect 25016 14684 25072 14740
rect 24808 14580 24864 14636
rect 24912 14580 24968 14636
rect 25016 14580 25072 14636
rect 24808 14476 24864 14532
rect 24912 14476 24968 14532
rect 25016 14476 25072 14532
rect 26852 14912 26908 14968
rect 18228 10592 18284 10648
rect 23492 10444 23548 10468
rect 23492 10412 23548 10444
rect 24808 10076 24864 10132
rect 24912 10076 24968 10132
rect 25016 10076 25072 10132
rect 24808 9972 24864 10028
rect 24912 9972 24968 10028
rect 25016 9972 25072 10028
rect 24808 9868 24864 9924
rect 24912 9868 24968 9924
rect 25016 9868 25072 9924
rect 22260 9512 22316 9568
rect 20838 7812 20894 7828
rect 20838 7772 20894 7812
rect 20942 7812 20998 7828
rect 20942 7772 20998 7812
rect 21046 7812 21102 7828
rect 21046 7772 21102 7812
rect 20838 7668 20894 7724
rect 20942 7668 20998 7724
rect 21046 7668 21102 7724
rect 20838 7564 20894 7620
rect 20942 7564 20998 7620
rect 21046 7564 21102 7620
rect 7700 3392 7756 3448
rect 12740 3392 12796 3448
rect 16868 5516 16924 5524
rect 16868 5468 16924 5516
rect 16972 5516 17028 5524
rect 16972 5468 17028 5516
rect 17076 5516 17132 5524
rect 17076 5468 17132 5516
rect 16868 5364 16924 5420
rect 16972 5364 17028 5420
rect 17076 5364 17132 5420
rect 16868 5260 16924 5316
rect 16972 5260 17028 5316
rect 17076 5260 17132 5316
rect 15204 4832 15260 4888
rect 12898 3164 12954 3220
rect 12898 3108 12954 3116
rect 12898 3060 12954 3108
rect 13002 3164 13058 3220
rect 13002 3108 13058 3116
rect 13002 3060 13058 3108
rect 13106 3164 13162 3220
rect 13106 3108 13162 3116
rect 13106 3060 13162 3108
rect 12898 2956 12954 3012
rect 13002 2956 13058 3012
rect 13106 2956 13162 3012
rect 15428 4112 15484 4168
rect 24808 5516 24864 5524
rect 24808 5468 24864 5516
rect 24912 5516 24968 5524
rect 24912 5468 24968 5516
rect 25016 5516 25072 5524
rect 25016 5468 25072 5516
rect 24808 5364 24864 5420
rect 24912 5364 24968 5420
rect 25016 5364 25072 5420
rect 24808 5260 24864 5316
rect 24912 5260 24968 5316
rect 25016 5260 25072 5316
rect 21364 4832 21420 4888
rect 20468 3444 20524 3448
rect 20468 3392 20524 3444
rect 20838 3164 20894 3220
rect 20838 3108 20894 3116
rect 20838 3060 20894 3108
rect 20942 3164 20998 3220
rect 20942 3108 20998 3116
rect 20942 3060 20998 3108
rect 21046 3164 21102 3220
rect 21046 3108 21102 3116
rect 21046 3060 21102 3108
rect 20838 2956 20894 3012
rect 20942 2956 20998 3012
rect 21046 2956 21102 3012
rect 28778 12380 28834 12436
rect 28882 12380 28938 12436
rect 28986 12380 29042 12436
rect 28778 12276 28834 12332
rect 28882 12276 28938 12332
rect 28986 12276 29042 12332
rect 28778 12172 28834 12228
rect 28882 12172 28938 12228
rect 28986 12172 29042 12228
rect 28778 7812 28834 7828
rect 28778 7772 28834 7812
rect 28882 7812 28938 7828
rect 28882 7772 28938 7812
rect 28986 7812 29042 7828
rect 28986 7772 29042 7812
rect 28778 7668 28834 7724
rect 28882 7668 28938 7724
rect 28986 7668 29042 7724
rect 28778 7564 28834 7620
rect 28882 7564 28938 7620
rect 28986 7564 29042 7620
rect 28778 3164 28834 3220
rect 28778 3108 28834 3116
rect 28778 3060 28834 3108
rect 28882 3164 28938 3220
rect 28882 3108 28938 3116
rect 28882 3060 28938 3108
rect 28986 3164 29042 3220
rect 28986 3108 29042 3116
rect 28986 3060 29042 3108
rect 28778 2956 28834 3012
rect 28882 2956 28938 3012
rect 28986 2956 29042 3012
<< metal5 >>
rect 4324 18388 18524 18404
rect 4324 18332 4340 18388
rect 4396 18332 18452 18388
rect 18508 18332 18524 18388
rect 4324 18316 18524 18332
rect 6340 17308 17628 17324
rect 6340 17252 6356 17308
rect 6412 17252 17556 17308
rect 17612 17252 17628 17308
rect 6340 17236 17628 17252
rect 1060 17044 32876 17072
rect 1060 16988 4958 17044
rect 5014 16988 5062 17044
rect 5118 16988 5166 17044
rect 5222 16988 12898 17044
rect 12954 16988 13002 17044
rect 13058 16988 13106 17044
rect 13162 16988 20838 17044
rect 20894 16988 20942 17044
rect 20998 16988 21046 17044
rect 21102 16988 28778 17044
rect 28834 16988 28882 17044
rect 28938 16988 28986 17044
rect 29042 16988 32876 17044
rect 1060 16940 32876 16988
rect 1060 16884 4958 16940
rect 5014 16884 5062 16940
rect 5118 16884 5166 16940
rect 5222 16884 12898 16940
rect 12954 16884 13002 16940
rect 13058 16884 13106 16940
rect 13162 16884 20838 16940
rect 20894 16884 20942 16940
rect 20998 16884 21046 16940
rect 21102 16884 28778 16940
rect 28834 16884 28882 16940
rect 28938 16884 28986 16940
rect 29042 16884 32876 16940
rect 1060 16836 32876 16884
rect 1060 16780 4958 16836
rect 5014 16780 5062 16836
rect 5118 16780 5166 16836
rect 5222 16780 12898 16836
rect 12954 16780 13002 16836
rect 13058 16780 13106 16836
rect 13162 16780 20838 16836
rect 20894 16780 20942 16836
rect 20998 16780 21046 16836
rect 21102 16780 28778 16836
rect 28834 16780 28882 16836
rect 28938 16780 28986 16836
rect 29042 16780 32876 16836
rect 1060 16752 32876 16780
rect 13284 16588 23116 16604
rect 13284 16532 13300 16588
rect 13356 16532 23044 16588
rect 23100 16532 23116 16588
rect 13284 16516 23116 16532
rect 2532 16408 10124 16424
rect 2532 16352 2548 16408
rect 2604 16352 10052 16408
rect 10108 16352 10124 16408
rect 2532 16336 10124 16352
rect 4772 16228 18412 16244
rect 4772 16172 4788 16228
rect 4844 16172 18340 16228
rect 18396 16172 18412 16228
rect 4772 16156 18412 16172
rect 11156 16048 23788 16064
rect 11156 15992 11172 16048
rect 11228 15992 23716 16048
rect 23772 15992 23788 16048
rect 11156 15976 23788 15992
rect 12500 15508 27708 15524
rect 12500 15452 12516 15508
rect 12572 15452 27636 15508
rect 27692 15452 27708 15508
rect 12500 15436 27708 15452
rect 15075 15328 24684 15344
rect 15075 15272 18564 15328
rect 18620 15272 24612 15328
rect 24668 15272 24684 15328
rect 15075 15256 24684 15272
rect 15075 15164 15163 15256
rect 3764 15148 15163 15164
rect 3764 15092 3780 15148
rect 3836 15092 12740 15148
rect 12796 15092 15163 15148
rect 3764 15076 15163 15092
rect 15412 15148 18972 15164
rect 15412 15092 15428 15148
rect 15484 15092 18900 15148
rect 18956 15092 18972 15148
rect 15412 15076 18972 15092
rect 12164 14968 26924 14984
rect 12164 14912 12180 14968
rect 12236 14912 26852 14968
rect 26908 14912 26924 14968
rect 12164 14896 26924 14912
rect 1060 14740 32876 14768
rect 1060 14684 8928 14740
rect 8984 14684 9032 14740
rect 9088 14684 9136 14740
rect 9192 14684 16868 14740
rect 16924 14684 16972 14740
rect 17028 14684 17076 14740
rect 17132 14684 24808 14740
rect 24864 14684 24912 14740
rect 24968 14684 25016 14740
rect 25072 14684 32876 14740
rect 1060 14636 32876 14684
rect 1060 14580 8928 14636
rect 8984 14580 9032 14636
rect 9088 14580 9136 14636
rect 9192 14580 16868 14636
rect 16924 14580 16972 14636
rect 17028 14580 17076 14636
rect 17132 14580 24808 14636
rect 24864 14580 24912 14636
rect 24968 14580 25016 14636
rect 25072 14580 32876 14636
rect 1060 14532 32876 14580
rect 1060 14476 8928 14532
rect 8984 14476 9032 14532
rect 9088 14476 9136 14532
rect 9192 14476 16868 14532
rect 16924 14476 16972 14532
rect 17028 14476 17076 14532
rect 17132 14476 24808 14532
rect 24864 14476 24912 14532
rect 24968 14476 25016 14532
rect 25072 14476 32876 14532
rect 1060 14448 32876 14476
rect 14628 14068 20540 14084
rect 14628 14012 14644 14068
rect 14700 14012 20468 14068
rect 20524 14012 20540 14068
rect 14628 13996 20540 14012
rect 16644 12808 18860 12824
rect 16644 12752 16660 12808
rect 16716 12752 18788 12808
rect 18844 12752 18860 12808
rect 16644 12736 18860 12752
rect 1060 12436 32876 12464
rect 1060 12380 4958 12436
rect 5014 12380 5062 12436
rect 5118 12380 5166 12436
rect 5222 12380 12898 12436
rect 12954 12380 13002 12436
rect 13058 12380 13106 12436
rect 13162 12380 20838 12436
rect 20894 12380 20942 12436
rect 20998 12380 21046 12436
rect 21102 12380 28778 12436
rect 28834 12380 28882 12436
rect 28938 12380 28986 12436
rect 29042 12380 32876 12436
rect 1060 12332 32876 12380
rect 1060 12276 4958 12332
rect 5014 12276 5062 12332
rect 5118 12276 5166 12332
rect 5222 12276 12898 12332
rect 12954 12276 13002 12332
rect 13058 12276 13106 12332
rect 13162 12276 20838 12332
rect 20894 12276 20942 12332
rect 20998 12276 21046 12332
rect 21102 12276 28778 12332
rect 28834 12276 28882 12332
rect 28938 12276 28986 12332
rect 29042 12276 32876 12332
rect 1060 12228 32876 12276
rect 1060 12172 4958 12228
rect 5014 12172 5062 12228
rect 5118 12172 5166 12228
rect 5222 12172 12898 12228
rect 12954 12172 13002 12228
rect 13058 12172 13106 12228
rect 13162 12172 20838 12228
rect 20894 12172 20942 12228
rect 20998 12172 21046 12228
rect 21102 12172 28778 12228
rect 28834 12172 28882 12228
rect 28938 12172 28986 12228
rect 29042 12172 32876 12228
rect 1060 12144 32876 12172
rect 14068 11728 17292 11744
rect 14068 11672 14084 11728
rect 14140 11672 17220 11728
rect 17276 11672 17292 11728
rect 14068 11656 17292 11672
rect 11604 11548 18076 11564
rect 11604 11492 11620 11548
rect 11676 11492 18004 11548
rect 18060 11492 18076 11548
rect 11604 11476 18076 11492
rect 8244 10648 18300 10664
rect 8244 10592 8260 10648
rect 8316 10592 18228 10648
rect 18284 10592 18300 10648
rect 8244 10576 18300 10592
rect 13284 10468 23564 10484
rect 13284 10412 13300 10468
rect 13356 10412 23492 10468
rect 23548 10412 23564 10468
rect 13284 10396 23564 10412
rect 1060 10132 32876 10160
rect 1060 10076 8928 10132
rect 8984 10076 9032 10132
rect 9088 10076 9136 10132
rect 9192 10076 16868 10132
rect 16924 10076 16972 10132
rect 17028 10076 17076 10132
rect 17132 10076 24808 10132
rect 24864 10076 24912 10132
rect 24968 10076 25016 10132
rect 25072 10076 32876 10132
rect 1060 10028 32876 10076
rect 1060 9972 8928 10028
rect 8984 9972 9032 10028
rect 9088 9972 9136 10028
rect 9192 9972 16868 10028
rect 16924 9972 16972 10028
rect 17028 9972 17076 10028
rect 17132 9972 24808 10028
rect 24864 9972 24912 10028
rect 24968 9972 25016 10028
rect 25072 9972 32876 10028
rect 1060 9924 32876 9972
rect 1060 9868 8928 9924
rect 8984 9868 9032 9924
rect 9088 9868 9136 9924
rect 9192 9868 16868 9924
rect 16924 9868 16972 9924
rect 17028 9868 17076 9924
rect 17132 9868 24808 9924
rect 24864 9868 24912 9924
rect 24968 9868 25016 9924
rect 25072 9868 32876 9924
rect 1060 9840 32876 9868
rect 5332 9568 22332 9584
rect 5332 9512 5348 9568
rect 5404 9512 22260 9568
rect 22316 9512 22332 9568
rect 5332 9496 22332 9512
rect 1060 7828 32876 7856
rect 1060 7772 4958 7828
rect 5014 7772 5062 7828
rect 5118 7772 5166 7828
rect 5222 7772 12898 7828
rect 12954 7772 13002 7828
rect 13058 7772 13106 7828
rect 13162 7772 20838 7828
rect 20894 7772 20942 7828
rect 20998 7772 21046 7828
rect 21102 7772 28778 7828
rect 28834 7772 28882 7828
rect 28938 7772 28986 7828
rect 29042 7772 32876 7828
rect 1060 7724 32876 7772
rect 1060 7668 4958 7724
rect 5014 7668 5062 7724
rect 5118 7668 5166 7724
rect 5222 7668 12898 7724
rect 12954 7668 13002 7724
rect 13058 7668 13106 7724
rect 13162 7668 20838 7724
rect 20894 7668 20942 7724
rect 20998 7668 21046 7724
rect 21102 7668 28778 7724
rect 28834 7668 28882 7724
rect 28938 7668 28986 7724
rect 29042 7668 32876 7724
rect 1060 7620 32876 7668
rect 1060 7564 4958 7620
rect 5014 7564 5062 7620
rect 5118 7564 5166 7620
rect 5222 7564 12898 7620
rect 12954 7564 13002 7620
rect 13058 7564 13106 7620
rect 13162 7564 20838 7620
rect 20894 7564 20942 7620
rect 20998 7564 21046 7620
rect 21102 7564 28778 7620
rect 28834 7564 28882 7620
rect 28938 7564 28986 7620
rect 29042 7564 32876 7620
rect 1060 7536 32876 7564
rect 1060 5524 32876 5552
rect 1060 5468 8928 5524
rect 8984 5468 9032 5524
rect 9088 5468 9136 5524
rect 9192 5468 16868 5524
rect 16924 5468 16972 5524
rect 17028 5468 17076 5524
rect 17132 5468 24808 5524
rect 24864 5468 24912 5524
rect 24968 5468 25016 5524
rect 25072 5468 32876 5524
rect 1060 5420 32876 5468
rect 1060 5364 8928 5420
rect 8984 5364 9032 5420
rect 9088 5364 9136 5420
rect 9192 5364 16868 5420
rect 16924 5364 16972 5420
rect 17028 5364 17076 5420
rect 17132 5364 24808 5420
rect 24864 5364 24912 5420
rect 24968 5364 25016 5420
rect 25072 5364 32876 5420
rect 1060 5316 32876 5364
rect 1060 5260 8928 5316
rect 8984 5260 9032 5316
rect 9088 5260 9136 5316
rect 9192 5260 16868 5316
rect 16924 5260 16972 5316
rect 17028 5260 17076 5316
rect 17132 5260 24808 5316
rect 24864 5260 24912 5316
rect 24968 5260 25016 5316
rect 25072 5260 32876 5316
rect 1060 5232 32876 5260
rect 15188 4888 21436 4904
rect 15188 4832 15204 4888
rect 15260 4832 21364 4888
rect 21420 4832 21436 4888
rect 15188 4816 21436 4832
rect 6676 4168 15500 4184
rect 6676 4112 6692 4168
rect 6748 4112 7028 4168
rect 7084 4112 15428 4168
rect 15484 4112 15500 4168
rect 6676 4096 15500 4112
rect 1524 3988 8444 4004
rect 1524 3932 1540 3988
rect 1596 3932 8372 3988
rect 8428 3932 8444 3988
rect 1524 3916 8444 3932
rect 6788 3448 20540 3464
rect 6788 3392 6804 3448
rect 6860 3392 7700 3448
rect 7756 3392 12740 3448
rect 12796 3392 20468 3448
rect 20524 3392 20540 3448
rect 6788 3376 20540 3392
rect 1060 3220 32876 3248
rect 1060 3164 4958 3220
rect 5014 3164 5062 3220
rect 5118 3164 5166 3220
rect 5222 3164 12898 3220
rect 12954 3164 13002 3220
rect 13058 3164 13106 3220
rect 13162 3164 20838 3220
rect 20894 3164 20942 3220
rect 20998 3164 21046 3220
rect 21102 3164 28778 3220
rect 28834 3164 28882 3220
rect 28938 3164 28986 3220
rect 29042 3164 32876 3220
rect 1060 3116 32876 3164
rect 1060 3060 4958 3116
rect 5014 3060 5062 3116
rect 5118 3060 5166 3116
rect 5222 3060 12898 3116
rect 12954 3060 13002 3116
rect 13058 3060 13106 3116
rect 13162 3060 20838 3116
rect 20894 3060 20942 3116
rect 20998 3060 21046 3116
rect 21102 3060 28778 3116
rect 28834 3060 28882 3116
rect 28938 3060 28986 3116
rect 29042 3060 32876 3116
rect 1060 3012 32876 3060
rect 1060 2956 4958 3012
rect 5014 2956 5062 3012
rect 5118 2956 5166 3012
rect 5222 2956 12898 3012
rect 12954 2956 13002 3012
rect 13058 2956 13106 3012
rect 13162 2956 20838 3012
rect 20894 2956 20942 3012
rect 20998 2956 21046 3012
rect 21102 2956 28778 3012
rect 28834 2956 28882 3012
rect 28938 2956 28986 3012
rect 29042 2956 32876 3012
rect 1060 2928 32876 2956
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__335__I pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 13328 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__I0
timestamp 1654395037
transform 1 0 16576 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__342__A1
timestamp 1654395037
transform -1 0 7728 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__342__A2
timestamp 1654395037
transform -1 0 7504 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__344__A1
timestamp 1654395037
transform 1 0 6272 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__344__A2
timestamp 1654395037
transform 1 0 6048 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__A1
timestamp 1654395037
transform 1 0 3808 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__A2
timestamp 1654395037
transform 1 0 4816 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__390__A1
timestamp 1654395037
transform -1 0 9744 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__404__A1
timestamp 1654395037
transform 1 0 12768 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__A1
timestamp 1654395037
transform -1 0 9744 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__A1
timestamp 1654395037
transform 1 0 9296 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__440__I
timestamp 1654395037
transform 1 0 25760 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__486__I
timestamp 1654395037
transform 1 0 12768 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__496__A1
timestamp 1654395037
transform -1 0 2240 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__499__A1
timestamp 1654395037
transform -1 0 6720 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__502__A1
timestamp 1654395037
transform 1 0 3696 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__513__A1
timestamp 1654395037
transform -1 0 10864 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__514__A1
timestamp 1654395037
transform 1 0 8848 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__519__A1
timestamp 1654395037
transform 1 0 19264 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__520__A1
timestamp 1654395037
transform -1 0 15344 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__524__I
timestamp 1654395037
transform -1 0 16912 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__529__I
timestamp 1654395037
transform 1 0 11424 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__547__A1
timestamp 1654395037
transform 1 0 21168 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__562__B2
timestamp 1654395037
transform 1 0 17360 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__564__A1
timestamp 1654395037
transform 1 0 20496 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__568__A1
timestamp 1654395037
transform 1 0 24752 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__577__A1
timestamp 1654395037
transform 1 0 23744 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__584__B2
timestamp 1654395037
transform -1 0 21616 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__590__A1
timestamp 1654395037
transform 1 0 24528 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__594__B2
timestamp 1654395037
transform -1 0 24976 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__595__A1
timestamp 1654395037
transform 1 0 26320 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__599__A1
timestamp 1654395037
transform 1 0 27440 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__600__A2
timestamp 1654395037
transform 1 0 26096 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__602__A1
timestamp 1654395037
transform 1 0 24752 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__604__A1
timestamp 1654395037
transform 1 0 22960 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__605__A2
timestamp 1654395037
transform 1 0 23520 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__634__I
timestamp 1654395037
transform 1 0 18816 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__646__I
timestamp 1654395037
transform 1 0 19712 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__663__CLK
timestamp 1654395037
transform 1 0 26096 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__664__CLK
timestamp 1654395037
transform 1 0 26432 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__665__CLK
timestamp 1654395037
transform 1 0 25984 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__666__CLK
timestamp 1654395037
transform 1 0 19936 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__667__CLK
timestamp 1654395037
transform 1 0 19600 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__668__CLK
timestamp 1654395037
transform 1 0 21168 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__669__CLK
timestamp 1654395037
transform 1 0 20384 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__670__CLK
timestamp 1654395037
transform 1 0 16800 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__671__CLK
timestamp 1654395037
transform 1 0 17248 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__672__CLK
timestamp 1654395037
transform 1 0 13888 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__673__CLK
timestamp 1654395037
transform 1 0 9072 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__674__CLK
timestamp 1654395037
transform 1 0 25200 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__675__CLK
timestamp 1654395037
transform 1 0 20944 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__676__CLK
timestamp 1654395037
transform 1 0 21840 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__677__CLK
timestamp 1654395037
transform 1 0 25424 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__678__CLK
timestamp 1654395037
transform 1 0 24304 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__679__CLK
timestamp 1654395037
transform 1 0 25648 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__680__CLK
timestamp 1654395037
transform 1 0 25872 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__681__CLK
timestamp 1654395037
transform 1 0 17248 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__682__CLK
timestamp 1654395037
transform 1 0 13440 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__683__CLK
timestamp 1654395037
transform 1 0 13216 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__684__CLK
timestamp 1654395037
transform 1 0 14672 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__685__CLK
timestamp 1654395037
transform 1 0 10304 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__686__I
timestamp 1654395037
transform 1 0 4928 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1654395037
transform 1 0 3696 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1654395037
transform 1 0 6608 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1654395037
transform -1 0 5040 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1654395037
transform 1 0 8064 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1654395037
transform 1 0 3696 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1654395037
transform -1 0 1568 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1654395037
transform -1 0 1568 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1654395037
transform 1 0 1344 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1654395037
transform -1 0 6384 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1654395037
transform 1 0 12656 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1654395037
transform -1 0 12992 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1654395037
transform 1 0 17248 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1654395037
transform 1 0 23744 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1654395037
transform 1 0 23968 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1654395037
transform -1 0 24640 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1654395037
transform 1 0 28112 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1654395037
transform 1 0 30688 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1654395037
transform -1 0 32592 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1654395037
transform 1 0 1568 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1654395037
transform -1 0 32144 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1654395037
transform -1 0 31920 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1654395037
transform -1 0 31920 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1654395037
transform -1 0 31920 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1654395037
transform -1 0 31920 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1654395037
transform -1 0 31920 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1654395037
transform 1 0 2016 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1654395037
transform 1 0 2016 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1654395037
transform 1 0 2688 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1654395037
transform 1 0 3136 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1654395037
transform 1 0 2912 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1654395037
transform 1 0 3360 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1654395037
transform 1 0 4480 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1654395037
transform -1 0 6160 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1654395037
transform 1 0 26208 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1654395037
transform 1 0 9744 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_ringosc.dstage\[0\].id.delaybuf1_I
timestamp 1654395037
transform 1 0 4704 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_ringosc.dstage\[0\].id.delayen1_EN
timestamp 1654395037
transform 1 0 4032 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_ringosc.dstage\[0\].id.delayenb0_I
timestamp 1654395037
transform 1 0 4816 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_ringosc.dstage\[0\].id.delayenb1_I
timestamp 1654395037
transform 1 0 5040 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_ringosc.dstage\[0\].id.trim1bar_I
timestamp 1654395037
transform -1 0 1680 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 4928 0 1 784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1654395037
transform 1 0 5264 0 1 784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 9184 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_103 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 12656 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_107
timestamp 1654395037
transform 1 0 13104 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1654395037
transform 1 0 20608 0 1 784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_201 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 23632 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1654395037
transform 1 0 24528 0 1 784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_212
timestamp 1654395037
transform 1 0 24864 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_216
timestamp 1654395037
transform 1 0 25312 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_226 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 26432 0 1 784
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_242
timestamp 1654395037
transform 1 0 28224 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1654395037
transform 1 0 28448 0 1 784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_247 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 28784 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_279
timestamp 1654395037
transform 1 0 32368 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_2
timestamp 1654395037
transform 1 0 1344 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_4
timestamp 1654395037
transform 1 0 1568 0 -1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_69
timestamp 1654395037
transform 1 0 8848 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_73
timestamp 1654395037
transform 1 0 9296 0 -1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_146
timestamp 1654395037
transform 1 0 17472 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_148
timestamp 1654395037
transform 1 0 17696 0 -1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_209
timestamp 1654395037
transform 1 0 24528 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_215
timestamp 1654395037
transform 1 0 25200 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_247
timestamp 1654395037
transform 1 0 28784 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_263
timestamp 1654395037
transform 1 0 30576 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_271
timestamp 1654395037
transform 1 0 31472 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_49
timestamp 1654395037
transform 1 0 6608 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1654395037
transform 1 0 12880 0 1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_167
timestamp 1654395037
transform 1 0 19824 0 1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1654395037
transform 1 0 20832 0 1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_223
timestamp 1654395037
transform 1 0 26096 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_239
timestamp 1654395037
transform 1 0 27888 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1654395037
transform 1 0 28784 0 1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_250
timestamp 1654395037
transform 1 0 29120 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_266
timestamp 1654395037
transform 1 0 30912 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_274
timestamp 1654395037
transform 1 0 31808 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_278
timestamp 1654395037
transform 1 0 32256 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_280
timestamp 1654395037
transform 1 0 32480 0 1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1654395037
transform 1 0 8960 0 -1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_105
timestamp 1654395037
transform 1 0 12880 0 -1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_122
timestamp 1654395037
transform 1 0 14784 0 -1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_139
timestamp 1654395037
transform 1 0 16688 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1654395037
transform 1 0 16912 0 -1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1654395037
transform 1 0 24864 0 -1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_227
timestamp 1654395037
transform 1 0 26544 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_259
timestamp 1654395037
transform 1 0 30128 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_275
timestamp 1654395037
transform 1 0 31920 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_279
timestamp 1654395037
transform 1 0 32368 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_69
timestamp 1654395037
transform 1 0 8848 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_71
timestamp 1654395037
transform 1 0 9072 0 1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_181
timestamp 1654395037
transform 1 0 21392 0 1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_224
timestamp 1654395037
transform 1 0 26208 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_240
timestamp 1654395037
transform 1 0 28000 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_250
timestamp 1654395037
transform 1 0 29120 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_266
timestamp 1654395037
transform 1 0 30912 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_274
timestamp 1654395037
transform 1 0 31808 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_278
timestamp 1654395037
transform 1 0 32256 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_280
timestamp 1654395037
transform 1 0 32480 0 1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_14
timestamp 1654395037
transform 1 0 2688 0 -1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_23
timestamp 1654395037
transform 1 0 3696 0 -1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1654395037
transform 1 0 8960 0 -1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_73
timestamp 1654395037
transform 1 0 9296 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_140
timestamp 1654395037
transform 1 0 16800 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_150
timestamp 1654395037
transform 1 0 17920 0 -1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_227
timestamp 1654395037
transform 1 0 26544 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_259
timestamp 1654395037
transform 1 0 30128 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_267
timestamp 1654395037
transform 1 0 31024 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_271
timestamp 1654395037
transform 1 0 31472 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_49
timestamp 1654395037
transform 1 0 6608 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_51
timestamp 1654395037
transform 1 0 6832 0 1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_99
timestamp 1654395037
transform 1 0 12208 0 1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_108
timestamp 1654395037
transform 1 0 13216 0 1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_163
timestamp 1654395037
transform 1 0 19376 0 1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_174
timestamp 1654395037
transform 1 0 20608 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1654395037
transform 1 0 20832 0 1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_185
timestamp 1654395037
transform 1 0 21840 0 1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_228
timestamp 1654395037
transform 1 0 26656 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_244
timestamp 1654395037
transform 1 0 28448 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_250
timestamp 1654395037
transform 1 0 29120 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_266
timestamp 1654395037
transform 1 0 30912 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_274
timestamp 1654395037
transform 1 0 31808 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_278
timestamp 1654395037
transform 1 0 32256 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_280
timestamp 1654395037
transform 1 0 32480 0 1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_8
timestamp 1654395037
transform 1 0 2016 0 -1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_7_73
timestamp 1654395037
transform 1 0 9296 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_81
timestamp 1654395037
transform 1 0 10192 0 -1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_144
timestamp 1654395037
transform 1 0 17248 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_154
timestamp 1654395037
transform 1 0 18368 0 -1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_7_167
timestamp 1654395037
transform 1 0 19824 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_169
timestamp 1654395037
transform 1 0 20048 0 -1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_233
timestamp 1654395037
transform 1 0 27216 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_265
timestamp 1654395037
transform 1 0 30800 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_54
timestamp 1654395037
transform 1 0 7168 0 1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_59
timestamp 1654395037
transform 1 0 7728 0 1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_8_79
timestamp 1654395037
transform 1 0 9968 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_81
timestamp 1654395037
transform 1 0 10192 0 1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_116
timestamp 1654395037
transform 1 0 14112 0 1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_135
timestamp 1654395037
transform 1 0 16240 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_157
timestamp 1654395037
transform 1 0 18704 0 1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1654395037
transform 1 0 20384 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1654395037
transform 1 0 20832 0 1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_179
timestamp 1654395037
transform 1 0 21168 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_201
timestamp 1654395037
transform 1 0 23632 0 1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_225
timestamp 1654395037
transform 1 0 26320 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_241
timestamp 1654395037
transform 1 0 28112 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_8_245
timestamp 1654395037
transform 1 0 28560 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1654395037
transform 1 0 28784 0 1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_250
timestamp 1654395037
transform 1 0 29120 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_266
timestamp 1654395037
transform 1 0 30912 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_274
timestamp 1654395037
transform 1 0 31808 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_8_278
timestamp 1654395037
transform 1 0 32256 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_280
timestamp 1654395037
transform 1 0 32480 0 1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_14
timestamp 1654395037
transform 1 0 2688 0 -1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_36
timestamp 1654395037
transform 1 0 5152 0 -1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_51
timestamp 1654395037
transform 1 0 6832 0 -1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_58
timestamp 1654395037
transform 1 0 7616 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1654395037
transform 1 0 8960 0 -1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_107
timestamp 1654395037
transform 1 0 13104 0 -1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_170
timestamp 1654395037
transform 1 0 20160 0 -1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_9_179
timestamp 1654395037
transform 1 0 21168 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_181
timestamp 1654395037
transform 1 0 21392 0 -1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1654395037
transform 1 0 24864 0 -1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_232
timestamp 1654395037
transform 1 0 27104 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_264
timestamp 1654395037
transform 1 0 30688 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_280
timestamp 1654395037
transform 1 0 32480 0 -1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_25
timestamp 1654395037
transform 1 0 3920 0 1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1654395037
transform 1 0 4928 0 1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_10_51
timestamp 1654395037
transform 1 0 6832 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_53
timestamp 1654395037
transform 1 0 7056 0 1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_10_74
timestamp 1654395037
transform 1 0 9408 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_88
timestamp 1654395037
transform 1 0 10976 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_116
timestamp 1654395037
transform 1 0 14112 0 1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_125
timestamp 1654395037
transform 1 0 15120 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_129
timestamp 1654395037
transform 1 0 15568 0 1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_170
timestamp 1654395037
transform 1 0 20160 0 1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_179
timestamp 1654395037
transform 1 0 21168 0 1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_10_186
timestamp 1654395037
transform 1 0 21952 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_194
timestamp 1654395037
transform 1 0 22848 0 1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_201
timestamp 1654395037
transform 1 0 23632 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_239
timestamp 1654395037
transform 1 0 27888 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1654395037
transform 1 0 28784 0 1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_250
timestamp 1654395037
transform 1 0 29120 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_266
timestamp 1654395037
transform 1 0 30912 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_10_270
timestamp 1654395037
transform 1 0 31360 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_272
timestamp 1654395037
transform 1 0 31584 0 1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_8
timestamp 1654395037
transform 1 0 2016 0 -1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_28
timestamp 1654395037
transform 1 0 4256 0 -1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_37
timestamp 1654395037
transform 1 0 5264 0 -1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_52
timestamp 1654395037
transform 1 0 6944 0 -1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_11_69
timestamp 1654395037
transform 1 0 8848 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_81
timestamp 1654395037
transform 1 0 10192 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_135
timestamp 1654395037
transform 1 0 16240 0 -1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_144
timestamp 1654395037
transform 1 0 17248 0 -1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_240
timestamp 1654395037
transform 1 0 28000 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_272
timestamp 1654395037
transform 1 0 31584 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_280
timestamp 1654395037
transform 1 0 32480 0 -1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_94
timestamp 1654395037
transform 1 0 11648 0 1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_135
timestamp 1654395037
transform 1 0 16240 0 1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_151
timestamp 1654395037
transform 1 0 18032 0 1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_164
timestamp 1654395037
transform 1 0 19488 0 1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_187
timestamp 1654395037
transform 1 0 22064 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_195
timestamp 1654395037
transform 1 0 22960 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_199
timestamp 1654395037
transform 1 0 23408 0 1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_202
timestamp 1654395037
transform 1 0 23744 0 1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_219
timestamp 1654395037
transform 1 0 25648 0 1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1654395037
transform 1 0 28336 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1654395037
transform 1 0 28784 0 1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_250
timestamp 1654395037
transform 1 0 29120 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_266
timestamp 1654395037
transform 1 0 30912 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_274
timestamp 1654395037
transform 1 0 31808 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_12_278
timestamp 1654395037
transform 1 0 32256 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_280
timestamp 1654395037
transform 1 0 32480 0 1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_2
timestamp 1654395037
transform 1 0 1344 0 -1 11760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_13_34
timestamp 1654395037
transform 1 0 4928 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_13_99
timestamp 1654395037
transform 1 0 12208 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_13_139
timestamp 1654395037
transform 1 0 16688 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1654395037
transform 1 0 16912 0 -1 11760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_168
timestamp 1654395037
transform 1 0 19936 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_13_176
timestamp 1654395037
transform 1 0 20832 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1654395037
transform 1 0 24864 0 -1 11760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_238
timestamp 1654395037
transform 1 0 27776 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_270
timestamp 1654395037
transform 1 0 31360 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_13_278
timestamp 1654395037
transform 1 0 32256 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_280
timestamp 1654395037
transform 1 0 32480 0 -1 11760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_14_6
timestamp 1654395037
transform 1 0 1792 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_14_33
timestamp 1654395037
transform 1 0 4816 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_56
timestamp 1654395037
transform 1 0 7392 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_14_64
timestamp 1654395037
transform 1 0 8288 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_66
timestamp 1654395037
transform 1 0 8512 0 1 11760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_103
timestamp 1654395037
transform 1 0 12656 0 1 11760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_14_120
timestamp 1654395037
transform 1 0 14560 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_122
timestamp 1654395037
transform 1 0 14784 0 1 11760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_14_179
timestamp 1654395037
transform 1 0 21168 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_191
timestamp 1654395037
transform 1 0 22512 0 1 11760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_206
timestamp 1654395037
transform 1 0 24192 0 1 11760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_237
timestamp 1654395037
transform 1 0 27664 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_241
timestamp 1654395037
transform 1 0 28112 0 1 11760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_267
timestamp 1654395037
transform 1 0 31024 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_14_271
timestamp 1654395037
transform 1 0 31472 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_2
timestamp 1654395037
transform 1 0 1344 0 -1 13328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_47
timestamp 1654395037
transform 1 0 6384 0 -1 13328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_15_73
timestamp 1654395037
transform 1 0 9296 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_104
timestamp 1654395037
transform 1 0 12768 0 -1 13328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_15_140
timestamp 1654395037
transform 1 0 16800 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_15_157
timestamp 1654395037
transform 1 0 18704 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_159
timestamp 1654395037
transform 1 0 18928 0 -1 13328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_186
timestamp 1654395037
transform 1 0 21952 0 -1 13328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_15_242
timestamp 1654395037
transform 1 0 28224 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_267
timestamp 1654395037
transform 1 0 31024 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_275
timestamp 1654395037
transform 1 0 31920 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_15_279
timestamp 1654395037
transform 1 0 32368 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1654395037
transform 1 0 4928 0 1 13328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_16_67
timestamp 1654395037
transform 1 0 8624 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_69
timestamp 1654395037
transform 1 0 8848 0 1 13328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1654395037
transform 1 0 12880 0 1 13328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_108
timestamp 1654395037
transform 1 0 13216 0 1 13328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_16_133
timestamp 1654395037
transform 1 0 16016 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_230
timestamp 1654395037
transform 1 0 26880 0 1 13328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_16_245
timestamp 1654395037
transform 1 0 28560 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1654395037
transform 1 0 28784 0 1 13328
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_273
timestamp 1654395037
transform 1 0 31696 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_37
timestamp 1654395037
transform 1 0 5264 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_45
timestamp 1654395037
transform 1 0 6160 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_49
timestamp 1654395037
transform 1 0 6608 0 -1 14896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_79
timestamp 1654395037
transform 1 0 9968 0 -1 14896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_109
timestamp 1654395037
transform 1 0 13328 0 -1 14896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_144
timestamp 1654395037
transform 1 0 17248 0 -1 14896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_17_175
timestamp 1654395037
transform 1 0 20720 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_17_210
timestamp 1654395037
transform 1 0 24640 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1654395037
transform 1 0 24864 0 -1 14896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_276
timestamp 1654395037
transform 1 0 32032 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_280
timestamp 1654395037
transform 1 0 32480 0 -1 14896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_8
timestamp 1654395037
transform 1 0 2016 0 1 14896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_18_41
timestamp 1654395037
transform 1 0 5712 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_89
timestamp 1654395037
transform 1 0 11088 0 1 14896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1654395037
transform 1 0 12880 0 1 14896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_108
timestamp 1654395037
transform 1 0 13216 0 1 14896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_18_162
timestamp 1654395037
transform 1 0 19264 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_18_175
timestamp 1654395037
transform 1 0 20720 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_202
timestamp 1654395037
transform 1 0 23744 0 1 14896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_230
timestamp 1654395037
transform 1 0 26880 0 1 14896
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_8
timestamp 1654395037
transform 1 0 2016 0 -1 16464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_38
timestamp 1654395037
transform 1 0 5376 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_19_46
timestamp 1654395037
transform 1 0 6272 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_127
timestamp 1654395037
transform 1 0 15344 0 -1 16464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_136
timestamp 1654395037
transform 1 0 16352 0 -1 16464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_152
timestamp 1654395037
transform 1 0 18144 0 -1 16464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_201
timestamp 1654395037
transform 1 0 23632 0 -1 16464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_210
timestamp 1654395037
transform 1 0 24640 0 -1 16464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_246
timestamp 1654395037
transform 1 0 28672 0 -1 16464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_274
timestamp 1654395037
transform 1 0 31808 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_19_278
timestamp 1654395037
transform 1 0 32256 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_280
timestamp 1654395037
transform 1 0 32480 0 -1 16464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_20_33
timestamp 1654395037
transform 1 0 4816 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_37
timestamp 1654395037
transform 1 0 5264 0 1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_20_41
timestamp 1654395037
transform 1 0 5712 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_83
timestamp 1654395037
transform 1 0 10416 0 1 16464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_127
timestamp 1654395037
transform 1 0 15344 0 1 16464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_153
timestamp 1654395037
transform 1 0 18256 0 1 16464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1654395037
transform 1 0 20832 0 1 16464
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_20_193
timestamp 1654395037
transform 1 0 22736 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_20_246
timestamp 1654395037
transform 1 0 28672 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_273
timestamp 1654395037
transform 1 0 31696 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_25
timestamp 1654395037
transform 1 0 3920 0 -1 18032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1654395037
transform 1 0 16912 0 -1 18032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_206
timestamp 1654395037
transform 1 0 24192 0 -1 18032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_21_272
timestamp 1654395037
transform 1 0 31584 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_274
timestamp 1654395037
transform 1 0 31808 0 -1 18032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_21_277
timestamp 1654395037
transform 1 0 32144 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_22_22
timestamp 1654395037
transform 1 0 3584 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_22_32
timestamp 1654395037
transform 1 0 4704 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1654395037
transform 1 0 4928 0 1 18032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_37
timestamp 1654395037
transform 1 0 5264 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_22_41
timestamp 1654395037
transform 1 0 5712 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_183
timestamp 1654395037
transform 1 0 21616 0 1 18032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_22_206
timestamp 1654395037
transform 1 0 24192 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_218
timestamp 1654395037
transform 1 0 25536 0 1 18032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_22_243
timestamp 1654395037
transform 1 0 28336 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_247
timestamp 1654395037
transform 1 0 28784 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_22_255
timestamp 1654395037
transform 1 0 29680 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_257
timestamp 1654395037
transform 1 0 29904 0 1 18032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_22_266
timestamp 1654395037
transform 1 0 30912 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_268
timestamp 1654395037
transform 1 0 31136 0 1 18032
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 1120 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1654395037
transform -1 0 32816 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1654395037
transform 1 0 1120 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1654395037
transform -1 0 32816 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1654395037
transform 1 0 1120 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1654395037
transform -1 0 32816 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1654395037
transform 1 0 1120 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1654395037
transform -1 0 32816 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1654395037
transform 1 0 1120 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1654395037
transform -1 0 32816 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1654395037
transform 1 0 1120 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1654395037
transform -1 0 32816 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1654395037
transform 1 0 1120 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1654395037
transform -1 0 32816 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1654395037
transform 1 0 1120 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1654395037
transform -1 0 32816 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1654395037
transform 1 0 1120 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1654395037
transform -1 0 32816 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1654395037
transform 1 0 1120 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1654395037
transform -1 0 32816 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1654395037
transform 1 0 1120 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1654395037
transform -1 0 32816 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1654395037
transform 1 0 1120 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1654395037
transform -1 0 32816 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1654395037
transform 1 0 1120 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1654395037
transform -1 0 32816 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1654395037
transform 1 0 1120 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1654395037
transform -1 0 32816 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1654395037
transform 1 0 1120 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1654395037
transform -1 0 32816 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1654395037
transform 1 0 1120 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1654395037
transform -1 0 32816 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1654395037
transform 1 0 1120 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1654395037
transform -1 0 32816 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1654395037
transform 1 0 1120 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1654395037
transform -1 0 32816 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1654395037
transform 1 0 1120 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1654395037
transform -1 0 32816 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1654395037
transform 1 0 1120 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1654395037
transform -1 0 32816 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1654395037
transform 1 0 1120 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1654395037
transform -1 0 32816 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1654395037
transform 1 0 1120 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1654395037
transform -1 0 32816 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1654395037
transform 1 0 1120 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1654395037
transform -1 0 32816 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_46
timestamp 1654395037
transform 1 0 5040 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_47
timestamp 1654395037
transform 1 0 8960 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_48
timestamp 1654395037
transform 1 0 12880 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_49
timestamp 1654395037
transform 1 0 16800 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_50
timestamp 1654395037
transform 1 0 20720 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_51
timestamp 1654395037
transform 1 0 24640 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_52
timestamp 1654395037
transform 1 0 28560 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_53
timestamp 1654395037
transform 1 0 9072 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_54
timestamp 1654395037
transform 1 0 17024 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_55
timestamp 1654395037
transform 1 0 24976 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_56
timestamp 1654395037
transform 1 0 5040 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_57
timestamp 1654395037
transform 1 0 12992 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_58
timestamp 1654395037
transform 1 0 20944 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_59
timestamp 1654395037
transform 1 0 28896 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_60
timestamp 1654395037
transform 1 0 9072 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_61
timestamp 1654395037
transform 1 0 17024 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_62
timestamp 1654395037
transform 1 0 24976 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_63
timestamp 1654395037
transform 1 0 5040 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_64
timestamp 1654395037
transform 1 0 12992 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_65
timestamp 1654395037
transform 1 0 20944 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_66
timestamp 1654395037
transform 1 0 28896 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_67
timestamp 1654395037
transform 1 0 9072 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_68
timestamp 1654395037
transform 1 0 17024 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_69
timestamp 1654395037
transform 1 0 24976 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_70
timestamp 1654395037
transform 1 0 5040 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_71
timestamp 1654395037
transform 1 0 12992 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_72
timestamp 1654395037
transform 1 0 20944 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_73
timestamp 1654395037
transform 1 0 28896 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_74
timestamp 1654395037
transform 1 0 9072 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_75
timestamp 1654395037
transform 1 0 17024 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_76
timestamp 1654395037
transform 1 0 24976 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_77
timestamp 1654395037
transform 1 0 5040 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_78
timestamp 1654395037
transform 1 0 12992 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_79
timestamp 1654395037
transform 1 0 20944 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_80
timestamp 1654395037
transform 1 0 28896 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_81
timestamp 1654395037
transform 1 0 9072 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_82
timestamp 1654395037
transform 1 0 17024 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_83
timestamp 1654395037
transform 1 0 24976 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_84
timestamp 1654395037
transform 1 0 5040 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_85
timestamp 1654395037
transform 1 0 12992 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_86
timestamp 1654395037
transform 1 0 20944 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_87
timestamp 1654395037
transform 1 0 28896 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_88
timestamp 1654395037
transform 1 0 9072 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_89
timestamp 1654395037
transform 1 0 17024 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_90
timestamp 1654395037
transform 1 0 24976 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_91
timestamp 1654395037
transform 1 0 5040 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_92
timestamp 1654395037
transform 1 0 12992 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_93
timestamp 1654395037
transform 1 0 20944 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_94
timestamp 1654395037
transform 1 0 28896 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_95
timestamp 1654395037
transform 1 0 9072 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_96
timestamp 1654395037
transform 1 0 17024 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_97
timestamp 1654395037
transform 1 0 24976 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_98
timestamp 1654395037
transform 1 0 5040 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_99
timestamp 1654395037
transform 1 0 12992 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_100
timestamp 1654395037
transform 1 0 20944 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_101
timestamp 1654395037
transform 1 0 28896 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_102
timestamp 1654395037
transform 1 0 9072 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_103
timestamp 1654395037
transform 1 0 17024 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_104
timestamp 1654395037
transform 1 0 24976 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_105
timestamp 1654395037
transform 1 0 5040 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_106
timestamp 1654395037
transform 1 0 12992 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_107
timestamp 1654395037
transform 1 0 20944 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_108
timestamp 1654395037
transform 1 0 28896 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_109
timestamp 1654395037
transform 1 0 9072 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110
timestamp 1654395037
transform 1 0 17024 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1654395037
transform 1 0 24976 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1654395037
transform 1 0 5040 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1654395037
transform 1 0 12992 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1654395037
transform 1 0 20944 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1654395037
transform 1 0 28896 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1654395037
transform 1 0 9072 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1654395037
transform 1 0 17024 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1654395037
transform 1 0 24976 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1654395037
transform 1 0 5040 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1654395037
transform 1 0 12992 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1654395037
transform 1 0 20944 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1654395037
transform 1 0 28896 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1654395037
transform 1 0 9072 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1654395037
transform 1 0 17024 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1654395037
transform 1 0 24976 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1654395037
transform 1 0 5040 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1654395037
transform 1 0 8960 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1654395037
transform 1 0 12880 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1654395037
transform 1 0 16800 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1654395037
transform 1 0 20720 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1654395037
transform 1 0 24640 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1654395037
transform 1 0 28560 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _318_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 12320 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _319_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 26544 0 -1 3920
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _320_
timestamp 1654395037
transform -1 0 19824 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _321_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 10864 0 1 7056
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _322_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 12096 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _323_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 10192 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _324_
timestamp 1654395037
transform -1 0 9072 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _325_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 20608 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _326_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 13552 0 -1 5488
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _327_
timestamp 1654395037
transform 1 0 9856 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _328_
timestamp 1654395037
transform -1 0 10304 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _329_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 24976 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _330_
timestamp 1654395037
transform 1 0 10528 0 -1 3920
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _331_
timestamp 1654395037
transform 1 0 8288 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _332_
timestamp 1654395037
transform 1 0 4256 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _333_
timestamp 1654395037
transform 1 0 10976 0 1 784
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _334_
timestamp 1654395037
transform 1 0 6496 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _335_
timestamp 1654395037
transform 1 0 13552 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _336_
timestamp 1654395037
transform 1 0 14224 0 1 784
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _337_
timestamp 1654395037
transform 1 0 10304 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _338_
timestamp 1654395037
transform 1 0 18816 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _339_
timestamp 1654395037
transform -1 0 20944 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _340_
timestamp 1654395037
transform 1 0 19824 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _341_
timestamp 1654395037
transform -1 0 8848 0 -1 2352
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _342_
timestamp 1654395037
transform -1 0 7056 0 -1 7056
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _343_
timestamp 1654395037
transform -1 0 2912 0 1 2352
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _344_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 4592 0 -1 3920
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _345_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 3360 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _346_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 4928 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _347_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 1680 0 -1 2352
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _348_
timestamp 1654395037
transform 1 0 4928 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _349_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 2240 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _350_
timestamp 1654395037
transform 1 0 1344 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _351_
timestamp 1654395037
transform -1 0 6608 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _352_
timestamp 1654395037
transform -1 0 8848 0 1 3920
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _353_
timestamp 1654395037
transform -1 0 7168 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _354_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 4928 0 -1 2352
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _355_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 7504 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _356_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 9072 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _357_
timestamp 1654395037
transform 1 0 5264 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _358_
timestamp 1654395037
transform -1 0 9856 0 -1 3920
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _359_
timestamp 1654395037
transform -1 0 5040 0 1 2352
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _360_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 7056 0 1 2352
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _361_
timestamp 1654395037
transform 1 0 7504 0 -1 5488
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _362_
timestamp 1654395037
transform 1 0 8064 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _363_
timestamp 1654395037
transform -1 0 5712 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _364_
timestamp 1654395037
transform 1 0 5376 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _365_
timestamp 1654395037
transform -1 0 8064 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _366_
timestamp 1654395037
transform -1 0 6048 0 -1 3920
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _367_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 1344 0 1 3920
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _368_
timestamp 1654395037
transform -1 0 8064 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _369_
timestamp 1654395037
transform -1 0 7840 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _370_
timestamp 1654395037
transform -1 0 6608 0 1 2352
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _371_
timestamp 1654395037
transform 1 0 1344 0 -1 5488
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _372_
timestamp 1654395037
transform -1 0 3136 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _373_
timestamp 1654395037
transform -1 0 5040 0 1 3920
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _374_
timestamp 1654395037
transform -1 0 2688 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _375_
timestamp 1654395037
transform -1 0 3696 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _376_
timestamp 1654395037
transform 1 0 2688 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _377_
timestamp 1654395037
transform -1 0 8400 0 -1 7056
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _378_
timestamp 1654395037
transform -1 0 6272 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _379_
timestamp 1654395037
transform -1 0 8400 0 1 5488
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _380_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 7504 0 -1 5488
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _381_
timestamp 1654395037
transform -1 0 4256 0 -1 8624
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _382_
timestamp 1654395037
transform 1 0 2128 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _383_
timestamp 1654395037
transform 1 0 1344 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _384_
timestamp 1654395037
transform 1 0 3920 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _385_
timestamp 1654395037
transform -1 0 6608 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _386_
timestamp 1654395037
transform 1 0 3920 0 -1 7056
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _387_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 3920 0 1 7056
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _388_
timestamp 1654395037
transform 1 0 5376 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _389_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 5264 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _390_
timestamp 1654395037
transform 1 0 9744 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _391_
timestamp 1654395037
transform 1 0 17696 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _392_
timestamp 1654395037
transform -1 0 10640 0 -1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _393_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 9632 0 1 8624
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _394_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 24976 0 -1 7056
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _395_
timestamp 1654395037
transform -1 0 7168 0 1 7056
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _396_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 3360 0 1 3920
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _397_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 3584 0 1 5488
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _398_
timestamp 1654395037
transform 1 0 10528 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _399_
timestamp 1654395037
transform 1 0 12208 0 1 7056
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _400_
timestamp 1654395037
transform -1 0 17920 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _401_
timestamp 1654395037
transform -1 0 15232 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _402_
timestamp 1654395037
transform 1 0 10640 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _403_
timestamp 1654395037
transform 1 0 14336 0 -1 10192
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _404_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 11760 0 -1 13328
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _405_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 14336 0 -1 10192
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _406_
timestamp 1654395037
transform -1 0 12096 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _407_
timestamp 1654395037
transform 1 0 12320 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _408_
timestamp 1654395037
transform 1 0 11088 0 1 10192
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _409_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 19824 0 1 11760
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _410_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 12208 0 1 10192
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _411_
timestamp 1654395037
transform 1 0 14000 0 1 10192
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _412_
timestamp 1654395037
transform 1 0 9744 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _413_
timestamp 1654395037
transform 1 0 10640 0 -1 13328
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _414_
timestamp 1654395037
transform 1 0 5152 0 -1 11760
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _415_
timestamp 1654395037
transform -1 0 11760 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _416_
timestamp 1654395037
transform -1 0 9408 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _417_
timestamp 1654395037
transform 1 0 5264 0 -1 8624
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _418_
timestamp 1654395037
transform -1 0 7616 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _419_
timestamp 1654395037
transform 1 0 6048 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _420_
timestamp 1654395037
transform 1 0 10752 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _421_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 6496 0 -1 11760
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _422_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 11760 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _423_
timestamp 1654395037
transform 1 0 13216 0 1 11760
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _424_
timestamp 1654395037
transform 1 0 13216 0 1 10192
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _425_
timestamp 1654395037
transform -1 0 14784 0 -1 11760
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _426_
timestamp 1654395037
transform 1 0 18592 0 -1 11760
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _427_
timestamp 1654395037
transform 1 0 21168 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _428_
timestamp 1654395037
transform 1 0 17248 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _429_
timestamp 1654395037
transform -1 0 14224 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _430_
timestamp 1654395037
transform 1 0 12432 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _431_
timestamp 1654395037
transform -1 0 15792 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _432_
timestamp 1654395037
transform 1 0 15232 0 -1 11760
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _433_
timestamp 1654395037
transform 1 0 16352 0 1 10192
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _434_
timestamp 1654395037
transform 1 0 16352 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _435_
timestamp 1654395037
transform 1 0 13216 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _436_
timestamp 1654395037
transform -1 0 15120 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _437_
timestamp 1654395037
transform -1 0 16240 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _438_
timestamp 1654395037
transform 1 0 15344 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _439_
timestamp 1654395037
transform 1 0 15568 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _440_
timestamp 1654395037
transform -1 0 24752 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _441_
timestamp 1654395037
transform -1 0 24192 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _442_
timestamp 1654395037
transform 1 0 8624 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _443_
timestamp 1654395037
transform 1 0 7952 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _444_
timestamp 1654395037
transform 1 0 11088 0 -1 11760
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _445_
timestamp 1654395037
transform 1 0 9296 0 1 10192
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _446_
timestamp 1654395037
transform 1 0 19600 0 1 10192
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _447_
timestamp 1654395037
transform 1 0 21392 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _448_
timestamp 1654395037
transform 1 0 7056 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _449_
timestamp 1654395037
transform -1 0 12208 0 -1 11760
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _450_
timestamp 1654395037
transform 1 0 9296 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _451_
timestamp 1654395037
transform 1 0 4368 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _452_
timestamp 1654395037
transform 1 0 8064 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _453_
timestamp 1654395037
transform 1 0 7168 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _454_
timestamp 1654395037
transform -1 0 8960 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _455_
timestamp 1654395037
transform 1 0 8400 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _456_
timestamp 1654395037
transform 1 0 11760 0 -1 10192
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _457_
timestamp 1654395037
transform -1 0 12992 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _458_
timestamp 1654395037
transform 1 0 13216 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _459_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 13664 0 -1 3920
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _460_
timestamp 1654395037
transform -1 0 13776 0 1 3920
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _461_
timestamp 1654395037
transform -1 0 12992 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _462_
timestamp 1654395037
transform 1 0 12320 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _463_
timestamp 1654395037
transform -1 0 13664 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _464_
timestamp 1654395037
transform 1 0 14000 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _465_
timestamp 1654395037
transform -1 0 12992 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _466_
timestamp 1654395037
transform 1 0 13328 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _467_
timestamp 1654395037
transform -1 0 16016 0 -1 5488
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _468_
timestamp 1654395037
transform -1 0 14672 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _469_
timestamp 1654395037
transform 1 0 15792 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _470_
timestamp 1654395037
transform -1 0 15792 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _471_
timestamp 1654395037
transform 1 0 15904 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _472_
timestamp 1654395037
transform 1 0 13664 0 1 2352
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _473_
timestamp 1654395037
transform 1 0 14896 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _474_
timestamp 1654395037
transform 1 0 17024 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _475_
timestamp 1654395037
transform 1 0 16016 0 -1 5488
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _476_
timestamp 1654395037
transform -1 0 22400 0 -1 5488
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _477_
timestamp 1654395037
transform -1 0 25872 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _478_
timestamp 1654395037
transform -1 0 24080 0 -1 5488
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _479_
timestamp 1654395037
transform -1 0 26432 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _480_
timestamp 1654395037
transform 1 0 19824 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _481_
timestamp 1654395037
transform -1 0 21840 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _482_
timestamp 1654395037
transform 1 0 6944 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _483_
timestamp 1654395037
transform 1 0 5264 0 1 11760
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _484_
timestamp 1654395037
transform 1 0 1680 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _485_
timestamp 1654395037
transform 1 0 10416 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _486_
timestamp 1654395037
transform -1 0 12208 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _487_
timestamp 1654395037
transform 1 0 19936 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _488_
timestamp 1654395037
transform 1 0 18032 0 1 13328
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _489_
timestamp 1654395037
transform -1 0 21952 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _490_
timestamp 1654395037
transform -1 0 9072 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _491_
timestamp 1654395037
transform -1 0 10752 0 1 13328
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _492_
timestamp 1654395037
transform 1 0 6832 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _493_
timestamp 1654395037
transform -1 0 6160 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _494_
timestamp 1654395037
transform 1 0 11984 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _495_
timestamp 1654395037
transform 1 0 12656 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _496_
timestamp 1654395037
transform 1 0 2016 0 1 13328
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _497_
timestamp 1654395037
transform 1 0 2576 0 1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _498_
timestamp 1654395037
transform -1 0 8176 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _499_
timestamp 1654395037
transform 1 0 6720 0 -1 13328
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _500_
timestamp 1654395037
transform -1 0 8624 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _501_
timestamp 1654395037
transform 1 0 6160 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _502_
timestamp 1654395037
transform 1 0 2240 0 -1 18032
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _503_
timestamp 1654395037
transform 1 0 17920 0 -1 13328
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _504_
timestamp 1654395037
transform 1 0 15792 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _505_
timestamp 1654395037
transform -1 0 14224 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _506_
timestamp 1654395037
transform -1 0 7168 0 -1 18032
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _507_
timestamp 1654395037
transform -1 0 20160 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _508_
timestamp 1654395037
transform 1 0 12880 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _509_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 13440 0 -1 14896
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _510_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 11984 0 1 11760
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _511_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 15344 0 -1 16464
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _512_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 14224 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _513_
timestamp 1654395037
transform 1 0 11424 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _514_
timestamp 1654395037
transform 1 0 10864 0 -1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _515_
timestamp 1654395037
transform -1 0 12768 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _516_
timestamp 1654395037
transform -1 0 11872 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _517_
timestamp 1654395037
transform 1 0 3248 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _518_
timestamp 1654395037
transform 1 0 18368 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _519_
timestamp 1654395037
transform -1 0 19264 0 -1 16464
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _520_
timestamp 1654395037
transform 1 0 14224 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _521_
timestamp 1654395037
transform 1 0 17920 0 1 11760
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _522_
timestamp 1654395037
transform -1 0 21280 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _523_
timestamp 1654395037
transform -1 0 16352 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _524_
timestamp 1654395037
transform -1 0 17024 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _525_
timestamp 1654395037
transform 1 0 9856 0 1 18032
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _526_
timestamp 1654395037
transform 1 0 15680 0 1 18032
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _527_
timestamp 1654395037
transform -1 0 18816 0 1 18032
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _528_
timestamp 1654395037
transform -1 0 16800 0 1 18032
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _529_
timestamp 1654395037
transform 1 0 11200 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _530_
timestamp 1654395037
transform 1 0 10640 0 -1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _531_
timestamp 1654395037
transform 1 0 11872 0 1 14896
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _532_
timestamp 1654395037
transform 1 0 27664 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _533_
timestamp 1654395037
transform 1 0 11760 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _534_
timestamp 1654395037
transform 1 0 27664 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _535_
timestamp 1654395037
transform 1 0 11200 0 -1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _536_
timestamp 1654395037
transform 1 0 11648 0 1 13328
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _537_
timestamp 1654395037
transform 1 0 24304 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _538_
timestamp 1654395037
transform -1 0 22288 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _539_
timestamp 1654395037
transform -1 0 22512 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _540_
timestamp 1654395037
transform 1 0 20160 0 1 13328
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _541_
timestamp 1654395037
transform 1 0 16464 0 -1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _542_
timestamp 1654395037
transform -1 0 10976 0 1 18032
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _543_
timestamp 1654395037
transform 1 0 17696 0 1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _544_
timestamp 1654395037
transform 1 0 15456 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _545_
timestamp 1654395037
transform 1 0 17696 0 1 18032
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _546_
timestamp 1654395037
transform -1 0 11536 0 1 18032
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _547_
timestamp 1654395037
transform 1 0 21392 0 -1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _548_
timestamp 1654395037
transform 1 0 17248 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _549_
timestamp 1654395037
transform -1 0 18256 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _550_
timestamp 1654395037
transform -1 0 19488 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _551_
timestamp 1654395037
transform 1 0 21952 0 -1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _552_
timestamp 1654395037
transform 1 0 13888 0 1 13328
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _553_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 14448 0 -1 14896
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _554_
timestamp 1654395037
transform 1 0 22848 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _555_
timestamp 1654395037
transform 1 0 17808 0 1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _556_
timestamp 1654395037
transform 1 0 21168 0 1 13328
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _557_
timestamp 1654395037
transform 1 0 13328 0 1 13328
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _558_
timestamp 1654395037
transform 1 0 15792 0 -1 13328
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _559_
timestamp 1654395037
transform 1 0 14896 0 1 13328
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _560_
timestamp 1654395037
transform -1 0 22064 0 1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _561_
timestamp 1654395037
transform 1 0 8960 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _562_
timestamp 1654395037
transform 1 0 18256 0 -1 14896
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _563_
timestamp 1654395037
transform 1 0 19040 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _564_
timestamp 1654395037
transform -1 0 20832 0 1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _565_
timestamp 1654395037
transform 1 0 19600 0 -1 14896
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _566_
timestamp 1654395037
transform -1 0 20496 0 1 14896
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _567_
timestamp 1654395037
transform 1 0 2128 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _568_
timestamp 1654395037
transform -1 0 25760 0 -1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _569_
timestamp 1654395037
transform 1 0 20944 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _570_
timestamp 1654395037
transform -1 0 23520 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _571_
timestamp 1654395037
transform 1 0 23744 0 1 13328
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _572_
timestamp 1654395037
transform 1 0 21616 0 1 14896
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _573_
timestamp 1654395037
transform 1 0 23072 0 -1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _574_
timestamp 1654395037
transform -1 0 17248 0 1 11760
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _575_
timestamp 1654395037
transform 1 0 15120 0 1 14896
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _576_
timestamp 1654395037
transform 1 0 15904 0 1 14896
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _577_
timestamp 1654395037
transform -1 0 26320 0 -1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _578_
timestamp 1654395037
transform 1 0 17248 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _579_
timestamp 1654395037
transform -1 0 6608 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _580_
timestamp 1654395037
transform 1 0 21728 0 1 13328
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _581_
timestamp 1654395037
transform 1 0 22512 0 -1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _582_
timestamp 1654395037
transform 1 0 21840 0 -1 14896
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _583_
timestamp 1654395037
transform -1 0 29680 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _584_
timestamp 1654395037
transform 1 0 22400 0 1 14896
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _585_
timestamp 1654395037
transform -1 0 17808 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _586_
timestamp 1654395037
transform -1 0 18592 0 -1 18032
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _587_
timestamp 1654395037
transform -1 0 18032 0 -1 18032
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _588_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 16240 0 1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _589_
timestamp 1654395037
transform 1 0 23184 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _590_
timestamp 1654395037
transform -1 0 26880 0 1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _591_
timestamp 1654395037
transform 1 0 25200 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _592_
timestamp 1654395037
transform -1 0 24528 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _593_
timestamp 1654395037
transform -1 0 32032 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _594_
timestamp 1654395037
transform 1 0 24976 0 1 14896
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _595_
timestamp 1654395037
transform -1 0 27104 0 -1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _596_
timestamp 1654395037
transform -1 0 25200 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _597_
timestamp 1654395037
transform 1 0 23520 0 -1 14896
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _598_
timestamp 1654395037
transform 1 0 27104 0 -1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _599_
timestamp 1654395037
transform -1 0 27776 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _600_
timestamp 1654395037
transform 1 0 25984 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _601_
timestamp 1654395037
transform 1 0 26992 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _602_
timestamp 1654395037
transform -1 0 24864 0 1 11760
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _603_
timestamp 1654395037
transform 1 0 25200 0 1 13328
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _604_
timestamp 1654395037
transform -1 0 22960 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _605_
timestamp 1654395037
transform -1 0 23520 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _606_
timestamp 1654395037
transform 1 0 23856 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _607_
timestamp 1654395037
transform -1 0 8400 0 1 7056
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _608_
timestamp 1654395037
transform -1 0 19376 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _609_
timestamp 1654395037
transform 1 0 19488 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _610_
timestamp 1654395037
transform 1 0 18480 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _611_
timestamp 1654395037
transform -1 0 25872 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _612_
timestamp 1654395037
transform -1 0 23632 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _613_
timestamp 1654395037
transform 1 0 25872 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _614_
timestamp 1654395037
transform -1 0 27216 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _615_
timestamp 1654395037
transform 1 0 25872 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _616_
timestamp 1654395037
transform -1 0 25984 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _617_
timestamp 1654395037
transform 1 0 20160 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _618_
timestamp 1654395037
transform -1 0 21616 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _619_
timestamp 1654395037
transform 1 0 17696 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _620_
timestamp 1654395037
transform 1 0 19600 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _621_
timestamp 1654395037
transform -1 0 19600 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _622_
timestamp 1654395037
transform -1 0 18032 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _623_
timestamp 1654395037
transform 1 0 18032 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _624_
timestamp 1654395037
transform -1 0 20944 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _625_
timestamp 1654395037
transform -1 0 19376 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _626_
timestamp 1654395037
transform -1 0 18816 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _627_
timestamp 1654395037
transform -1 0 17920 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _628_
timestamp 1654395037
transform 1 0 14224 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _629_
timestamp 1654395037
transform -1 0 17360 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _630_
timestamp 1654395037
transform 1 0 14896 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _631_
timestamp 1654395037
transform 1 0 19712 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _632_
timestamp 1654395037
transform -1 0 18704 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _633_
timestamp 1654395037
transform -1 0 18144 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _634_
timestamp 1654395037
transform 1 0 19040 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _635_
timestamp 1654395037
transform -1 0 20160 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _636_
timestamp 1654395037
transform -1 0 18816 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _637_
timestamp 1654395037
transform 1 0 21280 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _638_
timestamp 1654395037
transform 1 0 22960 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _639_
timestamp 1654395037
transform -1 0 20160 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _640_
timestamp 1654395037
transform -1 0 19488 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _641_
timestamp 1654395037
transform 1 0 20272 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _642_
timestamp 1654395037
transform -1 0 20944 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _643_
timestamp 1654395037
transform 1 0 19152 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _644_
timestamp 1654395037
transform -1 0 22288 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _645_
timestamp 1654395037
transform 1 0 23520 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _646_
timestamp 1654395037
transform -1 0 19712 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _647_
timestamp 1654395037
transform 1 0 21616 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _648_
timestamp 1654395037
transform -1 0 22960 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _649_
timestamp 1654395037
transform 1 0 23632 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _650_
timestamp 1654395037
transform 1 0 22960 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _651_
timestamp 1654395037
transform 1 0 22960 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _652_
timestamp 1654395037
transform -1 0 25648 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _653_
timestamp 1654395037
transform -1 0 22960 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _654_
timestamp 1654395037
transform -1 0 18368 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _655_
timestamp 1654395037
transform 1 0 17808 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _656_
timestamp 1654395037
transform -1 0 19040 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _657_
timestamp 1654395037
transform -1 0 10528 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _658_
timestamp 1654395037
transform 1 0 9184 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _659_
timestamp 1654395037
transform 1 0 10528 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _660_
timestamp 1654395037
transform 1 0 12208 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _661_
timestamp 1654395037
transform -1 0 11872 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _662_
timestamp 1654395037
transform 1 0 10864 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _663_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 20160 0 -1 7056
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _664_
timestamp 1654395037
transform -1 0 25760 0 1 5488
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _665_
timestamp 1654395037
transform -1 0 25312 0 1 3920
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _666_
timestamp 1654395037
transform 1 0 17248 0 -1 3920
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _667_
timestamp 1654395037
transform -1 0 18928 0 1 2352
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _668_
timestamp 1654395037
transform 1 0 15792 0 1 3920
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _669_
timestamp 1654395037
transform 1 0 14896 0 1 5488
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _670_
timestamp 1654395037
transform 1 0 12992 0 -1 7056
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _671_
timestamp 1654395037
transform 1 0 13216 0 -1 8624
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _672_
timestamp 1654395037
transform 1 0 9296 0 -1 8624
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _673_
timestamp 1654395037
transform 1 0 5264 0 1 10192
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _674_
timestamp 1654395037
transform 1 0 21056 0 -1 11760
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _675_
timestamp 1654395037
transform 1 0 15680 0 1 8624
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _676_
timestamp 1654395037
transform 1 0 17360 0 -1 10192
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _677_
timestamp 1654395037
transform 1 0 21168 0 -1 10192
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _678_
timestamp 1654395037
transform 1 0 18480 0 -1 2352
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _679_
timestamp 1654395037
transform 1 0 21056 0 -1 3920
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _680_
timestamp 1654395037
transform 1 0 21168 0 1 2352
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _681_
timestamp 1654395037
transform 1 0 13216 0 -1 2352
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _682_
timestamp 1654395037
transform 1 0 9408 0 -1 2352
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _683_
timestamp 1654395037
transform -1 0 12880 0 1 2352
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _684_
timestamp 1654395037
transform 1 0 9744 0 -1 5488
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _685_
timestamp 1654395037
transform 1 0 8400 0 1 5488
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _686_
timestamp 1654395037
transform -1 0 4928 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  input1
timestamp 1654395037
transform 1 0 3248 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1654395037
transform -1 0 5936 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1654395037
transform -1 0 6608 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1654395037
transform -1 0 4928 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1654395037
transform -1 0 3696 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1654395037
transform 1 0 1344 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1654395037
transform 1 0 1344 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1654395037
transform 1 0 1344 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1654395037
transform 1 0 9184 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1654395037
transform 1 0 11536 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1654395037
transform -1 0 15680 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1654395037
transform 1 0 17024 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1654395037
transform 1 0 20944 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1654395037
transform -1 0 22848 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1654395037
transform 1 0 24864 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1654395037
transform -1 0 27440 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1654395037
transform -1 0 30688 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1654395037
transform -1 0 32592 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1654395037
transform 1 0 1344 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1654395037
transform -1 0 31920 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1654395037
transform -1 0 32592 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1654395037
transform -1 0 32592 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1654395037
transform -1 0 32592 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1654395037
transform -1 0 32592 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1654395037
transform -1 0 32592 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1654395037
transform 1 0 1344 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1654395037
transform 1 0 1344 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1654395037
transform 1 0 1344 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1654395037
transform 1 0 2016 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1654395037
transform 1 0 1344 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1654395037
transform 1 0 1344 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1654395037
transform 1 0 3808 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1654395037
transform 1 0 6384 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1654395037
transform -1 0 26208 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1654395037
transform -1 0 9744 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output36 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 4480 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output37 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 1344 0 1 784
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  rebuffer1
timestamp 1654395037
transform 1 0 12208 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  rebuffer2
timestamp 1654395037
transform -1 0 16688 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[0\].id.delaybuf0
timestamp 1654395037
transform -1 0 22848 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp 1654395037
transform -1 0 4704 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[0\].id.delayen0 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 2352 0 -1 11760
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[0\].id.delayen1
timestamp 1654395037
transform 1 0 2128 0 -1 10192
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[0\].id.delayenb0
timestamp 1654395037
transform 1 0 1344 0 1 10192
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[0\].id.delayenb1
timestamp 1654395037
transform 1 0 1792 0 1 8624
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  ringosc.dstage\[0\].id.delayint0 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 4256 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[0\].id.trim0bar
timestamp 1654395037
transform -1 0 4928 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[0\].id.trim1bar
timestamp 1654395037
transform 1 0 1344 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[1\].id.delaybuf0
timestamp 1654395037
transform -1 0 4816 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1654395037
transform 1 0 1904 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[1\].id.delayen0
timestamp 1654395037
transform 1 0 2576 0 1 13328
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[1\].id.delayen1
timestamp 1654395037
transform -1 0 6384 0 -1 13328
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[1\].id.delayenb0
timestamp 1654395037
transform 1 0 2576 0 -1 13328
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[1\].id.delayenb1
timestamp 1654395037
transform -1 0 4144 0 1 11760
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  ringosc.dstage\[1\].id.delayint0
timestamp 1654395037
transform 1 0 3920 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[1\].id.trim0bar
timestamp 1654395037
transform 1 0 1456 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[1\].id.trim1bar
timestamp 1654395037
transform -1 0 5712 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[2\].id.delaybuf0
timestamp 1654395037
transform -1 0 5264 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1654395037
transform 1 0 4144 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[2\].id.delayen0
timestamp 1654395037
transform 1 0 3136 0 1 14896
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[2\].id.delayen1
timestamp 1654395037
transform 1 0 2800 0 -1 16464
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[2\].id.delayenb0
timestamp 1654395037
transform 1 0 2016 0 -1 14896
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[2\].id.delayenb1
timestamp 1654395037
transform 1 0 2240 0 1 16464
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  ringosc.dstage\[2\].id.delayint0
timestamp 1654395037
transform 1 0 4704 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[2\].id.trim0bar
timestamp 1654395037
transform -1 0 5712 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[2\].id.trim1bar
timestamp 1654395037
transform -1 0 3248 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[3\].id.delaybuf0
timestamp 1654395037
transform 1 0 5936 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1654395037
transform -1 0 9968 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[3\].id.delayen0
timestamp 1654395037
transform 1 0 8512 0 1 14896
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[3\].id.delayen1
timestamp 1654395037
transform 1 0 6608 0 1 14896
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[3\].id.delayenb0
timestamp 1654395037
transform 1 0 7168 0 -1 14896
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[3\].id.delayenb1
timestamp 1654395037
transform 1 0 6944 0 -1 16464
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  ringosc.dstage\[3\].id.delayint0
timestamp 1654395037
transform 1 0 10416 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[3\].id.trim0bar
timestamp 1654395037
transform 1 0 6720 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[3\].id.trim1bar
timestamp 1654395037
transform 1 0 6496 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[4\].id.delaybuf0
timestamp 1654395037
transform 1 0 9296 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1654395037
transform -1 0 10640 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[4\].id.delayen0
timestamp 1654395037
transform 1 0 8512 0 1 16464
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[4\].id.delayen1
timestamp 1654395037
transform 1 0 7056 0 1 18032
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[4\].id.delayenb0
timestamp 1654395037
transform 1 0 7168 0 -1 18032
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[4\].id.delayenb1
timestamp 1654395037
transform 1 0 6608 0 1 16464
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  ringosc.dstage\[4\].id.delayint0
timestamp 1654395037
transform 1 0 9296 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[4\].id.trim0bar
timestamp 1654395037
transform 1 0 6160 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[4\].id.trim1bar
timestamp 1654395037
transform 1 0 5712 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[5\].id.delaybuf0
timestamp 1654395037
transform 1 0 10528 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1654395037
transform -1 0 16016 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[5\].id.delayen0
timestamp 1654395037
transform 1 0 13216 0 1 16464
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[5\].id.delayen1
timestamp 1654395037
transform 1 0 13104 0 1 18032
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[5\].id.delayenb0
timestamp 1654395037
transform 1 0 12768 0 -1 18032
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[5\].id.delayenb1
timestamp 1654395037
transform 1 0 10864 0 -1 18032
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  ringosc.dstage\[5\].id.delayint0
timestamp 1654395037
transform 1 0 14672 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[5\].id.trim0bar
timestamp 1654395037
transform 1 0 10416 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[5\].id.trim1bar
timestamp 1654395037
transform 1 0 9968 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[6\].id.delaybuf0
timestamp 1654395037
transform 1 0 17024 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1654395037
transform -1 0 21168 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[6\].id.delayen0
timestamp 1654395037
transform 1 0 19488 0 -1 16464
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[6\].id.delayen1
timestamp 1654395037
transform 1 0 18816 0 1 18032
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[6\].id.delayenb0
timestamp 1654395037
transform -1 0 20272 0 1 16464
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[6\].id.delayenb1
timestamp 1654395037
transform -1 0 20496 0 -1 18032
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  ringosc.dstage\[6\].id.delayint0
timestamp 1654395037
transform 1 0 21168 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[6\].id.trim0bar
timestamp 1654395037
transform -1 0 21616 0 1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[6\].id.trim1bar
timestamp 1654395037
transform -1 0 23296 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[7\].id.delaybuf0
timestamp 1654395037
transform 1 0 22064 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1654395037
transform 1 0 23968 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[7\].id.delayen0
timestamp 1654395037
transform -1 0 27104 0 -1 18032
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[7\].id.delayen1
timestamp 1654395037
transform -1 0 26768 0 1 16464
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[7\].id.delayenb0
timestamp 1654395037
transform 1 0 22288 0 -1 18032
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[7\].id.delayenb1
timestamp 1654395037
transform 1 0 22960 0 1 16464
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  ringosc.dstage\[7\].id.delayint0
timestamp 1654395037
transform 1 0 24304 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[7\].id.trim0bar
timestamp 1654395037
transform 1 0 21728 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[7\].id.trim1bar
timestamp 1654395037
transform -1 0 23744 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[8\].id.delaybuf0
timestamp 1654395037
transform 1 0 26096 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1654395037
transform 1 0 27440 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[8\].id.delayen0
timestamp 1654395037
transform 1 0 29008 0 -1 18032
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[8\].id.delayen1
timestamp 1654395037
transform 1 0 26768 0 1 16464
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[8\].id.delayenb0
timestamp 1654395037
transform 1 0 27104 0 -1 18032
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[8\].id.delayenb1
timestamp 1654395037
transform -1 0 28224 0 -1 16464
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  ringosc.dstage\[8\].id.delayint0
timestamp 1654395037
transform 1 0 31024 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[8\].id.trim0bar
timestamp 1654395037
transform 1 0 25648 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[8\].id.trim1bar
timestamp 1654395037
transform -1 0 28672 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[9\].id.delaybuf0
timestamp 1654395037
transform -1 0 31584 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1654395037
transform -1 0 31360 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[9\].id.delayen0
timestamp 1654395037
transform 1 0 28784 0 -1 16464
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[9\].id.delayen1
timestamp 1654395037
transform 1 0 26992 0 1 14896
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[9\].id.delayenb0
timestamp 1654395037
transform 1 0 29120 0 1 14896
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[9\].id.delayenb1
timestamp 1654395037
transform 1 0 29120 0 1 16464
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  ringosc.dstage\[9\].id.delayint0
timestamp 1654395037
transform 1 0 31024 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[9\].id.trim0bar
timestamp 1654395037
transform 1 0 28112 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[9\].id.trim1bar
timestamp 1654395037
transform -1 0 31808 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[10\].id.delaybuf0
timestamp 1654395037
transform 1 0 30912 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1654395037
transform -1 0 31696 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[10\].id.delayen0
timestamp 1654395037
transform 1 0 29120 0 1 11760
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[10\].id.delayen1
timestamp 1654395037
transform 1 0 29008 0 -1 14896
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[10\].id.delayenb0
timestamp 1654395037
transform 1 0 28448 0 -1 13328
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[10\].id.delayenb1
timestamp 1654395037
transform 1 0 29120 0 1 13328
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  ringosc.dstage\[10\].id.delayint0
timestamp 1654395037
transform 1 0 30352 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[10\].id.trim0bar
timestamp 1654395037
transform 1 0 28112 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[10\].id.trim1bar
timestamp 1654395037
transform 1 0 28560 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[11\].id.delaybuf0
timestamp 1654395037
transform -1 0 28896 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1654395037
transform -1 0 27440 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  ringosc.dstage\[11\].id.delayen0 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 25200 0 -1 11760
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[11\].id.delayen1
timestamp 1654395037
transform 1 0 25200 0 -1 13328
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  ringosc.dstage\[11\].id.delayenb0
timestamp 1654395037
transform 1 0 25760 0 1 10192
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.dstage\[11\].id.delayenb1
timestamp 1654395037
transform 1 0 24864 0 1 11760
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  ringosc.dstage\[11\].id.delayint0
timestamp 1654395037
transform 1 0 27104 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[11\].id.trim0bar
timestamp 1654395037
transform 1 0 25200 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.dstage\[11\].id.trim1bar
timestamp 1654395037
transform -1 0 28224 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  ringosc.ibufp00
timestamp 1654395037
transform -1 0 22960 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_8  ringosc.ibufp01 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 23520 0 -1 8624
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  ringosc.ibufp10
timestamp 1654395037
transform -1 0 2800 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  ringosc.ibufp11 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 2688 0 -1 8624
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  ringosc.iss.ctrlen0
timestamp 1654395037
transform 1 0 24192 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1654395037
transform -1 0 28336 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  ringosc.iss.delayen0
timestamp 1654395037
transform 1 0 24080 0 1 8624
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.iss.delayen1
timestamp 1654395037
transform 1 0 25984 0 1 8624
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  ringosc.iss.delayenb0
timestamp 1654395037
transform 1 0 25200 0 -1 8624
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  ringosc.iss.delayenb1
timestamp 1654395037
transform 1 0 25648 0 -1 10192
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.iss.delayint0
timestamp 1654395037
transform -1 0 28000 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  ringosc.iss.reseten0_38 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 26096 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  ringosc.iss.reseten0
timestamp 1654395037
transform 1 0 23744 0 1 7056
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  ringosc.iss.trim1bar
timestamp 1654395037
transform 1 0 24752 0 1 10192
box -86 -86 534 870
<< labels >>
flabel metal4 s 4930 724 5250 18876 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 12870 724 13190 18876 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 20810 724 21130 18876 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 28750 724 29070 18876 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 1060 2928 32876 3248 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 1060 7536 32876 7856 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 1060 12144 32876 12464 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 1060 16752 32876 17072 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 8900 724 9220 18876 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 16840 724 17160 18876 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 24780 724 25100 18876 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 1060 5232 32876 5552 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 1060 9840 32876 10160 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 1060 14448 32876 14768 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal3 s 0 616 800 728 0 FreeSans 448 0 0 0 clockp[0]
port 2 nsew signal tristate
flabel metal3 s 0 1848 800 1960 0 FreeSans 448 0 0 0 clockp[1]
port 3 nsew signal tristate
flabel metal3 s 0 10584 800 10696 0 FreeSans 448 0 0 0 dco
port 4 nsew signal input
flabel metal3 s 0 3080 800 3192 0 FreeSans 448 0 0 0 div[0]
port 5 nsew signal input
flabel metal3 s 0 4312 800 4424 0 FreeSans 448 0 0 0 div[1]
port 6 nsew signal input
flabel metal3 s 0 5544 800 5656 0 FreeSans 448 0 0 0 div[2]
port 7 nsew signal input
flabel metal3 s 0 6776 800 6888 0 FreeSans 448 0 0 0 div[3]
port 8 nsew signal input
flabel metal3 s 0 8008 800 8120 0 FreeSans 448 0 0 0 div[4]
port 9 nsew signal input
flabel metal3 s 0 9240 800 9352 0 FreeSans 448 0 0 0 enable
port 10 nsew signal input
flabel metal3 s 0 11816 800 11928 0 FreeSans 448 0 0 0 ext_trim[0]
port 11 nsew signal input
flabel metal2 s 9016 19200 9128 20000 0 FreeSans 448 90 0 0 ext_trim[10]
port 12 nsew signal input
flabel metal2 s 11592 19200 11704 20000 0 FreeSans 448 90 0 0 ext_trim[11]
port 13 nsew signal input
flabel metal2 s 14168 19200 14280 20000 0 FreeSans 448 90 0 0 ext_trim[12]
port 14 nsew signal input
flabel metal2 s 16856 19200 16968 20000 0 FreeSans 448 90 0 0 ext_trim[13]
port 15 nsew signal input
flabel metal2 s 19432 19200 19544 20000 0 FreeSans 448 90 0 0 ext_trim[14]
port 16 nsew signal input
flabel metal2 s 22120 19200 22232 20000 0 FreeSans 448 90 0 0 ext_trim[15]
port 17 nsew signal input
flabel metal2 s 24696 19200 24808 20000 0 FreeSans 448 90 0 0 ext_trim[16]
port 18 nsew signal input
flabel metal2 s 27272 19200 27384 20000 0 FreeSans 448 90 0 0 ext_trim[17]
port 19 nsew signal input
flabel metal2 s 29960 19200 30072 20000 0 FreeSans 448 90 0 0 ext_trim[18]
port 20 nsew signal input
flabel metal2 s 32536 19200 32648 20000 0 FreeSans 448 90 0 0 ext_trim[19]
port 21 nsew signal input
flabel metal3 s 0 13048 800 13160 0 FreeSans 448 0 0 0 ext_trim[1]
port 22 nsew signal input
flabel metal3 s 33200 18200 34000 18312 0 FreeSans 448 0 0 0 ext_trim[20]
port 23 nsew signal input
flabel metal3 s 33200 14840 34000 14952 0 FreeSans 448 0 0 0 ext_trim[21]
port 24 nsew signal input
flabel metal3 s 33200 11592 34000 11704 0 FreeSans 448 0 0 0 ext_trim[22]
port 25 nsew signal input
flabel metal3 s 33200 8232 34000 8344 0 FreeSans 448 0 0 0 ext_trim[23]
port 26 nsew signal input
flabel metal3 s 33200 4872 34000 4984 0 FreeSans 448 0 0 0 ext_trim[24]
port 27 nsew signal input
flabel metal3 s 33200 1624 34000 1736 0 FreeSans 448 0 0 0 ext_trim[25]
port 28 nsew signal input
flabel metal3 s 0 14280 800 14392 0 FreeSans 448 0 0 0 ext_trim[2]
port 29 nsew signal input
flabel metal3 s 0 15512 800 15624 0 FreeSans 448 0 0 0 ext_trim[3]
port 30 nsew signal input
flabel metal3 s 0 16744 800 16856 0 FreeSans 448 0 0 0 ext_trim[4]
port 31 nsew signal input
flabel metal3 s 0 17976 800 18088 0 FreeSans 448 0 0 0 ext_trim[5]
port 32 nsew signal input
flabel metal3 s 0 19208 800 19320 0 FreeSans 448 0 0 0 ext_trim[6]
port 33 nsew signal input
flabel metal2 s 1176 19200 1288 20000 0 FreeSans 448 90 0 0 ext_trim[7]
port 34 nsew signal input
flabel metal2 s 3752 19200 3864 20000 0 FreeSans 448 90 0 0 ext_trim[8]
port 35 nsew signal input
flabel metal2 s 6328 19200 6440 20000 0 FreeSans 448 90 0 0 ext_trim[9]
port 36 nsew signal input
flabel metal2 s 25480 0 25592 800 0 FreeSans 448 90 0 0 osc
port 37 nsew signal input
flabel metal2 s 8456 0 8568 800 0 FreeSans 448 90 0 0 resetb
port 38 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 34000 20000
<< end >>
