magic
tech gf180mcuD
magscale 1 10
timestamp 1655304105
<< error_p >>
rect -808 -255 -797 -209
rect -594 -255 -583 -209
rect -380 -255 -369 -209
rect -166 -255 -155 -209
rect 53 -255 64 -209
rect 267 -255 278 -209
rect 481 -255 492 -209
rect 695 -255 706 -209
<< nwell >>
rect -1128 -486 1121 486
<< mvpmos >>
rect -810 -176 -700 224
rect -596 -176 -486 224
rect -382 -176 -272 224
rect -168 -176 -58 224
rect 51 -176 161 224
rect 265 -176 375 224
rect 479 -176 589 224
rect 693 -176 803 224
<< mvpdiff >>
rect -898 211 -810 224
rect -898 -163 -885 211
rect -839 -163 -810 211
rect -898 -176 -810 -163
rect -700 211 -596 224
rect -700 -163 -671 211
rect -625 -163 -596 211
rect -700 -176 -596 -163
rect -486 211 -382 224
rect -486 -163 -457 211
rect -411 -163 -382 211
rect -486 -176 -382 -163
rect -272 211 -168 224
rect -272 -163 -243 211
rect -197 -163 -168 211
rect -272 -176 -168 -163
rect -58 211 51 224
rect -58 -163 -29 211
rect 17 -163 51 211
rect -58 -176 51 -163
rect 161 211 265 224
rect 161 -163 190 211
rect 236 -163 265 211
rect 161 -176 265 -163
rect 375 211 479 224
rect 375 -163 404 211
rect 450 -163 479 211
rect 375 -176 479 -163
rect 589 211 693 224
rect 589 -163 618 211
rect 664 -163 693 211
rect 589 -176 693 -163
rect 803 211 891 224
rect 803 -163 832 211
rect 878 -163 891 211
rect 803 -176 891 -163
<< mvpdiffc >>
rect -885 -163 -839 211
rect -671 -163 -625 211
rect -457 -163 -411 211
rect -243 -163 -197 211
rect -29 -163 17 211
rect 190 -163 236 211
rect 404 -163 450 211
rect 618 -163 664 211
rect 832 -163 878 211
<< mvnsubdiff >>
rect -1042 387 1035 400
rect -1042 341 -880 387
rect 880 341 1035 387
rect -1042 328 1035 341
rect -1042 284 -970 328
rect -1042 -284 -1029 284
rect -983 -284 -970 284
rect 963 284 1035 328
rect -1042 -328 -970 -284
rect 963 -284 976 284
rect 1022 -284 1035 284
rect 963 -328 1035 -284
rect -1042 -400 1035 -328
<< mvnsubdiffcont >>
rect -880 341 880 387
rect -1029 -284 -983 284
rect 976 -284 1022 284
<< polysilicon >>
rect -810 224 -700 268
rect -596 224 -486 268
rect -382 224 -272 268
rect -168 224 -58 268
rect 51 224 161 268
rect 265 224 375 268
rect 479 224 589 268
rect 693 224 803 268
rect -810 -209 -700 -176
rect -810 -255 -797 -209
rect -713 -255 -700 -209
rect -810 -268 -700 -255
rect -596 -209 -486 -176
rect -596 -255 -583 -209
rect -499 -255 -486 -209
rect -596 -268 -486 -255
rect -382 -209 -272 -176
rect -382 -255 -369 -209
rect -285 -255 -272 -209
rect -382 -268 -272 -255
rect -168 -209 -58 -176
rect -168 -255 -155 -209
rect -71 -255 -58 -209
rect -168 -268 -58 -255
rect 51 -209 161 -176
rect 51 -255 64 -209
rect 148 -255 161 -209
rect 51 -268 161 -255
rect 265 -209 375 -176
rect 265 -255 278 -209
rect 362 -255 375 -209
rect 265 -268 375 -255
rect 479 -209 589 -176
rect 479 -255 492 -209
rect 576 -255 589 -209
rect 479 -268 589 -255
rect 693 -209 803 -176
rect 693 -255 706 -209
rect 790 -255 803 -209
rect 693 -268 803 -255
<< polycontact >>
rect -797 -255 -713 -209
rect -583 -255 -499 -209
rect -369 -255 -285 -209
rect -155 -255 -71 -209
rect 64 -255 148 -209
rect 278 -255 362 -209
rect 492 -255 576 -209
rect 706 -255 790 -209
<< metal1 >>
rect -1029 341 -880 387
rect 880 341 1022 387
rect -1029 284 -983 341
rect 976 284 1022 341
rect -885 211 -839 222
rect -885 -174 -839 -163
rect -671 211 -625 222
rect -671 -174 -625 -163
rect -457 211 -411 222
rect -457 -174 -411 -163
rect -243 211 -197 222
rect -243 -174 -197 -163
rect -29 211 17 222
rect -29 -174 17 -163
rect 190 211 236 222
rect 190 -174 236 -163
rect 404 211 450 222
rect 404 -174 450 -163
rect 618 211 664 222
rect 618 -174 664 -163
rect 832 211 878 222
rect 832 -174 878 -163
rect -808 -255 -797 -209
rect -713 -255 -702 -209
rect -594 -255 -583 -209
rect -499 -255 -488 -209
rect -380 -255 -369 -209
rect -285 -255 -274 -209
rect -166 -255 -155 -209
rect -71 -255 -60 -209
rect 53 -255 64 -209
rect 148 -255 159 -209
rect 267 -255 278 -209
rect 362 -255 373 -209
rect 481 -255 492 -209
rect 576 -255 587 -209
rect 695 -255 706 -209
rect 790 -255 801 -209
rect -1029 -341 -983 -284
rect 976 -341 1022 -284
rect -1029 -387 1022 -341
<< properties >>
string FIXED_BBOX -960 -364 960 364
string gencell pmos_6p0
string library gf180mcu
string parameters w 2 l 0.5 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.5 wmin 0.3 full_metal 1 compatible {pmos_3p3 pmos_6p0}
<< end >>
