magic
tech gf180mcuD
magscale 1 10
timestamp 1655307388
<< nwell >>
rect 1353 -110 1490 561
rect 1353 -418 2231 -110
rect 1353 -1211 1490 -418
<< metal1 >>
rect 526 385 3034 685
rect 744 -884 883 385
rect 1072 288 1124 300
rect 1072 -872 1124 -860
rect 946 -996 958 -944
rect 1032 -996 1044 -944
rect 946 -1019 1044 -996
rect 1242 -1112 1614 385
rect 1727 309 1779 310
rect 1706 297 1779 309
rect 1706 223 1727 297
rect 1706 209 1779 223
rect 2237 297 2310 310
rect 2289 223 2310 297
rect 2237 210 2310 223
rect 2400 219 2706 385
rect 1841 111 1853 167
rect 2154 111 2166 167
rect 2400 41 2625 219
rect 2696 41 2706 219
rect 2400 -2 2706 41
rect 2808 -62 3008 6
rect 2364 -77 3008 -62
rect 2364 -226 2379 -77
rect 2543 -194 3008 -77
rect 2543 -226 2561 -194
rect 2364 -243 2561 -226
rect 1869 -325 2420 -317
rect 1869 -406 1883 -325
rect 2058 -329 2420 -325
rect 2058 -406 2421 -329
rect 1869 -414 2421 -406
rect 1722 -693 1774 -681
rect 1722 -879 1774 -867
rect 1942 -693 1994 -681
rect 1942 -879 1994 -867
rect 1813 -998 1826 -946
rect 1900 -998 1913 -946
rect 1813 -999 1913 -998
rect 589 -1184 789 -1168
rect 589 -1352 604 -1184
rect 773 -1352 789 -1184
rect 2284 -1304 2421 -414
rect 2595 -484 2608 -425
rect 2751 -484 2767 -425
rect 2824 -540 2876 -528
rect 589 -1568 789 -1352
rect 1072 -1490 1087 -1438
rect 1201 -1490 1214 -1438
rect 877 -2015 1021 -1541
rect 1243 -1571 1297 -1559
rect 1295 -1915 1297 -1571
rect 1243 -1927 1297 -1915
rect 1401 -2015 1625 -1320
rect 1825 -1474 1837 -1422
rect 1951 -1474 1963 -1422
rect 1743 -1543 1795 -1531
rect 1993 -1543 2045 -1531
rect 1993 -1850 2045 -1837
rect 1743 -1930 1795 -1917
rect 2171 -2015 2421 -1304
rect 2514 -580 2566 -568
rect 2514 -1926 2566 -1914
rect 2824 -1926 2876 -1914
rect 607 -2315 3034 -2015
<< via1 >>
rect 1072 -860 1124 288
rect 958 -996 1032 -944
rect 1727 223 1779 297
rect 2237 223 2289 297
rect 1853 111 2154 167
rect 2625 41 2696 219
rect 2379 -226 2543 -77
rect 1883 -406 2058 -325
rect 1722 -867 1774 -693
rect 1942 -867 1994 -693
rect 1826 -998 1900 -946
rect 604 -1352 773 -1184
rect 2608 -484 2751 -425
rect 1087 -1490 1201 -1438
rect 1243 -1915 1295 -1571
rect 1837 -1474 1951 -1422
rect 1743 -1917 1795 -1543
rect 1993 -1837 2045 -1543
rect 2514 -1914 2566 -580
rect 2824 -1914 2876 -540
<< metal2 >>
rect 2242 313 2359 333
rect 1070 303 1126 304
rect 1725 303 1781 313
rect 1070 297 1781 303
rect 1070 288 1727 297
rect 1070 -860 1072 288
rect 1124 224 1727 288
rect 1124 -707 1126 224
rect 1725 223 1727 224
rect 1779 223 1781 297
rect 1725 207 1781 223
rect 2235 297 2359 313
rect 2235 223 2237 297
rect 2289 223 2359 297
rect 2235 207 2359 223
rect 2242 190 2359 207
rect 2622 219 2698 236
rect 1841 167 2166 170
rect 1841 111 1853 167
rect 2154 111 2166 167
rect 1841 109 2166 111
rect 1847 -175 1921 109
rect 2242 52 2318 190
rect 1719 -249 1921 -175
rect 1992 -24 2318 52
rect 2622 41 2625 219
rect 2696 41 2698 219
rect 2622 33 2698 41
rect 1719 -465 1793 -249
rect 1992 -322 2068 -24
rect 2364 -77 2561 -62
rect 2364 -97 2379 -77
rect 2128 -226 2379 -97
rect 2543 -226 2561 -77
rect 1869 -325 2070 -322
rect 1869 -406 1883 -325
rect 2058 -406 2070 -325
rect 1869 -408 2070 -406
rect 2128 -422 2257 -226
rect 2364 -243 2561 -226
rect 2622 -239 2696 33
rect 2622 -317 2889 -239
rect 2128 -425 2764 -422
rect 2128 -465 2608 -425
rect 1719 -484 2608 -465
rect 2751 -484 2764 -425
rect 1719 -486 2764 -484
rect 1719 -539 2257 -486
rect 1720 -693 1776 -680
rect 1720 -707 1722 -693
rect 1124 -855 1722 -707
rect 1124 -860 1126 -855
rect 1070 -876 1126 -860
rect 1720 -867 1722 -855
rect 1774 -867 1776 -693
rect 1720 -880 1776 -867
rect 1940 -687 1996 -680
rect 2128 -687 2257 -539
rect 2822 -540 2889 -317
rect 1940 -693 2257 -687
rect 1940 -867 1942 -693
rect 1994 -853 2257 -693
rect 1994 -867 1996 -853
rect 1940 -880 1996 -867
rect 946 -944 1044 -942
rect 946 -996 958 -944
rect 1032 -996 1044 -944
rect 946 -998 1044 -996
rect 1813 -946 1913 -944
rect 1813 -998 1826 -946
rect 1900 -998 1913 -946
rect 589 -1184 789 -1168
rect 589 -1352 604 -1184
rect 773 -1236 789 -1184
rect 961 -1236 1026 -998
rect 1813 -1000 1913 -998
rect 1832 -1236 1907 -1000
rect 773 -1305 1907 -1236
rect 773 -1352 789 -1305
rect 589 -1368 789 -1352
rect 961 -1421 1026 -1305
rect 1832 -1420 1907 -1305
rect 961 -1438 1215 -1421
rect 961 -1486 1087 -1438
rect 1072 -1490 1087 -1486
rect 1201 -1486 1215 -1438
rect 1825 -1422 1963 -1420
rect 1825 -1474 1837 -1422
rect 1951 -1474 1963 -1422
rect 1825 -1476 1963 -1474
rect 1201 -1490 1214 -1486
rect 1072 -1492 1214 -1490
rect 1741 -1543 1797 -1527
rect 1241 -1571 1297 -1555
rect 1241 -1915 1243 -1571
rect 1295 -1634 1297 -1571
rect 1741 -1634 1743 -1543
rect 1295 -1846 1743 -1634
rect 1295 -1915 1297 -1846
rect 1241 -1931 1297 -1915
rect 1741 -1917 1743 -1846
rect 1795 -1912 1797 -1543
rect 1991 -1543 2047 -1527
rect 1991 -1837 1993 -1543
rect 2045 -1557 2047 -1543
rect 2128 -1557 2257 -853
rect 2045 -1805 2257 -1557
rect 2512 -580 2568 -564
rect 2045 -1837 2047 -1805
rect 1991 -1853 2047 -1837
rect 2512 -1912 2514 -580
rect 1795 -1914 2514 -1912
rect 2566 -1914 2568 -580
rect 1795 -1917 2568 -1914
rect 1741 -1985 2568 -1917
rect 2822 -1914 2824 -540
rect 2876 -1914 2889 -540
rect 2822 -1926 2889 -1914
rect 2822 -1930 2878 -1926
use nmos_6p0_L3YBEV  X6 primitives
timestamp 1655307388
transform 1 0 2695 0 1 -1203
box -364 -932 364 932
use pmos_6p0_9YEQN4  XM1 primitives
timestamp 1655307388
transform 1 0 985 0 1 -325
box -378 -886 368 886
use nmos_6p0_BJPB5U  XM3 primitives
timestamp 1655307388
transform 1 0 1144 0 1 -1704
box -334 -432 334 432
use pmos_6p0_9859UL  XM5 primitives
timestamp 1655307388
transform 1 0 2008 0 1 226
box -518 -336 518 336
use nmos_6p0_BJPB5U  nmos_6p0_BJPB5U_0
timestamp 1655307388
transform 1 0 1894 0 1 -1706
box -334 -432 334 432
use pmos_6p0_UXEQNM  pmos_6p0_UXEQNM_0 primitives
timestamp 1655307388
transform 1 0 1863 0 1 -804
box -378 -386 368 386
<< labels >>
flabel metal1 577 445 777 645 0 FreeSans 1280 0 0 0 VDD
port 0 nsew
flabel metal1 639 -2288 839 -2088 0 FreeSans 1280 0 0 0 VSS
port 1 nsew
flabel metal1 2808 -194 3008 6 0 FreeSans 1280 0 0 0 Vout
port 3 nsew
flabel metal1 589 -1568 789 -1368 0 FreeSans 1280 0 0 0 Vin
port 2 nsew
<< end >>
