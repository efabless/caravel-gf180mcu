magic
tech gf180mcuC
magscale 1 10
timestamp 1670447232
<< fillblock >>
rect 0 4545 18699 8998
rect 0 0 8380 4545
use font_2D  font_2D_0 alpha
timestamp 1654634570
transform 1 0 5197 0 1 4980
box 0 648 864 864
use font_44  font_4A_0 alpha
timestamp 1654634570
transform 1 0 271 0 1 324
box 0 0 648 1512
use font_4B  font_4B_0 alpha
timestamp 1654634570
transform 1 0 6334 0 1 2739
box 0 0 648 1512
use font_6C  font_6C_0 alpha
timestamp 1654634570
transform 1 0 5567 0 1 7107
box 0 0 216 1512
use font_6C  font_6C_1
timestamp 1654634570
transform 1 0 3907 0 1 4990
box 0 0 216 1512
use font_6C  font_6C_2
timestamp 1654634570
transform 1 0 7120 0 1 4975
box 0 0 216 1512
use font_6C  font_6C_3
timestamp 1654634570
transform 1 0 10152 0 1 4965
box 0 0 216 1512
use font_6C  font_6C_4
timestamp 1654634570
transform 1 0 14929 0 1 7113
box 0 0 216 1512
use font_6E  font_6E_0 alpha
timestamp 1654634570
transform 1 0 2957 0 1 2748
box 0 0 648 1080
use font_43  font_6E_1
timestamp 1654634570
transform 1 0 1993 0 1 315
box 0 0 648 1080
use font_6E  font_6E_2
timestamp 1654634570
transform 1 0 13605 0 1 4983
box 0 0 648 1080
use font_6F  font_6F_0 alpha
timestamp 1654634570
transform 1 0 1308 0 1 5018
box 0 0 648 1080
use font_6F  font_6F_1
timestamp 1654634570
transform 1 0 2159 0 1 5008
box 0 0 648 1080
use font_6F  font_6F_2
timestamp 1654634570
transform 1 0 374 0 1 2776
box 0 0 648 1080
use font_6F  font_6F_3
timestamp 1654634570
transform 1 0 7560 0 1 4965
box 0 0 648 1080
use font_6F  font_6F_4
timestamp 1654634570
transform 1 0 11902 0 1 4992
box 0 0 648 1080
use font_28  font_28_0 alpha
timestamp 1654634570
transform 1 0 8569 0 1 7131
box 0 0 432 1512
use font_29  font_29_0 alpha
timestamp 1654634570
transform 1 0 10069 0 1 7113
box 0 0 432 1512
use font_30  font_30_0 alpha
timestamp 1654634570
transform 1 0 5352 0 1 332
box 0 0 648 1512
use font_32  font_32_0 alpha
timestamp 1654634570
transform 1 0 4482 0 1 323
box 0 0 648 1512
use font_32  font_32_1
timestamp 1654634570
transform 1 0 6232 0 1 324
box 0 0 648 1512
use font_32  font_32_2
timestamp 1654634570
transform 1 0 7120 0 1 332
box 0 0 648 1512
use font_43  font_43_0 alpha
timestamp 1654634570
transform 1 0 383 0 1 7116
box 0 0 648 1512
use font_44  font_44_0 alpha
timestamp 1654634570
transform 1 0 5474 0 1 2739
box 0 0 648 1512
use font_45  font_45_0 alpha
timestamp 1654634570
transform 1 0 11459 0 1 7113
box 0 0 648 1512
use font_46  font_46_0 alpha
timestamp 1654634570
transform 1 0 7336 0 1 7125
box 0 0 648 1512
use font_46  font_46_1
timestamp 1654634570
transform 1 0 11050 0 1 4956
box 0 0 648 1512
use font_47  font_47_0 alpha
timestamp 1654634570
transform 1 0 6456 0 1 7125
box 0 0 648 1512
use font_47  font_47_1
timestamp 1654634570
transform 1 0 468 0 1 5001
box 0 0 648 1512
use font_47  font_47_2
timestamp 1654634570
transform 1 0 6260 0 1 5001
box 0 0 648 1512
use font_50  font_50_0 alpha
timestamp 1654634570
transform 1 0 4613 0 1 2757
box 0 0 648 1512
use font_61  font_61_0 alpha
timestamp 1654634570
transform 1 0 1235 0 1 7107
box 0 0 648 1080
use font_61  font_61_1
timestamp 1654634570
transform 1 0 2966 0 1 7107
box 0 0 648 1080
use font_61  font_61_2
timestamp 1654634570
transform 1 0 9282 0 1 4984
box 0 0 648 1080
use font_61  font_61_3
timestamp 1654634570
transform 1 0 13189 0 1 7103
box 0 0 648 1080
use font_62  font_62_0 alpha
timestamp 1654634570
transform 1 0 8421 0 1 4984
box 0 0 648 1512
use font_62  font_62_1
timestamp 1654634570
transform 1 0 14059 0 1 7113
box 0 0 648 1512
use font_63  font_63_0 alpha
timestamp 1654634570
transform 1 0 9209 0 1 7301
box 0 0 648 1080
use font_64  font_64_0 alpha
timestamp 1654634570
transform 1 0 14484 0 1 5001
box 0 0 648 1512
use font_65  font_65_0 alpha
timestamp 1654634570
transform 1 0 4706 0 1 7125
box 0 0 648 1080
use font_65  font_65_1
timestamp 1654634570
transform 1 0 4347 0 1 4990
box 0 0 648 1080
use font_65  font_65_2
timestamp 1654634570
transform 1 0 16861 0 1 4992
box 0 0 648 1080
use font_65  font_65_3
timestamp 1654634570
transform 1 0 2105 0 1 2767
box 0 0 648 1080
use font_65  font_65_5
timestamp 1654634570
transform 1 0 15359 0 1 7113
box 0 0 648 1080
use font_66  font_66_0 alpha
timestamp 1654634570
transform 1 0 12319 0 1 7113
box 0 0 648 1512
use font_67  font_67_0 alpha
timestamp 1654634570
transform 1 0 3038 0 1 4999
box 0 -432 648 1080
use font_69  font_69_0 alpha
timestamp 1654634570
transform 1 0 16206 0 1 5001
box 0 0 432 1512
use font_70  font_70_0 alpha
timestamp 1654634570
transform 1 0 1235 0 1 2785
box 0 -432 648 1080
use font_72  font_72_0 alpha
timestamp 1654634570
transform 1 0 2096 0 1 7107
box 0 0 648 1080
use font_72  font_72_1
timestamp 1654634570
transform 1 0 15345 0 1 4992
box 0 0 648 1080
use font_73  font_73_0 alpha
timestamp 1654634570
transform 1 0 17731 0 1 5001
box 0 0 648 1080
use font_73  font_73_1
timestamp 1654634570
transform 1 0 16229 0 1 7121
box 0 0 648 1080
use font_73  font_73_2
timestamp 1654634570
transform 1 0 17089 0 1 7121
box 0 0 648 1080
use font_45  font_45_1 alpha
timestamp 1654634570
transform 1 0 1132 0 1 315
box 0 0 648 1080
use font_75  font_75_0
timestamp 1654634570
transform 1 0 12763 0 1 5001
box 0 0 648 1080
use font_76  font_76_0 alpha
timestamp 1654634570
transform 1 0 3874 0 1 7107
box 0 0 648 1080
<< end >>
