magic
tech gf180mcuC
magscale 1 5
timestamp 1670147979
<< obsm1 >>
rect 112 754 8424 5585
<< metal2 >>
rect 280 6100 336 6500
rect 504 6100 560 6500
rect 728 6100 784 6500
rect 952 6100 1008 6500
rect 1176 6100 1232 6500
rect 1400 6100 1456 6500
rect 1624 6100 1680 6500
rect 1848 6100 1904 6500
rect 2072 6100 2128 6500
rect 2296 6100 2352 6500
rect 2520 6100 2576 6500
rect 2744 6100 2800 6500
rect 2968 6100 3024 6500
rect 3192 6100 3248 6500
rect 3416 6100 3472 6500
rect 3640 6100 3696 6500
rect 3864 6100 3920 6500
rect 4088 6100 4144 6500
rect 4312 6100 4368 6500
rect 4536 6100 4592 6500
rect 4760 6100 4816 6500
rect 4984 6100 5040 6500
rect 5208 6100 5264 6500
rect 5432 6100 5488 6500
rect 5656 6100 5712 6500
rect 5880 6100 5936 6500
rect 6104 6100 6160 6500
rect 6328 6100 6384 6500
rect 6552 6100 6608 6500
rect 6776 6100 6832 6500
rect 7000 6100 7056 6500
rect 7224 6100 7280 6500
rect 7448 6100 7504 6500
rect 7672 6100 7728 6500
rect 7896 6100 7952 6500
rect 8120 6100 8176 6500
rect 280 0 336 400
rect 504 0 560 400
rect 728 0 784 400
rect 952 0 1008 400
rect 1176 0 1232 400
rect 1400 0 1456 400
rect 1624 0 1680 400
rect 1848 0 1904 400
rect 2072 0 2128 400
rect 2296 0 2352 400
rect 2520 0 2576 400
rect 2744 0 2800 400
rect 2968 0 3024 400
rect 3192 0 3248 400
rect 3416 0 3472 400
rect 3640 0 3696 400
rect 3864 0 3920 400
rect 4088 0 4144 400
rect 4312 0 4368 400
rect 4536 0 4592 400
rect 4760 0 4816 400
rect 4984 0 5040 400
rect 5208 0 5264 400
rect 5432 0 5488 400
rect 5656 0 5712 400
rect 5880 0 5936 400
rect 6104 0 6160 400
rect 6328 0 6384 400
rect 6552 0 6608 400
rect 6776 0 6832 400
rect 7000 0 7056 400
rect 7224 0 7280 400
rect 7448 0 7504 400
rect 7672 0 7728 400
rect 7896 0 7952 400
rect 8120 0 8176 400
<< obsm2 >>
rect 366 6070 474 6100
rect 590 6070 698 6100
rect 814 6070 922 6100
rect 1038 6070 1146 6100
rect 1262 6070 1370 6100
rect 1486 6070 1594 6100
rect 1710 6070 1818 6100
rect 1934 6070 2042 6100
rect 2158 6070 2266 6100
rect 2382 6070 2490 6100
rect 2606 6070 2714 6100
rect 2830 6070 2938 6100
rect 3054 6070 3162 6100
rect 3278 6070 3386 6100
rect 3502 6070 3610 6100
rect 3726 6070 3834 6100
rect 3950 6070 4058 6100
rect 4174 6070 4282 6100
rect 4398 6070 4506 6100
rect 4622 6070 4730 6100
rect 4846 6070 4954 6100
rect 5070 6070 5178 6100
rect 5294 6070 5402 6100
rect 5518 6070 5626 6100
rect 5742 6070 5850 6100
rect 5966 6070 6074 6100
rect 6190 6070 6298 6100
rect 6414 6070 6522 6100
rect 6638 6070 6746 6100
rect 6862 6070 6970 6100
rect 7086 6070 7194 6100
rect 7310 6070 7418 6100
rect 7534 6070 7642 6100
rect 7758 6070 7866 6100
rect 7982 6070 8090 6100
rect 8206 6070 8410 6100
rect 294 430 8410 6070
rect 366 400 474 430
rect 590 400 698 430
rect 814 400 922 430
rect 1038 400 1146 430
rect 1262 400 1370 430
rect 1486 400 1594 430
rect 1710 400 1818 430
rect 1934 400 2042 430
rect 2158 400 2266 430
rect 2382 400 2490 430
rect 2606 400 2714 430
rect 2830 400 2938 430
rect 3054 400 3162 430
rect 3278 400 3386 430
rect 3502 400 3610 430
rect 3726 400 3834 430
rect 3950 400 4058 430
rect 4174 400 4282 430
rect 4398 400 4506 430
rect 4622 400 4730 430
rect 4846 400 4954 430
rect 5070 400 5178 430
rect 5294 400 5402 430
rect 5518 400 5626 430
rect 5742 400 5850 430
rect 5966 400 6074 430
rect 6190 400 6298 430
rect 6414 400 6522 430
rect 6638 400 6746 430
rect 6862 400 6970 430
rect 7086 400 7194 430
rect 7310 400 7418 430
rect 7534 400 7642 430
rect 7758 400 7866 430
rect 7982 400 8090 430
rect 8206 400 8410 430
<< metal3 >>
rect 0 5320 400 5376
rect 8100 5320 8500 5376
rect 0 3192 400 3248
rect 8100 3192 8500 3248
rect 0 1064 400 1120
rect 8100 1064 8500 1120
<< obsm3 >>
rect 289 5406 8415 5502
rect 430 5290 8070 5406
rect 289 3278 8415 5290
rect 430 3162 8070 3278
rect 289 1150 8415 3162
rect 430 1034 8070 1150
rect 289 770 8415 1034
<< metal4 >>
rect 1061 754 1221 5518
rect 2090 754 2250 5518
rect 3119 754 3279 5518
rect 4148 754 4308 5518
rect 5177 754 5337 5518
rect 6206 754 6366 5518
rect 7235 754 7395 5518
rect 8264 754 8424 5518
<< labels >>
rlabel metal4 s 1061 754 1221 5518 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 3119 754 3279 5518 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 5177 754 5337 5518 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 7235 754 7395 5518 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 2090 754 2250 5518 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 4148 754 4308 5518 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 6206 754 6366 5518 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 8264 754 8424 5518 6 VSS
port 2 nsew ground bidirectional
rlabel metal2 s 280 0 336 400 6 mgmt_gpio_in[0]
port 3 nsew signal input
rlabel metal2 s 2520 0 2576 400 6 mgmt_gpio_in[10]
port 4 nsew signal input
rlabel metal2 s 2744 0 2800 400 6 mgmt_gpio_in[11]
port 5 nsew signal input
rlabel metal2 s 2968 0 3024 400 6 mgmt_gpio_in[12]
port 6 nsew signal input
rlabel metal2 s 3192 0 3248 400 6 mgmt_gpio_in[13]
port 7 nsew signal input
rlabel metal2 s 3416 0 3472 400 6 mgmt_gpio_in[14]
port 8 nsew signal input
rlabel metal2 s 3640 0 3696 400 6 mgmt_gpio_in[15]
port 9 nsew signal input
rlabel metal2 s 3864 0 3920 400 6 mgmt_gpio_in[16]
port 10 nsew signal input
rlabel metal2 s 4088 0 4144 400 6 mgmt_gpio_in[17]
port 11 nsew signal input
rlabel metal2 s 504 0 560 400 6 mgmt_gpio_in[1]
port 12 nsew signal input
rlabel metal2 s 728 0 784 400 6 mgmt_gpio_in[2]
port 13 nsew signal input
rlabel metal2 s 952 0 1008 400 6 mgmt_gpio_in[3]
port 14 nsew signal input
rlabel metal2 s 1176 0 1232 400 6 mgmt_gpio_in[4]
port 15 nsew signal input
rlabel metal2 s 1400 0 1456 400 6 mgmt_gpio_in[5]
port 16 nsew signal input
rlabel metal2 s 1624 0 1680 400 6 mgmt_gpio_in[6]
port 17 nsew signal input
rlabel metal2 s 1848 0 1904 400 6 mgmt_gpio_in[7]
port 18 nsew signal input
rlabel metal2 s 2072 0 2128 400 6 mgmt_gpio_in[8]
port 19 nsew signal input
rlabel metal2 s 2296 0 2352 400 6 mgmt_gpio_in[9]
port 20 nsew signal input
rlabel metal2 s 280 6100 336 6500 6 mgmt_gpio_in_buf[0]
port 21 nsew signal output
rlabel metal2 s 2520 6100 2576 6500 6 mgmt_gpio_in_buf[10]
port 22 nsew signal output
rlabel metal2 s 2744 6100 2800 6500 6 mgmt_gpio_in_buf[11]
port 23 nsew signal output
rlabel metal2 s 2968 6100 3024 6500 6 mgmt_gpio_in_buf[12]
port 24 nsew signal output
rlabel metal2 s 3192 6100 3248 6500 6 mgmt_gpio_in_buf[13]
port 25 nsew signal output
rlabel metal2 s 3416 6100 3472 6500 6 mgmt_gpio_in_buf[14]
port 26 nsew signal output
rlabel metal2 s 3640 6100 3696 6500 6 mgmt_gpio_in_buf[15]
port 27 nsew signal output
rlabel metal2 s 3864 6100 3920 6500 6 mgmt_gpio_in_buf[16]
port 28 nsew signal output
rlabel metal2 s 4088 6100 4144 6500 6 mgmt_gpio_in_buf[17]
port 29 nsew signal output
rlabel metal2 s 504 6100 560 6500 6 mgmt_gpio_in_buf[1]
port 30 nsew signal output
rlabel metal2 s 728 6100 784 6500 6 mgmt_gpio_in_buf[2]
port 31 nsew signal output
rlabel metal2 s 952 6100 1008 6500 6 mgmt_gpio_in_buf[3]
port 32 nsew signal output
rlabel metal2 s 1176 6100 1232 6500 6 mgmt_gpio_in_buf[4]
port 33 nsew signal output
rlabel metal2 s 1400 6100 1456 6500 6 mgmt_gpio_in_buf[5]
port 34 nsew signal output
rlabel metal2 s 1624 6100 1680 6500 6 mgmt_gpio_in_buf[6]
port 35 nsew signal output
rlabel metal2 s 1848 6100 1904 6500 6 mgmt_gpio_in_buf[7]
port 36 nsew signal output
rlabel metal2 s 2072 6100 2128 6500 6 mgmt_gpio_in_buf[8]
port 37 nsew signal output
rlabel metal2 s 2296 6100 2352 6500 6 mgmt_gpio_in_buf[9]
port 38 nsew signal output
rlabel metal3 s 0 1064 400 1120 6 mgmt_gpio_oeb[0]
port 39 nsew signal input
rlabel metal3 s 0 3192 400 3248 6 mgmt_gpio_oeb[1]
port 40 nsew signal input
rlabel metal3 s 0 5320 400 5376 6 mgmt_gpio_oeb[2]
port 41 nsew signal input
rlabel metal3 s 8100 1064 8500 1120 6 mgmt_gpio_oeb_buf[0]
port 42 nsew signal output
rlabel metal3 s 8100 3192 8500 3248 6 mgmt_gpio_oeb_buf[1]
port 43 nsew signal output
rlabel metal3 s 8100 5320 8500 5376 6 mgmt_gpio_oeb_buf[2]
port 44 nsew signal output
rlabel metal2 s 4312 6100 4368 6500 6 mgmt_gpio_out[0]
port 45 nsew signal input
rlabel metal2 s 6552 6100 6608 6500 6 mgmt_gpio_out[10]
port 46 nsew signal input
rlabel metal2 s 6776 6100 6832 6500 6 mgmt_gpio_out[11]
port 47 nsew signal input
rlabel metal2 s 7000 6100 7056 6500 6 mgmt_gpio_out[12]
port 48 nsew signal input
rlabel metal2 s 7224 6100 7280 6500 6 mgmt_gpio_out[13]
port 49 nsew signal input
rlabel metal2 s 7448 6100 7504 6500 6 mgmt_gpio_out[14]
port 50 nsew signal input
rlabel metal2 s 7672 6100 7728 6500 6 mgmt_gpio_out[15]
port 51 nsew signal input
rlabel metal2 s 7896 6100 7952 6500 6 mgmt_gpio_out[16]
port 52 nsew signal input
rlabel metal2 s 8120 6100 8176 6500 6 mgmt_gpio_out[17]
port 53 nsew signal input
rlabel metal2 s 4536 6100 4592 6500 6 mgmt_gpio_out[1]
port 54 nsew signal input
rlabel metal2 s 4760 6100 4816 6500 6 mgmt_gpio_out[2]
port 55 nsew signal input
rlabel metal2 s 4984 6100 5040 6500 6 mgmt_gpio_out[3]
port 56 nsew signal input
rlabel metal2 s 5208 6100 5264 6500 6 mgmt_gpio_out[4]
port 57 nsew signal input
rlabel metal2 s 5432 6100 5488 6500 6 mgmt_gpio_out[5]
port 58 nsew signal input
rlabel metal2 s 5656 6100 5712 6500 6 mgmt_gpio_out[6]
port 59 nsew signal input
rlabel metal2 s 5880 6100 5936 6500 6 mgmt_gpio_out[7]
port 60 nsew signal input
rlabel metal2 s 6104 6100 6160 6500 6 mgmt_gpio_out[8]
port 61 nsew signal input
rlabel metal2 s 6328 6100 6384 6500 6 mgmt_gpio_out[9]
port 62 nsew signal input
rlabel metal2 s 4312 0 4368 400 6 mgmt_gpio_out_buf[0]
port 63 nsew signal output
rlabel metal2 s 6552 0 6608 400 6 mgmt_gpio_out_buf[10]
port 64 nsew signal output
rlabel metal2 s 6776 0 6832 400 6 mgmt_gpio_out_buf[11]
port 65 nsew signal output
rlabel metal2 s 7000 0 7056 400 6 mgmt_gpio_out_buf[12]
port 66 nsew signal output
rlabel metal2 s 7224 0 7280 400 6 mgmt_gpio_out_buf[13]
port 67 nsew signal output
rlabel metal2 s 7448 0 7504 400 6 mgmt_gpio_out_buf[14]
port 68 nsew signal output
rlabel metal2 s 7672 0 7728 400 6 mgmt_gpio_out_buf[15]
port 69 nsew signal output
rlabel metal2 s 7896 0 7952 400 6 mgmt_gpio_out_buf[16]
port 70 nsew signal output
rlabel metal2 s 8120 0 8176 400 6 mgmt_gpio_out_buf[17]
port 71 nsew signal output
rlabel metal2 s 4536 0 4592 400 6 mgmt_gpio_out_buf[1]
port 72 nsew signal output
rlabel metal2 s 4760 0 4816 400 6 mgmt_gpio_out_buf[2]
port 73 nsew signal output
rlabel metal2 s 4984 0 5040 400 6 mgmt_gpio_out_buf[3]
port 74 nsew signal output
rlabel metal2 s 5208 0 5264 400 6 mgmt_gpio_out_buf[4]
port 75 nsew signal output
rlabel metal2 s 5432 0 5488 400 6 mgmt_gpio_out_buf[5]
port 76 nsew signal output
rlabel metal2 s 5656 0 5712 400 6 mgmt_gpio_out_buf[6]
port 77 nsew signal output
rlabel metal2 s 5880 0 5936 400 6 mgmt_gpio_out_buf[7]
port 78 nsew signal output
rlabel metal2 s 6104 0 6160 400 6 mgmt_gpio_out_buf[8]
port 79 nsew signal output
rlabel metal2 s 6328 0 6384 400 6 mgmt_gpio_out_buf[9]
port 80 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 8500 6500
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 165610
string GDS_FILE ../gds/mprj_io_buffer.gds
string GDS_START 36318
<< end >>

