magic
tech gf180mcuD
magscale 1 10
timestamp 1655307388
<< pwell >>
rect -364 -932 364 932
<< mvnmos >>
rect -100 -724 100 676
<< mvndiff >>
rect -188 663 -100 676
rect -188 -711 -175 663
rect -129 -711 -100 663
rect -188 -724 -100 -711
rect 100 663 188 676
rect 100 -711 129 663
rect 175 -711 188 663
rect 100 -724 188 -711
<< mvndiffc >>
rect -175 -711 -129 663
rect 129 -711 175 663
<< mvpsubdiff >>
rect -332 828 332 900
rect -332 784 -260 828
rect -332 -784 -319 784
rect -273 -784 -260 784
rect 260 784 332 828
rect -332 -828 -260 -784
rect 260 -784 273 784
rect 319 -784 332 784
rect 260 -828 332 -784
rect -332 -841 332 -828
rect -332 -887 -216 -841
rect 216 -887 332 -841
rect -332 -900 332 -887
<< mvpsubdiffcont >>
rect -319 -784 -273 784
rect 273 -784 319 784
rect -216 -887 216 -841
<< polysilicon >>
rect -100 755 100 768
rect -100 709 -87 755
rect 87 709 100 755
rect -100 676 100 709
rect -100 -768 100 -724
<< polycontact >>
rect -87 709 87 755
<< metal1 >>
rect -319 841 319 887
rect -319 784 -273 841
rect 273 784 319 841
rect -98 709 -87 755
rect 87 709 98 755
rect -175 663 -129 674
rect -175 -722 -129 -711
rect 129 663 175 674
rect 129 -722 175 -711
rect -319 -841 -273 -784
rect 273 -841 319 -784
rect -319 -887 -216 -841
rect 216 -887 319 -841
<< properties >>
string FIXED_BBOX -296 -864 296 864
string gencell nmos_6p0
string library gf180mcu
string parameters w 7.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.6 wmin 0.3 full_metal 1 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
