magic
tech micross
timestamp 1679504633
<< rdl >>
tri -3494 13040 -1177 13449 se
rect -1177 13040 1177 13449
tri 1177 13040 3494 13449 sw
tri -5705 12235 -3494 13040 se
rect -3494 12235 3494 13040
tri 3494 12235 5705 13040 sw
tri -7743 11059 -5705 12235 se
rect -5705 11059 5705 12235
tri 5705 11059 7743 12235 sw
tri -9546 9546 -7743 11059 se
rect -7743 9546 7743 11059
tri 7743 9546 9546 11059 sw
tri -11059 7743 -9546 9546 se
rect -9546 7743 9546 9546
tri 9546 7743 11349 9546 sw
tri -12235 5705 -11059 7743 se
rect -11059 5705 11349 7743
tri 11349 5705 13387 7743 sw
tri -13040 3494 -12235 5705 se
rect -12235 3494 13387 5705
tri 13387 3494 15598 5705 sw
tri -13449 1177 -13040 3494 se
rect -13040 1177 15598 3494
tri 15598 1177 17915 3494 sw
rect -13449 0 17915 1177
tri 17915 0 19092 1177 sw
rect -13449 -1177 9546 0
tri -13449 -3494 -13040 -1177 ne
rect -13040 -3494 9546 -1177
tri -13040 -5705 -12235 -3494 ne
rect -12235 -5705 9546 -3494
tri -12235 -7743 -11059 -5705 ne
rect -11059 -7743 9546 -5705
tri -11059 -9546 -9546 -7743 ne
rect -9546 -9546 9546 -7743
tri 9546 -9546 19092 0 nw
tri -9546 -11059 -7743 -9546 ne
rect -7743 -11059 7743 -9546
tri 7743 -11059 9546 -9546 nw
tri -7743 -12235 -5705 -11059 ne
rect -5705 -12235 5705 -11059
tri 5705 -12235 7743 -11059 nw
tri -5705 -13040 -3494 -12235 ne
rect -3494 -13040 3494 -12235
tri 3494 -13040 5705 -12235 nw
tri -3494 -13449 -1177 -13040 ne
rect -1177 -13449 1177 -13040
tri 1177 -13449 3494 -13040 nw
<< pi2 >>
tri -1910 10833 0 11000 se
tri 0 10833 1910 11000 sw
tri -3762 10337 -1910 10833 se
rect -1910 10337 1910 10833
tri 1910 10337 3762 10833 sw
tri -5500 9526 -3762 10337 se
rect -3762 9526 3762 10337
tri 3762 9526 5500 10337 sw
tri -7071 8426 -5500 9526 se
rect -5500 8426 5500 9526
tri 5500 8426 7071 9526 sw
tri -8426 7071 -7071 8426 se
rect -7071 7071 7071 8426
tri 7071 7071 8426 8426 sw
tri -9526 5500 -8426 7071 se
rect -8426 5500 8426 7071
tri 8426 5500 9526 7071 sw
tri -10337 3762 -9526 5500 se
rect -9526 3762 9526 5500
tri 9526 3762 10337 5500 sw
tri -10833 1910 -10337 3762 se
rect -10337 1910 10337 3762
tri 10337 1910 10833 3762 sw
tri -11000 0 -10833 1910 se
tri -11000 -1910 -10833 0 ne
rect -10833 -1910 10833 1910
tri 10833 0 11000 1910 sw
tri 10833 -1910 11000 0 nw
tri -10833 -3762 -10337 -1910 ne
rect -10337 -3762 10337 -1910
tri 10337 -3762 10833 -1910 nw
tri -10337 -5500 -9526 -3762 ne
rect -9526 -5500 9526 -3762
tri 9526 -5500 10337 -3762 nw
tri -9526 -7071 -8426 -5500 ne
rect -8426 -7071 8426 -5500
tri 8426 -7071 9526 -5500 nw
tri -8426 -8426 -7071 -7071 ne
rect -7071 -8426 7071 -7071
tri 7071 -8426 8426 -7071 nw
tri -7071 -9526 -5500 -8426 ne
rect -5500 -9526 5500 -8426
tri 5500 -9526 7071 -8426 nw
tri -5500 -10337 -3762 -9526 ne
rect -3762 -10337 3762 -9526
tri 3762 -10337 5500 -9526 nw
tri -3762 -10833 -1910 -10337 ne
rect -1910 -10833 1910 -10337
tri 1910 -10833 3762 -10337 nw
tri -1910 -11000 0 -10833 ne
tri 0 -11000 1910 -10833 nw
<< ubm >>
tri -2171 12310 0 12500 se
tri 0 12310 2171 12500 sw
tri -4275 11746 -2171 12310 se
rect -2171 11746 2171 12310
tri 2171 11746 4275 12310 sw
tri -6250 10825 -4275 11746 se
rect -4275 10825 4275 11746
tri 4275 10825 6250 11746 sw
tri -8035 9576 -6250 10825 se
rect -6250 9576 6250 10825
tri 6250 9576 8035 10825 sw
tri -9576 8035 -8035 9576 se
rect -8035 8035 8035 9576
tri 8035 8035 9576 9576 sw
tri -10825 6250 -9576 8035 se
rect -9576 6250 9576 8035
tri 9576 6250 10825 8035 sw
tri -11746 4275 -10825 6250 se
rect -10825 4275 10825 6250
tri 10825 4275 11746 6250 sw
tri -12310 2171 -11746 4275 se
rect -11746 2171 11746 4275
tri 11746 2171 12310 4275 sw
tri -12500 0 -12310 2171 se
tri -12500 -2171 -12310 0 ne
rect -12310 -2171 12310 2171
tri 12310 0 12500 2171 sw
tri 12310 -2171 12500 0 nw
tri -12310 -4275 -11746 -2171 ne
rect -11746 -4275 11746 -2171
tri 11746 -4275 12310 -2171 nw
tri -11746 -6250 -10825 -4275 ne
rect -10825 -6250 10825 -4275
tri 10825 -6250 11746 -4275 nw
tri -10825 -8035 -9576 -6250 ne
rect -9576 -8035 9576 -6250
tri 9576 -8035 10825 -6250 nw
tri -9576 -9576 -8035 -8035 ne
rect -8035 -9576 8035 -8035
tri 8035 -9576 9576 -8035 nw
tri -8035 -10825 -6250 -9576 ne
rect -6250 -10825 6250 -9576
tri 6250 -10825 8035 -9576 nw
tri -6250 -11746 -4275 -10825 ne
rect -4275 -11746 4275 -10825
tri 4275 -11746 6250 -10825 nw
tri -4275 -12310 -2171 -11746 ne
rect -2171 -12310 2171 -11746
tri 2171 -12310 4275 -11746 nw
tri -2171 -12500 0 -12310 ne
tri 0 -12500 2171 -12310 nw
<< properties >>
string FIXED_BBOX -13500 -13500 13500 13500
<< end >>
