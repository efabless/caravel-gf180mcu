magic
tech gf180mcuC
magscale 6 5
timestamp 1654634570
<< metal5 >>
rect 108 648 216 756
rect 0 540 216 648
rect 108 108 216 540
rect 0 0 324 108
<< properties >>
string FIXED_BBOX 0 0 432 756
<< end >>
