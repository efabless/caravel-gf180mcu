magic
tech gf180mcuD
magscale 1 10
timestamp 1670521662
<< metal5 >>
rect -3396 7367 3918 7615
rect -2505 1541 -2244 7367
rect -1286 -56 -1074 7233
rect 151 1510 412 7367
rect 1394 -56 1606 7243
rect 2835 1482 3096 7367
rect 4074 -56 4286 7244
rect -3458 -294 4286 -56
use mim_2p0fF_8KW78G  XC1 primitives
array 0 2 2680 0 2 2480
timestamp 1670521662
transform 1 0 -2294 0 1 1179
box -1220 -1120 1220 1120
<< labels >>
flabel metal5 s -3430 -269 -3230 -69 0 FreeSans 1280 0 0 0 VSS
port 1 nsew
flabel metal5 s -3367 7398 -3167 7598 0 FreeSans 1280 0 0 0 In
port 0 nsew
<< end >>
