VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_core
  CLASS BLOCK ;
  FOREIGN caravel_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 3170.000 BY 4360.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 14.080 17.440 24.080 4345.520 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 14.080 17.440 3155.520 27.440 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 14.080 4335.520 3155.520 4345.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3145.520 17.440 3155.520 4345.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 106.080 5.440 109.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 106.080 4282.880 109.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 186.080 5.440 189.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 186.080 4282.880 189.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 266.080 5.440 269.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 266.080 4282.880 269.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 346.080 5.440 349.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 346.080 4282.880 349.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 426.080 5.440 429.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 426.080 4282.880 429.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 506.080 5.440 509.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 506.080 4282.880 509.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 586.080 5.440 589.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 586.080 4282.880 589.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 666.080 5.440 669.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 666.080 4282.880 669.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 746.080 5.440 749.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 746.080 4282.880 749.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 826.080 5.440 829.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 826.080 4282.880 829.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 906.080 5.440 909.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 906.080 4282.880 909.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 986.080 5.440 989.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 986.080 4282.880 989.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1066.080 5.440 1069.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1066.080 4282.880 1069.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1146.080 5.440 1149.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1146.080 4282.880 1149.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1226.080 5.440 1229.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1226.080 4282.880 1229.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1306.080 5.440 1309.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1306.080 4282.880 1309.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1386.080 5.440 1389.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1386.080 4282.880 1389.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1466.080 5.440 1469.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1466.080 4282.880 1469.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 5.440 1549.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1546.080 4282.880 1549.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1626.080 5.440 1629.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1626.080 4282.880 1629.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1706.080 5.440 1709.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1706.080 4282.880 1709.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1786.080 5.440 1789.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1786.080 4282.880 1789.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1866.080 5.440 1869.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1866.080 4282.880 1869.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1946.080 5.440 1949.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1946.080 4282.880 1949.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2026.080 5.440 2029.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2026.080 4282.880 2029.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2106.080 5.440 2109.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2106.080 4282.880 2109.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2186.080 5.440 2189.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2186.080 4282.880 2189.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2266.080 5.440 2269.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2266.080 4282.880 2269.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2346.080 5.440 2349.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2346.080 4282.880 2349.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2426.080 5.440 2429.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2426.080 4282.880 2429.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2506.080 5.440 2509.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2506.080 4282.880 2509.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2586.080 5.440 2589.080 219.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2586.080 984.710 2589.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2586.080 4282.880 2589.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2666.080 5.440 2669.080 219.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2666.080 984.710 2669.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2666.080 4282.880 2669.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2746.080 5.440 2749.080 219.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2746.080 984.710 2749.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2746.080 4282.880 2749.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2826.080 5.440 2829.080 219.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2826.080 984.710 2829.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2826.080 4282.880 2829.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2906.080 5.440 2909.080 86.730 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2906.080 144.725 2909.080 219.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2906.080 984.710 2909.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2906.080 4282.880 2909.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2986.080 5.440 2989.080 219.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2986.080 984.710 2989.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2986.080 4282.880 2989.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3099.080 5.440 3102.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3126.620 5.440 3129.620 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 36.080 5.440 39.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.940 5.440 63.940 4357.520 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 56.590 3167.520 59.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 116.590 2896.355 119.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 176.590 3167.520 179.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 236.590 2549.760 239.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 296.590 2549.760 299.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 356.590 2549.760 359.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 416.590 2549.760 419.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 476.590 2549.760 479.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 536.590 2549.760 539.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 596.590 2549.760 599.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 656.590 2549.760 659.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 716.590 2549.760 719.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 776.590 2549.760 779.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 836.590 2549.760 839.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 896.590 601.540 899.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 956.590 601.540 959.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1016.590 3167.520 1019.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1076.590 1561.540 1079.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1136.590 3167.520 1139.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1196.590 3167.520 1199.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1256.590 3167.520 1259.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1316.590 93.140 1319.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1376.590 93.140 1379.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1436.590 93.140 1439.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1496.590 93.140 1499.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1556.590 93.140 1559.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1616.590 93.140 1619.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1676.590 93.140 1679.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1736.590 93.140 1739.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1796.590 93.140 1799.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1856.590 93.140 1859.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1916.590 93.140 1919.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1976.590 93.140 1979.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2036.590 93.140 2039.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2096.590 93.140 2099.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2156.590 93.140 2159.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2216.590 93.140 2219.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2276.590 93.140 2279.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2336.590 93.140 2339.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2396.590 93.140 2399.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2456.590 93.140 2459.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2516.590 93.140 2519.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2576.590 93.140 2579.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2636.590 93.140 2639.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2696.590 93.140 2699.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2756.590 93.140 2759.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2816.590 93.140 2819.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2876.590 93.140 2879.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2936.590 93.140 2939.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2996.590 93.140 2999.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3056.590 93.140 3059.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3116.590 93.140 3119.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3176.590 93.140 3179.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3236.590 93.140 3239.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3296.590 93.140 3299.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3356.590 93.140 3359.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3416.590 93.140 3419.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3476.590 93.140 3479.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3536.590 93.140 3539.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3596.590 93.140 3599.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3656.590 93.140 3659.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3716.590 93.140 3719.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3776.590 93.140 3779.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3836.590 93.140 3839.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3896.590 93.140 3899.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3956.590 93.140 3959.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4016.590 93.140 4019.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4076.590 93.140 4079.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4136.590 93.140 4139.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4196.590 93.140 4199.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4256.590 93.140 4259.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4316.590 3167.520 4319.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 672.460 896.590 1081.540 899.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 672.460 956.590 1081.540 959.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1152.460 896.590 2549.760 899.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1152.460 956.590 2549.760 959.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1632.460 1076.590 2121.040 1079.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2191.960 1076.590 3167.520 1079.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2966.995 116.590 3167.520 119.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 236.590 3167.520 239.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 296.590 3167.520 299.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 356.590 3167.520 359.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 416.590 3167.520 419.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 476.590 3167.520 479.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 536.590 3167.520 539.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 596.590 3167.520 599.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 656.590 3167.520 659.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 716.590 3167.520 719.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 776.590 3167.520 779.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 836.590 3167.520 839.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 896.590 3167.520 899.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 956.590 3167.520 959.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1316.590 3167.520 1319.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1376.590 3167.520 1379.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1436.590 3167.520 1439.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1496.590 3167.520 1499.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1556.590 3167.520 1559.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1616.590 3167.520 1619.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1676.590 3167.520 1679.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1736.590 3167.520 1739.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1796.590 3167.520 1799.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1856.590 3167.520 1859.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1916.590 3167.520 1919.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1976.590 3167.520 1979.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2036.590 3167.520 2039.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2096.590 3167.520 2099.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2156.590 3167.520 2159.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2216.590 3167.520 2219.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2276.590 3167.520 2279.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2336.590 3167.520 2339.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2396.590 3167.520 2399.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2456.590 3167.520 2459.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2516.590 3167.520 2519.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2576.590 3167.520 2579.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2636.590 3167.520 2639.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2696.590 3167.520 2699.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2756.590 3167.520 2759.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2816.590 3167.520 2819.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2876.590 3167.520 2879.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2936.590 3167.520 2939.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2996.590 3167.520 2999.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3056.590 3167.520 3059.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3116.590 3167.520 3119.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3176.590 3167.520 3179.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3236.590 3167.520 3239.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3296.590 3167.520 3299.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3356.590 3167.520 3359.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3416.590 3167.520 3419.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3476.590 3167.520 3479.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3536.590 3167.520 3539.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3596.590 3167.520 3599.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3656.590 3167.520 3659.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3716.590 3167.520 3719.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3776.590 3167.520 3779.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3836.590 3167.520 3839.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3896.590 3167.520 3899.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3956.590 3167.520 3959.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 4016.590 3167.520 4019.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 4076.590 3167.520 4079.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 4136.590 3167.520 4139.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 4196.590 3167.520 4199.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 4256.590 3167.520 4259.590 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2331.080 5.440 2334.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2331.080 4282.880 2334.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2880.580 5.440 2883.580 219.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2880.580 984.710 2883.580 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2880.580 4282.880 2883.580 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2163.080 5.440 2166.080 1031.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2163.080 1123.280 2166.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2163.080 4282.880 2166.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1916.380 5.440 1919.380 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1916.380 4282.880 1919.380 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1359.380 5.440 1362.380 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1359.380 4282.880 1362.380 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1116.480 5.440 1119.480 891.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1116.480 983.280 1119.480 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1116.480 4282.880 1119.480 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 864.780 5.440 867.780 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 864.780 4282.880 867.780 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 556.280 5.440 559.280 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 556.280 4282.880 559.280 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 306.580 5.440 309.580 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 306.580 4282.880 309.580 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 566.620 62.420 569.620 572.620 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1023.770 58.500 1025.270 576.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1480.730 58.500 1482.230 576.540 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 2.080 5.440 12.080 4357.520 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 5.440 3167.520 15.440 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4347.520 3167.520 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3157.520 5.440 3167.520 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 128.080 5.440 131.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 128.080 4282.880 131.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 208.080 5.440 211.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 208.080 4282.880 211.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 288.080 5.440 291.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 288.080 4282.880 291.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 368.080 5.440 371.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 368.080 4282.880 371.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 448.080 5.440 451.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 448.080 4282.880 451.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 528.080 5.440 531.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 528.080 4282.880 531.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 608.080 5.440 611.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 608.080 4282.880 611.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 688.080 5.440 691.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 688.080 4282.880 691.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 768.080 5.440 771.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 768.080 4282.880 771.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 848.080 5.440 851.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 848.080 4282.880 851.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 928.080 5.440 931.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 928.080 4282.880 931.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1008.080 5.440 1011.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1008.080 4282.880 1011.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1088.080 5.440 1091.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1088.080 4282.880 1091.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1168.080 5.440 1171.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1168.080 4282.880 1171.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1248.080 5.440 1251.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1248.080 4282.880 1251.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1328.080 5.440 1331.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1328.080 4282.880 1331.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1408.080 5.440 1411.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1408.080 4282.880 1411.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1488.080 5.440 1491.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1488.080 4282.880 1491.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1568.080 5.440 1571.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1568.080 4282.880 1571.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1648.080 5.440 1651.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1648.080 4282.880 1651.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1728.080 5.440 1731.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1728.080 4282.880 1731.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1808.080 5.440 1811.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1808.080 4282.880 1811.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1888.080 5.440 1891.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1888.080 4282.880 1891.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1968.080 5.440 1971.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1968.080 4282.880 1971.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2048.080 5.440 2051.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2048.080 4282.880 2051.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2128.080 5.440 2131.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2128.080 4282.880 2131.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2208.080 5.440 2211.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2208.080 4282.880 2211.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2288.080 5.440 2291.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2288.080 4282.880 2291.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2368.080 5.440 2371.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2368.080 4282.880 2371.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2448.080 5.440 2451.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2448.080 4282.880 2451.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2528.080 5.440 2531.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2528.080 4282.880 2531.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2608.080 5.440 2611.080 219.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2608.080 984.710 2611.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2608.080 4282.880 2611.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2688.080 5.440 2691.080 219.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2688.080 984.710 2691.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2688.080 4282.880 2691.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2768.080 5.440 2771.080 219.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2768.080 984.710 2771.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2768.080 4282.880 2771.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2848.080 5.440 2851.080 219.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2848.080 984.710 2851.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2848.080 4282.880 2851.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2928.080 5.440 2931.080 86.730 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2928.080 144.725 2931.080 219.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2928.080 984.710 2931.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2928.080 4282.880 2931.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3008.080 5.440 3011.080 219.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3008.080 984.710 3011.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3008.080 4282.880 3011.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3108.080 5.440 3111.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 3135.620 5.440 3138.620 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 45.080 5.440 48.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 69.940 5.440 72.940 4357.520 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 86.590 2896.855 89.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 146.590 2896.355 149.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 206.590 3167.520 209.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 266.590 2549.760 269.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 326.590 2549.760 329.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 386.590 2549.760 389.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 446.590 2549.760 449.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 506.590 2549.760 509.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 566.590 2549.760 569.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 626.590 2549.760 629.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 686.590 2549.760 689.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 746.590 2549.760 749.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 806.590 2549.760 809.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 866.590 2549.760 869.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 926.590 601.540 929.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 986.590 3167.520 989.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1046.590 1561.540 1049.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1106.590 1561.540 1109.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1166.590 3167.520 1169.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1226.590 3167.520 1229.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1286.590 93.140 1289.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1346.590 93.140 1349.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1406.590 93.140 1409.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1466.590 93.140 1469.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1526.590 93.140 1529.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1586.590 93.140 1589.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1646.590 93.140 1649.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1706.590 93.140 1709.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1766.590 93.140 1769.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1826.590 93.140 1829.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1886.590 93.140 1889.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 1946.590 93.140 1949.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2006.590 93.140 2009.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2066.590 93.140 2069.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2126.590 93.140 2129.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2186.590 93.140 2189.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2246.590 93.140 2249.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2306.590 93.140 2309.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2366.590 93.140 2369.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2426.590 93.140 2429.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2486.590 93.140 2489.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2546.590 93.140 2549.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2606.590 93.140 2609.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2666.590 93.140 2669.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2726.590 93.140 2729.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2786.590 93.140 2789.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2846.590 93.140 2849.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2906.590 93.140 2909.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 2966.590 93.140 2969.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3026.590 93.140 3029.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3086.590 93.140 3089.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3146.590 93.140 3149.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3206.590 93.140 3209.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3266.590 93.140 3269.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3326.590 93.140 3329.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3386.590 93.140 3389.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3446.590 93.140 3449.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3506.590 93.140 3509.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3566.590 93.140 3569.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3626.590 93.140 3629.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3686.590 93.140 3689.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3746.590 93.140 3749.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3806.590 93.140 3809.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3866.590 93.140 3869.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3926.590 93.140 3929.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 3986.590 93.140 3989.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4046.590 93.140 4049.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4106.590 93.140 4109.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4166.590 93.140 4169.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4226.590 93.140 4229.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.080 4286.590 3167.520 4289.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 672.460 926.590 1081.540 929.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1152.460 926.590 2549.760 929.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1632.460 1046.590 2121.040 1049.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1632.460 1106.590 2121.040 1109.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2191.960 1046.590 3167.520 1049.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2191.960 1106.590 3167.520 1109.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2966.995 86.590 3167.520 89.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2966.995 146.590 3167.520 149.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 266.590 3167.520 269.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 326.590 3167.520 329.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 386.590 3167.520 389.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 446.590 3167.520 449.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 506.590 3167.520 509.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 566.590 3167.520 569.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 626.590 3167.520 629.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 686.590 3167.520 689.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 746.590 3167.520 749.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 806.590 3167.520 809.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 866.590 3167.520 869.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3054.560 926.590 3167.520 929.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1286.590 3167.520 1289.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1346.590 3167.520 1349.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1406.590 3167.520 1409.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1466.590 3167.520 1469.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1526.590 3167.520 1529.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1586.590 3167.520 1589.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1646.590 3167.520 1649.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1706.590 3167.520 1709.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1766.590 3167.520 1769.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1826.590 3167.520 1829.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1886.590 3167.520 1889.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 1946.590 3167.520 1949.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2006.590 3167.520 2009.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2066.590 3167.520 2069.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2126.590 3167.520 2129.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2186.590 3167.520 2189.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2246.590 3167.520 2249.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2306.590 3167.520 2309.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2366.590 3167.520 2369.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2426.590 3167.520 2429.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2486.590 3167.520 2489.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2546.590 3167.520 2549.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2606.590 3167.520 2609.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2666.590 3167.520 2669.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2726.590 3167.520 2729.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2786.590 3167.520 2789.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2846.590 3167.520 2849.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2906.590 3167.520 2909.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 2966.590 3167.520 2969.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3026.590 3167.520 3029.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3086.590 3167.520 3089.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3146.590 3167.520 3149.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3206.590 3167.520 3209.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3266.590 3167.520 3269.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3326.590 3167.520 3329.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3386.590 3167.520 3389.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3446.590 3167.520 3449.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3506.590 3167.520 3509.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3566.590 3167.520 3569.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3626.590 3167.520 3629.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3686.590 3167.520 3689.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3746.590 3167.520 3749.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3806.590 3167.520 3809.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3866.590 3167.520 3869.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3926.590 3167.520 3929.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 3986.590 3167.520 3989.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 4046.590 3167.520 4049.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 4106.590 3167.520 4109.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 4166.590 3167.520 4169.590 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3076.860 4226.590 3167.520 4229.590 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2353.080 5.440 2356.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2353.080 4282.880 2356.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2892.580 5.440 2895.580 219.050 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2892.580 984.710 2895.580 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2892.580 4282.880 2895.580 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2170.080 5.440 2173.080 1031.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2170.080 1123.280 2173.080 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2170.080 4282.880 2173.080 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1923.380 5.440 1926.380 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1923.380 4282.880 1926.380 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1366.380 5.440 1369.380 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1366.380 4282.880 1369.380 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1123.480 5.440 1126.480 891.720 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1123.480 983.280 1126.480 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1123.480 4282.880 1126.480 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 871.780 5.440 874.780 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 871.780 4282.880 874.780 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 563.280 5.440 566.280 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 563.280 4282.880 566.280 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 313.580 5.440 316.580 1266.320 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 313.580 4282.880 316.580 4357.520 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1026.010 58.500 1027.510 576.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1482.970 58.500 1484.470 576.540 ;
    END
  END VSS
  PIN clock_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 790.860 -4.000 791.240 4.000 ;
    END
  END clock_core
  PIN const_one[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.965 -4.000 451.345 4.000 ;
    END
  END const_one[0]
  PIN const_one[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1275.965 -4.220 1276.345 4.000 ;
    END
  END const_one[1]
  PIN const_zero[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2163.670 -4.010 2164.050 4.000 ;
    END
  END const_zero[0]
  PIN const_zero[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1888.670 -4.010 1889.050 4.000 ;
    END
  END const_zero[1]
  PIN const_zero[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1613.670 -4.010 1614.050 4.000 ;
    END
  END const_zero[2]
  PIN const_zero[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1338.665 -4.000 1339.055 4.000 ;
    END
  END const_zero[3]
  PIN const_zero[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 725.965 -4.050 726.345 4.000 ;
    END
  END const_zero[4]
  PIN const_zero[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 455.330 -4.000 455.710 4.000 ;
    END
  END const_zero[5]
  PIN const_zero[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2373.360 -4.010 2373.740 4.000 ;
    END
  END const_zero[6]
  PIN const_zero[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2375.965 -4.010 2376.345 4.000 ;
    END
  END const_zero[7]
  PIN const_zero[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2380.330 -4.010 2380.710 4.000 ;
    END
  END const_zero[8]
  PIN const_zero[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2438.670 -4.010 2439.050 4.000 ;
    END
  END const_zero[9]
  PIN flash_clk_frame
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1614.400 -4.000 1614.780 4.000 ;
    END
  END flash_clk_frame
  PIN flash_clk_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1615.130 -4.000 1615.510 4.000 ;
    END
  END flash_clk_oe
  PIN flash_csb_frame
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1339.400 -4.000 1339.780 4.000 ;
    END
  END flash_csb_frame
  PIN flash_csb_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1340.130 -4.000 1340.510 4.000 ;
    END
  END flash_csb_oe
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1890.855 -4.000 1891.235 4.000 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1889.400 -4.000 1889.780 4.000 ;
    END
  END flash_io0_do
  PIN flash_io0_ie
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1831.385 -4.000 1831.765 4.000 ;
    END
  END flash_io0_ie
  PIN flash_io0_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1890.130 -4.000 1890.510 4.000 ;
    END
  END flash_io0_oe
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2165.860 -4.000 2166.240 4.000 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2164.400 -4.000 2164.780 4.000 ;
    END
  END flash_io1_do
  PIN flash_io1_ie
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2106.385 -4.000 2106.765 4.000 ;
    END
  END flash_io1_ie
  PIN flash_io1_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2165.130 -4.000 2165.510 4.000 ;
    END
  END flash_io1_oe
  PIN gpio_drive_select_core[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2377.110 -4.000 2377.490 4.000 ;
    END
  END gpio_drive_select_core[0]
  PIN gpio_drive_select_core[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2377.820 -4.000 2378.200 4.000 ;
    END
  END gpio_drive_select_core[1]
  PIN gpio_in_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2440.860 -4.000 2441.240 4.000 ;
    END
  END gpio_in_core
  PIN gpio_inenb_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2381.385 -4.000 2381.765 4.000 ;
    END
  END gpio_inenb_core
  PIN gpio_out_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2439.400 -4.000 2439.780 4.000 ;
    END
  END gpio_out_core
  PIN gpio_outenb_core
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2440.130 -4.000 2440.510 4.000 ;
    END
  END gpio_outenb_core
  PIN mprj_io_drive_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 97.110 3174.000 97.490 ;
    END
  END mprj_io_drive_sel[0]
  PIN mprj_io_drive_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1172.110 3174.000 1172.490 ;
    END
  END mprj_io_drive_sel[10]
  PIN mprj_io_drive_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1172.820 3174.000 1173.200 ;
    END
  END mprj_io_drive_sel[11]
  PIN mprj_io_drive_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1387.110 3174.000 1387.490 ;
    END
  END mprj_io_drive_sel[12]
  PIN mprj_io_drive_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1387.820 3174.000 1388.200 ;
    END
  END mprj_io_drive_sel[13]
  PIN mprj_io_drive_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2247.110 3174.000 2247.490 ;
    END
  END mprj_io_drive_sel[14]
  PIN mprj_io_drive_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2247.820 3174.000 2248.200 ;
    END
  END mprj_io_drive_sel[15]
  PIN mprj_io_drive_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2462.110 3174.000 2462.490 ;
    END
  END mprj_io_drive_sel[16]
  PIN mprj_io_drive_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2462.820 3174.000 2463.200 ;
    END
  END mprj_io_drive_sel[17]
  PIN mprj_io_drive_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2677.110 3174.000 2677.490 ;
    END
  END mprj_io_drive_sel[18]
  PIN mprj_io_drive_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2677.820 3174.000 2678.200 ;
    END
  END mprj_io_drive_sel[19]
  PIN mprj_io_drive_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 97.820 3174.000 98.200 ;
    END
  END mprj_io_drive_sel[1]
  PIN mprj_io_drive_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2892.110 3174.000 2892.490 ;
    END
  END mprj_io_drive_sel[20]
  PIN mprj_io_drive_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2892.820 3174.000 2893.200 ;
    END
  END mprj_io_drive_sel[21]
  PIN mprj_io_drive_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3107.110 3174.000 3107.490 ;
    END
  END mprj_io_drive_sel[22]
  PIN mprj_io_drive_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3107.820 3174.000 3108.200 ;
    END
  END mprj_io_drive_sel[23]
  PIN mprj_io_drive_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3322.110 3174.000 3322.490 ;
    END
  END mprj_io_drive_sel[24]
  PIN mprj_io_drive_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3322.820 3174.000 3323.200 ;
    END
  END mprj_io_drive_sel[25]
  PIN mprj_io_drive_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3752.110 3174.000 3752.490 ;
    END
  END mprj_io_drive_sel[26]
  PIN mprj_io_drive_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3752.820 3174.000 3753.200 ;
    END
  END mprj_io_drive_sel[27]
  PIN mprj_io_drive_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 4182.110 3174.000 4182.490 ;
    END
  END mprj_io_drive_sel[28]
  PIN mprj_io_drive_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 4182.820 3174.000 4183.200 ;
    END
  END mprj_io_drive_sel[29]
  PIN mprj_io_drive_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 312.110 3174.000 312.490 ;
    END
  END mprj_io_drive_sel[2]
  PIN mprj_io_drive_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2982.510 4356.000 2982.890 4364.000 ;
    END
  END mprj_io_drive_sel[30]
  PIN mprj_io_drive_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2981.800 4356.000 2982.180 4364.000 ;
    END
  END mprj_io_drive_sel[31]
  PIN mprj_io_drive_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2432.510 4356.000 2432.890 4364.000 ;
    END
  END mprj_io_drive_sel[32]
  PIN mprj_io_drive_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2431.800 4356.000 2432.180 4364.000 ;
    END
  END mprj_io_drive_sel[33]
  PIN mprj_io_drive_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2157.510 4356.000 2157.890 4364.000 ;
    END
  END mprj_io_drive_sel[34]
  PIN mprj_io_drive_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2156.800 4356.000 2157.180 4364.000 ;
    END
  END mprj_io_drive_sel[35]
  PIN mprj_io_drive_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1882.510 4356.000 1882.890 4364.000 ;
    END
  END mprj_io_drive_sel[36]
  PIN mprj_io_drive_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1881.800 4356.000 1882.180 4364.000 ;
    END
  END mprj_io_drive_sel[37]
  PIN mprj_io_drive_sel[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1332.510 4356.000 1332.890 4364.000 ;
    END
  END mprj_io_drive_sel[38]
  PIN mprj_io_drive_sel[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1331.800 4356.000 1332.180 4364.000 ;
    END
  END mprj_io_drive_sel[39]
  PIN mprj_io_drive_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 312.820 3174.000 313.200 ;
    END
  END mprj_io_drive_sel[3]
  PIN mprj_io_drive_sel[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1057.510 4356.000 1057.890 4364.000 ;
    END
  END mprj_io_drive_sel[40]
  PIN mprj_io_drive_sel[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1056.800 4356.000 1057.180 4364.000 ;
    END
  END mprj_io_drive_sel[41]
  PIN mprj_io_drive_sel[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 782.510 4356.000 782.890 4364.000 ;
    END
  END mprj_io_drive_sel[42]
  PIN mprj_io_drive_sel[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 781.800 4356.000 782.180 4364.000 ;
    END
  END mprj_io_drive_sel[43]
  PIN mprj_io_drive_sel[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 507.510 4356.000 507.890 4364.000 ;
    END
  END mprj_io_drive_sel[44]
  PIN mprj_io_drive_sel[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 506.800 4356.000 507.180 4364.000 ;
    END
  END mprj_io_drive_sel[45]
  PIN mprj_io_drive_sel[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 232.510 4356.000 232.890 4364.000 ;
    END
  END mprj_io_drive_sel[46]
  PIN mprj_io_drive_sel[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.800 4356.000 232.180 4364.000 ;
    END
  END mprj_io_drive_sel[47]
  PIN mprj_io_drive_sel[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 4237.510 4.000 4237.890 ;
    END
  END mprj_io_drive_sel[48]
  PIN mprj_io_drive_sel[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 4236.800 4.000 4237.180 ;
    END
  END mprj_io_drive_sel[49]
  PIN mprj_io_drive_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 527.110 3174.000 527.490 ;
    END
  END mprj_io_drive_sel[4]
  PIN mprj_io_drive_sel[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3417.510 4.000 3417.890 ;
    END
  END mprj_io_drive_sel[50]
  PIN mprj_io_drive_sel[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3416.800 4.000 3417.180 ;
    END
  END mprj_io_drive_sel[51]
  PIN mprj_io_drive_sel[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3212.510 4.000 3212.890 ;
    END
  END mprj_io_drive_sel[52]
  PIN mprj_io_drive_sel[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3211.800 4.000 3212.180 ;
    END
  END mprj_io_drive_sel[53]
  PIN mprj_io_drive_sel[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3007.510 4.000 3007.890 ;
    END
  END mprj_io_drive_sel[54]
  PIN mprj_io_drive_sel[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3006.800 4.000 3007.180 ;
    END
  END mprj_io_drive_sel[55]
  PIN mprj_io_drive_sel[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2802.510 4.000 2802.890 ;
    END
  END mprj_io_drive_sel[56]
  PIN mprj_io_drive_sel[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2801.800 4.000 2802.180 ;
    END
  END mprj_io_drive_sel[57]
  PIN mprj_io_drive_sel[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2597.510 4.000 2597.890 ;
    END
  END mprj_io_drive_sel[58]
  PIN mprj_io_drive_sel[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2596.800 4.000 2597.180 ;
    END
  END mprj_io_drive_sel[59]
  PIN mprj_io_drive_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 527.820 3174.000 528.200 ;
    END
  END mprj_io_drive_sel[5]
  PIN mprj_io_drive_sel[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2392.510 4.000 2392.890 ;
    END
  END mprj_io_drive_sel[60]
  PIN mprj_io_drive_sel[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2391.800 4.000 2392.180 ;
    END
  END mprj_io_drive_sel[61]
  PIN mprj_io_drive_sel[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2187.510 4.000 2187.890 ;
    END
  END mprj_io_drive_sel[62]
  PIN mprj_io_drive_sel[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2186.800 4.000 2187.180 ;
    END
  END mprj_io_drive_sel[63]
  PIN mprj_io_drive_sel[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1572.510 4.000 1572.890 ;
    END
  END mprj_io_drive_sel[64]
  PIN mprj_io_drive_sel[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1571.800 4.000 1572.180 ;
    END
  END mprj_io_drive_sel[65]
  PIN mprj_io_drive_sel[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1367.510 4.000 1367.890 ;
    END
  END mprj_io_drive_sel[66]
  PIN mprj_io_drive_sel[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1366.800 4.000 1367.180 ;
    END
  END mprj_io_drive_sel[67]
  PIN mprj_io_drive_sel[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1162.510 4.000 1162.890 ;
    END
  END mprj_io_drive_sel[68]
  PIN mprj_io_drive_sel[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1161.800 4.000 1162.180 ;
    END
  END mprj_io_drive_sel[69]
  PIN mprj_io_drive_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 742.110 3174.000 742.490 ;
    END
  END mprj_io_drive_sel[6]
  PIN mprj_io_drive_sel[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 957.510 4.000 957.890 ;
    END
  END mprj_io_drive_sel[70]
  PIN mprj_io_drive_sel[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 956.800 4.000 957.180 ;
    END
  END mprj_io_drive_sel[71]
  PIN mprj_io_drive_sel[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 752.510 4.000 752.890 ;
    END
  END mprj_io_drive_sel[72]
  PIN mprj_io_drive_sel[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 751.800 4.000 752.180 ;
    END
  END mprj_io_drive_sel[73]
  PIN mprj_io_drive_sel[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 547.510 4.000 547.890 ;
    END
  END mprj_io_drive_sel[74]
  PIN mprj_io_drive_sel[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 546.800 4.000 547.180 ;
    END
  END mprj_io_drive_sel[75]
  PIN mprj_io_drive_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 742.820 3174.000 743.200 ;
    END
  END mprj_io_drive_sel[7]
  PIN mprj_io_drive_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 957.110 3174.000 957.490 ;
    END
  END mprj_io_drive_sel[8]
  PIN mprj_io_drive_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 957.820 3174.000 958.200 ;
    END
  END mprj_io_drive_sel[9]
  PIN mprj_io_ie[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 101.385 3174.000 101.765 ;
    END
  END mprj_io_ie[0]
  PIN mprj_io_ie[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2896.385 3174.000 2896.765 ;
    END
  END mprj_io_ie[10]
  PIN mprj_io_ie[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3111.385 3174.000 3111.765 ;
    END
  END mprj_io_ie[11]
  PIN mprj_io_ie[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3326.385 3174.000 3326.765 ;
    END
  END mprj_io_ie[12]
  PIN mprj_io_ie[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3756.385 3174.000 3756.765 ;
    END
  END mprj_io_ie[13]
  PIN mprj_io_ie[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 4186.385 3174.000 4186.765 ;
    END
  END mprj_io_ie[14]
  PIN mprj_io_ie[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2978.235 4356.000 2978.615 4364.000 ;
    END
  END mprj_io_ie[15]
  PIN mprj_io_ie[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2428.235 4356.000 2428.615 4364.000 ;
    END
  END mprj_io_ie[16]
  PIN mprj_io_ie[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2153.235 4356.000 2153.615 4364.000 ;
    END
  END mprj_io_ie[17]
  PIN mprj_io_ie[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1878.235 4356.000 1878.615 4364.000 ;
    END
  END mprj_io_ie[18]
  PIN mprj_io_ie[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1328.235 4356.000 1328.615 4364.000 ;
    END
  END mprj_io_ie[19]
  PIN mprj_io_ie[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 316.385 3174.000 316.765 ;
    END
  END mprj_io_ie[1]
  PIN mprj_io_ie[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1053.235 4356.000 1053.615 4364.000 ;
    END
  END mprj_io_ie[20]
  PIN mprj_io_ie[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 778.235 4356.000 778.615 4364.000 ;
    END
  END mprj_io_ie[21]
  PIN mprj_io_ie[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 503.235 4356.000 503.615 4364.000 ;
    END
  END mprj_io_ie[22]
  PIN mprj_io_ie[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.235 4356.000 228.615 4364.000 ;
    END
  END mprj_io_ie[23]
  PIN mprj_io_ie[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 4233.235 4.000 4233.615 ;
    END
  END mprj_io_ie[24]
  PIN mprj_io_ie[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3413.235 4.000 3413.615 ;
    END
  END mprj_io_ie[25]
  PIN mprj_io_ie[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3208.235 4.000 3208.615 ;
    END
  END mprj_io_ie[26]
  PIN mprj_io_ie[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3003.235 4.000 3003.615 ;
    END
  END mprj_io_ie[27]
  PIN mprj_io_ie[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2798.235 4.000 2798.615 ;
    END
  END mprj_io_ie[28]
  PIN mprj_io_ie[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2593.235 4.000 2593.615 ;
    END
  END mprj_io_ie[29]
  PIN mprj_io_ie[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 531.385 3174.000 531.765 ;
    END
  END mprj_io_ie[2]
  PIN mprj_io_ie[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2388.235 4.000 2388.615 ;
    END
  END mprj_io_ie[30]
  PIN mprj_io_ie[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2183.235 4.000 2183.615 ;
    END
  END mprj_io_ie[31]
  PIN mprj_io_ie[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1568.235 4.000 1568.615 ;
    END
  END mprj_io_ie[32]
  PIN mprj_io_ie[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1363.235 4.000 1363.615 ;
    END
  END mprj_io_ie[33]
  PIN mprj_io_ie[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1158.235 4.000 1158.615 ;
    END
  END mprj_io_ie[34]
  PIN mprj_io_ie[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 953.235 4.000 953.615 ;
    END
  END mprj_io_ie[35]
  PIN mprj_io_ie[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 748.235 4.000 748.615 ;
    END
  END mprj_io_ie[36]
  PIN mprj_io_ie[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 543.235 4.000 543.615 ;
    END
  END mprj_io_ie[37]
  PIN mprj_io_ie[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 746.385 3174.000 746.765 ;
    END
  END mprj_io_ie[3]
  PIN mprj_io_ie[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 961.385 3174.000 961.765 ;
    END
  END mprj_io_ie[4]
  PIN mprj_io_ie[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1176.385 3174.000 1176.765 ;
    END
  END mprj_io_ie[5]
  PIN mprj_io_ie[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1391.385 3174.000 1391.765 ;
    END
  END mprj_io_ie[6]
  PIN mprj_io_ie[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2251.385 3174.000 2251.765 ;
    END
  END mprj_io_ie[7]
  PIN mprj_io_ie[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2466.385 3174.000 2466.765 ;
    END
  END mprj_io_ie[8]
  PIN mprj_io_ie[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2681.385 3174.000 2681.765 ;
    END
  END mprj_io_ie[9]
  PIN mprj_io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 160.860 3174.000 161.240 ;
    END
  END mprj_io_in[0]
  PIN mprj_io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2955.860 3174.000 2956.240 ;
    END
  END mprj_io_in[10]
  PIN mprj_io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3170.860 3174.000 3171.240 ;
    END
  END mprj_io_in[11]
  PIN mprj_io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3385.860 3174.000 3386.240 ;
    END
  END mprj_io_in[12]
  PIN mprj_io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3815.860 3174.000 3816.240 ;
    END
  END mprj_io_in[13]
  PIN mprj_io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 4245.860 3174.000 4246.240 ;
    END
  END mprj_io_in[14]
  PIN mprj_io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2918.760 4356.000 2919.140 4364.000 ;
    END
  END mprj_io_in[15]
  PIN mprj_io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2368.760 4356.000 2369.140 4364.000 ;
    END
  END mprj_io_in[16]
  PIN mprj_io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2093.760 4356.000 2094.140 4364.000 ;
    END
  END mprj_io_in[17]
  PIN mprj_io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1818.760 4356.000 1819.140 4364.000 ;
    END
  END mprj_io_in[18]
  PIN mprj_io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1268.760 4356.000 1269.140 4364.000 ;
    END
  END mprj_io_in[19]
  PIN mprj_io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 375.860 3174.000 376.240 ;
    END
  END mprj_io_in[1]
  PIN mprj_io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 993.760 4356.000 994.140 4364.000 ;
    END
  END mprj_io_in[20]
  PIN mprj_io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 718.760 4356.000 719.140 4364.000 ;
    END
  END mprj_io_in[21]
  PIN mprj_io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 443.760 4356.000 444.140 4364.000 ;
    END
  END mprj_io_in[22]
  PIN mprj_io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.760 4356.000 169.140 4364.000 ;
    END
  END mprj_io_in[23]
  PIN mprj_io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 4173.760 4.000 4174.140 ;
    END
  END mprj_io_in[24]
  PIN mprj_io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3353.760 4.000 3354.140 ;
    END
  END mprj_io_in[25]
  PIN mprj_io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3148.760 4.000 3149.140 ;
    END
  END mprj_io_in[26]
  PIN mprj_io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2943.760 4.000 2944.140 ;
    END
  END mprj_io_in[27]
  PIN mprj_io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2738.760 4.000 2739.140 ;
    END
  END mprj_io_in[28]
  PIN mprj_io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2533.760 4.000 2534.140 ;
    END
  END mprj_io_in[29]
  PIN mprj_io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 590.860 3174.000 591.240 ;
    END
  END mprj_io_in[2]
  PIN mprj_io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2328.760 4.000 2329.140 ;
    END
  END mprj_io_in[30]
  PIN mprj_io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2123.760 4.000 2124.140 ;
    END
  END mprj_io_in[31]
  PIN mprj_io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1508.760 4.000 1509.140 ;
    END
  END mprj_io_in[32]
  PIN mprj_io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1303.760 4.000 1304.140 ;
    END
  END mprj_io_in[33]
  PIN mprj_io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1098.760 4.000 1099.140 ;
    END
  END mprj_io_in[34]
  PIN mprj_io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 893.760 4.000 894.140 ;
    END
  END mprj_io_in[35]
  PIN mprj_io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 688.760 4.000 689.140 ;
    END
  END mprj_io_in[36]
  PIN mprj_io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 483.760 4.000 484.140 ;
    END
  END mprj_io_in[37]
  PIN mprj_io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 805.860 3174.000 806.240 ;
    END
  END mprj_io_in[3]
  PIN mprj_io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1020.860 3174.000 1021.240 ;
    END
  END mprj_io_in[4]
  PIN mprj_io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1235.860 3174.000 1236.240 ;
    END
  END mprj_io_in[5]
  PIN mprj_io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1450.860 3174.000 1451.240 ;
    END
  END mprj_io_in[6]
  PIN mprj_io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2310.860 3174.000 2311.240 ;
    END
  END mprj_io_in[7]
  PIN mprj_io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2525.860 3174.000 2526.240 ;
    END
  END mprj_io_in[8]
  PIN mprj_io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2740.860 3174.000 2741.240 ;
    END
  END mprj_io_in[9]
  PIN mprj_io_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 160.130 3174.000 160.510 ;
    END
  END mprj_io_oe[0]
  PIN mprj_io_oe[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2955.130 3174.000 2955.510 ;
    END
  END mprj_io_oe[10]
  PIN mprj_io_oe[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3170.130 3174.000 3170.510 ;
    END
  END mprj_io_oe[11]
  PIN mprj_io_oe[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3385.130 3174.000 3385.510 ;
    END
  END mprj_io_oe[12]
  PIN mprj_io_oe[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3815.130 3174.000 3815.510 ;
    END
  END mprj_io_oe[13]
  PIN mprj_io_oe[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 4245.130 3174.000 4245.510 ;
    END
  END mprj_io_oe[14]
  PIN mprj_io_oe[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2919.490 4356.000 2919.870 4364.000 ;
    END
  END mprj_io_oe[15]
  PIN mprj_io_oe[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2369.490 4356.000 2369.870 4364.000 ;
    END
  END mprj_io_oe[16]
  PIN mprj_io_oe[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2094.490 4356.000 2094.870 4364.000 ;
    END
  END mprj_io_oe[17]
  PIN mprj_io_oe[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1819.490 4356.000 1819.870 4364.000 ;
    END
  END mprj_io_oe[18]
  PIN mprj_io_oe[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1269.490 4356.000 1269.870 4364.000 ;
    END
  END mprj_io_oe[19]
  PIN mprj_io_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 375.130 3174.000 375.510 ;
    END
  END mprj_io_oe[1]
  PIN mprj_io_oe[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 994.490 4356.000 994.870 4364.000 ;
    END
  END mprj_io_oe[20]
  PIN mprj_io_oe[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 719.490 4356.000 719.870 4364.000 ;
    END
  END mprj_io_oe[21]
  PIN mprj_io_oe[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 444.490 4356.000 444.870 4364.000 ;
    END
  END mprj_io_oe[22]
  PIN mprj_io_oe[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 169.490 4356.000 169.870 4364.000 ;
    END
  END mprj_io_oe[23]
  PIN mprj_io_oe[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 4174.490 4.000 4174.870 ;
    END
  END mprj_io_oe[24]
  PIN mprj_io_oe[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3354.490 4.000 3354.870 ;
    END
  END mprj_io_oe[25]
  PIN mprj_io_oe[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3149.490 4.000 3149.870 ;
    END
  END mprj_io_oe[26]
  PIN mprj_io_oe[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2944.490 4.000 2944.870 ;
    END
  END mprj_io_oe[27]
  PIN mprj_io_oe[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2739.490 4.000 2739.870 ;
    END
  END mprj_io_oe[28]
  PIN mprj_io_oe[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2534.490 4.000 2534.870 ;
    END
  END mprj_io_oe[29]
  PIN mprj_io_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 590.130 3174.000 590.510 ;
    END
  END mprj_io_oe[2]
  PIN mprj_io_oe[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2329.490 4.000 2329.870 ;
    END
  END mprj_io_oe[30]
  PIN mprj_io_oe[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2124.490 4.000 2124.870 ;
    END
  END mprj_io_oe[31]
  PIN mprj_io_oe[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1509.490 4.000 1509.870 ;
    END
  END mprj_io_oe[32]
  PIN mprj_io_oe[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1304.490 4.000 1304.870 ;
    END
  END mprj_io_oe[33]
  PIN mprj_io_oe[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1099.490 4.000 1099.870 ;
    END
  END mprj_io_oe[34]
  PIN mprj_io_oe[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 894.490 4.000 894.870 ;
    END
  END mprj_io_oe[35]
  PIN mprj_io_oe[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 689.490 4.000 689.870 ;
    END
  END mprj_io_oe[36]
  PIN mprj_io_oe[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 484.490 4.000 484.870 ;
    END
  END mprj_io_oe[37]
  PIN mprj_io_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 805.130 3174.000 805.510 ;
    END
  END mprj_io_oe[3]
  PIN mprj_io_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1020.130 3174.000 1020.510 ;
    END
  END mprj_io_oe[4]
  PIN mprj_io_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1235.130 3174.000 1235.510 ;
    END
  END mprj_io_oe[5]
  PIN mprj_io_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1450.130 3174.000 1450.510 ;
    END
  END mprj_io_oe[6]
  PIN mprj_io_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2310.130 3174.000 2310.510 ;
    END
  END mprj_io_oe[7]
  PIN mprj_io_oe[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2525.130 3174.000 2525.510 ;
    END
  END mprj_io_oe[8]
  PIN mprj_io_oe[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2740.130 3174.000 2740.510 ;
    END
  END mprj_io_oe[9]
  PIN mprj_io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 159.400 3174.000 159.780 ;
    END
  END mprj_io_out[0]
  PIN mprj_io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2954.400 3174.000 2954.780 ;
    END
  END mprj_io_out[10]
  PIN mprj_io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3169.400 3174.000 3169.780 ;
    END
  END mprj_io_out[11]
  PIN mprj_io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3384.400 3174.000 3384.780 ;
    END
  END mprj_io_out[12]
  PIN mprj_io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3814.400 3174.000 3814.780 ;
    END
  END mprj_io_out[13]
  PIN mprj_io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 4244.400 3174.000 4244.780 ;
    END
  END mprj_io_out[14]
  PIN mprj_io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2920.220 4356.000 2920.600 4364.000 ;
    END
  END mprj_io_out[15]
  PIN mprj_io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2370.220 4356.000 2370.600 4364.000 ;
    END
  END mprj_io_out[16]
  PIN mprj_io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2095.220 4356.000 2095.600 4364.000 ;
    END
  END mprj_io_out[17]
  PIN mprj_io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1820.220 4356.000 1820.600 4364.000 ;
    END
  END mprj_io_out[18]
  PIN mprj_io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1270.220 4356.000 1270.600 4364.000 ;
    END
  END mprj_io_out[19]
  PIN mprj_io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 374.400 3174.000 374.780 ;
    END
  END mprj_io_out[1]
  PIN mprj_io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 995.220 4356.000 995.600 4364.000 ;
    END
  END mprj_io_out[20]
  PIN mprj_io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 720.220 4356.000 720.600 4364.000 ;
    END
  END mprj_io_out[21]
  PIN mprj_io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 445.220 4356.000 445.600 4364.000 ;
    END
  END mprj_io_out[22]
  PIN mprj_io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 170.220 4356.000 170.600 4364.000 ;
    END
  END mprj_io_out[23]
  PIN mprj_io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 4175.220 4.000 4175.600 ;
    END
  END mprj_io_out[24]
  PIN mprj_io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3355.220 4.000 3355.600 ;
    END
  END mprj_io_out[25]
  PIN mprj_io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3150.220 4.000 3150.600 ;
    END
  END mprj_io_out[26]
  PIN mprj_io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2945.220 4.000 2945.600 ;
    END
  END mprj_io_out[27]
  PIN mprj_io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2740.220 4.000 2740.600 ;
    END
  END mprj_io_out[28]
  PIN mprj_io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2535.220 4.000 2535.600 ;
    END
  END mprj_io_out[29]
  PIN mprj_io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 589.400 3174.000 589.780 ;
    END
  END mprj_io_out[2]
  PIN mprj_io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2330.220 4.000 2330.600 ;
    END
  END mprj_io_out[30]
  PIN mprj_io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2125.220 4.000 2125.600 ;
    END
  END mprj_io_out[31]
  PIN mprj_io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1510.220 4.000 1510.600 ;
    END
  END mprj_io_out[32]
  PIN mprj_io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1305.220 4.000 1305.600 ;
    END
  END mprj_io_out[33]
  PIN mprj_io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1100.220 4.000 1100.600 ;
    END
  END mprj_io_out[34]
  PIN mprj_io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 895.220 4.000 895.600 ;
    END
  END mprj_io_out[35]
  PIN mprj_io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 690.220 4.000 690.600 ;
    END
  END mprj_io_out[36]
  PIN mprj_io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 485.220 4.000 485.600 ;
    END
  END mprj_io_out[37]
  PIN mprj_io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 804.400 3174.000 804.780 ;
    END
  END mprj_io_out[3]
  PIN mprj_io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1019.400 3174.000 1019.780 ;
    END
  END mprj_io_out[4]
  PIN mprj_io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1234.400 3174.000 1234.780 ;
    END
  END mprj_io_out[5]
  PIN mprj_io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1449.400 3174.000 1449.780 ;
    END
  END mprj_io_out[6]
  PIN mprj_io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2309.400 3174.000 2309.780 ;
    END
  END mprj_io_out[7]
  PIN mprj_io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2524.400 3174.000 2524.780 ;
    END
  END mprj_io_out[8]
  PIN mprj_io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2739.400 3174.000 2739.780 ;
    END
  END mprj_io_out[9]
  PIN mprj_io_pulldown_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 100.330 3174.000 100.710 ;
    END
  END mprj_io_pulldown_sel[0]
  PIN mprj_io_pulldown_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2895.330 3174.000 2895.710 ;
    END
  END mprj_io_pulldown_sel[10]
  PIN mprj_io_pulldown_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3110.330 3174.000 3110.710 ;
    END
  END mprj_io_pulldown_sel[11]
  PIN mprj_io_pulldown_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3325.330 3174.000 3325.710 ;
    END
  END mprj_io_pulldown_sel[12]
  PIN mprj_io_pulldown_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3755.330 3174.000 3755.710 ;
    END
  END mprj_io_pulldown_sel[13]
  PIN mprj_io_pulldown_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 4185.330 3174.000 4185.710 ;
    END
  END mprj_io_pulldown_sel[14]
  PIN mprj_io_pulldown_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2979.290 4356.000 2979.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[15]
  PIN mprj_io_pulldown_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2429.290 4356.000 2429.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[16]
  PIN mprj_io_pulldown_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2154.290 4356.000 2154.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[17]
  PIN mprj_io_pulldown_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1879.290 4356.000 1879.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[18]
  PIN mprj_io_pulldown_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1329.290 4356.000 1329.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[19]
  PIN mprj_io_pulldown_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 315.330 3174.000 315.710 ;
    END
  END mprj_io_pulldown_sel[1]
  PIN mprj_io_pulldown_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1054.290 4356.000 1054.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[20]
  PIN mprj_io_pulldown_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 779.290 4356.000 779.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[21]
  PIN mprj_io_pulldown_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 504.290 4356.000 504.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[22]
  PIN mprj_io_pulldown_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 229.290 4356.000 229.670 4364.000 ;
    END
  END mprj_io_pulldown_sel[23]
  PIN mprj_io_pulldown_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 4234.290 4.000 4234.670 ;
    END
  END mprj_io_pulldown_sel[24]
  PIN mprj_io_pulldown_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3414.290 4.000 3414.670 ;
    END
  END mprj_io_pulldown_sel[25]
  PIN mprj_io_pulldown_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3209.290 4.000 3209.670 ;
    END
  END mprj_io_pulldown_sel[26]
  PIN mprj_io_pulldown_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3004.290 4.000 3004.670 ;
    END
  END mprj_io_pulldown_sel[27]
  PIN mprj_io_pulldown_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2799.290 4.000 2799.670 ;
    END
  END mprj_io_pulldown_sel[28]
  PIN mprj_io_pulldown_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2594.290 4.000 2594.670 ;
    END
  END mprj_io_pulldown_sel[29]
  PIN mprj_io_pulldown_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 530.330 3174.000 530.710 ;
    END
  END mprj_io_pulldown_sel[2]
  PIN mprj_io_pulldown_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2389.290 4.000 2389.670 ;
    END
  END mprj_io_pulldown_sel[30]
  PIN mprj_io_pulldown_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2184.290 4.000 2184.670 ;
    END
  END mprj_io_pulldown_sel[31]
  PIN mprj_io_pulldown_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1569.290 4.000 1569.670 ;
    END
  END mprj_io_pulldown_sel[32]
  PIN mprj_io_pulldown_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1364.290 4.000 1364.670 ;
    END
  END mprj_io_pulldown_sel[33]
  PIN mprj_io_pulldown_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1159.290 4.000 1159.670 ;
    END
  END mprj_io_pulldown_sel[34]
  PIN mprj_io_pulldown_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 954.290 4.000 954.670 ;
    END
  END mprj_io_pulldown_sel[35]
  PIN mprj_io_pulldown_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 749.290 4.000 749.670 ;
    END
  END mprj_io_pulldown_sel[36]
  PIN mprj_io_pulldown_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 544.290 4.000 544.670 ;
    END
  END mprj_io_pulldown_sel[37]
  PIN mprj_io_pulldown_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 745.330 3174.000 745.710 ;
    END
  END mprj_io_pulldown_sel[3]
  PIN mprj_io_pulldown_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 960.330 3174.000 960.710 ;
    END
  END mprj_io_pulldown_sel[4]
  PIN mprj_io_pulldown_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1175.330 3174.000 1175.710 ;
    END
  END mprj_io_pulldown_sel[5]
  PIN mprj_io_pulldown_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1390.330 3174.000 1390.710 ;
    END
  END mprj_io_pulldown_sel[6]
  PIN mprj_io_pulldown_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2250.330 3174.000 2250.710 ;
    END
  END mprj_io_pulldown_sel[7]
  PIN mprj_io_pulldown_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2465.330 3174.000 2465.710 ;
    END
  END mprj_io_pulldown_sel[8]
  PIN mprj_io_pulldown_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2680.330 3174.000 2680.710 ;
    END
  END mprj_io_pulldown_sel[9]
  PIN mprj_io_pullup_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 95.965 3174.000 96.345 ;
    END
  END mprj_io_pullup_sel[0]
  PIN mprj_io_pullup_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2890.965 3174.000 2891.345 ;
    END
  END mprj_io_pullup_sel[10]
  PIN mprj_io_pullup_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3105.965 3174.000 3106.345 ;
    END
  END mprj_io_pullup_sel[11]
  PIN mprj_io_pullup_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3320.965 3174.000 3321.345 ;
    END
  END mprj_io_pullup_sel[12]
  PIN mprj_io_pullup_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3750.965 3174.000 3751.345 ;
    END
  END mprj_io_pullup_sel[13]
  PIN mprj_io_pullup_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 4180.965 3174.000 4181.345 ;
    END
  END mprj_io_pullup_sel[14]
  PIN mprj_io_pullup_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2983.655 4356.000 2984.035 4364.000 ;
    END
  END mprj_io_pullup_sel[15]
  PIN mprj_io_pullup_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2433.655 4356.000 2434.035 4364.000 ;
    END
  END mprj_io_pullup_sel[16]
  PIN mprj_io_pullup_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2158.655 4356.000 2159.035 4364.000 ;
    END
  END mprj_io_pullup_sel[17]
  PIN mprj_io_pullup_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1883.655 4356.000 1884.035 4364.000 ;
    END
  END mprj_io_pullup_sel[18]
  PIN mprj_io_pullup_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1333.655 4356.000 1334.035 4364.000 ;
    END
  END mprj_io_pullup_sel[19]
  PIN mprj_io_pullup_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 310.965 3174.000 311.345 ;
    END
  END mprj_io_pullup_sel[1]
  PIN mprj_io_pullup_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1058.655 4356.000 1059.035 4364.000 ;
    END
  END mprj_io_pullup_sel[20]
  PIN mprj_io_pullup_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 783.655 4356.000 784.035 4364.000 ;
    END
  END mprj_io_pullup_sel[21]
  PIN mprj_io_pullup_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 508.655 4356.000 509.035 4364.000 ;
    END
  END mprj_io_pullup_sel[22]
  PIN mprj_io_pullup_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 233.655 4356.000 234.035 4364.000 ;
    END
  END mprj_io_pullup_sel[23]
  PIN mprj_io_pullup_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 4238.655 4.000 4239.035 ;
    END
  END mprj_io_pullup_sel[24]
  PIN mprj_io_pullup_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3418.655 4.000 3419.035 ;
    END
  END mprj_io_pullup_sel[25]
  PIN mprj_io_pullup_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3213.655 4.000 3214.035 ;
    END
  END mprj_io_pullup_sel[26]
  PIN mprj_io_pullup_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3008.655 4.000 3009.035 ;
    END
  END mprj_io_pullup_sel[27]
  PIN mprj_io_pullup_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2803.655 4.000 2804.035 ;
    END
  END mprj_io_pullup_sel[28]
  PIN mprj_io_pullup_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2598.655 4.000 2599.035 ;
    END
  END mprj_io_pullup_sel[29]
  PIN mprj_io_pullup_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 525.965 3174.000 526.345 ;
    END
  END mprj_io_pullup_sel[2]
  PIN mprj_io_pullup_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2393.655 4.000 2394.035 ;
    END
  END mprj_io_pullup_sel[30]
  PIN mprj_io_pullup_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2188.655 4.000 2189.035 ;
    END
  END mprj_io_pullup_sel[31]
  PIN mprj_io_pullup_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1573.655 4.000 1574.035 ;
    END
  END mprj_io_pullup_sel[32]
  PIN mprj_io_pullup_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1368.655 4.000 1369.035 ;
    END
  END mprj_io_pullup_sel[33]
  PIN mprj_io_pullup_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1163.655 4.000 1164.035 ;
    END
  END mprj_io_pullup_sel[34]
  PIN mprj_io_pullup_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 958.655 4.000 959.035 ;
    END
  END mprj_io_pullup_sel[35]
  PIN mprj_io_pullup_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 753.655 4.000 754.035 ;
    END
  END mprj_io_pullup_sel[36]
  PIN mprj_io_pullup_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 548.655 4.000 549.035 ;
    END
  END mprj_io_pullup_sel[37]
  PIN mprj_io_pullup_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 740.965 3174.000 741.345 ;
    END
  END mprj_io_pullup_sel[3]
  PIN mprj_io_pullup_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 955.965 3174.000 956.345 ;
    END
  END mprj_io_pullup_sel[4]
  PIN mprj_io_pullup_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1170.965 3174.000 1171.345 ;
    END
  END mprj_io_pullup_sel[5]
  PIN mprj_io_pullup_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1385.965 3174.000 1386.345 ;
    END
  END mprj_io_pullup_sel[6]
  PIN mprj_io_pullup_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2245.965 3174.000 2246.345 ;
    END
  END mprj_io_pullup_sel[7]
  PIN mprj_io_pullup_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2460.965 3174.000 2461.345 ;
    END
  END mprj_io_pullup_sel[8]
  PIN mprj_io_pullup_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2675.965 3174.000 2676.345 ;
    END
  END mprj_io_pullup_sel[9]
  PIN mprj_io_schmitt_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 93.360 3174.000 93.740 ;
    END
  END mprj_io_schmitt_sel[0]
  PIN mprj_io_schmitt_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2888.360 3174.000 2888.740 ;
    END
  END mprj_io_schmitt_sel[10]
  PIN mprj_io_schmitt_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3103.360 3174.000 3103.740 ;
    END
  END mprj_io_schmitt_sel[11]
  PIN mprj_io_schmitt_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3318.360 3174.000 3318.740 ;
    END
  END mprj_io_schmitt_sel[12]
  PIN mprj_io_schmitt_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3748.360 3174.000 3748.740 ;
    END
  END mprj_io_schmitt_sel[13]
  PIN mprj_io_schmitt_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 4178.360 3174.000 4178.740 ;
    END
  END mprj_io_schmitt_sel[14]
  PIN mprj_io_schmitt_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2986.260 4356.000 2986.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[15]
  PIN mprj_io_schmitt_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2436.260 4356.000 2436.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[16]
  PIN mprj_io_schmitt_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2161.260 4356.000 2161.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[17]
  PIN mprj_io_schmitt_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1886.260 4356.000 1886.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[18]
  PIN mprj_io_schmitt_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1336.260 4356.000 1336.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[19]
  PIN mprj_io_schmitt_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 308.360 3174.000 308.740 ;
    END
  END mprj_io_schmitt_sel[1]
  PIN mprj_io_schmitt_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1061.260 4356.000 1061.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[20]
  PIN mprj_io_schmitt_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 786.260 4356.000 786.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[21]
  PIN mprj_io_schmitt_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 511.260 4356.000 511.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[22]
  PIN mprj_io_schmitt_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 236.260 4356.000 236.640 4364.000 ;
    END
  END mprj_io_schmitt_sel[23]
  PIN mprj_io_schmitt_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 4241.260 4.000 4241.640 ;
    END
  END mprj_io_schmitt_sel[24]
  PIN mprj_io_schmitt_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3421.260 4.000 3421.640 ;
    END
  END mprj_io_schmitt_sel[25]
  PIN mprj_io_schmitt_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3216.260 4.000 3216.640 ;
    END
  END mprj_io_schmitt_sel[26]
  PIN mprj_io_schmitt_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3011.260 4.000 3011.640 ;
    END
  END mprj_io_schmitt_sel[27]
  PIN mprj_io_schmitt_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2806.260 4.000 2806.640 ;
    END
  END mprj_io_schmitt_sel[28]
  PIN mprj_io_schmitt_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2601.260 4.000 2601.640 ;
    END
  END mprj_io_schmitt_sel[29]
  PIN mprj_io_schmitt_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 523.360 3174.000 523.740 ;
    END
  END mprj_io_schmitt_sel[2]
  PIN mprj_io_schmitt_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2396.260 4.000 2396.640 ;
    END
  END mprj_io_schmitt_sel[30]
  PIN mprj_io_schmitt_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2191.260 4.000 2191.640 ;
    END
  END mprj_io_schmitt_sel[31]
  PIN mprj_io_schmitt_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1576.260 4.000 1576.640 ;
    END
  END mprj_io_schmitt_sel[32]
  PIN mprj_io_schmitt_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1371.260 4.000 1371.640 ;
    END
  END mprj_io_schmitt_sel[33]
  PIN mprj_io_schmitt_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1166.260 4.000 1166.640 ;
    END
  END mprj_io_schmitt_sel[34]
  PIN mprj_io_schmitt_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 961.260 4.000 961.640 ;
    END
  END mprj_io_schmitt_sel[35]
  PIN mprj_io_schmitt_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 756.260 4.000 756.640 ;
    END
  END mprj_io_schmitt_sel[36]
  PIN mprj_io_schmitt_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 551.260 4.000 551.640 ;
    END
  END mprj_io_schmitt_sel[37]
  PIN mprj_io_schmitt_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 738.360 3174.000 738.740 ;
    END
  END mprj_io_schmitt_sel[3]
  PIN mprj_io_schmitt_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 953.360 3174.000 953.740 ;
    END
  END mprj_io_schmitt_sel[4]
  PIN mprj_io_schmitt_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1168.360 3174.000 1168.740 ;
    END
  END mprj_io_schmitt_sel[5]
  PIN mprj_io_schmitt_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1383.360 3174.000 1383.740 ;
    END
  END mprj_io_schmitt_sel[6]
  PIN mprj_io_schmitt_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2243.360 3174.000 2243.740 ;
    END
  END mprj_io_schmitt_sel[7]
  PIN mprj_io_schmitt_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2458.360 3174.000 2458.740 ;
    END
  END mprj_io_schmitt_sel[8]
  PIN mprj_io_schmitt_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2673.360 3174.000 2673.740 ;
    END
  END mprj_io_schmitt_sel[9]
  PIN mprj_io_slew_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 158.670 3174.000 159.050 ;
    END
  END mprj_io_slew_sel[0]
  PIN mprj_io_slew_sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2953.670 3174.000 2954.050 ;
    END
  END mprj_io_slew_sel[10]
  PIN mprj_io_slew_sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3168.670 3174.000 3169.050 ;
    END
  END mprj_io_slew_sel[11]
  PIN mprj_io_slew_sel[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3383.670 3174.000 3384.050 ;
    END
  END mprj_io_slew_sel[12]
  PIN mprj_io_slew_sel[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 3813.670 3174.000 3814.050 ;
    END
  END mprj_io_slew_sel[13]
  PIN mprj_io_slew_sel[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 4243.670 3174.000 4244.050 ;
    END
  END mprj_io_slew_sel[14]
  PIN mprj_io_slew_sel[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2920.950 4356.000 2921.330 4364.000 ;
    END
  END mprj_io_slew_sel[15]
  PIN mprj_io_slew_sel[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2370.950 4356.000 2371.330 4364.000 ;
    END
  END mprj_io_slew_sel[16]
  PIN mprj_io_slew_sel[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2095.950 4356.000 2096.330 4364.000 ;
    END
  END mprj_io_slew_sel[17]
  PIN mprj_io_slew_sel[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1820.950 4356.000 1821.330 4364.000 ;
    END
  END mprj_io_slew_sel[18]
  PIN mprj_io_slew_sel[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1270.950 4356.000 1271.330 4364.000 ;
    END
  END mprj_io_slew_sel[19]
  PIN mprj_io_slew_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 373.670 3174.000 374.050 ;
    END
  END mprj_io_slew_sel[1]
  PIN mprj_io_slew_sel[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 995.950 4356.000 996.330 4364.000 ;
    END
  END mprj_io_slew_sel[20]
  PIN mprj_io_slew_sel[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 720.950 4356.000 721.330 4364.000 ;
    END
  END mprj_io_slew_sel[21]
  PIN mprj_io_slew_sel[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 445.950 4356.000 446.330 4364.000 ;
    END
  END mprj_io_slew_sel[22]
  PIN mprj_io_slew_sel[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 170.950 4356.000 171.330 4364.000 ;
    END
  END mprj_io_slew_sel[23]
  PIN mprj_io_slew_sel[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 4175.950 4.000 4176.330 ;
    END
  END mprj_io_slew_sel[24]
  PIN mprj_io_slew_sel[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3355.950 4.000 3356.330 ;
    END
  END mprj_io_slew_sel[25]
  PIN mprj_io_slew_sel[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 3150.950 4.000 3151.330 ;
    END
  END mprj_io_slew_sel[26]
  PIN mprj_io_slew_sel[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2945.950 4.000 2946.330 ;
    END
  END mprj_io_slew_sel[27]
  PIN mprj_io_slew_sel[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2740.950 4.000 2741.330 ;
    END
  END mprj_io_slew_sel[28]
  PIN mprj_io_slew_sel[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2535.950 4.000 2536.330 ;
    END
  END mprj_io_slew_sel[29]
  PIN mprj_io_slew_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 588.670 3174.000 589.050 ;
    END
  END mprj_io_slew_sel[2]
  PIN mprj_io_slew_sel[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2330.950 4.000 2331.330 ;
    END
  END mprj_io_slew_sel[30]
  PIN mprj_io_slew_sel[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 2125.950 4.000 2126.330 ;
    END
  END mprj_io_slew_sel[31]
  PIN mprj_io_slew_sel[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1510.950 4.000 1511.330 ;
    END
  END mprj_io_slew_sel[32]
  PIN mprj_io_slew_sel[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1305.950 4.000 1306.330 ;
    END
  END mprj_io_slew_sel[33]
  PIN mprj_io_slew_sel[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 1100.950 4.000 1101.330 ;
    END
  END mprj_io_slew_sel[34]
  PIN mprj_io_slew_sel[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 895.950 4.000 896.330 ;
    END
  END mprj_io_slew_sel[35]
  PIN mprj_io_slew_sel[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 690.950 4.000 691.330 ;
    END
  END mprj_io_slew_sel[36]
  PIN mprj_io_slew_sel[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT -4.000 485.950 4.000 486.330 ;
    END
  END mprj_io_slew_sel[37]
  PIN mprj_io_slew_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 803.670 3174.000 804.050 ;
    END
  END mprj_io_slew_sel[3]
  PIN mprj_io_slew_sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1018.670 3174.000 1019.050 ;
    END
  END mprj_io_slew_sel[4]
  PIN mprj_io_slew_sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1233.670 3174.000 1234.050 ;
    END
  END mprj_io_slew_sel[5]
  PIN mprj_io_slew_sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 1448.670 3174.000 1449.050 ;
    END
  END mprj_io_slew_sel[6]
  PIN mprj_io_slew_sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2308.670 3174.000 2309.050 ;
    END
  END mprj_io_slew_sel[7]
  PIN mprj_io_slew_sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2523.670 3174.000 2524.050 ;
    END
  END mprj_io_slew_sel[8]
  PIN mprj_io_slew_sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 3166.000 2738.670 3174.000 2739.050 ;
    END
  END mprj_io_slew_sel[9]
  PIN rstb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 515.860 -4.000 516.240 4.000 ;
    END
  END rstb
  OBS
      LAYER Metal1 ;
        RECT 22.490 26.470 3151.030 4353.850 ;
      LAYER Metal2 ;
        RECT 6.300 4355.700 168.460 4356.660 ;
        RECT 171.630 4355.700 227.935 4356.660 ;
        RECT 228.915 4355.700 228.990 4356.660 ;
        RECT 229.970 4355.700 231.500 4356.660 ;
        RECT 233.190 4355.700 233.355 4356.660 ;
        RECT 234.335 4355.700 235.960 4356.660 ;
        RECT 236.940 4355.700 443.460 4356.660 ;
        RECT 446.630 4355.700 502.935 4356.660 ;
        RECT 503.915 4355.700 503.990 4356.660 ;
        RECT 504.970 4355.700 506.500 4356.660 ;
        RECT 508.190 4355.700 508.355 4356.660 ;
        RECT 509.335 4355.700 510.960 4356.660 ;
        RECT 511.940 4355.700 718.460 4356.660 ;
        RECT 721.630 4355.700 777.935 4356.660 ;
        RECT 778.915 4355.700 778.990 4356.660 ;
        RECT 779.970 4355.700 781.500 4356.660 ;
        RECT 783.190 4355.700 783.355 4356.660 ;
        RECT 784.335 4355.700 785.960 4356.660 ;
        RECT 786.940 4355.700 993.460 4356.660 ;
        RECT 996.630 4355.700 1052.935 4356.660 ;
        RECT 1053.915 4355.700 1053.990 4356.660 ;
        RECT 1054.970 4355.700 1056.500 4356.660 ;
        RECT 1058.190 4355.700 1058.355 4356.660 ;
        RECT 1059.335 4355.700 1060.960 4356.660 ;
        RECT 1061.940 4355.700 1268.460 4356.660 ;
        RECT 1271.630 4355.700 1327.935 4356.660 ;
        RECT 1328.915 4355.700 1328.990 4356.660 ;
        RECT 1329.970 4355.700 1331.500 4356.660 ;
        RECT 1333.190 4355.700 1333.355 4356.660 ;
        RECT 1334.335 4355.700 1335.960 4356.660 ;
        RECT 1336.940 4355.700 1818.460 4356.660 ;
        RECT 1821.630 4355.700 1877.935 4356.660 ;
        RECT 1878.915 4355.700 1878.990 4356.660 ;
        RECT 1879.970 4355.700 1881.500 4356.660 ;
        RECT 1883.190 4355.700 1883.355 4356.660 ;
        RECT 1884.335 4355.700 1885.960 4356.660 ;
        RECT 1886.940 4355.700 2093.460 4356.660 ;
        RECT 2096.630 4355.700 2152.935 4356.660 ;
        RECT 2153.915 4355.700 2153.990 4356.660 ;
        RECT 2154.970 4355.700 2156.500 4356.660 ;
        RECT 2158.190 4355.700 2158.355 4356.660 ;
        RECT 2159.335 4355.700 2160.960 4356.660 ;
        RECT 2161.940 4355.700 2368.460 4356.660 ;
        RECT 2371.630 4355.700 2427.935 4356.660 ;
        RECT 2428.915 4355.700 2428.990 4356.660 ;
        RECT 2429.970 4355.700 2431.500 4356.660 ;
        RECT 2433.190 4355.700 2433.355 4356.660 ;
        RECT 2434.335 4355.700 2435.960 4356.660 ;
        RECT 2436.940 4355.700 2918.460 4356.660 ;
        RECT 2921.630 4355.700 2977.935 4356.660 ;
        RECT 2978.915 4355.700 2978.990 4356.660 ;
        RECT 2979.970 4355.700 2981.500 4356.660 ;
        RECT 2983.190 4355.700 2983.355 4356.660 ;
        RECT 2984.335 4355.700 2985.960 4356.660 ;
        RECT 2986.940 4355.700 3164.420 4356.660 ;
        RECT 6.300 4.300 3164.420 4355.700 ;
        RECT 6.300 3.500 450.665 4.300 ;
        RECT 451.645 3.500 455.030 4.300 ;
        RECT 456.010 3.500 515.560 4.300 ;
        RECT 516.540 3.500 725.665 4.300 ;
        RECT 726.645 3.500 790.560 4.300 ;
        RECT 791.540 3.500 1275.665 4.300 ;
        RECT 1276.645 3.500 1338.365 4.300 ;
        RECT 1340.810 3.500 1613.370 4.300 ;
        RECT 1615.810 3.500 1831.085 4.300 ;
        RECT 1832.065 3.500 1888.370 4.300 ;
        RECT 1891.535 3.500 2106.085 4.300 ;
        RECT 2107.065 3.500 2163.370 4.300 ;
        RECT 2166.540 3.500 2373.060 4.300 ;
        RECT 2374.040 3.500 2375.665 4.300 ;
        RECT 2376.645 3.500 2376.810 4.300 ;
        RECT 2378.500 3.500 2380.030 4.300 ;
        RECT 2381.010 3.500 2381.085 4.300 ;
        RECT 2382.065 3.500 2438.370 4.300 ;
        RECT 2441.540 3.500 3164.420 4.300 ;
      LAYER Metal3 ;
        RECT 1.210 4246.540 3168.390 4354.420 ;
        RECT 1.210 4243.370 3165.700 4246.540 ;
        RECT 1.210 4241.940 3168.390 4243.370 ;
        RECT 4.300 4240.960 3168.390 4241.940 ;
        RECT 1.210 4239.335 3168.390 4240.960 ;
        RECT 4.300 4238.355 3168.390 4239.335 ;
        RECT 1.210 4238.190 3168.390 4238.355 ;
        RECT 4.300 4236.500 3168.390 4238.190 ;
        RECT 1.210 4234.970 3168.390 4236.500 ;
        RECT 4.300 4233.990 3168.390 4234.970 ;
        RECT 1.210 4233.915 3168.390 4233.990 ;
        RECT 4.300 4232.935 3168.390 4233.915 ;
        RECT 1.210 4187.065 3168.390 4232.935 ;
        RECT 1.210 4186.085 3165.700 4187.065 ;
        RECT 1.210 4186.010 3168.390 4186.085 ;
        RECT 1.210 4185.030 3165.700 4186.010 ;
        RECT 1.210 4183.500 3168.390 4185.030 ;
        RECT 1.210 4181.810 3165.700 4183.500 ;
        RECT 1.210 4181.645 3168.390 4181.810 ;
        RECT 1.210 4180.665 3165.700 4181.645 ;
        RECT 1.210 4179.040 3168.390 4180.665 ;
        RECT 1.210 4178.060 3165.700 4179.040 ;
        RECT 1.210 4176.630 3168.390 4178.060 ;
        RECT 4.300 4173.460 3168.390 4176.630 ;
        RECT 1.210 3816.540 3168.390 4173.460 ;
        RECT 1.210 3813.370 3165.700 3816.540 ;
        RECT 1.210 3757.065 3168.390 3813.370 ;
        RECT 1.210 3756.085 3165.700 3757.065 ;
        RECT 1.210 3756.010 3168.390 3756.085 ;
        RECT 1.210 3755.030 3165.700 3756.010 ;
        RECT 1.210 3753.500 3168.390 3755.030 ;
        RECT 1.210 3751.810 3165.700 3753.500 ;
        RECT 1.210 3751.645 3168.390 3751.810 ;
        RECT 1.210 3750.665 3165.700 3751.645 ;
        RECT 1.210 3749.040 3168.390 3750.665 ;
        RECT 1.210 3748.060 3165.700 3749.040 ;
        RECT 1.210 3421.940 3168.390 3748.060 ;
        RECT 4.300 3420.960 3168.390 3421.940 ;
        RECT 1.210 3419.335 3168.390 3420.960 ;
        RECT 4.300 3418.355 3168.390 3419.335 ;
        RECT 1.210 3418.190 3168.390 3418.355 ;
        RECT 4.300 3416.500 3168.390 3418.190 ;
        RECT 1.210 3414.970 3168.390 3416.500 ;
        RECT 4.300 3413.990 3168.390 3414.970 ;
        RECT 1.210 3413.915 3168.390 3413.990 ;
        RECT 4.300 3412.935 3168.390 3413.915 ;
        RECT 1.210 3386.540 3168.390 3412.935 ;
        RECT 1.210 3383.370 3165.700 3386.540 ;
        RECT 1.210 3356.630 3168.390 3383.370 ;
        RECT 4.300 3353.460 3168.390 3356.630 ;
        RECT 1.210 3327.065 3168.390 3353.460 ;
        RECT 1.210 3326.085 3165.700 3327.065 ;
        RECT 1.210 3326.010 3168.390 3326.085 ;
        RECT 1.210 3325.030 3165.700 3326.010 ;
        RECT 1.210 3323.500 3168.390 3325.030 ;
        RECT 1.210 3321.810 3165.700 3323.500 ;
        RECT 1.210 3321.645 3168.390 3321.810 ;
        RECT 1.210 3320.665 3165.700 3321.645 ;
        RECT 1.210 3319.040 3168.390 3320.665 ;
        RECT 1.210 3318.060 3165.700 3319.040 ;
        RECT 1.210 3216.940 3168.390 3318.060 ;
        RECT 4.300 3215.960 3168.390 3216.940 ;
        RECT 1.210 3214.335 3168.390 3215.960 ;
        RECT 4.300 3213.355 3168.390 3214.335 ;
        RECT 1.210 3213.190 3168.390 3213.355 ;
        RECT 4.300 3211.500 3168.390 3213.190 ;
        RECT 1.210 3209.970 3168.390 3211.500 ;
        RECT 4.300 3208.990 3168.390 3209.970 ;
        RECT 1.210 3208.915 3168.390 3208.990 ;
        RECT 4.300 3207.935 3168.390 3208.915 ;
        RECT 1.210 3171.540 3168.390 3207.935 ;
        RECT 1.210 3168.370 3165.700 3171.540 ;
        RECT 1.210 3151.630 3168.390 3168.370 ;
        RECT 4.300 3148.460 3168.390 3151.630 ;
        RECT 1.210 3112.065 3168.390 3148.460 ;
        RECT 1.210 3111.085 3165.700 3112.065 ;
        RECT 1.210 3111.010 3168.390 3111.085 ;
        RECT 1.210 3110.030 3165.700 3111.010 ;
        RECT 1.210 3108.500 3168.390 3110.030 ;
        RECT 1.210 3106.810 3165.700 3108.500 ;
        RECT 1.210 3106.645 3168.390 3106.810 ;
        RECT 1.210 3105.665 3165.700 3106.645 ;
        RECT 1.210 3104.040 3168.390 3105.665 ;
        RECT 1.210 3103.060 3165.700 3104.040 ;
        RECT 1.210 3011.940 3168.390 3103.060 ;
        RECT 4.300 3010.960 3168.390 3011.940 ;
        RECT 1.210 3009.335 3168.390 3010.960 ;
        RECT 4.300 3008.355 3168.390 3009.335 ;
        RECT 1.210 3008.190 3168.390 3008.355 ;
        RECT 4.300 3006.500 3168.390 3008.190 ;
        RECT 1.210 3004.970 3168.390 3006.500 ;
        RECT 4.300 3003.990 3168.390 3004.970 ;
        RECT 1.210 3003.915 3168.390 3003.990 ;
        RECT 4.300 3002.935 3168.390 3003.915 ;
        RECT 1.210 2956.540 3168.390 3002.935 ;
        RECT 1.210 2953.370 3165.700 2956.540 ;
        RECT 1.210 2946.630 3168.390 2953.370 ;
        RECT 4.300 2943.460 3168.390 2946.630 ;
        RECT 1.210 2897.065 3168.390 2943.460 ;
        RECT 1.210 2896.085 3165.700 2897.065 ;
        RECT 1.210 2896.010 3168.390 2896.085 ;
        RECT 1.210 2895.030 3165.700 2896.010 ;
        RECT 1.210 2893.500 3168.390 2895.030 ;
        RECT 1.210 2891.810 3165.700 2893.500 ;
        RECT 1.210 2891.645 3168.390 2891.810 ;
        RECT 1.210 2890.665 3165.700 2891.645 ;
        RECT 1.210 2889.040 3168.390 2890.665 ;
        RECT 1.210 2888.060 3165.700 2889.040 ;
        RECT 1.210 2806.940 3168.390 2888.060 ;
        RECT 4.300 2805.960 3168.390 2806.940 ;
        RECT 1.210 2804.335 3168.390 2805.960 ;
        RECT 4.300 2803.355 3168.390 2804.335 ;
        RECT 1.210 2803.190 3168.390 2803.355 ;
        RECT 4.300 2801.500 3168.390 2803.190 ;
        RECT 1.210 2799.970 3168.390 2801.500 ;
        RECT 4.300 2798.990 3168.390 2799.970 ;
        RECT 1.210 2798.915 3168.390 2798.990 ;
        RECT 4.300 2797.935 3168.390 2798.915 ;
        RECT 1.210 2741.630 3168.390 2797.935 ;
        RECT 4.300 2741.540 3168.390 2741.630 ;
        RECT 4.300 2738.460 3165.700 2741.540 ;
        RECT 1.210 2738.370 3165.700 2738.460 ;
        RECT 1.210 2682.065 3168.390 2738.370 ;
        RECT 1.210 2681.085 3165.700 2682.065 ;
        RECT 1.210 2681.010 3168.390 2681.085 ;
        RECT 1.210 2680.030 3165.700 2681.010 ;
        RECT 1.210 2678.500 3168.390 2680.030 ;
        RECT 1.210 2676.810 3165.700 2678.500 ;
        RECT 1.210 2676.645 3168.390 2676.810 ;
        RECT 1.210 2675.665 3165.700 2676.645 ;
        RECT 1.210 2674.040 3168.390 2675.665 ;
        RECT 1.210 2673.060 3165.700 2674.040 ;
        RECT 1.210 2601.940 3168.390 2673.060 ;
        RECT 4.300 2600.960 3168.390 2601.940 ;
        RECT 1.210 2599.335 3168.390 2600.960 ;
        RECT 4.300 2598.355 3168.390 2599.335 ;
        RECT 1.210 2598.190 3168.390 2598.355 ;
        RECT 4.300 2596.500 3168.390 2598.190 ;
        RECT 1.210 2594.970 3168.390 2596.500 ;
        RECT 4.300 2593.990 3168.390 2594.970 ;
        RECT 1.210 2593.915 3168.390 2593.990 ;
        RECT 4.300 2592.935 3168.390 2593.915 ;
        RECT 1.210 2536.630 3168.390 2592.935 ;
        RECT 4.300 2533.460 3168.390 2536.630 ;
        RECT 1.210 2526.540 3168.390 2533.460 ;
        RECT 1.210 2523.370 3165.700 2526.540 ;
        RECT 1.210 2467.065 3168.390 2523.370 ;
        RECT 1.210 2466.085 3165.700 2467.065 ;
        RECT 1.210 2466.010 3168.390 2466.085 ;
        RECT 1.210 2465.030 3165.700 2466.010 ;
        RECT 1.210 2463.500 3168.390 2465.030 ;
        RECT 1.210 2461.810 3165.700 2463.500 ;
        RECT 1.210 2461.645 3168.390 2461.810 ;
        RECT 1.210 2460.665 3165.700 2461.645 ;
        RECT 1.210 2459.040 3168.390 2460.665 ;
        RECT 1.210 2458.060 3165.700 2459.040 ;
        RECT 1.210 2396.940 3168.390 2458.060 ;
        RECT 4.300 2395.960 3168.390 2396.940 ;
        RECT 1.210 2394.335 3168.390 2395.960 ;
        RECT 4.300 2393.355 3168.390 2394.335 ;
        RECT 1.210 2393.190 3168.390 2393.355 ;
        RECT 4.300 2391.500 3168.390 2393.190 ;
        RECT 1.210 2389.970 3168.390 2391.500 ;
        RECT 4.300 2388.990 3168.390 2389.970 ;
        RECT 1.210 2388.915 3168.390 2388.990 ;
        RECT 4.300 2387.935 3168.390 2388.915 ;
        RECT 1.210 2331.630 3168.390 2387.935 ;
        RECT 4.300 2328.460 3168.390 2331.630 ;
        RECT 1.210 2311.540 3168.390 2328.460 ;
        RECT 1.210 2308.370 3165.700 2311.540 ;
        RECT 1.210 2252.065 3168.390 2308.370 ;
        RECT 1.210 2251.085 3165.700 2252.065 ;
        RECT 1.210 2251.010 3168.390 2251.085 ;
        RECT 1.210 2250.030 3165.700 2251.010 ;
        RECT 1.210 2248.500 3168.390 2250.030 ;
        RECT 1.210 2246.810 3165.700 2248.500 ;
        RECT 1.210 2246.645 3168.390 2246.810 ;
        RECT 1.210 2245.665 3165.700 2246.645 ;
        RECT 1.210 2244.040 3168.390 2245.665 ;
        RECT 1.210 2243.060 3165.700 2244.040 ;
        RECT 1.210 2191.940 3168.390 2243.060 ;
        RECT 4.300 2190.960 3168.390 2191.940 ;
        RECT 1.210 2189.335 3168.390 2190.960 ;
        RECT 4.300 2188.355 3168.390 2189.335 ;
        RECT 1.210 2188.190 3168.390 2188.355 ;
        RECT 4.300 2186.500 3168.390 2188.190 ;
        RECT 1.210 2184.970 3168.390 2186.500 ;
        RECT 4.300 2183.990 3168.390 2184.970 ;
        RECT 1.210 2183.915 3168.390 2183.990 ;
        RECT 4.300 2182.935 3168.390 2183.915 ;
        RECT 1.210 2126.630 3168.390 2182.935 ;
        RECT 4.300 2123.460 3168.390 2126.630 ;
        RECT 1.210 1576.940 3168.390 2123.460 ;
        RECT 4.300 1575.960 3168.390 1576.940 ;
        RECT 1.210 1574.335 3168.390 1575.960 ;
        RECT 4.300 1573.355 3168.390 1574.335 ;
        RECT 1.210 1573.190 3168.390 1573.355 ;
        RECT 4.300 1571.500 3168.390 1573.190 ;
        RECT 1.210 1569.970 3168.390 1571.500 ;
        RECT 4.300 1568.990 3168.390 1569.970 ;
        RECT 1.210 1568.915 3168.390 1568.990 ;
        RECT 4.300 1567.935 3168.390 1568.915 ;
        RECT 1.210 1511.630 3168.390 1567.935 ;
        RECT 4.300 1508.460 3168.390 1511.630 ;
        RECT 1.210 1451.540 3168.390 1508.460 ;
        RECT 1.210 1448.370 3165.700 1451.540 ;
        RECT 1.210 1392.065 3168.390 1448.370 ;
        RECT 1.210 1391.085 3165.700 1392.065 ;
        RECT 1.210 1391.010 3168.390 1391.085 ;
        RECT 1.210 1390.030 3165.700 1391.010 ;
        RECT 1.210 1388.500 3168.390 1390.030 ;
        RECT 1.210 1386.810 3165.700 1388.500 ;
        RECT 1.210 1386.645 3168.390 1386.810 ;
        RECT 1.210 1385.665 3165.700 1386.645 ;
        RECT 1.210 1384.040 3168.390 1385.665 ;
        RECT 1.210 1383.060 3165.700 1384.040 ;
        RECT 1.210 1371.940 3168.390 1383.060 ;
        RECT 4.300 1370.960 3168.390 1371.940 ;
        RECT 1.210 1369.335 3168.390 1370.960 ;
        RECT 4.300 1368.355 3168.390 1369.335 ;
        RECT 1.210 1368.190 3168.390 1368.355 ;
        RECT 4.300 1366.500 3168.390 1368.190 ;
        RECT 1.210 1364.970 3168.390 1366.500 ;
        RECT 4.300 1363.990 3168.390 1364.970 ;
        RECT 1.210 1363.915 3168.390 1363.990 ;
        RECT 4.300 1362.935 3168.390 1363.915 ;
        RECT 1.210 1306.630 3168.390 1362.935 ;
        RECT 4.300 1303.460 3168.390 1306.630 ;
        RECT 1.210 1236.540 3168.390 1303.460 ;
        RECT 1.210 1233.370 3165.700 1236.540 ;
        RECT 1.210 1177.065 3168.390 1233.370 ;
        RECT 1.210 1176.085 3165.700 1177.065 ;
        RECT 1.210 1176.010 3168.390 1176.085 ;
        RECT 1.210 1175.030 3165.700 1176.010 ;
        RECT 1.210 1173.500 3168.390 1175.030 ;
        RECT 1.210 1171.810 3165.700 1173.500 ;
        RECT 1.210 1171.645 3168.390 1171.810 ;
        RECT 1.210 1170.665 3165.700 1171.645 ;
        RECT 1.210 1169.040 3168.390 1170.665 ;
        RECT 1.210 1168.060 3165.700 1169.040 ;
        RECT 1.210 1166.940 3168.390 1168.060 ;
        RECT 4.300 1165.960 3168.390 1166.940 ;
        RECT 1.210 1164.335 3168.390 1165.960 ;
        RECT 4.300 1163.355 3168.390 1164.335 ;
        RECT 1.210 1163.190 3168.390 1163.355 ;
        RECT 4.300 1161.500 3168.390 1163.190 ;
        RECT 1.210 1159.970 3168.390 1161.500 ;
        RECT 4.300 1158.990 3168.390 1159.970 ;
        RECT 1.210 1158.915 3168.390 1158.990 ;
        RECT 4.300 1157.935 3168.390 1158.915 ;
        RECT 1.210 1101.630 3168.390 1157.935 ;
        RECT 4.300 1098.460 3168.390 1101.630 ;
        RECT 1.210 1021.540 3168.390 1098.460 ;
        RECT 1.210 1018.370 3165.700 1021.540 ;
        RECT 1.210 962.065 3168.390 1018.370 ;
        RECT 1.210 961.940 3165.700 962.065 ;
        RECT 4.300 961.085 3165.700 961.940 ;
        RECT 4.300 961.010 3168.390 961.085 ;
        RECT 4.300 960.960 3165.700 961.010 ;
        RECT 1.210 960.030 3165.700 960.960 ;
        RECT 1.210 959.335 3168.390 960.030 ;
        RECT 4.300 958.500 3168.390 959.335 ;
        RECT 4.300 958.355 3165.700 958.500 ;
        RECT 1.210 958.190 3165.700 958.355 ;
        RECT 4.300 956.810 3165.700 958.190 ;
        RECT 4.300 956.645 3168.390 956.810 ;
        RECT 4.300 956.500 3165.700 956.645 ;
        RECT 1.210 955.665 3165.700 956.500 ;
        RECT 1.210 954.970 3168.390 955.665 ;
        RECT 4.300 954.040 3168.390 954.970 ;
        RECT 4.300 953.990 3165.700 954.040 ;
        RECT 1.210 953.915 3165.700 953.990 ;
        RECT 4.300 953.060 3165.700 953.915 ;
        RECT 4.300 952.935 3168.390 953.060 ;
        RECT 1.210 896.630 3168.390 952.935 ;
        RECT 4.300 893.460 3168.390 896.630 ;
        RECT 1.210 806.540 3168.390 893.460 ;
        RECT 1.210 803.370 3165.700 806.540 ;
        RECT 1.210 756.940 3168.390 803.370 ;
        RECT 4.300 755.960 3168.390 756.940 ;
        RECT 1.210 754.335 3168.390 755.960 ;
        RECT 4.300 753.355 3168.390 754.335 ;
        RECT 1.210 753.190 3168.390 753.355 ;
        RECT 4.300 751.500 3168.390 753.190 ;
        RECT 1.210 749.970 3168.390 751.500 ;
        RECT 4.300 748.990 3168.390 749.970 ;
        RECT 1.210 748.915 3168.390 748.990 ;
        RECT 4.300 747.935 3168.390 748.915 ;
        RECT 1.210 747.065 3168.390 747.935 ;
        RECT 1.210 746.085 3165.700 747.065 ;
        RECT 1.210 746.010 3168.390 746.085 ;
        RECT 1.210 745.030 3165.700 746.010 ;
        RECT 1.210 743.500 3168.390 745.030 ;
        RECT 1.210 741.810 3165.700 743.500 ;
        RECT 1.210 741.645 3168.390 741.810 ;
        RECT 1.210 740.665 3165.700 741.645 ;
        RECT 1.210 739.040 3168.390 740.665 ;
        RECT 1.210 738.060 3165.700 739.040 ;
        RECT 1.210 691.630 3168.390 738.060 ;
        RECT 4.300 688.460 3168.390 691.630 ;
        RECT 1.210 591.540 3168.390 688.460 ;
        RECT 1.210 588.370 3165.700 591.540 ;
        RECT 1.210 551.940 3168.390 588.370 ;
        RECT 4.300 550.960 3168.390 551.940 ;
        RECT 1.210 549.335 3168.390 550.960 ;
        RECT 4.300 548.355 3168.390 549.335 ;
        RECT 1.210 548.190 3168.390 548.355 ;
        RECT 4.300 546.500 3168.390 548.190 ;
        RECT 1.210 544.970 3168.390 546.500 ;
        RECT 4.300 543.990 3168.390 544.970 ;
        RECT 1.210 543.915 3168.390 543.990 ;
        RECT 4.300 542.935 3168.390 543.915 ;
        RECT 1.210 532.065 3168.390 542.935 ;
        RECT 1.210 531.085 3165.700 532.065 ;
        RECT 1.210 531.010 3168.390 531.085 ;
        RECT 1.210 530.030 3165.700 531.010 ;
        RECT 1.210 528.500 3168.390 530.030 ;
        RECT 1.210 526.810 3165.700 528.500 ;
        RECT 1.210 526.645 3168.390 526.810 ;
        RECT 1.210 525.665 3165.700 526.645 ;
        RECT 1.210 524.040 3168.390 525.665 ;
        RECT 1.210 523.060 3165.700 524.040 ;
        RECT 1.210 486.630 3168.390 523.060 ;
        RECT 4.300 483.460 3168.390 486.630 ;
        RECT 1.210 376.540 3168.390 483.460 ;
        RECT 1.210 373.370 3165.700 376.540 ;
        RECT 1.210 317.065 3168.390 373.370 ;
        RECT 1.210 316.085 3165.700 317.065 ;
        RECT 1.210 316.010 3168.390 316.085 ;
        RECT 1.210 315.030 3165.700 316.010 ;
        RECT 1.210 313.500 3168.390 315.030 ;
        RECT 1.210 311.810 3165.700 313.500 ;
        RECT 1.210 311.645 3168.390 311.810 ;
        RECT 1.210 310.665 3165.700 311.645 ;
        RECT 1.210 309.040 3168.390 310.665 ;
        RECT 1.210 308.060 3165.700 309.040 ;
        RECT 1.210 161.540 3168.390 308.060 ;
        RECT 1.210 158.370 3165.700 161.540 ;
        RECT 1.210 102.065 3168.390 158.370 ;
        RECT 1.210 101.085 3165.700 102.065 ;
        RECT 1.210 101.010 3168.390 101.085 ;
        RECT 1.210 100.030 3165.700 101.010 ;
        RECT 1.210 98.500 3168.390 100.030 ;
        RECT 1.210 96.810 3165.700 98.500 ;
        RECT 1.210 96.645 3168.390 96.810 ;
        RECT 1.210 95.665 3165.700 96.645 ;
        RECT 1.210 94.040 3168.390 95.665 ;
        RECT 1.210 93.060 3165.700 94.040 ;
        RECT 1.210 25.340 3168.390 93.060 ;
      LAYER Metal4 ;
        RECT 1.260 33.690 1.780 4332.630 ;
        RECT 12.380 33.690 13.780 4332.630 ;
        RECT 24.380 33.690 35.780 4332.630 ;
        RECT 39.380 33.690 44.780 4332.630 ;
        RECT 48.380 33.690 60.640 4332.630 ;
        RECT 64.240 33.690 69.640 4332.630 ;
        RECT 73.240 4282.580 105.780 4332.630 ;
        RECT 109.380 4282.580 127.780 4332.630 ;
        RECT 131.380 4282.580 185.780 4332.630 ;
        RECT 189.380 4282.580 207.780 4332.630 ;
        RECT 211.380 4282.580 265.780 4332.630 ;
        RECT 269.380 4282.580 287.780 4332.630 ;
        RECT 291.380 4282.580 306.280 4332.630 ;
        RECT 309.880 4282.580 313.280 4332.630 ;
        RECT 316.880 4282.580 345.780 4332.630 ;
        RECT 349.380 4282.580 367.780 4332.630 ;
        RECT 371.380 4282.580 425.780 4332.630 ;
        RECT 429.380 4282.580 447.780 4332.630 ;
        RECT 451.380 4282.580 505.780 4332.630 ;
        RECT 509.380 4282.580 527.780 4332.630 ;
        RECT 531.380 4282.580 555.980 4332.630 ;
        RECT 559.580 4282.580 562.980 4332.630 ;
        RECT 566.580 4282.580 585.780 4332.630 ;
        RECT 589.380 4282.580 607.780 4332.630 ;
        RECT 611.380 4282.580 665.780 4332.630 ;
        RECT 669.380 4282.580 687.780 4332.630 ;
        RECT 691.380 4282.580 745.780 4332.630 ;
        RECT 749.380 4282.580 767.780 4332.630 ;
        RECT 771.380 4282.580 825.780 4332.630 ;
        RECT 829.380 4282.580 847.780 4332.630 ;
        RECT 851.380 4282.580 864.480 4332.630 ;
        RECT 868.080 4282.580 871.480 4332.630 ;
        RECT 875.080 4282.580 905.780 4332.630 ;
        RECT 909.380 4282.580 927.780 4332.630 ;
        RECT 931.380 4282.580 985.780 4332.630 ;
        RECT 989.380 4282.580 1007.780 4332.630 ;
        RECT 1011.380 4282.580 1065.780 4332.630 ;
        RECT 1069.380 4282.580 1087.780 4332.630 ;
        RECT 1091.380 4282.580 1116.180 4332.630 ;
        RECT 1119.780 4282.580 1123.180 4332.630 ;
        RECT 1126.780 4282.580 1145.780 4332.630 ;
        RECT 1149.380 4282.580 1167.780 4332.630 ;
        RECT 1171.380 4282.580 1225.780 4332.630 ;
        RECT 1229.380 4282.580 1247.780 4332.630 ;
        RECT 1251.380 4282.580 1305.780 4332.630 ;
        RECT 1309.380 4282.580 1327.780 4332.630 ;
        RECT 1331.380 4282.580 1359.080 4332.630 ;
        RECT 1362.680 4282.580 1366.080 4332.630 ;
        RECT 1369.680 4282.580 1385.780 4332.630 ;
        RECT 1389.380 4282.580 1407.780 4332.630 ;
        RECT 1411.380 4282.580 1465.780 4332.630 ;
        RECT 1469.380 4282.580 1487.780 4332.630 ;
        RECT 1491.380 4282.580 1545.780 4332.630 ;
        RECT 1549.380 4282.580 1567.780 4332.630 ;
        RECT 1571.380 4282.580 1625.780 4332.630 ;
        RECT 1629.380 4282.580 1647.780 4332.630 ;
        RECT 1651.380 4282.580 1705.780 4332.630 ;
        RECT 1709.380 4282.580 1727.780 4332.630 ;
        RECT 1731.380 4282.580 1785.780 4332.630 ;
        RECT 1789.380 4282.580 1807.780 4332.630 ;
        RECT 1811.380 4282.580 1865.780 4332.630 ;
        RECT 1869.380 4282.580 1887.780 4332.630 ;
        RECT 1891.380 4282.580 1916.080 4332.630 ;
        RECT 1919.680 4282.580 1923.080 4332.630 ;
        RECT 1926.680 4282.580 1945.780 4332.630 ;
        RECT 1949.380 4282.580 1967.780 4332.630 ;
        RECT 1971.380 4282.580 2025.780 4332.630 ;
        RECT 2029.380 4282.580 2047.780 4332.630 ;
        RECT 2051.380 4282.580 2105.780 4332.630 ;
        RECT 2109.380 4282.580 2127.780 4332.630 ;
        RECT 2131.380 4282.580 2162.780 4332.630 ;
        RECT 2166.380 4282.580 2169.780 4332.630 ;
        RECT 2173.380 4282.580 2185.780 4332.630 ;
        RECT 2189.380 4282.580 2207.780 4332.630 ;
        RECT 2211.380 4282.580 2265.780 4332.630 ;
        RECT 2269.380 4282.580 2287.780 4332.630 ;
        RECT 2291.380 4282.580 2330.780 4332.630 ;
        RECT 2334.380 4282.580 2345.780 4332.630 ;
        RECT 2349.380 4282.580 2352.780 4332.630 ;
        RECT 2356.380 4282.580 2367.780 4332.630 ;
        RECT 2371.380 4282.580 2425.780 4332.630 ;
        RECT 2429.380 4282.580 2447.780 4332.630 ;
        RECT 2451.380 4282.580 2505.780 4332.630 ;
        RECT 2509.380 4282.580 2527.780 4332.630 ;
        RECT 2531.380 4282.580 2585.780 4332.630 ;
        RECT 2589.380 4282.580 2607.780 4332.630 ;
        RECT 2611.380 4282.580 2665.780 4332.630 ;
        RECT 2669.380 4282.580 2687.780 4332.630 ;
        RECT 2691.380 4282.580 2745.780 4332.630 ;
        RECT 2749.380 4282.580 2767.780 4332.630 ;
        RECT 2771.380 4282.580 2825.780 4332.630 ;
        RECT 2829.380 4282.580 2847.780 4332.630 ;
        RECT 2851.380 4282.580 2880.280 4332.630 ;
        RECT 2883.880 4282.580 2892.280 4332.630 ;
        RECT 2895.880 4282.580 2905.780 4332.630 ;
        RECT 2909.380 4282.580 2927.780 4332.630 ;
        RECT 2931.380 4282.580 2985.780 4332.630 ;
        RECT 2989.380 4282.580 3007.780 4332.630 ;
        RECT 3011.380 4282.580 3098.780 4332.630 ;
        RECT 73.240 1266.620 3098.780 4282.580 ;
        RECT 73.240 33.690 105.780 1266.620 ;
        RECT 109.380 33.690 127.780 1266.620 ;
        RECT 131.380 33.690 185.780 1266.620 ;
        RECT 189.380 33.690 207.780 1266.620 ;
        RECT 211.380 33.690 265.780 1266.620 ;
        RECT 269.380 33.690 287.780 1266.620 ;
        RECT 291.380 33.690 306.280 1266.620 ;
        RECT 309.880 33.690 313.280 1266.620 ;
        RECT 316.880 33.690 345.780 1266.620 ;
        RECT 349.380 33.690 367.780 1266.620 ;
        RECT 371.380 33.690 425.780 1266.620 ;
        RECT 429.380 33.690 447.780 1266.620 ;
        RECT 451.380 33.690 505.780 1266.620 ;
        RECT 509.380 33.690 527.780 1266.620 ;
        RECT 531.380 33.690 555.980 1266.620 ;
        RECT 559.580 33.690 562.980 1266.620 ;
        RECT 566.580 572.920 585.780 1266.620 ;
        RECT 569.920 62.120 585.780 572.920 ;
        RECT 566.580 33.690 585.780 62.120 ;
        RECT 589.380 33.690 607.780 1266.620 ;
        RECT 611.380 33.690 665.780 1266.620 ;
        RECT 669.380 33.690 687.780 1266.620 ;
        RECT 691.380 33.690 745.780 1266.620 ;
        RECT 749.380 33.690 767.780 1266.620 ;
        RECT 771.380 33.690 825.780 1266.620 ;
        RECT 829.380 33.690 847.780 1266.620 ;
        RECT 851.380 33.690 864.480 1266.620 ;
        RECT 868.080 33.690 871.480 1266.620 ;
        RECT 875.080 33.690 905.780 1266.620 ;
        RECT 909.380 33.690 927.780 1266.620 ;
        RECT 931.380 33.690 985.780 1266.620 ;
        RECT 989.380 33.690 1007.780 1266.620 ;
        RECT 1011.380 576.840 1065.780 1266.620 ;
        RECT 1011.380 58.200 1023.470 576.840 ;
        RECT 1025.570 58.200 1025.710 576.840 ;
        RECT 1027.810 58.200 1065.780 576.840 ;
        RECT 1011.380 33.690 1065.780 58.200 ;
        RECT 1069.380 33.690 1087.780 1266.620 ;
        RECT 1091.380 982.980 1116.180 1266.620 ;
        RECT 1119.780 982.980 1123.180 1266.620 ;
        RECT 1126.780 982.980 1145.780 1266.620 ;
        RECT 1091.380 892.020 1145.780 982.980 ;
        RECT 1091.380 33.690 1116.180 892.020 ;
        RECT 1119.780 33.690 1123.180 892.020 ;
        RECT 1126.780 33.690 1145.780 892.020 ;
        RECT 1149.380 33.690 1167.780 1266.620 ;
        RECT 1171.380 33.690 1225.780 1266.620 ;
        RECT 1229.380 33.690 1247.780 1266.620 ;
        RECT 1251.380 33.690 1305.780 1266.620 ;
        RECT 1309.380 33.690 1327.780 1266.620 ;
        RECT 1331.380 33.690 1359.080 1266.620 ;
        RECT 1362.680 33.690 1366.080 1266.620 ;
        RECT 1369.680 33.690 1385.780 1266.620 ;
        RECT 1389.380 33.690 1407.780 1266.620 ;
        RECT 1411.380 33.690 1465.780 1266.620 ;
        RECT 1469.380 576.840 1487.780 1266.620 ;
        RECT 1469.380 58.200 1480.430 576.840 ;
        RECT 1482.530 58.200 1482.670 576.840 ;
        RECT 1484.770 58.200 1487.780 576.840 ;
        RECT 1469.380 33.690 1487.780 58.200 ;
        RECT 1491.380 33.690 1545.780 1266.620 ;
        RECT 1549.380 33.690 1567.780 1266.620 ;
        RECT 1571.380 33.690 1625.780 1266.620 ;
        RECT 1629.380 33.690 1647.780 1266.620 ;
        RECT 1651.380 33.690 1705.780 1266.620 ;
        RECT 1709.380 33.690 1727.780 1266.620 ;
        RECT 1731.380 33.690 1785.780 1266.620 ;
        RECT 1789.380 33.690 1807.780 1266.620 ;
        RECT 1811.380 33.690 1865.780 1266.620 ;
        RECT 1869.380 33.690 1887.780 1266.620 ;
        RECT 1891.380 33.690 1916.080 1266.620 ;
        RECT 1919.680 33.690 1923.080 1266.620 ;
        RECT 1926.680 33.690 1945.780 1266.620 ;
        RECT 1949.380 33.690 1967.780 1266.620 ;
        RECT 1971.380 33.690 2025.780 1266.620 ;
        RECT 2029.380 33.690 2047.780 1266.620 ;
        RECT 2051.380 33.690 2105.780 1266.620 ;
        RECT 2109.380 33.690 2127.780 1266.620 ;
        RECT 2131.380 1122.980 2162.780 1266.620 ;
        RECT 2166.380 1122.980 2169.780 1266.620 ;
        RECT 2173.380 1122.980 2185.780 1266.620 ;
        RECT 2131.380 1032.020 2185.780 1122.980 ;
        RECT 2131.380 33.690 2162.780 1032.020 ;
        RECT 2166.380 33.690 2169.780 1032.020 ;
        RECT 2173.380 33.690 2185.780 1032.020 ;
        RECT 2189.380 33.690 2207.780 1266.620 ;
        RECT 2211.380 33.690 2265.780 1266.620 ;
        RECT 2269.380 33.690 2287.780 1266.620 ;
        RECT 2291.380 33.690 2330.780 1266.620 ;
        RECT 2334.380 33.690 2345.780 1266.620 ;
        RECT 2349.380 33.690 2352.780 1266.620 ;
        RECT 2356.380 33.690 2367.780 1266.620 ;
        RECT 2371.380 33.690 2425.780 1266.620 ;
        RECT 2429.380 33.690 2447.780 1266.620 ;
        RECT 2451.380 33.690 2505.780 1266.620 ;
        RECT 2509.380 33.690 2527.780 1266.620 ;
        RECT 2531.380 984.410 2585.780 1266.620 ;
        RECT 2589.380 984.410 2607.780 1266.620 ;
        RECT 2611.380 984.410 2665.780 1266.620 ;
        RECT 2669.380 984.410 2687.780 1266.620 ;
        RECT 2691.380 984.410 2745.780 1266.620 ;
        RECT 2749.380 984.410 2767.780 1266.620 ;
        RECT 2771.380 984.410 2825.780 1266.620 ;
        RECT 2829.380 984.410 2847.780 1266.620 ;
        RECT 2851.380 984.410 2880.280 1266.620 ;
        RECT 2883.880 984.410 2892.280 1266.620 ;
        RECT 2895.880 984.410 2905.780 1266.620 ;
        RECT 2909.380 984.410 2927.780 1266.620 ;
        RECT 2931.380 984.410 2985.780 1266.620 ;
        RECT 2989.380 984.410 3007.780 1266.620 ;
        RECT 3011.380 984.410 3098.780 1266.620 ;
        RECT 2531.380 219.350 3098.780 984.410 ;
        RECT 2531.380 33.690 2585.780 219.350 ;
        RECT 2589.380 33.690 2607.780 219.350 ;
        RECT 2611.380 33.690 2665.780 219.350 ;
        RECT 2669.380 33.690 2687.780 219.350 ;
        RECT 2691.380 33.690 2745.780 219.350 ;
        RECT 2749.380 33.690 2767.780 219.350 ;
        RECT 2771.380 33.690 2825.780 219.350 ;
        RECT 2829.380 33.690 2847.780 219.350 ;
        RECT 2851.380 33.690 2880.280 219.350 ;
        RECT 2883.880 33.690 2892.280 219.350 ;
        RECT 2895.880 144.425 2905.780 219.350 ;
        RECT 2909.380 144.425 2927.780 219.350 ;
        RECT 2931.380 144.425 2985.780 219.350 ;
        RECT 2895.880 87.030 2985.780 144.425 ;
        RECT 2895.880 33.690 2905.780 87.030 ;
        RECT 2909.380 33.690 2927.780 87.030 ;
        RECT 2931.380 33.690 2985.780 87.030 ;
        RECT 2989.380 33.690 3007.780 219.350 ;
        RECT 3011.380 33.690 3098.780 219.350 ;
        RECT 3102.380 33.690 3107.780 4332.630 ;
        RECT 3111.380 33.690 3126.320 4332.630 ;
        RECT 3129.920 33.690 3135.320 4332.630 ;
        RECT 3138.920 33.690 3145.220 4332.630 ;
        RECT 3155.820 33.690 3157.220 4332.630 ;
        RECT 3167.820 33.690 3168.340 4332.630 ;
      LAYER Metal5 ;
        RECT 1.180 4320.090 3168.420 4332.660 ;
        RECT 1.180 4316.090 1.580 4320.090 ;
        RECT 3168.020 4316.090 3168.420 4320.090 ;
        RECT 1.180 4290.090 3168.420 4316.090 ;
        RECT 1.180 4286.090 1.580 4290.090 ;
        RECT 3168.020 4286.090 3168.420 4290.090 ;
        RECT 1.180 4260.090 3168.420 4286.090 ;
        RECT 1.180 4256.090 1.580 4260.090 ;
        RECT 93.640 4256.090 3076.360 4260.090 ;
        RECT 3168.020 4256.090 3168.420 4260.090 ;
        RECT 1.180 4230.090 3168.420 4256.090 ;
        RECT 1.180 4226.090 1.580 4230.090 ;
        RECT 93.640 4226.090 3076.360 4230.090 ;
        RECT 3168.020 4226.090 3168.420 4230.090 ;
        RECT 1.180 4200.090 3168.420 4226.090 ;
        RECT 1.180 4196.090 1.580 4200.090 ;
        RECT 93.640 4196.090 3076.360 4200.090 ;
        RECT 3168.020 4196.090 3168.420 4200.090 ;
        RECT 1.180 4170.090 3168.420 4196.090 ;
        RECT 1.180 4166.090 1.580 4170.090 ;
        RECT 93.640 4166.090 3076.360 4170.090 ;
        RECT 3168.020 4166.090 3168.420 4170.090 ;
        RECT 1.180 4140.090 3168.420 4166.090 ;
        RECT 1.180 4136.090 1.580 4140.090 ;
        RECT 93.640 4136.090 3076.360 4140.090 ;
        RECT 3168.020 4136.090 3168.420 4140.090 ;
        RECT 1.180 4110.090 3168.420 4136.090 ;
        RECT 1.180 4106.090 1.580 4110.090 ;
        RECT 93.640 4106.090 3076.360 4110.090 ;
        RECT 3168.020 4106.090 3168.420 4110.090 ;
        RECT 1.180 4080.090 3168.420 4106.090 ;
        RECT 1.180 4076.090 1.580 4080.090 ;
        RECT 93.640 4076.090 3076.360 4080.090 ;
        RECT 3168.020 4076.090 3168.420 4080.090 ;
        RECT 1.180 4050.090 3168.420 4076.090 ;
        RECT 1.180 4046.090 1.580 4050.090 ;
        RECT 93.640 4046.090 3076.360 4050.090 ;
        RECT 3168.020 4046.090 3168.420 4050.090 ;
        RECT 1.180 4020.090 3168.420 4046.090 ;
        RECT 1.180 4016.090 1.580 4020.090 ;
        RECT 93.640 4016.090 3076.360 4020.090 ;
        RECT 3168.020 4016.090 3168.420 4020.090 ;
        RECT 1.180 3990.090 3168.420 4016.090 ;
        RECT 1.180 3986.090 1.580 3990.090 ;
        RECT 93.640 3986.090 3076.360 3990.090 ;
        RECT 3168.020 3986.090 3168.420 3990.090 ;
        RECT 1.180 3960.090 3168.420 3986.090 ;
        RECT 1.180 3956.090 1.580 3960.090 ;
        RECT 93.640 3956.090 3076.360 3960.090 ;
        RECT 3168.020 3956.090 3168.420 3960.090 ;
        RECT 1.180 3930.090 3168.420 3956.090 ;
        RECT 1.180 3926.090 1.580 3930.090 ;
        RECT 93.640 3926.090 3076.360 3930.090 ;
        RECT 3168.020 3926.090 3168.420 3930.090 ;
        RECT 1.180 3900.090 3168.420 3926.090 ;
        RECT 1.180 3896.090 1.580 3900.090 ;
        RECT 93.640 3896.090 3076.360 3900.090 ;
        RECT 3168.020 3896.090 3168.420 3900.090 ;
        RECT 1.180 3870.090 3168.420 3896.090 ;
        RECT 1.180 3866.090 1.580 3870.090 ;
        RECT 93.640 3866.090 3076.360 3870.090 ;
        RECT 3168.020 3866.090 3168.420 3870.090 ;
        RECT 1.180 3840.090 3168.420 3866.090 ;
        RECT 1.180 3836.090 1.580 3840.090 ;
        RECT 93.640 3836.090 3076.360 3840.090 ;
        RECT 3168.020 3836.090 3168.420 3840.090 ;
        RECT 1.180 3810.090 3168.420 3836.090 ;
        RECT 1.180 3806.090 1.580 3810.090 ;
        RECT 93.640 3806.090 3076.360 3810.090 ;
        RECT 3168.020 3806.090 3168.420 3810.090 ;
        RECT 1.180 3780.090 3168.420 3806.090 ;
        RECT 1.180 3776.090 1.580 3780.090 ;
        RECT 93.640 3776.090 3076.360 3780.090 ;
        RECT 3168.020 3776.090 3168.420 3780.090 ;
        RECT 1.180 3750.090 3168.420 3776.090 ;
        RECT 1.180 3746.090 1.580 3750.090 ;
        RECT 93.640 3746.090 3076.360 3750.090 ;
        RECT 3168.020 3746.090 3168.420 3750.090 ;
        RECT 1.180 3720.090 3168.420 3746.090 ;
        RECT 1.180 3716.090 1.580 3720.090 ;
        RECT 93.640 3716.090 3076.360 3720.090 ;
        RECT 3168.020 3716.090 3168.420 3720.090 ;
        RECT 1.180 3690.090 3168.420 3716.090 ;
        RECT 1.180 3686.090 1.580 3690.090 ;
        RECT 93.640 3686.090 3076.360 3690.090 ;
        RECT 3168.020 3686.090 3168.420 3690.090 ;
        RECT 1.180 3660.090 3168.420 3686.090 ;
        RECT 1.180 3656.090 1.580 3660.090 ;
        RECT 93.640 3656.090 3076.360 3660.090 ;
        RECT 3168.020 3656.090 3168.420 3660.090 ;
        RECT 1.180 3630.090 3168.420 3656.090 ;
        RECT 1.180 3626.090 1.580 3630.090 ;
        RECT 93.640 3626.090 3076.360 3630.090 ;
        RECT 3168.020 3626.090 3168.420 3630.090 ;
        RECT 1.180 3600.090 3168.420 3626.090 ;
        RECT 1.180 3596.090 1.580 3600.090 ;
        RECT 93.640 3596.090 3076.360 3600.090 ;
        RECT 3168.020 3596.090 3168.420 3600.090 ;
        RECT 1.180 3570.090 3168.420 3596.090 ;
        RECT 1.180 3566.090 1.580 3570.090 ;
        RECT 93.640 3566.090 3076.360 3570.090 ;
        RECT 3168.020 3566.090 3168.420 3570.090 ;
        RECT 1.180 3540.090 3168.420 3566.090 ;
        RECT 1.180 3536.090 1.580 3540.090 ;
        RECT 93.640 3536.090 3076.360 3540.090 ;
        RECT 3168.020 3536.090 3168.420 3540.090 ;
        RECT 1.180 3510.090 3168.420 3536.090 ;
        RECT 1.180 3506.090 1.580 3510.090 ;
        RECT 93.640 3506.090 3076.360 3510.090 ;
        RECT 3168.020 3506.090 3168.420 3510.090 ;
        RECT 1.180 3480.090 3168.420 3506.090 ;
        RECT 1.180 3476.090 1.580 3480.090 ;
        RECT 93.640 3476.090 3076.360 3480.090 ;
        RECT 3168.020 3476.090 3168.420 3480.090 ;
        RECT 1.180 3450.090 3168.420 3476.090 ;
        RECT 1.180 3446.090 1.580 3450.090 ;
        RECT 93.640 3446.090 3076.360 3450.090 ;
        RECT 3168.020 3446.090 3168.420 3450.090 ;
        RECT 1.180 3420.090 3168.420 3446.090 ;
        RECT 1.180 3416.090 1.580 3420.090 ;
        RECT 93.640 3416.090 3076.360 3420.090 ;
        RECT 3168.020 3416.090 3168.420 3420.090 ;
        RECT 1.180 3390.090 3168.420 3416.090 ;
        RECT 1.180 3386.090 1.580 3390.090 ;
        RECT 93.640 3386.090 3076.360 3390.090 ;
        RECT 3168.020 3386.090 3168.420 3390.090 ;
        RECT 1.180 3360.090 3168.420 3386.090 ;
        RECT 1.180 3356.090 1.580 3360.090 ;
        RECT 93.640 3356.090 3076.360 3360.090 ;
        RECT 3168.020 3356.090 3168.420 3360.090 ;
        RECT 1.180 3330.090 3168.420 3356.090 ;
        RECT 1.180 3326.090 1.580 3330.090 ;
        RECT 93.640 3326.090 3076.360 3330.090 ;
        RECT 3168.020 3326.090 3168.420 3330.090 ;
        RECT 1.180 3300.090 3168.420 3326.090 ;
        RECT 1.180 3296.090 1.580 3300.090 ;
        RECT 93.640 3296.090 3076.360 3300.090 ;
        RECT 3168.020 3296.090 3168.420 3300.090 ;
        RECT 1.180 3270.090 3168.420 3296.090 ;
        RECT 1.180 3266.090 1.580 3270.090 ;
        RECT 93.640 3266.090 3076.360 3270.090 ;
        RECT 3168.020 3266.090 3168.420 3270.090 ;
        RECT 1.180 3240.090 3168.420 3266.090 ;
        RECT 1.180 3236.090 1.580 3240.090 ;
        RECT 93.640 3236.090 3076.360 3240.090 ;
        RECT 3168.020 3236.090 3168.420 3240.090 ;
        RECT 1.180 3210.090 3168.420 3236.090 ;
        RECT 1.180 3206.090 1.580 3210.090 ;
        RECT 93.640 3206.090 3076.360 3210.090 ;
        RECT 3168.020 3206.090 3168.420 3210.090 ;
        RECT 1.180 3180.090 3168.420 3206.090 ;
        RECT 1.180 3176.090 1.580 3180.090 ;
        RECT 93.640 3176.090 3076.360 3180.090 ;
        RECT 3168.020 3176.090 3168.420 3180.090 ;
        RECT 1.180 3150.090 3168.420 3176.090 ;
        RECT 1.180 3146.090 1.580 3150.090 ;
        RECT 93.640 3146.090 3076.360 3150.090 ;
        RECT 3168.020 3146.090 3168.420 3150.090 ;
        RECT 1.180 3120.090 3168.420 3146.090 ;
        RECT 1.180 3116.090 1.580 3120.090 ;
        RECT 93.640 3116.090 3076.360 3120.090 ;
        RECT 3168.020 3116.090 3168.420 3120.090 ;
        RECT 1.180 3090.090 3168.420 3116.090 ;
        RECT 1.180 3086.090 1.580 3090.090 ;
        RECT 93.640 3086.090 3076.360 3090.090 ;
        RECT 3168.020 3086.090 3168.420 3090.090 ;
        RECT 1.180 3060.090 3168.420 3086.090 ;
        RECT 1.180 3056.090 1.580 3060.090 ;
        RECT 93.640 3056.090 3076.360 3060.090 ;
        RECT 3168.020 3056.090 3168.420 3060.090 ;
        RECT 1.180 3030.090 3168.420 3056.090 ;
        RECT 1.180 3026.090 1.580 3030.090 ;
        RECT 93.640 3026.090 3076.360 3030.090 ;
        RECT 3168.020 3026.090 3168.420 3030.090 ;
        RECT 1.180 3000.090 3168.420 3026.090 ;
        RECT 1.180 2996.090 1.580 3000.090 ;
        RECT 93.640 2996.090 3076.360 3000.090 ;
        RECT 3168.020 2996.090 3168.420 3000.090 ;
        RECT 1.180 2970.090 3168.420 2996.090 ;
        RECT 1.180 2966.090 1.580 2970.090 ;
        RECT 93.640 2966.090 3076.360 2970.090 ;
        RECT 3168.020 2966.090 3168.420 2970.090 ;
        RECT 1.180 2940.090 3168.420 2966.090 ;
        RECT 1.180 2936.090 1.580 2940.090 ;
        RECT 93.640 2936.090 3076.360 2940.090 ;
        RECT 3168.020 2936.090 3168.420 2940.090 ;
        RECT 1.180 2910.090 3168.420 2936.090 ;
        RECT 1.180 2906.090 1.580 2910.090 ;
        RECT 93.640 2906.090 3076.360 2910.090 ;
        RECT 3168.020 2906.090 3168.420 2910.090 ;
        RECT 1.180 2880.090 3168.420 2906.090 ;
        RECT 1.180 2876.090 1.580 2880.090 ;
        RECT 93.640 2876.090 3076.360 2880.090 ;
        RECT 3168.020 2876.090 3168.420 2880.090 ;
        RECT 1.180 2850.090 3168.420 2876.090 ;
        RECT 1.180 2846.090 1.580 2850.090 ;
        RECT 93.640 2846.090 3076.360 2850.090 ;
        RECT 3168.020 2846.090 3168.420 2850.090 ;
        RECT 1.180 2820.090 3168.420 2846.090 ;
        RECT 1.180 2816.090 1.580 2820.090 ;
        RECT 93.640 2816.090 3076.360 2820.090 ;
        RECT 3168.020 2816.090 3168.420 2820.090 ;
        RECT 1.180 2790.090 3168.420 2816.090 ;
        RECT 1.180 2786.090 1.580 2790.090 ;
        RECT 93.640 2786.090 3076.360 2790.090 ;
        RECT 3168.020 2786.090 3168.420 2790.090 ;
        RECT 1.180 2760.090 3168.420 2786.090 ;
        RECT 1.180 2756.090 1.580 2760.090 ;
        RECT 93.640 2756.090 3076.360 2760.090 ;
        RECT 3168.020 2756.090 3168.420 2760.090 ;
        RECT 1.180 2730.090 3168.420 2756.090 ;
        RECT 1.180 2726.090 1.580 2730.090 ;
        RECT 93.640 2726.090 3076.360 2730.090 ;
        RECT 3168.020 2726.090 3168.420 2730.090 ;
        RECT 1.180 2700.090 3168.420 2726.090 ;
        RECT 1.180 2696.090 1.580 2700.090 ;
        RECT 93.640 2696.090 3076.360 2700.090 ;
        RECT 3168.020 2696.090 3168.420 2700.090 ;
        RECT 1.180 2670.090 3168.420 2696.090 ;
        RECT 1.180 2666.090 1.580 2670.090 ;
        RECT 93.640 2666.090 3076.360 2670.090 ;
        RECT 3168.020 2666.090 3168.420 2670.090 ;
        RECT 1.180 2640.090 3168.420 2666.090 ;
        RECT 1.180 2636.090 1.580 2640.090 ;
        RECT 93.640 2636.090 3076.360 2640.090 ;
        RECT 3168.020 2636.090 3168.420 2640.090 ;
        RECT 1.180 2610.090 3168.420 2636.090 ;
        RECT 1.180 2606.090 1.580 2610.090 ;
        RECT 93.640 2606.090 3076.360 2610.090 ;
        RECT 3168.020 2606.090 3168.420 2610.090 ;
        RECT 1.180 2580.090 3168.420 2606.090 ;
        RECT 1.180 2576.090 1.580 2580.090 ;
        RECT 93.640 2576.090 3076.360 2580.090 ;
        RECT 3168.020 2576.090 3168.420 2580.090 ;
        RECT 1.180 2550.090 3168.420 2576.090 ;
        RECT 1.180 2546.090 1.580 2550.090 ;
        RECT 93.640 2546.090 3076.360 2550.090 ;
        RECT 3168.020 2546.090 3168.420 2550.090 ;
        RECT 1.180 2520.090 3168.420 2546.090 ;
        RECT 1.180 2516.090 1.580 2520.090 ;
        RECT 93.640 2516.090 3076.360 2520.090 ;
        RECT 3168.020 2516.090 3168.420 2520.090 ;
        RECT 1.180 2490.090 3168.420 2516.090 ;
        RECT 1.180 2486.090 1.580 2490.090 ;
        RECT 93.640 2486.090 3076.360 2490.090 ;
        RECT 3168.020 2486.090 3168.420 2490.090 ;
        RECT 1.180 2460.090 3168.420 2486.090 ;
        RECT 1.180 2456.090 1.580 2460.090 ;
        RECT 93.640 2456.090 3076.360 2460.090 ;
        RECT 3168.020 2456.090 3168.420 2460.090 ;
        RECT 1.180 2430.090 3168.420 2456.090 ;
        RECT 1.180 2426.090 1.580 2430.090 ;
        RECT 93.640 2426.090 3076.360 2430.090 ;
        RECT 3168.020 2426.090 3168.420 2430.090 ;
        RECT 1.180 2400.090 3168.420 2426.090 ;
        RECT 1.180 2396.090 1.580 2400.090 ;
        RECT 93.640 2396.090 3076.360 2400.090 ;
        RECT 3168.020 2396.090 3168.420 2400.090 ;
        RECT 1.180 2370.090 3168.420 2396.090 ;
        RECT 1.180 2366.090 1.580 2370.090 ;
        RECT 93.640 2366.090 3076.360 2370.090 ;
        RECT 3168.020 2366.090 3168.420 2370.090 ;
        RECT 1.180 2340.090 3168.420 2366.090 ;
        RECT 1.180 2336.090 1.580 2340.090 ;
        RECT 93.640 2336.090 3076.360 2340.090 ;
        RECT 3168.020 2336.090 3168.420 2340.090 ;
        RECT 1.180 2310.090 3168.420 2336.090 ;
        RECT 1.180 2306.090 1.580 2310.090 ;
        RECT 93.640 2306.090 3076.360 2310.090 ;
        RECT 3168.020 2306.090 3168.420 2310.090 ;
        RECT 1.180 2280.090 3168.420 2306.090 ;
        RECT 1.180 2276.090 1.580 2280.090 ;
        RECT 93.640 2276.090 3076.360 2280.090 ;
        RECT 3168.020 2276.090 3168.420 2280.090 ;
        RECT 1.180 2250.090 3168.420 2276.090 ;
        RECT 1.180 2246.090 1.580 2250.090 ;
        RECT 93.640 2246.090 3076.360 2250.090 ;
        RECT 3168.020 2246.090 3168.420 2250.090 ;
        RECT 1.180 2220.090 3168.420 2246.090 ;
        RECT 1.180 2216.090 1.580 2220.090 ;
        RECT 93.640 2216.090 3076.360 2220.090 ;
        RECT 3168.020 2216.090 3168.420 2220.090 ;
        RECT 1.180 2190.090 3168.420 2216.090 ;
        RECT 1.180 2186.090 1.580 2190.090 ;
        RECT 93.640 2186.090 3076.360 2190.090 ;
        RECT 3168.020 2186.090 3168.420 2190.090 ;
        RECT 1.180 2160.090 3168.420 2186.090 ;
        RECT 1.180 2156.090 1.580 2160.090 ;
        RECT 93.640 2156.090 3076.360 2160.090 ;
        RECT 3168.020 2156.090 3168.420 2160.090 ;
        RECT 1.180 2130.090 3168.420 2156.090 ;
        RECT 1.180 2126.090 1.580 2130.090 ;
        RECT 93.640 2126.090 3076.360 2130.090 ;
        RECT 3168.020 2126.090 3168.420 2130.090 ;
        RECT 1.180 2100.090 3168.420 2126.090 ;
        RECT 1.180 2096.090 1.580 2100.090 ;
        RECT 93.640 2096.090 3076.360 2100.090 ;
        RECT 3168.020 2096.090 3168.420 2100.090 ;
        RECT 1.180 2070.090 3168.420 2096.090 ;
        RECT 1.180 2066.090 1.580 2070.090 ;
        RECT 93.640 2066.090 3076.360 2070.090 ;
        RECT 3168.020 2066.090 3168.420 2070.090 ;
        RECT 1.180 2040.090 3168.420 2066.090 ;
        RECT 1.180 2036.090 1.580 2040.090 ;
        RECT 93.640 2036.090 3076.360 2040.090 ;
        RECT 3168.020 2036.090 3168.420 2040.090 ;
        RECT 1.180 2010.090 3168.420 2036.090 ;
        RECT 1.180 2006.090 1.580 2010.090 ;
        RECT 93.640 2006.090 3076.360 2010.090 ;
        RECT 3168.020 2006.090 3168.420 2010.090 ;
        RECT 1.180 1980.090 3168.420 2006.090 ;
        RECT 1.180 1976.090 1.580 1980.090 ;
        RECT 93.640 1976.090 3076.360 1980.090 ;
        RECT 3168.020 1976.090 3168.420 1980.090 ;
        RECT 1.180 1950.090 3168.420 1976.090 ;
        RECT 1.180 1946.090 1.580 1950.090 ;
        RECT 93.640 1946.090 3076.360 1950.090 ;
        RECT 3168.020 1946.090 3168.420 1950.090 ;
        RECT 1.180 1920.090 3168.420 1946.090 ;
        RECT 1.180 1916.090 1.580 1920.090 ;
        RECT 93.640 1916.090 3076.360 1920.090 ;
        RECT 3168.020 1916.090 3168.420 1920.090 ;
        RECT 1.180 1890.090 3168.420 1916.090 ;
        RECT 1.180 1886.090 1.580 1890.090 ;
        RECT 93.640 1886.090 3076.360 1890.090 ;
        RECT 3168.020 1886.090 3168.420 1890.090 ;
        RECT 1.180 1860.090 3168.420 1886.090 ;
        RECT 1.180 1856.090 1.580 1860.090 ;
        RECT 93.640 1856.090 3076.360 1860.090 ;
        RECT 3168.020 1856.090 3168.420 1860.090 ;
        RECT 1.180 1830.090 3168.420 1856.090 ;
        RECT 1.180 1826.090 1.580 1830.090 ;
        RECT 93.640 1826.090 3076.360 1830.090 ;
        RECT 3168.020 1826.090 3168.420 1830.090 ;
        RECT 1.180 1800.090 3168.420 1826.090 ;
        RECT 1.180 1796.090 1.580 1800.090 ;
        RECT 93.640 1796.090 3076.360 1800.090 ;
        RECT 3168.020 1796.090 3168.420 1800.090 ;
        RECT 1.180 1770.090 3168.420 1796.090 ;
        RECT 1.180 1766.090 1.580 1770.090 ;
        RECT 93.640 1766.090 3076.360 1770.090 ;
        RECT 3168.020 1766.090 3168.420 1770.090 ;
        RECT 1.180 1740.090 3168.420 1766.090 ;
        RECT 1.180 1736.090 1.580 1740.090 ;
        RECT 93.640 1736.090 3076.360 1740.090 ;
        RECT 3168.020 1736.090 3168.420 1740.090 ;
        RECT 1.180 1710.090 3168.420 1736.090 ;
        RECT 1.180 1706.090 1.580 1710.090 ;
        RECT 93.640 1706.090 3076.360 1710.090 ;
        RECT 3168.020 1706.090 3168.420 1710.090 ;
        RECT 1.180 1680.090 3168.420 1706.090 ;
        RECT 1.180 1676.090 1.580 1680.090 ;
        RECT 93.640 1676.090 3076.360 1680.090 ;
        RECT 3168.020 1676.090 3168.420 1680.090 ;
        RECT 1.180 1650.090 3168.420 1676.090 ;
        RECT 1.180 1646.090 1.580 1650.090 ;
        RECT 93.640 1646.090 3076.360 1650.090 ;
        RECT 3168.020 1646.090 3168.420 1650.090 ;
        RECT 1.180 1620.090 3168.420 1646.090 ;
        RECT 1.180 1616.090 1.580 1620.090 ;
        RECT 93.640 1616.090 3076.360 1620.090 ;
        RECT 3168.020 1616.090 3168.420 1620.090 ;
        RECT 1.180 1590.090 3168.420 1616.090 ;
        RECT 1.180 1586.090 1.580 1590.090 ;
        RECT 93.640 1586.090 3076.360 1590.090 ;
        RECT 3168.020 1586.090 3168.420 1590.090 ;
        RECT 1.180 1560.090 3168.420 1586.090 ;
        RECT 1.180 1556.090 1.580 1560.090 ;
        RECT 93.640 1556.090 3076.360 1560.090 ;
        RECT 3168.020 1556.090 3168.420 1560.090 ;
        RECT 1.180 1530.090 3168.420 1556.090 ;
        RECT 1.180 1526.090 1.580 1530.090 ;
        RECT 93.640 1526.090 3076.360 1530.090 ;
        RECT 3168.020 1526.090 3168.420 1530.090 ;
        RECT 1.180 1500.090 3168.420 1526.090 ;
        RECT 1.180 1496.090 1.580 1500.090 ;
        RECT 93.640 1496.090 3076.360 1500.090 ;
        RECT 3168.020 1496.090 3168.420 1500.090 ;
        RECT 1.180 1470.090 3168.420 1496.090 ;
        RECT 1.180 1466.090 1.580 1470.090 ;
        RECT 93.640 1466.090 3076.360 1470.090 ;
        RECT 3168.020 1466.090 3168.420 1470.090 ;
        RECT 1.180 1440.090 3168.420 1466.090 ;
        RECT 1.180 1436.090 1.580 1440.090 ;
        RECT 93.640 1436.090 3076.360 1440.090 ;
        RECT 3168.020 1436.090 3168.420 1440.090 ;
        RECT 1.180 1410.090 3168.420 1436.090 ;
        RECT 1.180 1406.090 1.580 1410.090 ;
        RECT 93.640 1406.090 3076.360 1410.090 ;
        RECT 3168.020 1406.090 3168.420 1410.090 ;
        RECT 1.180 1380.090 3168.420 1406.090 ;
        RECT 1.180 1376.090 1.580 1380.090 ;
        RECT 93.640 1376.090 3076.360 1380.090 ;
        RECT 3168.020 1376.090 3168.420 1380.090 ;
        RECT 1.180 1350.090 3168.420 1376.090 ;
        RECT 1.180 1346.090 1.580 1350.090 ;
        RECT 93.640 1346.090 3076.360 1350.090 ;
        RECT 3168.020 1346.090 3168.420 1350.090 ;
        RECT 1.180 1320.090 3168.420 1346.090 ;
        RECT 1.180 1316.090 1.580 1320.090 ;
        RECT 93.640 1316.090 3076.360 1320.090 ;
        RECT 3168.020 1316.090 3168.420 1320.090 ;
        RECT 1.180 1290.090 3168.420 1316.090 ;
        RECT 1.180 1286.090 1.580 1290.090 ;
        RECT 93.640 1286.090 3076.360 1290.090 ;
        RECT 3168.020 1286.090 3168.420 1290.090 ;
        RECT 1.180 1260.090 3168.420 1286.090 ;
        RECT 1.180 1256.090 1.580 1260.090 ;
        RECT 3168.020 1256.090 3168.420 1260.090 ;
        RECT 1.180 1230.090 3168.420 1256.090 ;
        RECT 1.180 1226.090 1.580 1230.090 ;
        RECT 3168.020 1226.090 3168.420 1230.090 ;
        RECT 1.180 1200.090 3168.420 1226.090 ;
        RECT 1.180 1196.090 1.580 1200.090 ;
        RECT 3168.020 1196.090 3168.420 1200.090 ;
        RECT 1.180 1170.090 3168.420 1196.090 ;
        RECT 1.180 1166.090 1.580 1170.090 ;
        RECT 3168.020 1166.090 3168.420 1170.090 ;
        RECT 1.180 1140.090 3168.420 1166.090 ;
        RECT 1.180 1136.090 1.580 1140.090 ;
        RECT 3168.020 1136.090 3168.420 1140.090 ;
        RECT 1.180 1110.090 3168.420 1136.090 ;
        RECT 1.180 1106.090 1.580 1110.090 ;
        RECT 1562.040 1106.090 1631.960 1110.090 ;
        RECT 2121.540 1106.090 2191.460 1110.090 ;
        RECT 3168.020 1106.090 3168.420 1110.090 ;
        RECT 1.180 1080.090 3168.420 1106.090 ;
        RECT 1.180 1076.090 1.580 1080.090 ;
        RECT 1562.040 1076.090 1631.960 1080.090 ;
        RECT 2121.540 1076.090 2191.460 1080.090 ;
        RECT 3168.020 1076.090 3168.420 1080.090 ;
        RECT 1.180 1050.090 3168.420 1076.090 ;
        RECT 1.180 1046.090 1.580 1050.090 ;
        RECT 1562.040 1046.090 1631.960 1050.090 ;
        RECT 2121.540 1046.090 2191.460 1050.090 ;
        RECT 3168.020 1046.090 3168.420 1050.090 ;
        RECT 1.180 1020.090 3168.420 1046.090 ;
        RECT 1.180 1016.090 1.580 1020.090 ;
        RECT 3168.020 1016.090 3168.420 1020.090 ;
        RECT 1.180 990.090 3168.420 1016.090 ;
        RECT 1.180 986.090 1.580 990.090 ;
        RECT 3168.020 986.090 3168.420 990.090 ;
        RECT 1.180 960.090 3168.420 986.090 ;
        RECT 1.180 956.090 1.580 960.090 ;
        RECT 602.040 956.090 671.960 960.090 ;
        RECT 1082.040 956.090 1151.960 960.090 ;
        RECT 2550.260 956.090 3054.060 960.090 ;
        RECT 3168.020 956.090 3168.420 960.090 ;
        RECT 1.180 930.090 3168.420 956.090 ;
        RECT 1.180 926.090 1.580 930.090 ;
        RECT 602.040 926.090 671.960 930.090 ;
        RECT 1082.040 926.090 1151.960 930.090 ;
        RECT 2550.260 926.090 3054.060 930.090 ;
        RECT 3168.020 926.090 3168.420 930.090 ;
        RECT 1.180 900.090 3168.420 926.090 ;
        RECT 1.180 896.090 1.580 900.090 ;
        RECT 602.040 896.090 671.960 900.090 ;
        RECT 1082.040 896.090 1151.960 900.090 ;
        RECT 2550.260 896.090 3054.060 900.090 ;
        RECT 3168.020 896.090 3168.420 900.090 ;
        RECT 1.180 870.090 3168.420 896.090 ;
        RECT 1.180 866.090 1.580 870.090 ;
        RECT 2550.260 866.090 3054.060 870.090 ;
        RECT 3168.020 866.090 3168.420 870.090 ;
        RECT 1.180 840.090 3168.420 866.090 ;
        RECT 1.180 836.090 1.580 840.090 ;
        RECT 2550.260 836.090 3054.060 840.090 ;
        RECT 3168.020 836.090 3168.420 840.090 ;
        RECT 1.180 810.090 3168.420 836.090 ;
        RECT 1.180 806.090 1.580 810.090 ;
        RECT 2550.260 806.090 3054.060 810.090 ;
        RECT 3168.020 806.090 3168.420 810.090 ;
        RECT 1.180 780.090 3168.420 806.090 ;
        RECT 1.180 776.090 1.580 780.090 ;
        RECT 2550.260 776.090 3054.060 780.090 ;
        RECT 3168.020 776.090 3168.420 780.090 ;
        RECT 1.180 750.090 3168.420 776.090 ;
        RECT 1.180 746.090 1.580 750.090 ;
        RECT 2550.260 746.090 3054.060 750.090 ;
        RECT 3168.020 746.090 3168.420 750.090 ;
        RECT 1.180 720.090 3168.420 746.090 ;
        RECT 1.180 716.090 1.580 720.090 ;
        RECT 2550.260 716.090 3054.060 720.090 ;
        RECT 3168.020 716.090 3168.420 720.090 ;
        RECT 1.180 690.090 3168.420 716.090 ;
        RECT 1.180 686.090 1.580 690.090 ;
        RECT 2550.260 686.090 3054.060 690.090 ;
        RECT 3168.020 686.090 3168.420 690.090 ;
        RECT 1.180 660.090 3168.420 686.090 ;
        RECT 1.180 656.090 1.580 660.090 ;
        RECT 2550.260 656.090 3054.060 660.090 ;
        RECT 3168.020 656.090 3168.420 660.090 ;
        RECT 1.180 630.090 3168.420 656.090 ;
        RECT 1.180 626.090 1.580 630.090 ;
        RECT 2550.260 626.090 3054.060 630.090 ;
        RECT 3168.020 626.090 3168.420 630.090 ;
        RECT 1.180 600.090 3168.420 626.090 ;
        RECT 1.180 596.090 1.580 600.090 ;
        RECT 2550.260 596.090 3054.060 600.090 ;
        RECT 3168.020 596.090 3168.420 600.090 ;
        RECT 1.180 570.090 3168.420 596.090 ;
        RECT 1.180 566.090 1.580 570.090 ;
        RECT 2550.260 566.090 3054.060 570.090 ;
        RECT 3168.020 566.090 3168.420 570.090 ;
        RECT 1.180 540.090 3168.420 566.090 ;
        RECT 1.180 536.090 1.580 540.090 ;
        RECT 2550.260 536.090 3054.060 540.090 ;
        RECT 3168.020 536.090 3168.420 540.090 ;
        RECT 1.180 510.090 3168.420 536.090 ;
        RECT 1.180 506.090 1.580 510.090 ;
        RECT 2550.260 506.090 3054.060 510.090 ;
        RECT 3168.020 506.090 3168.420 510.090 ;
        RECT 1.180 480.090 3168.420 506.090 ;
        RECT 1.180 476.090 1.580 480.090 ;
        RECT 2550.260 476.090 3054.060 480.090 ;
        RECT 3168.020 476.090 3168.420 480.090 ;
        RECT 1.180 450.090 3168.420 476.090 ;
        RECT 1.180 446.090 1.580 450.090 ;
        RECT 2550.260 446.090 3054.060 450.090 ;
        RECT 3168.020 446.090 3168.420 450.090 ;
        RECT 1.180 420.090 3168.420 446.090 ;
        RECT 1.180 416.090 1.580 420.090 ;
        RECT 2550.260 416.090 3054.060 420.090 ;
        RECT 3168.020 416.090 3168.420 420.090 ;
        RECT 1.180 390.090 3168.420 416.090 ;
        RECT 1.180 386.090 1.580 390.090 ;
        RECT 2550.260 386.090 3054.060 390.090 ;
        RECT 3168.020 386.090 3168.420 390.090 ;
        RECT 1.180 360.090 3168.420 386.090 ;
        RECT 1.180 356.090 1.580 360.090 ;
        RECT 2550.260 356.090 3054.060 360.090 ;
        RECT 3168.020 356.090 3168.420 360.090 ;
        RECT 1.180 330.090 3168.420 356.090 ;
        RECT 1.180 326.090 1.580 330.090 ;
        RECT 2550.260 326.090 3054.060 330.090 ;
        RECT 3168.020 326.090 3168.420 330.090 ;
        RECT 1.180 300.090 3168.420 326.090 ;
        RECT 1.180 296.090 1.580 300.090 ;
        RECT 2550.260 296.090 3054.060 300.090 ;
        RECT 3168.020 296.090 3168.420 300.090 ;
        RECT 1.180 270.090 3168.420 296.090 ;
        RECT 1.180 266.090 1.580 270.090 ;
        RECT 2550.260 266.090 3054.060 270.090 ;
        RECT 3168.020 266.090 3168.420 270.090 ;
        RECT 1.180 240.090 3168.420 266.090 ;
        RECT 1.180 236.090 1.580 240.090 ;
        RECT 2550.260 236.090 3054.060 240.090 ;
        RECT 3168.020 236.090 3168.420 240.090 ;
        RECT 1.180 210.090 3168.420 236.090 ;
        RECT 1.180 206.090 1.580 210.090 ;
        RECT 3168.020 206.090 3168.420 210.090 ;
        RECT 1.180 180.090 3168.420 206.090 ;
        RECT 1.180 176.090 1.580 180.090 ;
        RECT 3168.020 176.090 3168.420 180.090 ;
        RECT 1.180 150.090 3168.420 176.090 ;
        RECT 1.180 146.090 1.580 150.090 ;
        RECT 2896.855 146.090 2966.495 150.090 ;
        RECT 3168.020 146.090 3168.420 150.090 ;
        RECT 1.180 120.090 3168.420 146.090 ;
        RECT 1.180 116.090 1.580 120.090 ;
        RECT 2896.855 116.090 2966.495 120.090 ;
        RECT 3168.020 116.090 3168.420 120.090 ;
        RECT 1.180 95.010 3168.420 116.090 ;
  END
END caravel_core
END LIBRARY

