magic
tech gf180mcuC
magscale 1 10
timestamp 1655126753
<< metal1 >>
rect 1487 1786 1562 2040
rect 1805 1907 1880 2050
rect 1805 1847 1812 1907
rect 1872 1847 1880 1907
rect 1805 1826 1880 1847
rect 2831 1786 2906 2040
rect 3149 1907 3224 2050
rect 3149 1847 3156 1907
rect 3216 1847 3224 1907
rect 3149 1826 3224 1847
rect 3951 1786 4026 2040
rect 4269 1907 4344 2050
rect 4269 1847 4276 1907
rect 4336 1847 4344 1907
rect 4269 1826 4344 1847
rect 5295 1786 5370 2040
rect 5613 1907 5688 2050
rect 5613 1847 5620 1907
rect 5680 1847 5688 1907
rect 5613 1826 5688 1847
rect 6415 1786 6490 2040
rect 6733 1907 6808 2050
rect 6733 1847 6740 1907
rect 6800 1847 6808 1907
rect 6733 1826 6808 1847
rect 7759 1786 7834 2040
rect 8077 1907 8152 2050
rect 8077 1847 8084 1907
rect 8144 1847 8152 1907
rect 8077 1826 8152 1847
rect 8879 1786 8954 2040
rect 9197 1907 9272 2050
rect 9197 1847 9204 1907
rect 9264 1847 9272 1907
rect 9197 1826 9272 1847
rect 10223 1786 10298 2040
rect 10541 1907 10616 2050
rect 10541 1847 10548 1907
rect 10608 1847 10616 1907
rect 10541 1826 10616 1847
rect 11343 1786 11418 2040
rect 11661 1907 11736 2050
rect 11661 1847 11668 1907
rect 11728 1847 11736 1907
rect 11661 1826 11736 1847
rect 12687 1786 12762 2040
rect 13005 1907 13080 2050
rect 13005 1847 13012 1907
rect 13072 1847 13080 1907
rect 13005 1826 13080 1847
rect 13807 1786 13882 2040
rect 14125 1907 14200 2050
rect 14125 1847 14132 1907
rect 14192 1847 14200 1907
rect 14125 1826 14200 1847
rect 15151 1786 15226 2040
rect 15469 1907 15544 2050
rect 15469 1847 15476 1907
rect 15536 1847 15544 1907
rect 15469 1826 15544 1847
rect 16271 1786 16346 2040
rect 16589 1907 16664 2050
rect 16589 1847 16596 1907
rect 16656 1847 16664 1907
rect 16589 1826 16664 1847
rect 17615 1786 17690 2040
rect 17933 1907 18008 2050
rect 17933 1847 17940 1907
rect 18000 1847 18008 1907
rect 17933 1826 18008 1847
rect 18735 1786 18810 2040
rect 19053 1907 19128 2050
rect 19053 1847 19060 1907
rect 19120 1847 19128 1907
rect 19053 1826 19128 1847
rect 20079 1786 20154 2040
rect 20397 1907 20472 2050
rect 20397 1847 20404 1907
rect 20464 1847 20472 1907
rect 20397 1826 20472 1847
rect 1357 1714 1562 1786
rect 2701 1714 2906 1786
rect 3821 1714 4026 1786
rect 5165 1714 5370 1786
rect 6285 1714 6490 1786
rect 7629 1714 7834 1786
rect 8749 1714 8954 1786
rect 10093 1714 10298 1786
rect 11213 1714 11418 1786
rect 12557 1714 12762 1786
rect 13677 1714 13882 1786
rect 15021 1714 15226 1786
rect 16141 1714 16346 1786
rect 17485 1714 17690 1786
rect 18605 1714 18810 1786
rect 19949 1714 20154 1786
rect 1357 1695 1429 1714
rect 2701 1695 2773 1714
rect 3821 1695 3893 1714
rect 5165 1695 5237 1714
rect 6285 1695 6357 1714
rect 7629 1695 7701 1714
rect 8749 1695 8821 1714
rect 10093 1695 10165 1714
rect 11213 1695 11285 1714
rect 12557 1695 12629 1714
rect 13677 1695 13749 1714
rect 15021 1695 15093 1714
rect 16141 1695 16213 1714
rect 17485 1695 17557 1714
rect 18605 1695 18677 1714
rect 19949 1695 20021 1714
rect 1357 1030 1429 1049
rect 2701 1030 2773 1049
rect 3821 1030 3893 1049
rect 5165 1030 5237 1049
rect 6285 1030 6357 1049
rect 7629 1030 7701 1049
rect 8749 1030 8821 1049
rect 10093 1030 10165 1049
rect 11213 1030 11285 1049
rect 12557 1030 12629 1049
rect 13677 1030 13749 1049
rect 15021 1030 15093 1049
rect 16141 1030 16213 1049
rect 16711 1037 16771 1049
rect 1357 958 1562 1030
rect 2701 958 2906 1030
rect 3821 958 4026 1030
rect 5165 958 5370 1030
rect 6285 958 6490 1030
rect 7629 958 7834 1030
rect 8749 958 8954 1030
rect 10093 958 10298 1030
rect 11213 958 11418 1030
rect 12557 958 12762 1030
rect 13677 958 13882 1030
rect 15021 958 15226 1030
rect 16141 958 16346 1030
rect 16711 965 16771 977
rect 17485 1030 17557 1049
rect 18068 1032 18128 1044
rect 1487 704 1562 958
rect 1805 897 1880 918
rect 1805 837 1812 897
rect 1872 837 1880 897
rect 1805 694 1880 837
rect 2831 704 2906 958
rect 3149 897 3224 918
rect 3149 837 3156 897
rect 3216 837 3224 897
rect 3149 694 3224 837
rect 3951 704 4026 958
rect 4269 897 4344 918
rect 4269 837 4276 897
rect 4336 837 4344 897
rect 4269 694 4344 837
rect 5295 704 5370 958
rect 5613 897 5688 918
rect 5613 837 5620 897
rect 5680 837 5688 897
rect 5613 694 5688 837
rect 6415 704 6490 958
rect 6733 897 6808 918
rect 6733 837 6740 897
rect 6800 837 6808 897
rect 6733 694 6808 837
rect 7759 704 7834 958
rect 8077 897 8152 918
rect 8077 837 8084 897
rect 8144 837 8152 897
rect 8077 694 8152 837
rect 8879 704 8954 958
rect 9197 897 9272 918
rect 9197 837 9204 897
rect 9264 837 9272 897
rect 9197 694 9272 837
rect 10223 704 10298 958
rect 10541 897 10616 918
rect 10541 837 10548 897
rect 10608 837 10616 897
rect 10541 694 10616 837
rect 11343 704 11418 958
rect 11661 897 11736 918
rect 11661 837 11668 897
rect 11728 837 11736 897
rect 11661 694 11736 837
rect 12687 704 12762 958
rect 13005 897 13080 918
rect 13005 837 13012 897
rect 13072 837 13080 897
rect 13005 694 13080 837
rect 13807 704 13882 958
rect 14125 897 14200 918
rect 14125 837 14132 897
rect 14192 837 14200 897
rect 14125 694 14200 837
rect 15151 704 15226 958
rect 15469 897 15544 918
rect 15469 837 15476 897
rect 15536 837 15544 897
rect 15469 694 15544 837
rect 16271 704 16346 958
rect 16589 897 16664 918
rect 16589 837 16596 897
rect 16656 837 16664 897
rect 16589 694 16664 837
rect 16715 789 16768 965
rect 17485 958 17690 1030
rect 18068 960 18128 972
rect 18605 1030 18677 1049
rect 19183 1037 19243 1049
rect 16711 777 16771 789
rect 16711 705 16771 717
rect 17615 704 17690 958
rect 17933 897 18008 918
rect 17933 837 17940 897
rect 18000 837 18008 897
rect 17933 694 18008 837
rect 18072 784 18125 960
rect 18605 958 18810 1030
rect 19183 965 19243 977
rect 19949 1030 20021 1049
rect 20524 1032 20584 1044
rect 18068 772 18128 784
rect 18068 700 18128 712
rect 18735 704 18810 958
rect 19053 897 19128 918
rect 19053 837 19060 897
rect 19120 837 19128 897
rect 19053 694 19128 837
rect 19187 789 19240 965
rect 19949 958 20154 1030
rect 20524 960 20584 972
rect 19183 777 19243 789
rect 19183 705 19243 717
rect 20079 704 20154 958
rect 20397 897 20472 918
rect 20397 837 20404 897
rect 20464 837 20472 897
rect 20397 694 20472 837
rect 20529 784 20582 960
rect 20524 772 20584 784
rect 20524 700 20584 712
rect 1709 645 2002 648
rect 1997 531 2002 645
rect 1709 528 2002 531
<< via1 >>
rect 1707 2098 2000 2212
rect 10707 2098 11000 2212
rect 19707 2098 20000 2212
rect 1812 1847 1872 1907
rect 3156 1847 3216 1907
rect 4276 1847 4336 1907
rect 5620 1847 5680 1907
rect 6740 1847 6800 1907
rect 8084 1847 8144 1907
rect 9204 1847 9264 1907
rect 10548 1847 10608 1907
rect 11668 1847 11728 1907
rect 13012 1847 13072 1907
rect 14132 1847 14192 1907
rect 15476 1847 15536 1907
rect 16596 1847 16656 1907
rect 17940 1847 18000 1907
rect 19060 1847 19120 1907
rect 20404 1847 20464 1907
rect 6209 1312 6499 1432
rect 15209 1312 15499 1432
rect 16711 977 16771 1037
rect 1812 837 1872 897
rect 3156 837 3216 897
rect 4276 837 4336 897
rect 5620 837 5680 897
rect 6740 837 6800 897
rect 8084 837 8144 897
rect 9204 837 9264 897
rect 10548 837 10608 897
rect 11668 837 11728 897
rect 13012 837 13072 897
rect 14132 837 14192 897
rect 15476 837 15536 897
rect 16596 837 16656 897
rect 18068 972 18128 1032
rect 16711 717 16771 777
rect 17940 837 18000 897
rect 19183 977 19243 1037
rect 18068 712 18128 772
rect 19060 837 19120 897
rect 20524 972 20584 1032
rect 19183 717 19243 777
rect 20404 837 20464 897
rect 20524 712 20584 772
rect 1709 531 1997 645
rect 10709 531 10997 645
rect 19709 531 19997 645
<< metal2 >>
rect 1694 2302 2014 2313
rect 1694 2095 1707 2302
rect 1696 2002 1707 2095
rect 2000 2002 2014 2302
rect 10696 2302 11014 2313
rect 10696 2216 10707 2302
rect 10694 2095 10707 2216
rect 1696 1993 2014 2002
rect 10696 2002 10707 2095
rect 11000 2002 11014 2302
rect 19696 2302 20014 2313
rect 19696 2216 19707 2302
rect 19694 2095 19707 2216
rect 10696 1993 11014 2002
rect 19696 2002 19707 2095
rect 20000 2002 20014 2302
rect 19696 1993 20014 2002
rect 1051 1907 1893 1909
rect 1051 1847 1812 1907
rect 1872 1847 1893 1907
rect 1051 1845 1893 1847
rect 2338 1907 3237 1909
rect 2338 1847 3156 1907
rect 3216 1847 3237 1907
rect 2338 1845 3237 1847
rect 3313 1907 4357 1909
rect 3313 1847 4276 1907
rect 4336 1847 4357 1907
rect 3313 1845 4357 1847
rect 4740 1907 5701 1909
rect 4740 1847 5620 1907
rect 5680 1847 5701 1907
rect 4740 1845 5701 1847
rect 6067 1907 6821 1909
rect 6067 1847 6740 1907
rect 6800 1847 6821 1907
rect 6067 1845 6821 1847
rect 6944 1907 8165 1909
rect 6944 1847 8084 1907
rect 8144 1847 8165 1907
rect 6944 1845 8165 1847
rect 8400 1907 9287 1909
rect 8400 1847 9204 1907
rect 9264 1847 9287 1907
rect 8400 1845 9287 1847
rect 9744 1907 10627 1909
rect 9744 1847 10548 1907
rect 10608 1847 10627 1907
rect 9744 1845 10627 1847
rect 11200 1907 11747 1909
rect 11200 1847 11668 1907
rect 11728 1847 11747 1907
rect 11200 1845 11747 1847
rect 12544 1907 13091 1909
rect 12544 1847 13012 1907
rect 13072 1847 13091 1907
rect 12544 1845 13091 1847
rect 13625 1907 14211 1909
rect 13625 1847 14132 1907
rect 14192 1847 14211 1907
rect 13625 1845 14211 1847
rect 14978 1907 15553 1909
rect 14978 1847 15476 1907
rect 15536 1847 15553 1907
rect 14978 1845 15553 1847
rect 16257 1907 16771 1909
rect 16257 1847 16596 1907
rect 16656 1847 16771 1907
rect 16257 1845 16771 1847
rect 17602 1907 18126 1909
rect 17602 1847 17940 1907
rect 18000 1847 18126 1907
rect 17602 1845 18126 1847
rect 18723 1907 19241 1909
rect 18723 1847 19060 1907
rect 19120 1847 19241 1907
rect 18723 1845 19241 1847
rect 20066 1907 20582 1909
rect 20066 1847 20404 1907
rect 20464 1847 20582 1907
rect 20066 1845 20582 1847
rect 1051 1076 1107 1845
rect 0 1020 1107 1076
rect 0 0 56 1020
rect 672 897 1893 899
rect 672 837 1812 897
rect 1872 837 1893 897
rect 672 835 1893 837
rect 672 0 728 835
rect 2338 766 2394 1845
rect 1456 710 2394 766
rect 2542 897 3237 899
rect 2542 837 3156 897
rect 3216 837 3237 897
rect 2542 835 3237 837
rect 1456 0 1512 710
rect 1696 645 2013 648
rect 1696 531 1709 645
rect 1997 531 2013 645
rect 2542 608 2598 835
rect 3313 618 3369 1845
rect 3471 897 4357 899
rect 3471 837 4276 897
rect 4336 837 4357 897
rect 3471 835 4357 837
rect 1696 444 1719 531
rect 1993 444 2013 531
rect 1696 425 2013 444
rect 2128 552 2598 608
rect 2800 562 3369 618
rect 2128 0 2184 552
rect 2800 0 2856 562
rect 3472 0 3528 835
rect 4740 722 4796 1845
rect 4927 897 5701 899
rect 4927 837 5620 897
rect 5680 837 5701 897
rect 4927 835 5701 837
rect 4144 666 4796 722
rect 4144 0 4200 666
rect 4928 0 4984 835
rect 6067 659 6123 1845
rect 6196 1530 6513 1545
rect 6196 1240 6209 1530
rect 6499 1240 6513 1530
rect 6196 1225 6513 1240
rect 5600 603 6123 659
rect 6272 897 6821 899
rect 6272 837 6740 897
rect 6800 837 6821 897
rect 6272 835 6821 837
rect 5600 0 5656 603
rect 6272 0 6328 835
rect 6944 0 7000 1845
rect 7728 899 7784 900
rect 7728 897 8165 899
rect 7728 837 8084 897
rect 8144 837 8165 897
rect 7728 835 8165 837
rect 7728 0 7784 835
rect 8400 0 8456 1845
rect 8866 897 9293 899
rect 8866 837 9204 897
rect 9264 837 9293 897
rect 8866 835 9293 837
rect 9072 0 9128 835
rect 9744 0 9800 1845
rect 10210 897 10628 899
rect 10210 837 10548 897
rect 10608 837 10628 897
rect 10210 835 10628 837
rect 10416 0 10472 835
rect 10696 645 11013 648
rect 10696 531 10709 645
rect 10997 531 11013 645
rect 10696 444 10719 531
rect 10993 444 11013 531
rect 10696 425 11013 444
rect 11200 0 11256 1845
rect 11330 897 11929 899
rect 11330 837 11668 897
rect 11728 837 11929 897
rect 11330 835 11929 837
rect 11872 0 11928 835
rect 12544 0 12600 1845
rect 12674 897 13271 899
rect 12674 837 13012 897
rect 13072 878 13271 897
rect 13072 837 13272 878
rect 12674 835 13272 837
rect 13216 0 13272 835
rect 13625 609 13681 1845
rect 13794 897 14728 899
rect 13794 837 14132 897
rect 14192 837 14728 897
rect 13794 835 14728 837
rect 13625 553 14056 609
rect 14000 0 14056 553
rect 14672 0 14728 835
rect 14978 709 15034 1845
rect 15196 1530 15513 1545
rect 15196 1240 15209 1530
rect 15499 1240 15513 1530
rect 15196 1225 15513 1240
rect 16715 1039 16771 1845
rect 16697 1037 16790 1039
rect 16697 977 16711 1037
rect 16771 977 16790 1037
rect 18070 1034 18126 1845
rect 19185 1039 19241 1845
rect 19171 1037 19255 1039
rect 16697 975 16790 977
rect 18056 1032 18140 1034
rect 18056 972 18068 1032
rect 18128 972 18140 1032
rect 19171 977 19183 1037
rect 19243 977 19255 1037
rect 20526 1034 20582 1845
rect 19171 974 19255 977
rect 20512 1032 20596 1034
rect 18056 970 18140 972
rect 20512 972 20524 1032
rect 20584 972 20596 1032
rect 20512 970 20596 972
rect 15138 897 16073 899
rect 15138 837 15476 897
rect 15536 837 16073 897
rect 15138 835 16073 837
rect 16258 897 17528 899
rect 16258 837 16596 897
rect 16656 837 17528 897
rect 16258 835 17528 837
rect 17602 897 18400 899
rect 17602 837 17940 897
rect 18000 837 18400 897
rect 17602 835 18400 837
rect 18720 897 19792 899
rect 18720 837 19060 897
rect 19120 837 19792 897
rect 18720 835 19792 837
rect 20066 897 21672 899
rect 20066 837 20404 897
rect 20464 837 21672 897
rect 20066 835 21672 837
rect 14978 653 15400 709
rect 15344 0 15400 653
rect 16016 0 16072 835
rect 16688 777 16790 779
rect 16688 717 16711 777
rect 16771 717 16790 777
rect 16688 715 16790 717
rect 16688 0 16744 715
rect 17472 0 17528 835
rect 18056 772 18200 774
rect 18056 712 18068 772
rect 18128 712 18200 772
rect 18056 710 18200 712
rect 18144 0 18200 710
rect 18344 731 18400 835
rect 19171 777 19544 779
rect 18344 675 18872 731
rect 19171 717 19183 777
rect 19243 723 19544 777
rect 19243 717 19255 723
rect 19171 714 19255 717
rect 18816 0 18872 675
rect 19488 0 19544 723
rect 19736 767 19792 835
rect 20512 772 20596 774
rect 19736 711 20328 767
rect 19696 645 20013 648
rect 19696 531 19709 645
rect 19997 531 20013 645
rect 19696 444 19719 531
rect 19993 444 20013 531
rect 19696 425 20013 444
rect 20272 0 20328 711
rect 20512 712 20524 772
rect 20584 769 20596 772
rect 20584 713 21000 769
rect 20584 712 20596 713
rect 20512 710 20596 712
rect 20944 0 21000 713
rect 21616 0 21672 835
<< via2 >>
rect 1707 2212 2000 2302
rect 1707 2098 2000 2212
rect 1707 2002 2000 2098
rect 10707 2212 11000 2302
rect 10707 2098 11000 2212
rect 10707 2002 11000 2098
rect 19707 2212 20000 2302
rect 19707 2098 20000 2212
rect 19707 2002 20000 2098
rect 1719 531 1993 639
rect 1719 444 1993 531
rect 6209 1432 6499 1530
rect 6209 1312 6499 1432
rect 6209 1240 6499 1312
rect 10719 531 10993 639
rect 10719 444 10993 531
rect 15209 1432 15499 1530
rect 15209 1312 15499 1432
rect 15209 1240 15499 1312
rect 19719 531 19993 639
rect 19719 444 19993 531
<< metal3 >>
rect 1696 2302 2014 2313
rect 1696 2002 1707 2302
rect 2000 2002 2014 2302
rect 1696 1993 2014 2002
rect 10696 2302 11014 2313
rect 10696 2002 10707 2302
rect 11000 2002 11014 2302
rect 10696 1993 11014 2002
rect 19696 2302 20014 2313
rect 19696 2002 19707 2302
rect 20000 2002 20014 2302
rect 19696 1993 20014 2002
rect 6196 1530 6513 1545
rect 6196 1240 6209 1530
rect 6499 1240 6513 1530
rect 6196 1225 6513 1240
rect 15196 1530 15513 1545
rect 15196 1240 15209 1530
rect 15499 1240 15513 1530
rect 15196 1225 15513 1240
rect 1696 733 2013 745
rect 1696 437 1710 733
rect 2002 437 2013 733
rect 1696 425 2013 437
rect 10696 733 11013 745
rect 10696 437 10710 733
rect 11002 437 11013 733
rect 10696 425 11013 437
rect 19696 733 20013 745
rect 19696 437 19710 733
rect 20002 437 20013 733
rect 19696 425 20013 437
<< via3 >>
rect 1707 2002 2000 2302
rect 10707 2002 11000 2302
rect 19707 2002 20000 2302
rect 6209 1240 6499 1530
rect 15209 1240 15499 1530
rect 1710 639 2002 733
rect 1710 444 1719 639
rect 1719 444 1993 639
rect 1993 444 2002 639
rect 1710 437 2002 444
rect 10710 639 11002 733
rect 10710 444 10719 639
rect 10719 444 10993 639
rect 10993 444 11002 639
rect 10710 437 11002 444
rect 19710 639 20002 733
rect 19710 444 19719 639
rect 19719 444 19993 639
rect 19993 444 20002 639
rect 19710 437 20002 444
<< metal4 >>
rect 1696 2302 2013 2313
rect 1696 2002 1707 2302
rect 2000 2002 2013 2302
rect 1696 733 2013 2002
rect 10696 2302 11013 2313
rect 10696 2002 10707 2302
rect 11000 2002 11013 2302
rect 6196 1530 6513 1545
rect 6196 1240 6209 1530
rect 6499 1240 6513 1530
rect 6196 1225 6513 1240
rect 1696 433 1709 733
rect 2002 433 2013 733
rect 1696 425 2013 433
rect 10696 733 11013 2002
rect 19696 2302 20013 2313
rect 19696 2002 19707 2302
rect 20000 2002 20013 2302
rect 15196 1530 15513 1545
rect 15196 1240 15209 1530
rect 15499 1240 15513 1530
rect 15196 1225 15513 1240
rect 10696 433 10709 733
rect 11002 433 11013 733
rect 10696 425 11013 433
rect 19696 733 20013 2002
rect 19696 433 19709 733
rect 20002 433 20013 733
rect 19696 425 20013 433
<< via4 >>
rect 1707 2002 2000 2302
rect 10707 2002 11000 2302
rect 6209 1240 6499 1530
rect 1709 437 1710 733
rect 1710 437 2002 733
rect 1709 433 2002 437
rect 19707 2002 20000 2302
rect 15209 1240 15499 1530
rect 10709 437 10710 733
rect 10710 437 11002 733
rect 10709 433 11002 437
rect 19709 437 19710 733
rect 19710 437 20002 733
rect 19709 433 20002 437
<< metal5 >>
rect 741 2302 20916 2313
rect 741 2002 1707 2302
rect 2000 2002 10707 2302
rect 11000 2002 19707 2302
rect 20000 2002 20916 2302
rect 741 1993 20916 2002
rect 741 1530 20916 1545
rect 741 1240 6209 1530
rect 6499 1240 15209 1530
rect 15499 1240 20916 1530
rect 741 1225 20916 1240
rect 741 733 20916 745
rect 741 433 1709 733
rect 2002 433 10709 733
rect 11002 433 19709 733
rect 20002 433 20916 733
rect 741 425 20916 433
use gf180mcu_fd_sc_mcu7t5v0__endcap  gf180mcu_fd_sc_mcu7t5v0__endcap_0 $PDKPATH/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654792614
transform 1 0 889 0 -1 2156
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  gf180mcu_fd_sc_mcu7t5v0__endcap_1
timestamp 1654792614
transform 1 0 20601 0 -1 2156
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  gf180mcu_fd_sc_mcu7t5v0__endcap_2
timestamp 1654792614
transform 1 0 20601 0 1 588
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  gf180mcu_fd_sc_mcu7t5v0__endcap_3
timestamp 1654792614
transform 1 0 889 0 1 588
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_0 $PDKPATH/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654792614
transform 1 0 14329 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_1
timestamp 1654792614
transform 1 0 11865 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_2
timestamp 1654792614
transform 1 0 16793 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_3
timestamp 1654792614
transform 1 0 9401 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_4
timestamp 1654792614
transform 1 0 19257 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_5
timestamp 1654792614
transform 1 0 6937 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_7
timestamp 1654792614
transform 1 0 4473 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_8
timestamp 1654792614
transform 1 0 2009 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_9
timestamp 1654792614
transform 1 0 2009 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_10
timestamp 1654792614
transform 1 0 4473 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_11
timestamp 1654792614
transform 1 0 6937 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_12
timestamp 1654792614
transform 1 0 9401 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_13
timestamp 1654792614
transform 1 0 11865 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_14
timestamp 1654792614
transform 1 0 14329 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_15
timestamp 1654792614
transform 1 0 16793 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  gf180mcu_fd_sc_mcu7t5v0__fillcap_4_16
timestamp 1654792614
transform 1 0 19257 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_0 $PDKPATH/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654792614
transform 1 0 13209 0 1 588
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_1
timestamp 1654792614
transform 1 0 15673 0 1 588
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_2
timestamp 1654792614
transform 1 0 18137 0 1 588
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_4
timestamp 1654792614
transform 1 0 10745 0 1 588
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_5
timestamp 1654792614
transform 1 0 8281 0 1 588
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_6
timestamp 1654792614
transform 1 0 5817 0 1 588
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_7
timestamp 1654792614
transform 1 0 3353 0 1 588
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_8
timestamp 1654792614
transform 1 0 3353 0 -1 2156
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_9
timestamp 1654792614
transform 1 0 5817 0 -1 2156
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_10
timestamp 1654792614
transform 1 0 8281 0 -1 2156
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_11
timestamp 1654792614
transform 1 0 10745 0 -1 2156
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_12
timestamp 1654792614
transform 1 0 13209 0 -1 2156
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_13
timestamp 1654792614
transform 1 0 15673 0 -1 2156
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  gf180mcu_fd_sc_mcu7t5v0__filltie_14
timestamp 1654792614
transform 1 0 18137 0 -1 2156
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_0 $PDKPATH/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654792614
transform 1 0 14777 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_1
timestamp 1654792614
transform 1 0 13433 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_2
timestamp 1654792614
transform 1 0 17241 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_3
timestamp 1654792614
transform 1 0 15897 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_4
timestamp 1654792614
transform 1 0 19705 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_5
timestamp 1654792614
transform 1 0 18361 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_8
timestamp 1654792614
transform 1 0 1113 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_9
timestamp 1654792614
transform 1 0 2457 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_10
timestamp 1654792614
transform 1 0 12313 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_11
timestamp 1654792614
transform 1 0 10969 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_12
timestamp 1654792614
transform 1 0 9849 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_13
timestamp 1654792614
transform 1 0 8505 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_14
timestamp 1654792614
transform 1 0 7385 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_15
timestamp 1654792614
transform 1 0 6041 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_16
timestamp 1654792614
transform 1 0 4921 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_17
timestamp 1654792614
transform 1 0 3577 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_18
timestamp 1654792614
transform 1 0 2457 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_19
timestamp 1654792614
transform 1 0 1113 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_20
timestamp 1654792614
transform 1 0 3577 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_21
timestamp 1654792614
transform 1 0 4921 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_22
timestamp 1654792614
transform 1 0 6041 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_23
timestamp 1654792614
transform 1 0 7385 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_24
timestamp 1654792614
transform 1 0 8505 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_25
timestamp 1654792614
transform 1 0 9849 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_26
timestamp 1654792614
transform 1 0 10969 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_27
timestamp 1654792614
transform 1 0 12313 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_28
timestamp 1654792614
transform 1 0 13433 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_29
timestamp 1654792614
transform 1 0 14777 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_30
timestamp 1654792614
transform 1 0 15897 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_31
timestamp 1654792614
transform 1 0 17241 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_32
timestamp 1654792614
transform 1 0 18361 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  gf180mcu_fd_sc_mcu7t5v0__tieh_33
timestamp 1654792614
transform 1 0 19705 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_0 $PDKPATH/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654792614
transform 1 0 15225 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_1
timestamp 1654792614
transform 1 0 13881 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_2
timestamp 1654792614
transform 1 0 17689 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_3
timestamp 1654792614
transform 1 0 16345 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_4
timestamp 1654792614
transform 1 0 20153 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_5
timestamp 1654792614
transform 1 0 18809 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_8
timestamp 1654792614
transform 1 0 1561 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_9
timestamp 1654792614
transform 1 0 2905 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_10
timestamp 1654792614
transform 1 0 12761 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_11
timestamp 1654792614
transform 1 0 11417 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_12
timestamp 1654792614
transform 1 0 10297 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_13
timestamp 1654792614
transform 1 0 8953 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_14
timestamp 1654792614
transform 1 0 7833 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_15
timestamp 1654792614
transform 1 0 6489 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_16
timestamp 1654792614
transform 1 0 5369 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_17
timestamp 1654792614
transform 1 0 4025 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_18
timestamp 1654792614
transform 1 0 2905 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_19
timestamp 1654792614
transform 1 0 1561 0 1 588
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_20
timestamp 1654792614
transform 1 0 4025 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_21
timestamp 1654792614
transform 1 0 5369 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_22
timestamp 1654792614
transform 1 0 6489 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_23
timestamp 1654792614
transform 1 0 7833 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_24
timestamp 1654792614
transform 1 0 8953 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_25
timestamp 1654792614
transform 1 0 10297 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_26
timestamp 1654792614
transform 1 0 11417 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_27
timestamp 1654792614
transform 1 0 12761 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_28
timestamp 1654792614
transform 1 0 13881 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_29
timestamp 1654792614
transform 1 0 15225 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_30
timestamp 1654792614
transform 1 0 16345 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_31
timestamp 1654792614
transform 1 0 17689 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_32
timestamp 1654792614
transform 1 0 18809 0 -1 2156
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  gf180mcu_fd_sc_mcu7t5v0__tiel_33
timestamp 1654792614
transform 1 0 20153 0 -1 2156
box -86 -86 534 870
<< labels >>
flabel metal5 741 1225 880 1545 0 FreeSans 1600 0 0 0 VDD
port 32 nsew
flabel metal5 741 425 880 745 0 FreeSans 1600 0 0 0 VSS
port 33 nsew
flabel metal2 21616 0 21672 410 0 FreeSans 400 90 0 0 mask_rev[31]
port 24 nsew
flabel metal2 20944 0 21000 410 0 FreeSans 400 90 0 0 mask_rev[30]
port 23 nsew
flabel metal2 20272 0 20328 410 0 FreeSans 400 90 0 0 mask_rev[29]
port 21 nsew
flabel metal2 19488 0 19544 410 0 FreeSans 400 90 0 0 mask_rev[28]
port 20 nsew
flabel metal2 18816 0 18872 410 0 FreeSans 400 90 0 0 mask_rev[27]
port 19 nsew
flabel metal2 18144 0 18200 410 0 FreeSans 400 90 0 0 mask_rev[26]
port 18 nsew
flabel metal2 17472 0 17528 410 0 FreeSans 400 90 0 0 mask_rev[25]
port 17 nsew
flabel metal2 16688 0 16744 410 0 FreeSans 400 90 0 0 mask_rev[24]
port 16 nsew
flabel metal2 16016 0 16072 410 0 FreeSans 400 90 0 0 mask_rev[23]
port 15 nsew
flabel metal2 15344 0 15400 410 0 FreeSans 400 90 0 0 mask_rev[22]
port 14 nsew
flabel metal2 14672 0 14728 410 0 FreeSans 400 90 0 0 mask_rev[21]
port 13 nsew
flabel metal2 14000 0 14056 410 0 FreeSans 400 90 0 0 mask_rev[20]
port 12 nsew
flabel metal2 13216 0 13272 410 0 FreeSans 400 90 0 0 mask_rev[19]
port 10 nsew
flabel metal2 12544 0 12600 410 0 FreeSans 400 90 0 0 mask_rev[18]
port 9 nsew
flabel metal2 11872 0 11928 410 0 FreeSans 400 90 0 0 mask_rev[17]
port 8 nsew
flabel metal2 11200 0 11256 410 0 FreeSans 400 90 0 0 mask_rev[16]
port 7 nsew
flabel metal2 10416 0 10472 410 0 FreeSans 400 90 0 0 mask_rev[15]
port 6 nsew
flabel metal2 9744 0 9800 410 0 FreeSans 400 90 0 0 mask_rev[14]
port 5 nsew
flabel metal2 9072 0 9128 410 0 FreeSans 400 90 0 0 mask_rev[13]
port 4 nsew
flabel metal2 8400 0 8456 410 0 FreeSans 400 90 0 0 mask_rev[12]
port 3 nsew
flabel metal2 7728 0 7784 410 0 FreeSans 400 90 0 0 mask_rev[11]
port 2 nsew
flabel metal2 6944 0 7000 410 0 FreeSans 400 90 0 0 mask_rev[10]
port 1 nsew
flabel metal2 6272 0 6328 410 0 FreeSans 400 90 0 0 mask_rev[9]
port 31 nsew
flabel metal2 5600 0 5656 410 0 FreeSans 400 90 0 0 mask_rev[8]
port 30 nsew
flabel metal2 4928 0 4984 410 0 FreeSans 400 90 0 0 mask_rev[7]
port 29 nsew
flabel metal2 4144 0 4200 410 0 FreeSans 400 90 0 0 mask_rev[6]
port 28 nsew
flabel metal2 3472 0 3528 410 0 FreeSans 400 90 0 0 mask_rev[5]
port 27 nsew
flabel metal2 2800 0 2856 410 0 FreeSans 400 90 0 0 mask_rev[4]
port 26 nsew
flabel metal2 2128 0 2184 410 0 FreeSans 400 90 0 0 mask_rev[3]
port 25 nsew
flabel metal2 1456 0 1512 410 0 FreeSans 400 90 0 0 mask_rev[2]
port 22 nsew
flabel metal2 672 0 728 410 0 FreeSans 400 90 0 0 mask_rev[1]
port 11 nsew
flabel metal2 0 0 56 410 0 FreeSans 400 90 0 0 mask_rev[0]
port 0 nsew
<< end >>
