VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO open_source
  CLASS BLOCK ;
  FOREIGN open_source ;
  ORIGIN -1.880 -12.910 ;
  SIZE 70.695 BY 27.695 ;
  OBS
      LAYER Metal5 ;
        POLYGON 15.300 39.150 15.300 38.700 14.850 38.700 ;
        RECT 15.300 38.700 19.800 40.050 ;
        POLYGON 19.800 39.150 20.250 38.700 19.800 38.700 ;
        POLYGON 14.850 37.800 14.850 37.350 14.400 37.350 ;
        RECT 14.850 37.350 20.250 38.700 ;
        POLYGON 20.250 37.800 20.700 37.350 20.250 37.350 ;
        POLYGON 8.095 37.350 8.095 36.455 7.200 36.455 ;
        POLYGON 8.095 37.350 8.545 36.900 8.095 36.900 ;
        RECT 8.095 36.455 8.995 36.900 ;
        RECT 7.200 36.450 8.995 36.455 ;
        POLYGON 8.995 36.900 9.445 36.450 8.995 36.450 ;
        RECT 14.400 36.450 20.700 37.350 ;
        POLYGON 27.005 37.350 27.005 36.900 26.555 36.900 ;
        POLYGON 26.105 36.900 26.105 36.450 25.655 36.450 ;
        RECT 26.105 36.455 27.005 36.900 ;
        POLYGON 27.005 37.350 27.900 36.455 27.005 36.455 ;
        RECT 26.105 36.450 27.900 36.455 ;
        POLYGON 7.200 36.450 7.200 34.650 5.400 34.650 ;
        RECT 7.200 36.000 9.895 36.450 ;
        POLYGON 9.895 36.450 10.345 36.000 9.895 36.000 ;
        POLYGON 13.945 36.450 13.945 36.000 13.495 36.000 ;
        RECT 13.945 36.000 21.155 36.450 ;
        RECT 7.200 35.100 10.795 36.000 ;
        POLYGON 10.795 36.000 11.695 35.100 10.795 35.100 ;
        POLYGON 13.495 36.000 13.495 35.550 13.045 35.550 ;
        RECT 13.495 35.550 21.155 36.000 ;
        POLYGON 21.155 36.450 22.055 35.550 21.155 35.550 ;
        POLYGON 25.205 36.450 25.205 36.000 24.755 36.000 ;
        RECT 25.205 36.000 27.900 36.450 ;
        POLYGON 24.305 36.000 24.305 35.550 23.855 35.550 ;
        RECT 24.305 35.550 27.900 36.000 ;
        POLYGON 12.145 35.550 12.145 35.100 11.695 35.100 ;
        RECT 12.145 35.100 22.955 35.550 ;
        POLYGON 22.955 35.550 23.405 35.100 22.955 35.100 ;
        POLYGON 23.855 35.550 23.855 35.100 23.405 35.100 ;
        RECT 23.855 35.100 27.900 35.550 ;
        RECT 7.200 34.650 27.900 35.100 ;
        POLYGON 27.900 36.450 29.700 34.650 27.900 34.650 ;
        POLYGON 5.400 34.650 6.300 34.650 6.300 33.750 ;
        RECT 6.300 33.300 28.800 34.650 ;
        POLYGON 28.800 34.650 29.700 34.650 28.800 33.750 ;
        POLYGON 6.300 33.300 7.650 33.300 7.650 31.950 ;
        POLYGON 7.650 30.600 7.650 30.150 7.200 30.150 ;
        RECT 7.650 30.150 27.450 33.300 ;
        POLYGON 27.450 33.300 28.800 33.300 27.450 31.950 ;
        POLYGON 27.450 30.600 27.900 30.150 27.450 30.150 ;
        RECT 35.280 30.505 36.780 30.805 ;
        RECT 38.880 30.505 40.380 30.805 ;
        RECT 42.180 30.505 44.280 30.805 ;
        RECT 45.480 30.505 47.580 30.805 ;
        RECT 51.480 30.505 53.580 30.805 ;
        RECT 55.080 30.505 56.580 30.805 ;
        RECT 34.980 30.205 37.080 30.505 ;
        RECT 38.580 30.205 40.680 30.505 ;
        RECT 7.200 29.700 16.200 30.150 ;
        POLYGON 16.200 30.150 16.650 30.150 16.200 29.700 ;
        POLYGON 18.450 30.150 18.900 30.150 18.900 29.700 ;
        RECT 18.900 29.700 27.900 30.150 ;
        POLYGON 7.200 29.250 7.200 28.350 6.300 28.350 ;
        RECT 7.200 28.350 13.500 29.700 ;
        POLYGON 4.500 28.350 4.500 27.900 4.050 27.900 ;
        RECT 4.500 27.900 13.500 28.350 ;
        RECT 2.700 23.850 13.500 27.900 ;
        POLYGON 13.500 29.700 15.750 29.700 13.500 27.450 ;
        POLYGON 19.350 29.700 21.600 29.700 21.600 27.450 ;
        RECT 21.600 28.350 27.900 29.700 ;
        RECT 34.680 29.605 37.380 30.205 ;
        POLYGON 27.900 29.250 28.800 28.350 27.900 28.350 ;
        RECT 21.600 27.900 30.600 28.350 ;
        POLYGON 30.600 28.350 31.050 27.900 30.600 27.900 ;
        RECT 21.600 23.850 32.400 27.900 ;
        RECT 34.680 27.505 35.580 29.605 ;
        RECT 36.480 27.505 37.380 29.605 ;
        RECT 34.680 26.905 37.380 27.505 ;
        RECT 38.280 29.605 40.980 30.205 ;
        RECT 38.280 27.505 39.180 29.605 ;
        RECT 40.080 27.505 40.980 29.605 ;
        RECT 38.280 26.905 40.980 27.505 ;
        RECT 41.880 29.905 44.580 30.505 ;
        RECT 41.880 29.005 42.780 29.905 ;
        RECT 43.680 29.005 44.580 29.905 ;
        RECT 41.880 28.405 44.580 29.005 ;
        RECT 45.480 30.205 47.880 30.505 ;
        RECT 51.180 30.205 53.580 30.505 ;
        RECT 54.780 30.205 56.880 30.505 ;
        RECT 45.480 29.605 48.180 30.205 ;
        RECT 41.880 28.105 44.280 28.405 ;
        RECT 41.880 27.205 42.780 28.105 ;
        RECT 34.980 26.605 37.080 26.905 ;
        RECT 38.280 26.605 40.680 26.905 ;
        RECT 41.880 26.605 44.580 27.205 ;
        RECT 35.280 26.305 36.780 26.605 ;
        RECT 38.280 26.305 40.380 26.605 ;
        RECT 42.180 26.305 44.580 26.605 ;
        RECT 45.480 26.305 46.380 29.605 ;
        RECT 47.280 26.305 48.180 29.605 ;
        RECT 50.880 29.905 53.580 30.205 ;
        RECT 50.880 29.005 52.080 29.905 ;
        RECT 54.480 29.605 57.180 30.205 ;
        RECT 50.880 28.705 52.980 29.005 ;
        RECT 51.180 28.405 53.280 28.705 ;
        RECT 51.480 28.105 53.580 28.405 ;
        RECT 52.380 27.205 53.580 28.105 ;
        RECT 50.880 26.905 53.580 27.205 ;
        RECT 54.480 27.505 55.380 29.605 ;
        RECT 56.280 27.505 57.180 29.605 ;
        RECT 54.480 26.905 57.180 27.505 ;
        RECT 58.080 27.505 58.980 30.805 ;
        RECT 59.880 27.505 60.780 30.805 ;
        RECT 58.080 26.905 60.780 27.505 ;
        RECT 61.680 30.505 63.780 30.805 ;
        RECT 65.880 30.505 67.380 30.805 ;
        RECT 69.180 30.505 71.280 30.805 ;
        RECT 61.680 30.205 64.080 30.505 ;
        RECT 65.580 30.205 67.680 30.505 ;
        RECT 61.680 29.605 64.380 30.205 ;
        RECT 50.880 26.605 53.280 26.905 ;
        RECT 54.780 26.605 56.880 26.905 ;
        RECT 58.380 26.605 60.480 26.905 ;
        RECT 50.880 26.305 52.980 26.605 ;
        RECT 55.080 26.305 56.580 26.605 ;
        RECT 58.680 26.305 60.180 26.605 ;
        RECT 61.680 26.305 62.580 29.605 ;
        RECT 63.480 29.005 64.380 29.605 ;
        RECT 65.280 29.605 67.980 30.205 ;
        RECT 65.280 27.505 66.180 29.605 ;
        RECT 67.080 29.005 67.980 29.605 ;
        RECT 68.880 29.905 71.580 30.505 ;
        RECT 68.880 29.005 69.780 29.905 ;
        RECT 70.680 29.005 71.580 29.905 ;
        RECT 68.880 28.405 71.580 29.005 ;
        RECT 68.880 28.105 71.280 28.405 ;
        RECT 67.080 27.505 67.980 28.105 ;
        RECT 65.280 26.905 67.980 27.505 ;
        RECT 68.880 27.205 69.780 28.105 ;
        RECT 65.580 26.605 67.680 26.905 ;
        RECT 68.880 26.605 71.580 27.205 ;
        RECT 65.880 26.305 67.380 26.605 ;
        RECT 69.180 26.305 71.580 26.605 ;
        RECT 38.280 24.505 39.180 26.305 ;
        RECT 50.880 24.505 51.780 26.305 ;
        RECT 38.280 24.205 40.380 24.505 ;
        RECT 41.880 24.205 44.280 24.505 ;
        RECT 45.480 24.205 47.580 24.505 ;
        RECT 49.680 24.205 51.780 24.505 ;
        RECT 38.280 23.905 40.680 24.205 ;
        POLYGON 4.050 23.850 4.500 23.850 4.500 23.400 ;
        RECT 4.500 23.400 13.500 23.850 ;
        POLYGON 5.850 23.400 6.750 23.400 6.750 22.500 ;
        RECT 6.750 22.050 13.500 23.400 ;
        POLYGON 13.500 23.850 15.300 22.050 13.500 22.050 ;
        RECT 6.750 21.600 15.300 22.050 ;
        POLYGON 6.750 21.600 7.200 21.600 7.200 21.150 ;
        RECT 7.200 21.150 15.300 21.600 ;
        RECT 7.200 20.700 14.850 21.150 ;
        POLYGON 14.850 21.150 15.300 21.150 14.850 20.700 ;
        POLYGON 21.600 23.850 21.600 22.050 19.800 22.050 ;
        RECT 21.600 23.400 30.600 23.850 ;
        POLYGON 30.600 23.850 31.050 23.850 30.600 23.400 ;
        RECT 21.600 22.050 28.350 23.400 ;
        POLYGON 28.350 23.400 29.250 23.400 28.350 22.500 ;
        RECT 38.280 23.305 40.980 23.905 ;
        RECT 41.880 23.605 44.580 24.205 ;
        RECT 19.800 21.600 28.350 22.050 ;
        RECT 19.800 21.150 27.900 21.600 ;
        POLYGON 27.900 21.600 28.350 21.600 27.900 21.150 ;
        POLYGON 19.800 21.150 20.250 21.150 20.250 20.700 ;
        RECT 20.250 20.700 27.900 21.150 ;
        POLYGON 7.200 20.700 7.650 20.700 7.650 20.250 ;
        POLYGON 7.650 20.250 7.650 19.800 7.200 19.800 ;
        RECT 7.650 19.800 14.850 20.700 ;
        POLYGON 7.200 19.350 7.200 18.450 6.300 18.450 ;
        RECT 7.200 18.900 14.400 19.800 ;
        POLYGON 14.400 19.800 14.850 19.800 14.400 19.350 ;
        RECT 20.250 19.800 27.450 20.700 ;
        POLYGON 27.450 20.700 27.900 20.700 27.450 20.250 ;
        POLYGON 27.450 20.250 27.900 19.800 27.450 19.800 ;
        RECT 38.280 20.005 39.180 23.305 ;
        RECT 40.080 20.005 40.980 23.305 ;
        RECT 43.680 22.705 44.580 23.605 ;
        RECT 41.880 21.805 44.580 22.705 ;
        RECT 41.880 20.905 42.780 21.805 ;
        RECT 43.680 20.905 44.580 21.805 ;
        RECT 41.880 20.305 44.580 20.905 ;
        RECT 42.180 20.005 44.580 20.305 ;
        RECT 45.480 23.905 47.880 24.205 ;
        RECT 49.380 23.905 51.780 24.205 ;
        RECT 45.480 23.305 48.180 23.905 ;
        RECT 45.480 20.005 46.380 23.305 ;
        RECT 47.280 22.705 48.180 23.305 ;
        RECT 49.080 23.305 51.780 23.905 ;
        RECT 49.080 21.205 49.980 23.305 ;
        RECT 50.880 21.205 51.780 23.305 ;
        RECT 49.080 20.605 51.780 21.205 ;
        RECT 52.680 21.205 53.580 24.505 ;
        RECT 54.480 21.205 55.380 24.505 ;
        RECT 56.280 21.205 57.180 24.505 ;
        RECT 58.080 24.205 60.480 24.505 ;
        RECT 61.680 24.205 63.780 24.505 ;
        RECT 65.580 24.205 67.680 24.505 ;
        RECT 58.080 23.605 60.780 24.205 ;
        RECT 59.880 22.705 60.780 23.605 ;
        RECT 58.380 22.405 60.780 22.705 ;
        RECT 52.680 20.605 57.180 21.205 ;
        RECT 58.080 21.805 60.780 22.405 ;
        RECT 58.080 20.905 58.980 21.805 ;
        RECT 59.880 20.905 60.780 21.805 ;
        RECT 49.380 20.305 51.780 20.605 ;
        RECT 52.980 20.305 56.880 20.605 ;
        RECT 58.080 20.305 60.780 20.905 ;
        RECT 49.680 20.005 51.780 20.305 ;
        RECT 53.280 20.005 54.480 20.305 ;
        RECT 55.380 20.005 56.580 20.305 ;
        RECT 58.380 20.005 60.780 20.305 ;
        RECT 61.680 23.905 64.080 24.205 ;
        RECT 61.680 23.305 64.380 23.905 ;
        RECT 61.680 20.005 62.580 23.305 ;
        RECT 63.480 22.705 64.380 23.305 ;
        RECT 65.280 23.605 67.980 24.205 ;
        RECT 65.280 22.705 66.180 23.605 ;
        RECT 67.080 22.705 67.980 23.605 ;
        RECT 65.280 21.805 67.980 22.705 ;
        RECT 65.280 20.905 66.180 21.805 ;
        RECT 65.280 20.305 67.980 20.905 ;
        RECT 65.580 20.005 67.980 20.305 ;
        POLYGON 20.250 19.800 20.700 19.800 20.700 19.350 ;
        RECT 7.200 18.450 13.950 18.900 ;
        POLYGON 13.950 18.900 14.400 18.900 13.950 18.450 ;
        RECT 20.700 18.900 27.900 19.800 ;
        POLYGON 20.700 18.900 21.150 18.900 21.150 18.450 ;
        RECT 21.150 18.450 27.900 18.900 ;
        POLYGON 27.900 19.350 28.800 18.450 27.900 18.450 ;
        POLYGON 6.300 18.000 6.300 17.100 5.400 17.100 ;
        RECT 6.300 17.550 13.950 18.450 ;
        RECT 6.300 17.100 13.500 17.550 ;
        POLYGON 13.500 17.550 13.950 17.550 13.500 17.100 ;
        RECT 21.150 17.550 28.800 18.450 ;
        POLYGON 21.150 17.550 21.600 17.550 21.600 17.100 ;
        RECT 21.600 17.100 28.800 17.550 ;
        POLYGON 28.800 18.000 29.700 17.100 28.800 17.100 ;
        POLYGON 5.400 17.100 8.100 17.100 8.100 14.400 ;
        RECT 8.100 16.650 13.500 17.100 ;
        RECT 8.100 16.200 13.170 16.650 ;
        POLYGON 13.170 16.650 13.500 16.650 13.170 16.320 ;
        RECT 21.600 16.650 27.000 17.100 ;
        POLYGON 21.600 16.650 21.930 16.650 21.930 16.320 ;
        RECT 8.100 15.750 10.800 16.200 ;
        POLYGON 10.800 16.200 11.250 16.200 10.800 15.750 ;
        POLYGON 11.575 16.200 12.025 16.200 12.025 15.750 ;
        RECT 12.025 15.870 13.170 16.200 ;
        RECT 12.025 15.750 12.600 15.870 ;
        RECT 8.100 15.300 9.900 15.750 ;
        POLYGON 9.900 15.750 10.350 15.750 9.900 15.300 ;
        POLYGON 12.025 15.750 12.475 15.750 12.475 15.300 ;
        RECT 12.475 15.300 12.600 15.750 ;
        POLYGON 12.600 15.870 13.170 15.870 12.600 15.300 ;
        RECT 21.930 16.200 27.000 16.650 ;
        RECT 21.930 15.870 22.625 16.200 ;
        POLYGON 21.930 15.870 22.500 15.870 22.500 15.300 ;
        RECT 22.500 15.300 22.625 15.870 ;
        POLYGON 22.625 16.200 23.525 16.200 22.625 15.300 ;
        POLYGON 23.850 16.200 24.300 16.200 24.300 15.750 ;
        RECT 24.300 15.750 27.000 16.200 ;
        POLYGON 24.750 15.750 25.200 15.750 25.200 15.300 ;
        RECT 25.200 15.300 27.000 15.750 ;
        RECT 8.100 14.400 8.550 15.300 ;
        POLYGON 8.550 15.300 9.450 15.300 8.550 14.400 ;
        POLYGON 25.650 15.300 26.550 15.300 26.550 14.400 ;
        RECT 26.550 14.400 27.000 15.300 ;
        POLYGON 27.000 17.100 29.700 17.100 27.000 14.400 ;
  END
END open_source
END LIBRARY

