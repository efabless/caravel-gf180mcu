magic
tech micross
timestamp 1679504633
<< pi1 >>
tri 53750 505270 54280 505800 se
rect 54280 505270 57220 505800
tri 57220 505270 57750 505800 sw
rect 53750 502330 57750 505270
tri 53750 501800 54280 502330 ne
rect 54280 501800 57220 502330
tri 57220 501800 57750 502330 nw
tri 81250 505270 81780 505800 se
rect 81780 505270 84720 505800
tri 84720 505270 85250 505800 sw
rect 81250 502330 85250 505270
tri 81250 501800 81780 502330 ne
rect 81780 501800 84720 502330
tri 84720 501800 85250 502330 nw
tri 108750 505270 109280 505800 se
rect 109280 505270 112220 505800
tri 112220 505270 112750 505800 sw
rect 108750 502330 112750 505270
tri 108750 501800 109280 502330 ne
rect 109280 501800 112220 502330
tri 112220 501800 112750 502330 nw
tri 136250 505270 136780 505800 se
rect 136780 505270 139720 505800
tri 139720 505270 140250 505800 sw
rect 136250 502330 140250 505270
tri 136250 501800 136780 502330 ne
rect 136780 501800 139720 502330
tri 139720 501800 140250 502330 nw
tri 163750 505270 164280 505800 se
rect 164280 505270 167220 505800
tri 167220 505270 167750 505800 sw
rect 163750 502330 167750 505270
tri 163750 501800 164280 502330 ne
rect 164280 501800 167220 502330
tri 167220 501800 167750 502330 nw
tri 191250 505270 191780 505800 se
rect 191780 505270 194720 505800
tri 194720 505270 195250 505800 sw
rect 191250 502330 195250 505270
tri 191250 501800 191780 502330 ne
rect 191780 501800 194720 502330
tri 194720 501800 195250 502330 nw
tri 218750 505270 219280 505800 se
rect 219280 505270 222220 505800
tri 222220 505270 222750 505800 sw
rect 218750 502330 222750 505270
tri 218750 501800 219280 502330 ne
rect 219280 501800 222220 502330
tri 222220 501800 222750 502330 nw
tri 246250 505270 246780 505800 se
rect 246780 505270 249720 505800
tri 249720 505270 250250 505800 sw
rect 246250 502330 250250 505270
tri 246250 501800 246780 502330 ne
rect 246780 501800 249720 502330
tri 249720 501800 250250 502330 nw
tri 273750 505270 274280 505800 se
rect 274280 505270 277220 505800
tri 277220 505270 277750 505800 sw
rect 273750 502330 277750 505270
tri 273750 501800 274280 502330 ne
rect 274280 501800 277220 502330
tri 277220 501800 277750 502330 nw
tri 301250 505270 301780 505800 se
rect 301780 505270 304720 505800
tri 304720 505270 305250 505800 sw
rect 301250 502330 305250 505270
tri 301250 501800 301780 502330 ne
rect 301780 501800 304720 502330
tri 304720 501800 305250 502330 nw
tri 328750 505270 329280 505800 se
rect 329280 505270 332220 505800
tri 332220 505270 332750 505800 sw
rect 328750 502330 332750 505270
tri 328750 501800 329280 502330 ne
rect 329280 501800 332220 502330
tri 332220 501800 332750 502330 nw
tri 1200 457720 1730 458250 se
rect 1730 457720 4670 458250
tri 4670 457720 5200 458250 sw
rect 1200 454780 5200 457720
tri 1200 454250 1730 454780 ne
rect 1730 454250 4670 454780
tri 4670 454250 5200 454780 nw
tri 382800 458220 383330 458750 se
rect 383330 458220 386270 458750
tri 386270 458220 386800 458750 sw
rect 382800 455280 386800 458220
tri 382800 454750 383330 455280 ne
rect 383330 454750 386270 455280
tri 386270 454750 386800 455280 nw
tri 1200 437220 1730 437750 se
rect 1730 437220 4670 437750
tri 4670 437220 5200 437750 sw
rect 1200 434280 5200 437220
tri 1200 433750 1730 434280 ne
rect 1730 433750 4670 434280
tri 4670 433750 5200 434280 nw
tri 382800 436720 383330 437250 se
rect 383330 436720 386270 437250
tri 386270 436720 386800 437250 sw
rect 382800 433780 386800 436720
tri 382800 433250 383330 433780 ne
rect 383330 433250 386270 433780
tri 386270 433250 386800 433780 nw
tri 1200 416720 1730 417250 se
rect 1730 416720 4670 417250
tri 4670 416720 5200 417250 sw
rect 1200 413780 5200 416720
tri 1200 413250 1730 413780 ne
rect 1730 413250 4670 413780
tri 4670 413250 5200 413780 nw
tri 382800 415220 383330 415750 se
rect 383330 415220 386270 415750
tri 386270 415220 386800 415750 sw
rect 382800 412280 386800 415220
tri 382800 411750 383330 412280 ne
rect 383330 411750 386270 412280
tri 386270 411750 386800 412280 nw
tri 1200 396220 1730 396750 se
rect 1730 396220 4670 396750
tri 4670 396220 5200 396750 sw
rect 1200 393280 5200 396220
tri 1200 392750 1730 393280 ne
rect 1730 392750 4670 393280
tri 4670 392750 5200 393280 nw
tri 382800 393720 383330 394250 se
rect 383330 393720 386270 394250
tri 386270 393720 386800 394250 sw
rect 382800 390780 386800 393720
tri 382800 390250 383330 390780 ne
rect 383330 390250 386270 390780
tri 386270 390250 386800 390780 nw
tri 1200 375720 1730 376250 se
rect 1730 375720 4670 376250
tri 4670 375720 5200 376250 sw
rect 1200 372780 5200 375720
tri 1200 372250 1730 372780 ne
rect 1730 372250 4670 372780
tri 4670 372250 5200 372780 nw
tri 382800 372220 383330 372750 se
rect 383330 372220 386270 372750
tri 386270 372220 386800 372750 sw
rect 382800 369280 386800 372220
tri 382800 368750 383330 369280 ne
rect 383330 368750 386270 369280
tri 386270 368750 386800 369280 nw
tri 1200 355220 1730 355750 se
rect 1730 355220 4670 355750
tri 4670 355220 5200 355750 sw
rect 1200 352280 5200 355220
tri 1200 351750 1730 352280 ne
rect 1730 351750 4670 352280
tri 4670 351750 5200 352280 nw
tri 382800 350720 383330 351250 se
rect 383330 350720 386270 351250
tri 386270 350720 386800 351250 sw
rect 382800 347780 386800 350720
tri 382800 347250 383330 347780 ne
rect 383330 347250 386270 347780
tri 386270 347250 386800 347780 nw
tri 1200 334720 1730 335250 se
rect 1730 334720 4670 335250
tri 4670 334720 5200 335250 sw
rect 1200 331780 5200 334720
tri 1200 331250 1730 331780 ne
rect 1730 331250 4670 331780
tri 4670 331250 5200 331780 nw
tri 382800 329220 383330 329750 se
rect 383330 329220 386270 329750
tri 386270 329220 386800 329750 sw
rect 382800 326280 386800 329220
tri 382800 325750 383330 326280 ne
rect 383330 325750 386270 326280
tri 386270 325750 386800 326280 nw
tri 1200 314220 1730 314750 se
rect 1730 314220 4670 314750
tri 4670 314220 5200 314750 sw
rect 1200 311280 5200 314220
tri 1200 310750 1730 311280 ne
rect 1730 310750 4670 311280
tri 4670 310750 5200 311280 nw
tri 382800 307720 383330 308250 se
rect 383330 307720 386270 308250
tri 386270 307720 386800 308250 sw
rect 382800 304780 386800 307720
tri 382800 304250 383330 304780 ne
rect 383330 304250 386270 304780
tri 386270 304250 386800 304780 nw
tri 1200 293720 1730 294250 se
rect 1730 293720 4670 294250
tri 4670 293720 5200 294250 sw
rect 1200 290780 5200 293720
tri 1200 290250 1730 290780 ne
rect 1730 290250 4670 290780
tri 4670 290250 5200 290780 nw
tri 382800 286220 383330 286750 se
rect 383330 286220 386270 286750
tri 386270 286220 386800 286750 sw
rect 382800 283280 386800 286220
tri 382800 282750 383330 283280 ne
rect 383330 282750 386270 283280
tri 386270 282750 386800 283280 nw
tri 1200 273220 1730 273750 se
rect 1730 273220 4670 273750
tri 4670 273220 5200 273750 sw
rect 1200 270280 5200 273220
tri 1200 269750 1730 270280 ne
rect 1730 269750 4670 270280
tri 4670 269750 5200 270280 nw
tri 382800 264720 383330 265250 se
rect 383330 264720 386270 265250
tri 386270 264720 386800 265250 sw
rect 382800 261780 386800 264720
tri 382800 261250 383330 261780 ne
rect 383330 261250 386270 261780
tri 386270 261250 386800 261780 nw
tri 1200 252720 1730 253250 se
rect 1730 252720 4670 253250
tri 4670 252720 5200 253250 sw
rect 1200 249780 5200 252720
tri 1200 249250 1730 249780 ne
rect 1730 249250 4670 249780
tri 4670 249250 5200 249780 nw
tri 382800 243220 383330 243750 se
rect 383330 243220 386270 243750
tri 386270 243220 386800 243750 sw
rect 382800 240280 386800 243220
tri 382800 239750 383330 240280 ne
rect 383330 239750 386270 240280
tri 386270 239750 386800 240280 nw
tri 1200 232220 1730 232750 se
rect 1730 232220 4670 232750
tri 4670 232220 5200 232750 sw
rect 1200 229280 5200 232220
tri 1200 228750 1730 229280 ne
rect 1730 228750 4670 229280
tri 4670 228750 5200 229280 nw
tri 382800 221720 383330 222250 se
rect 383330 221720 386270 222250
tri 386270 221720 386800 222250 sw
rect 382800 218780 386800 221720
tri 382800 218250 383330 218780 ne
rect 383330 218250 386270 218780
tri 386270 218250 386800 218780 nw
tri 1200 211720 1730 212250 se
rect 1730 211720 4670 212250
tri 4670 211720 5200 212250 sw
rect 1200 208780 5200 211720
tri 1200 208250 1730 208780 ne
rect 1730 208250 4670 208780
tri 4670 208250 5200 208780 nw
tri 382800 200220 383330 200750 se
rect 383330 200220 386270 200750
tri 386270 200220 386800 200750 sw
rect 382800 197280 386800 200220
tri 382800 196750 383330 197280 ne
rect 383330 196750 386270 197280
tri 386270 196750 386800 197280 nw
tri 1200 191220 1730 191750 se
rect 1730 191220 4670 191750
tri 4670 191220 5200 191750 sw
rect 1200 188280 5200 191220
tri 1200 187750 1730 188280 ne
rect 1730 187750 4670 188280
tri 4670 187750 5200 188280 nw
tri 382800 178720 383330 179250 se
rect 383330 178720 386270 179250
tri 386270 178720 386800 179250 sw
rect 382800 175780 386800 178720
tri 382800 175250 383330 175780 ne
rect 383330 175250 386270 175780
tri 386270 175250 386800 175780 nw
tri 1200 170720 1730 171250 se
rect 1730 170720 4670 171250
tri 4670 170720 5200 171250 sw
rect 1200 167780 5200 170720
tri 1200 167250 1730 167780 ne
rect 1730 167250 4670 167780
tri 4670 167250 5200 167780 nw
tri 382800 157220 383330 157750 se
rect 383330 157220 386270 157750
tri 386270 157220 386800 157750 sw
rect 382800 154280 386800 157220
tri 382800 153750 383330 154280 ne
rect 383330 153750 386270 154280
tri 386270 153750 386800 154280 nw
tri 1200 150220 1730 150750 se
rect 1730 150220 4670 150750
tri 4670 150220 5200 150750 sw
rect 1200 147280 5200 150220
tri 1200 146750 1730 147280 ne
rect 1730 146750 4670 147280
tri 4670 146750 5200 147280 nw
tri 382800 135720 383330 136250 se
rect 383330 135720 386270 136250
tri 386270 135720 386800 136250 sw
rect 382800 132780 386800 135720
tri 382800 132250 383330 132780 ne
rect 383330 132250 386270 132780
tri 386270 132250 386800 132780 nw
tri 1200 129720 1730 130250 se
rect 1730 129720 4670 130250
tri 4670 129720 5200 130250 sw
rect 1200 126780 5200 129720
tri 1200 126250 1730 126780 ne
rect 1730 126250 4670 126780
tri 4670 126250 5200 126780 nw
tri 382800 114220 383330 114750 se
rect 383330 114220 386270 114750
tri 386270 114220 386800 114750 sw
rect 382800 111280 386800 114220
tri 382800 110750 383330 111280 ne
rect 383330 110750 386270 111280
tri 386270 110750 386800 111280 nw
tri 1200 109220 1730 109750 se
rect 1730 109220 4670 109750
tri 4670 109220 5200 109750 sw
rect 1200 106280 5200 109220
tri 1200 105750 1730 106280 ne
rect 1730 105750 4670 106280
tri 4670 105750 5200 106280 nw
tri 382800 92720 383330 93250 se
rect 383330 92720 386270 93250
tri 386270 92720 386800 93250 sw
rect 382800 89780 386800 92720
tri 382800 89250 383330 89780 ne
rect 383330 89250 386270 89780
tri 386270 89250 386800 89780 nw
tri 1200 88720 1730 89250 se
rect 1730 88720 4670 89250
tri 4670 88720 5200 89250 sw
rect 1200 85780 5200 88720
tri 1200 85250 1730 85780 ne
rect 1730 85250 4670 85780
tri 4670 85250 5200 85780 nw
tri 382800 71220 383330 71750 se
rect 383330 71220 386270 71750
tri 386270 71220 386800 71750 sw
tri 1200 68220 1730 68750 se
rect 1730 68220 4670 68750
tri 4670 68220 5200 68750 sw
rect 1200 65280 5200 68220
rect 382800 68280 386800 71220
tri 382800 67750 383330 68280 ne
rect 383330 67750 386270 68280
tri 386270 67750 386800 68280 nw
tri 1200 64750 1730 65280 ne
rect 1730 64750 4670 65280
tri 4670 64750 5200 65280 nw
tri 382800 49720 383330 50250 se
rect 383330 49720 386270 50250
tri 386270 49720 386800 50250 sw
tri 1200 47720 1730 48250 se
rect 1730 47720 4670 48250
tri 4670 47720 5200 48250 sw
rect 1200 44780 5200 47720
rect 382800 46780 386800 49720
tri 382800 46250 383330 46780 ne
rect 383330 46250 386270 46780
tri 386270 46250 386800 46780 nw
tri 1200 44250 1730 44780 ne
rect 1730 44250 4670 44780
tri 4670 44250 5200 44780 nw
tri 54250 4670 54780 5200 se
rect 54780 4670 57720 5200
tri 57720 4670 58250 5200 sw
rect 54250 1730 58250 4670
tri 54250 1200 54780 1730 ne
rect 54780 1200 57720 1730
tri 57720 1200 58250 1730 nw
tri 81750 4670 82280 5200 se
rect 82280 4670 85220 5200
tri 85220 4670 85750 5200 sw
rect 81750 1730 85750 4670
tri 81750 1200 82280 1730 ne
rect 82280 1200 85220 1730
tri 85220 1200 85750 1730 nw
tri 109250 4670 109780 5200 se
rect 109780 4670 112720 5200
tri 112720 4670 113250 5200 sw
rect 109250 1730 113250 4670
tri 109250 1200 109780 1730 ne
rect 109780 1200 112720 1730
tri 112720 1200 113250 1730 nw
tri 136750 4670 137280 5200 se
rect 137280 4670 140220 5200
tri 140220 4670 140750 5200 sw
rect 136750 1730 140750 4670
tri 136750 1200 137280 1730 ne
rect 137280 1200 140220 1730
tri 140220 1200 140750 1730 nw
tri 164250 4670 164780 5200 se
rect 164780 4670 167720 5200
tri 167720 4670 168250 5200 sw
rect 164250 1730 168250 4670
tri 164250 1200 164780 1730 ne
rect 164780 1200 167720 1730
tri 167720 1200 168250 1730 nw
tri 191750 4670 192280 5200 se
rect 192280 4670 195220 5200
tri 195220 4670 195750 5200 sw
rect 191750 1730 195750 4670
tri 191750 1200 192280 1730 ne
rect 192280 1200 195220 1730
tri 195220 1200 195750 1730 nw
tri 219250 4670 219780 5200 se
rect 219780 4670 222720 5200
tri 222720 4670 223250 5200 sw
rect 219250 1730 223250 4670
tri 219250 1200 219780 1730 ne
rect 219780 1200 222720 1730
tri 222720 1200 223250 1730 nw
tri 246750 4670 247280 5200 se
rect 247280 4670 250220 5200
tri 250220 4670 250750 5200 sw
rect 246750 1730 250750 4670
tri 246750 1200 247280 1730 ne
rect 247280 1200 250220 1730
tri 250220 1200 250750 1730 nw
tri 274250 4670 274780 5200 se
rect 274780 4670 277720 5200
tri 277720 4670 278250 5200 sw
rect 274250 1730 278250 4670
tri 274250 1200 274780 1730 ne
rect 274780 1200 277720 1730
tri 277720 1200 278250 1730 nw
tri 301750 4670 302280 5200 se
rect 302280 4670 305220 5200
tri 305220 4670 305750 5200 sw
rect 301750 1730 305750 4670
tri 301750 1200 302280 1730 ne
rect 302280 1200 305220 1730
tri 305220 1200 305750 1730 nw
tri 329250 4670 329780 5200 se
rect 329780 4670 332720 5200
tri 332720 4670 333250 5200 sw
rect 329250 1730 333250 4670
tri 329250 1200 329780 1730 ne
rect 329780 1200 332720 1730
tri 332720 1200 333250 1730 nw
<< rdl >>
tri 52906 506249 53457 506800 se
rect 53457 506249 58043 506800
tri 58043 506249 58594 506800 sw
tri 80785 506628 80957 506800 se
rect 80957 506628 85543 506800
tri 85543 506628 85715 506800 sw
tri 80422 506265 80785 506628 se
rect 80785 506265 85715 506628
tri 52750 506093 52906 506249 se
rect 52906 506093 58594 506249
tri 58594 506093 58750 506249 sw
rect 52750 501507 58750 506093
tri 52750 500956 53301 501507 ne
rect 53301 501263 58506 501507
tri 58506 501263 58750 501507 nw
tri 80250 506093 80422 506265 se
rect 80422 506138 85715 506265
tri 85715 506138 86205 506628 sw
tri 108284 506627 108457 506800 se
rect 108457 506627 113043 506800
tri 113043 506627 113216 506800 sw
tri 107923 506266 108284 506627 se
rect 108284 506266 113216 506627
rect 80422 506093 86205 506138
tri 86205 506093 86250 506138 sw
rect 80250 501507 86250 506093
tri 107750 506093 107923 506266 se
rect 107923 506098 113216 506266
tri 113216 506098 113745 506627 sw
tri 135783 506626 135957 506800 se
rect 135957 506626 140543 506800
tri 140543 506626 140717 506800 sw
tri 135424 506267 135783 506626 se
rect 135783 506267 140717 506626
rect 107923 506093 113745 506098
tri 113745 506093 113750 506098 sw
tri 80250 501335 80422 501507 ne
rect 80422 501462 86250 501507
tri 86250 501462 88582 503696 sw
rect 107750 501507 113750 506093
tri 135250 506093 135424 506267 se
rect 135424 506093 140717 506267
tri 140717 506093 141250 506626 sw
tri 163278 506621 163457 506800 se
rect 163457 506621 168043 506800
tri 162929 506272 163278 506621 se
rect 163278 506272 168043 506621
rect 80422 501335 88582 501462
rect 53301 500956 58500 501263
tri 58500 501257 58506 501263 nw
tri 53301 500800 53457 500956 ne
rect 53457 500800 58500 500956
tri 80422 500800 80957 501335 ne
rect 80957 500800 88582 501335
tri 88582 500800 89273 501462 sw
tri 107750 501334 107923 501507 ne
rect 107923 501502 113750 501507
tri 113750 501502 116091 503716 sw
rect 135250 503685 141250 506093
tri 162750 506093 162929 506272 se
rect 162929 506093 168043 506272
tri 168043 506093 168750 506800 sw
tri 190406 506249 190957 506800 se
rect 190957 506249 195543 506800
tri 195543 506249 196094 506800 sw
tri 218213 506556 218457 506800 se
rect 218457 506556 223043 506800
tri 223043 506556 223287 506800 sw
tri 245768 506611 245957 506800 se
rect 245957 506611 250543 506800
tri 250543 506611 250732 506800 sw
tri 273278 506621 273457 506800 se
rect 273457 506621 278043 506800
tri 278043 506621 278222 506800 sw
tri 300781 506624 300957 506800 se
rect 300957 506624 305543 506800
tri 305543 506624 305719 506800 sw
tri 141250 503685 141326 503755 sw
rect 135250 501507 141326 503685
rect 107923 501334 116091 501502
tri 107923 500800 108457 501334 ne
rect 108457 501333 116091 501334
tri 116091 501333 116270 501502 sw
tri 135250 501333 135424 501507 ne
rect 135424 501333 141326 501507
rect 108457 500800 116270 501333
tri 116270 500800 116833 501333 sw
tri 135424 500800 135957 501333 ne
rect 135957 500800 141326 501333
tri 141326 500800 144456 503685 sw
rect 162750 501917 168750 506093
tri 190250 506093 190406 506249 se
rect 190406 506093 196094 506249
tri 196094 506093 196250 506249 sw
tri 168750 501917 171000 503855 sw
rect 162750 501507 171000 501917
tri 162750 501328 162929 501507 ne
rect 162929 501328 171000 501507
tri 162929 500800 163457 501328 ne
rect 163457 500800 171000 501328
rect 190250 501507 196250 506093
tri 217750 506093 218213 506556 se
rect 218213 506337 223287 506556
tri 223287 506337 223506 506556 sw
rect 218213 506093 223506 506337
tri 223506 506093 223750 506337 sw
tri 190250 500956 190801 501507 ne
rect 190801 501263 196006 501507
tri 196006 501263 196250 501507 nw
tri 217000 501574 217750 502774 se
rect 217750 501574 223750 506093
tri 245250 506093 245768 506611 se
rect 245768 506282 250732 506611
tri 250732 506282 251061 506611 sw
rect 245768 506093 251061 506282
tri 251061 506093 251250 506282 sw
rect 217000 501507 223750 501574
rect 217000 501263 223506 501507
tri 223506 501263 223750 501507 nw
rect 190801 500956 196000 501263
tri 196000 501257 196006 501263 nw
tri 190801 500800 190957 500956 ne
rect 190957 500800 196000 500956
tri 54483 500737 54500 500800 ne
rect 54500 490172 58500 500800
tri 83490 500737 83556 500800 ne
rect 83556 500737 89273 500800
tri 89273 500737 89339 500800 sw
tri 111012 500737 111079 500800 ne
rect 111079 500737 116833 500800
tri 116833 500737 116900 500800 sw
tri 138554 500737 138622 500800 ne
rect 138622 500737 144456 500800
tri 144456 500737 144524 500800 sw
tri 166167 500737 166240 500800 ne
rect 166240 500737 171000 500800
tri 191983 500737 192000 500800 ne
tri 83556 498199 86205 500737 ne
rect 86205 498199 89339 500737
tri 89339 498199 91988 500737 sw
tri 111079 498245 113715 500737 ne
rect 113715 500643 116900 500737
tri 116900 500643 117000 500737 sw
rect 113715 498245 117000 500643
tri 117000 498245 119536 500643 sw
tri 138622 498245 141326 500737 ne
rect 141326 499377 144524 500737
tri 144524 499377 146000 500737 sw
tri 166240 500083 167000 500737 ne
rect 141326 498245 146000 499377
tri 113715 498217 113745 498245 ne
rect 113745 498217 119536 498245
tri 119536 498217 119565 498245 sw
tri 113745 498199 113764 498217 ne
rect 113764 498199 119565 498217
tri 119565 498199 119584 498217 sw
tri 141326 498199 141375 498245 ne
rect 141375 498199 146000 498245
tri 86205 492658 91988 498199 ne
tri 91988 494354 96000 498199 sw
tri 113764 497623 114373 498199 ne
rect 114373 497623 119584 498199
tri 119584 497623 120194 498199 sw
tri 141375 497623 142000 498199 ne
tri 114373 495139 117000 497623 ne
rect 117000 496861 120194 497623
tri 120194 496861 121000 497623 sw
rect 91988 492658 96000 494354
tri 91988 492646 92000 492658 ne
tri 58500 490172 60156 491828 sw
tri 54500 484516 60156 490172 ne
tri 60156 484516 65812 490172 sw
tri 60156 478860 65812 484516 ne
tri 65812 481328 69000 484516 sw
rect 65812 478860 69000 481328
tri 69000 478860 71468 481328 sw
tri 65812 475672 69000 478860 ne
rect 69000 478500 71468 478860
tri 71468 478500 71828 478860 sw
tri 69000 475672 71828 478500 nw
tri 724 459067 907 459250 se
rect 907 459067 5493 459250
tri 5493 459067 5676 459250 sw
tri 383 458726 724 459067 se
rect 724 458967 5676 459067
tri 5676 458967 5776 459067 sw
rect 724 458726 5776 458967
tri 200 458543 383 458726 se
rect 383 458543 5776 458726
tri 5776 458543 6200 458967 sw
rect 200 456352 6200 458543
rect 200 455500 6201 456352
tri 6201 455500 7224 456352 sw
rect 200 453957 82328 455500
tri 200 453774 383 453957 ne
rect 383 453774 82328 453957
tri 383 453250 907 453774 ne
rect 907 453533 82328 453774
tri 82328 453533 84295 455500 sw
rect 92000 453533 96000 492658
rect 117000 476500 121000 496861
tri 96000 453533 96795 454328 sw
rect 142000 453533 146000 498199
rect 167000 476500 171000 500737
tri 146000 453533 146795 454328 sw
rect 907 453250 84295 453533
tri 3675 451500 5776 453250 ne
rect 5776 451500 84295 453250
tri 84295 451500 86328 453533 sw
rect 92000 452672 96795 453533
tri 96795 452672 97656 453533 sw
rect 142000 452672 146795 453533
tri 146795 452672 147656 453533 sw
tri 92000 451500 93172 452672 ne
rect 93172 451500 97656 452672
tri 80672 445844 86328 451500 ne
tri 86328 445844 91984 451500 sw
tri 93172 447016 97656 451500 ne
tri 97656 447016 103312 452672 sw
tri 142000 447016 147656 452672 ne
tri 147656 447016 153312 452672 sw
tri 97656 445844 98828 447016 ne
rect 98828 445844 103312 447016
tri 86328 440188 91984 445844 ne
tri 91984 441828 96000 445844 sw
rect 91984 440188 96000 441828
tri 98828 441360 103312 445844 ne
tri 103312 441360 108968 447016 sw
tri 147656 441360 153312 447016 ne
tri 153312 441360 158968 447016 sw
tri 91984 440172 92000 440188 ne
tri 729 438572 907 438750 se
rect 907 438572 5493 438750
tri 5493 438572 5671 438750 sw
tri 378 438221 729 438572 se
rect 729 438221 5671 438572
tri 200 438043 378 438221 se
rect 378 438043 5671 438221
tri 5671 438043 6200 438572 sw
rect 200 435559 6200 438043
tri 6200 435559 6459 435785 sw
rect 200 433457 6459 435559
tri 200 433279 378 433457 ne
rect 378 433279 6459 433457
tri 378 432750 907 433279 ne
rect 907 432750 6459 433279
tri 3594 430248 6459 432750 ne
tri 6459 430500 12251 435559 sw
rect 6459 430248 71000 430500
tri 6459 426500 10749 430248 ne
rect 10749 426500 71000 430248
tri 727 418070 907 418250 se
rect 907 418070 5493 418250
tri 5493 418070 5673 418250 sw
tri 380 417723 727 418070 se
rect 727 417723 5673 418070
tri 200 417543 380 417723 se
rect 380 417543 5673 417723
tri 5673 417543 6200 418070 sw
rect 200 412957 6200 417543
rect 92000 415172 96000 440188
tri 103312 435704 108968 441360 ne
tri 108968 435704 114624 441360 sw
tri 153312 435704 158968 441360 ne
tri 158968 435704 164624 441360 sw
tri 108968 430048 114624 435704 ne
tri 114624 431328 119000 435704 sw
tri 158968 431328 163344 435704 ne
rect 163344 431328 164624 435704
tri 164624 431328 169000 435704 sw
rect 114624 430048 119000 431328
tri 119000 430048 120280 431328 sw
tri 163344 430048 164624 431328 ne
rect 164624 430048 169000 431328
tri 169000 430048 170280 431328 sw
tri 114624 425672 119000 430048 ne
rect 119000 428500 120280 430048
tri 120280 428500 121828 430048 sw
tri 119000 425672 121828 428500 nw
tri 164624 425672 169000 430048 ne
rect 169000 428500 170280 430048
tri 170280 428500 171828 430048 sw
tri 169000 425672 171828 428500 nw
tri 96000 415172 97656 416828 sw
tri 92000 414827 92345 415172 ne
rect 92345 414827 97656 415172
tri 200 412777 380 412957 ne
rect 380 412777 6200 412957
tri 380 412250 907 412777 ne
rect 907 412411 6200 412777
tri 6200 412411 8276 414827 sw
tri 92345 412411 94761 414827 ne
rect 94761 412411 97656 414827
rect 907 412250 8276 412411
tri 3141 409326 5654 412250 ne
rect 5654 410500 8276 412250
tri 8276 410500 9918 412411 sw
tri 94761 410500 96672 412411 ne
rect 96672 410500 97656 412411
tri 97656 410500 102328 415172 sw
rect 5654 409326 84828 410500
tri 84828 409326 86002 410500 sw
tri 96672 409516 97656 410500 ne
rect 97656 409516 139828 410500
tri 139828 409516 140812 410500 sw
tri 97656 409326 97846 409516 ne
rect 97846 409326 140812 409516
tri 5654 406500 8082 409326 ne
rect 8082 406500 86002 409326
tri 86002 406500 88828 409326 sw
tri 97846 406500 100672 409326 ne
rect 100672 406500 140812 409326
tri 140812 406500 143828 409516 sw
tri 83172 404328 85344 406500 ne
rect 85344 404328 88828 406500
tri 88828 404328 91000 406500 sw
tri 138172 404328 140344 406500 ne
rect 140344 404328 143828 406500
tri 143828 404328 146000 406500 sw
tri 85344 400844 88828 404328 ne
rect 88828 402156 91000 404328
tri 91000 402156 93172 404328 sw
tri 140344 402156 142516 404328 ne
rect 142516 402156 146000 404328
rect 88828 400844 93172 402156
tri 93172 400844 94484 402156 sw
tri 142516 400844 143828 402156 ne
rect 143828 400844 146000 402156
tri 146000 400844 149484 404328 sw
tri 3176 397750 5596 400500 se
rect 5596 397750 77260 400500
tri 77260 397750 80353 400500 sw
tri 88828 397750 91922 400844 ne
rect 91922 400500 94484 400844
tri 94484 400500 94828 400844 sw
tri 143828 400500 144172 400844 ne
rect 144172 400500 149484 400844
rect 91922 397750 129828 400500
tri 200 397043 907 397750 se
rect 907 397043 80353 397750
rect 200 396500 80353 397043
tri 80353 396500 81760 397750 sw
tri 91922 396500 93172 397750 ne
rect 93172 396500 129828 397750
tri 129828 396500 133828 400500 sw
tri 144172 396500 148172 400500 ne
rect 148172 396500 149484 400500
rect 200 392457 6200 396500
tri 6200 395132 7404 396500 nw
tri 75740 395132 77279 396500 ne
rect 77279 395132 81760 396500
tri 200 392280 377 392457 ne
rect 377 392280 5670 392457
tri 377 391927 730 392280 ne
rect 730 391927 5670 392280
tri 5670 391927 6200 392457 nw
tri 77279 391927 80884 395132 ne
rect 80884 391927 81760 395132
tri 730 391750 907 391927 ne
rect 907 391750 5493 391927
tri 5493 391750 5670 391927 nw
tri 80884 391750 81083 391927 ne
rect 81083 391750 81760 391927
tri 81760 391750 87103 396500 sw
tri 128172 391750 132922 396500 ne
rect 132922 391750 133828 396500
tri 81083 391149 81760 391750 ne
rect 81760 391149 87103 391750
tri 87103 391149 87780 391750 sw
tri 81760 390844 82103 391149 ne
rect 82103 390844 87780 391149
tri 87780 390844 88123 391149 sw
tri 132922 390844 133828 391750 ne
tri 133828 390844 139484 396500 sw
tri 148172 395188 149484 396500 ne
tri 149484 395188 155140 400844 sw
tri 187000 399328 192000 404328 se
rect 192000 402672 196000 500800
rect 217000 500800 223043 501263
tri 223043 500800 223506 501263 nw
tri 243281 500800 245250 503255 se
rect 245250 501507 251250 506093
tri 272750 506093 273278 506621 se
rect 273278 506272 278222 506621
tri 278222 506272 278571 506621 sw
rect 273278 506093 278571 506272
tri 278571 506093 278750 506272 sw
rect 245250 501318 251061 501507
tri 251061 501318 251250 501507 nw
tri 270958 501318 272750 503389 se
rect 272750 501507 278750 506093
tri 300250 506093 300781 506624 se
rect 300781 506269 305719 506624
tri 305719 506269 306074 506624 sw
tri 328278 506621 328457 506800 se
rect 328457 506621 333043 506800
tri 327929 506272 328278 506621 se
rect 328278 506272 333043 506621
rect 300781 506093 306074 506269
tri 306074 506093 306250 506269 sw
rect 272750 501328 278571 501507
tri 278571 501328 278750 501507 nw
rect 272750 501318 278043 501328
rect 245250 500800 250543 501318
tri 250543 500800 251061 501318 nw
tri 270510 500800 270958 501318 se
rect 270958 500800 278043 501318
tri 278043 500800 278571 501328 nw
tri 297868 500800 300250 503452 se
rect 300250 501507 306250 506093
rect 300250 501331 306074 501507
tri 306074 501331 306250 501507 nw
tri 327750 506093 327929 506272 se
rect 327929 506093 333043 506272
tri 333043 506093 333750 506800 sw
rect 327750 501917 333750 506093
tri 333750 501917 336000 503855 sw
rect 327750 501507 336000 501917
rect 300250 500800 305543 501331
tri 305543 500800 306074 501331 nw
tri 327750 501328 327929 501507 ne
rect 327929 501328 336000 501507
tri 327929 500800 328457 501328 ne
rect 328457 500800 336000 501328
rect 217000 500799 221233 500800
tri 221233 500799 221234 500800 nw
rect 243281 500799 248408 500800
tri 270509 500799 270510 500800 se
rect 270510 500799 275798 500800
tri 275798 500799 275799 500800 nw
rect 297868 500799 303243 500800
rect 217000 500637 221132 500799
tri 221132 500638 221233 500799 nw
tri 243152 500639 243281 500799 se
rect 243281 500639 248278 500799
rect 217000 476500 221000 500637
tri 221000 500426 221132 500637 nw
tri 242814 500217 243152 500638 se
rect 243152 500637 248278 500639
tri 248278 500638 248408 500799 nw
tri 270369 500638 270509 500799 se
rect 270509 500638 275658 500799
tri 275658 500638 275798 500799 nw
tri 297723 500638 297868 500799 se
rect 297868 500638 303098 500799
tri 303098 500638 303243 500799 nw
tri 331167 500638 331355 500800 ne
rect 331355 500638 336000 500800
rect 270369 500637 275658 500638
rect 243152 500217 247941 500637
tri 247941 500217 248278 500637 nw
tri 270257 500508 270369 500637 se
rect 270369 500508 275546 500637
tri 275546 500508 275658 500637 nw
tri 270005 500217 270257 500508 se
rect 270257 500217 272289 500508
tri 242000 499203 242814 500217 se
rect 242814 499203 247128 500217
tri 247128 499203 247941 500217 nw
tri 269127 499203 270005 500217 se
rect 270005 499203 272289 500217
tri 241422 453750 242000 454328 se
rect 242000 453750 246000 499203
tri 246000 497797 247128 499203 nw
tri 267911 497798 269127 499202 se
rect 269127 497798 272289 499203
tri 267000 496745 267911 497797 se
rect 267911 496745 272289 497798
tri 272289 496745 275546 500508 nw
rect 267000 496744 272289 496745
rect 267000 476500 271000 496744
tri 271000 495255 272289 496744 nw
tri 292347 494652 297723 500638 se
tri 297723 494652 303098 500638 nw
tri 331355 500083 332000 500638 ne
tri 292000 494266 292347 494652 se
rect 292347 494266 297376 494652
tri 297376 494266 297723 494652 nw
tri 331938 494266 332000 494328 se
rect 332000 494266 336000 500638
tri 286344 461172 292000 466828 se
rect 292000 465172 296000 494266
tri 296000 492734 297376 494266 nw
tri 330406 492734 331938 494266 se
rect 331938 492734 336000 494266
tri 326344 488672 330406 492734 se
rect 330406 492672 336000 492734
rect 330406 488672 332000 492672
tri 332000 488672 336000 492672 nw
tri 320688 483016 326344 488672 se
tri 326344 483016 332000 488672 nw
tri 316172 478500 320688 483016 se
rect 320688 478500 321828 483016
tri 321828 478500 326344 483016 nw
tri 316172 475672 319000 478500 ne
tri 319000 475672 321828 478500 nw
tri 292000 461172 296000 465172 nw
tri 284922 459750 286344 461172 se
rect 286344 459750 290578 461172
tri 290578 459750 292000 461172 nw
tri 280688 455516 284922 459750 se
rect 284922 455516 286344 459750
tri 286344 455516 290578 459750 nw
tri 381927 459170 382507 459750 se
rect 382507 459170 387093 459750
tri 387093 459170 387673 459750 sw
tri 381800 459043 381927 459170 se
rect 381927 459043 387673 459170
tri 387673 459043 387800 459170 sw
tri 280672 455500 280688 455516 se
rect 280688 455500 286328 455516
tri 286328 455500 286344 455516 nw
rect 381800 455500 387800 459043
tri 253922 453750 255672 455500 se
rect 255672 453750 284578 455500
tri 284578 453750 286328 455500 nw
tri 291422 453750 293172 455500 se
rect 293172 454457 387800 455500
rect 293172 453877 387220 454457
tri 387220 453877 387800 454457 nw
rect 293172 453750 387093 453877
tri 387093 453750 387220 453877 nw
tri 237516 449844 241422 453750 se
rect 241422 452672 246000 453750
rect 241422 449844 243172 452672
tri 243172 449844 246000 452672 nw
tri 250016 449844 253922 453750 se
rect 253922 451500 282328 453750
tri 282328 451500 284578 453750 nw
tri 289172 451500 291422 453750 se
rect 291422 451500 385567 453750
tri 385567 451500 386121 453750 nw
rect 253922 449844 255672 451500
tri 255672 449844 257328 451500 nw
tri 287516 449844 289172 451500 se
rect 289172 449844 293172 451500
tri 293172 449844 294828 451500 nw
tri 236344 448672 237516 449844 se
rect 237516 448672 242000 449844
tri 242000 448672 243172 449844 nw
tri 248844 448672 250016 449844 se
tri 231860 444188 236344 448672 se
rect 236344 444188 237516 448672
tri 237516 444188 242000 448672 nw
tri 244360 444188 248844 448672 se
rect 248844 444188 250016 448672
tri 250016 444188 255672 449844 nw
tri 281860 444188 287516 449844 se
tri 287516 444188 293172 449844 nw
tri 230688 443016 231860 444188 se
rect 231860 443016 236344 444188
tri 236344 443016 237516 444188 nw
tri 225032 437360 230688 443016 se
tri 230688 437360 236344 443016 nw
tri 242000 441828 244360 444188 se
rect 244360 441828 247656 444188
tri 247656 441828 250016 444188 nw
tri 279500 441828 281860 444188 se
tri 219376 431704 225032 437360 se
tri 225032 431704 230688 437360 nw
tri 216172 428500 219376 431704 se
rect 219376 428500 221828 431704
tri 221828 428500 225032 431704 nw
tri 216172 425672 219000 428500 ne
tri 219000 425672 221828 428500 nw
tri 241922 416750 242000 416828 se
rect 242000 416750 246000 441828
tri 246000 440172 247656 441828 nw
tri 277844 440172 279500 441828 se
rect 279500 440172 281860 441828
tri 276204 438532 277844 440172 se
rect 277844 438532 281860 440172
tri 281860 438532 287516 444188 nw
tri 328566 440894 330672 443000 se
rect 330672 440894 379823 443000
tri 379823 440894 381947 443000 sw
tri 326204 438532 328566 440894 se
rect 328566 439000 381947 440894
rect 328566 438532 331018 439000
tri 275922 438250 276204 438532 se
rect 276204 438250 281578 438532
tri 281578 438250 281860 438532 nw
tri 325922 438250 326204 438532 se
rect 326204 438250 331018 438532
tri 270548 432876 275922 438250 se
rect 275922 432876 276204 438250
tri 276204 432876 281578 438250 nw
tri 325362 437690 325922 438250 se
rect 325922 437690 331018 438250
tri 331018 437690 332328 439000 nw
tri 378177 437690 379498 439000 ne
rect 379498 438532 381947 439000
tri 381947 438532 384329 440894 sw
rect 379498 438250 384329 438532
tri 384329 438250 384614 438532 sw
rect 379498 437715 387093 438250
tri 387093 437715 387628 438250 sw
rect 379498 437690 387628 437715
tri 325016 437344 325362 437690 se
rect 325362 437344 330672 437690
tri 330672 437344 331018 437690 nw
tri 379498 437344 379847 437690 ne
rect 379847 437543 387628 437690
tri 387628 437543 387800 437715 sw
rect 379847 437344 387800 437543
tri 320548 432876 325016 437344 se
rect 325016 432876 325578 437344
tri 269922 432250 270548 432876 se
rect 270548 432250 275578 432876
tri 275578 432250 276204 432876 nw
tri 319922 432250 320548 432876 se
rect 320548 432250 325578 432876
tri 325578 432250 330672 437344 nw
tri 379847 435407 381800 437344 ne
rect 381800 432957 387800 437344
tri 381800 432810 381947 432957 ne
rect 381947 432810 387628 432957
tri 381947 432422 382335 432810 ne
rect 382335 432785 387628 432810
tri 387628 432785 387800 432957 nw
rect 382335 432422 387265 432785
tri 387265 432422 387628 432785 nw
tri 382335 432250 382507 432422 ne
rect 382507 432250 387093 432422
tri 387093 432250 387265 432422 nw
tri 266172 428500 269922 432250 se
rect 269922 428500 271828 432250
tri 271828 428500 275578 432250 nw
tri 319360 431688 319922 432250 se
rect 319922 431688 325016 432250
tri 325016 431688 325578 432250 nw
tri 316172 428500 319360 431688 se
rect 319360 428500 321828 431688
tri 321828 428500 325016 431688 nw
tri 266172 425672 269000 428500 ne
tri 269000 425672 271828 428500 nw
tri 316172 425672 319000 428500 ne
tri 319000 425672 321828 428500 nw
tri 236344 411172 241922 416750 se
rect 241922 415172 246000 416750
tri 382332 416575 382507 416750 se
rect 382507 416575 387093 416750
tri 387093 416575 387268 416750 sw
rect 241922 411172 242000 415172
tri 242000 411172 246000 415172 nw
tri 381800 416043 382332 416575 se
rect 382332 416218 387268 416575
tri 387268 416218 387625 416575 sw
rect 382332 416043 387625 416218
tri 387625 416043 387800 416218 sw
tri 378980 411179 381800 413732 se
rect 381800 411457 387800 416043
rect 381800 411282 387625 411457
tri 387625 411282 387800 411457 nw
rect 381800 411179 387522 411282
tri 387522 411179 387625 411282 nw
tri 378972 411172 378980 411179 se
rect 378980 411172 387093 411179
tri 235922 410750 236344 411172 se
rect 236344 410750 241578 411172
tri 241578 410750 242000 411172 nw
tri 378506 410750 378972 411172 se
rect 378972 410750 387093 411172
tri 387093 410750 387522 411179 nw
tri 230688 405516 235922 410750 se
rect 235922 405516 236344 410750
tri 236344 405516 241578 410750 nw
tri 378229 410500 378506 410750 se
rect 378506 410500 384191 410750
tri 384191 410500 384467 410750 nw
tri 243188 405516 248172 410500 se
rect 248172 406500 379771 410500
tri 379771 406500 384191 410500 nw
tri 230672 405500 230688 405516 se
rect 230688 405500 236328 405516
tri 236328 405500 236344 405516 nw
tri 243172 405500 243188 405516 se
rect 243188 405500 248172 405516
rect 192000 399328 192656 402672
tri 192656 399328 196000 402672 nw
tri 205016 399844 210672 405500 se
rect 210672 401500 232328 405500
tri 232328 401500 236328 405500 nw
tri 242516 404844 243172 405500 se
rect 243172 404844 248172 405500
tri 248172 404844 249828 406500 nw
tri 239172 401500 242516 404844 se
rect 242516 401500 243828 404844
tri 210672 399844 212328 401500 nw
tri 238172 400500 239172 401500 se
rect 239172 400500 243828 401500
tri 243828 400500 248172 404844 nw
tri 237516 399844 238172 400500 se
rect 238172 399844 243172 400500
tri 243172 399844 243828 400500 nw
tri 252516 399844 253172 400500 se
rect 253172 399844 379873 400500
tri 379873 399844 380481 400500 sw
tri 204500 399328 205016 399844 se
rect 205016 399328 206078 399844
rect 187000 397750 191078 399328
tri 191078 397750 192656 399328 nw
tri 202922 397750 204500 399328 se
rect 204500 397750 206078 399328
tri 149484 390844 153828 395188 ne
rect 153828 390844 155140 395188
tri 82103 385798 87780 390844 ne
rect 87780 385798 88123 390844
tri 88123 385798 93800 390844 sw
tri 87780 385188 88466 385798 ne
rect 88466 385188 93800 385798
tri 93800 385188 94486 385798 sw
tri 133828 385188 139484 390844 ne
tri 139484 388328 142000 390844 sw
tri 153828 389532 155140 390844 ne
tri 155140 389532 160796 395188 sw
tri 155140 388328 156344 389532 ne
rect 156344 388328 160796 389532
rect 139484 385188 142000 388328
tri 142000 385188 145140 388328 sw
tri 156344 385188 159484 388328 ne
rect 159484 385188 160796 388328
tri 88466 382672 91296 385188 ne
rect 91296 382672 94486 385188
tri 94486 382672 97316 385188 sw
tri 139484 382672 142000 385188 ne
rect 142000 384328 145140 385188
tri 145140 384328 146000 385188 sw
tri 91296 380500 93740 382672 ne
rect 93740 380500 97316 382672
tri 97316 380500 99760 382672 sw
tri 2998 377250 5521 380500 se
rect 5521 377250 71000 380500
tri 93740 380447 93800 380500 ne
rect 93800 380447 121000 380500
tri 200 376543 907 377250 se
rect 907 376543 71000 377250
rect 200 376500 71000 376543
tri 93800 376500 98240 380447 ne
rect 98240 376500 121000 380447
rect 200 371957 6200 376500
tri 6200 374853 7479 376500 nw
tri 200 371763 394 371957 ne
rect 394 371763 5687 371957
tri 394 371444 713 371763 ne
rect 713 371444 5687 371763
tri 5687 371444 6200 371957 nw
tri 713 371250 907 371444 ne
rect 907 371250 5493 371444
tri 5493 371250 5687 371444 nw
tri 200 356043 907 356750 se
rect 907 356043 5493 356750
tri 5493 356043 6200 356750 sw
rect 200 355528 6200 356043
rect 200 355500 6206 355528
tri 6206 355500 6576 355528 sw
rect 200 351907 94828 355500
tri 94828 351907 98421 355500 sw
rect 200 351516 98421 351907
rect 200 351457 6200 351516
tri 6212 351500 6424 351516 ne
rect 6424 351500 98421 351516
tri 98421 351500 98828 351907 sw
tri 200 350750 907 351457 ne
rect 907 350750 5493 351457
tri 5493 350750 6200 351457 nw
tri 93172 350750 93922 351500 ne
rect 93922 350750 98828 351500
tri 93922 345844 98828 350750 ne
tri 98828 345844 104484 351500 sw
tri 98828 340188 104484 345844 ne
tri 104484 340188 110140 345844 sw
tri 104484 336250 108422 340188 ne
rect 108422 336250 110140 340188
tri 722 336065 907 336250 se
rect 907 336065 5493 336250
tri 5493 336065 5678 336250 sw
tri 108422 336065 108607 336250 ne
rect 108607 336065 110140 336250
tri 385 335728 722 336065 se
rect 722 335728 5678 336065
tri 200 335543 385 335728 se
rect 385 335543 5678 335728
tri 5678 335543 6200 336065 sw
rect 200 332970 6200 335543
tri 108607 334532 110140 336065 ne
tri 110140 334532 115796 340188 sw
tri 110140 333378 111294 334532 ne
rect 111294 333378 115796 334532
tri 6200 332970 6699 333378 sw
tri 111294 332970 111702 333378 ne
rect 111702 332970 115796 333378
rect 200 330957 6699 332970
tri 200 330772 385 330957 ne
rect 385 330772 6699 330957
tri 385 330250 907 330772 ne
rect 907 330500 6699 330772
tri 6699 330500 9714 332970 sw
tri 111702 330500 114172 332970 ne
rect 114172 331328 115796 332970
tri 115796 331328 119000 334532 sw
rect 114172 330500 119000 331328
rect 907 330250 71000 330500
tri 3706 327800 6699 330250 ne
rect 6699 327800 71000 330250
tri 114172 328876 115796 330500 ne
rect 115796 328876 119000 330500
tri 119000 328876 121452 331328 sw
rect 142000 330500 146000 384328
tri 159484 383876 160796 385188 ne
tri 160796 383876 166452 389532 sw
tri 160796 378220 166452 383876 ne
tri 166452 378500 171828 383876 sw
rect 166452 378220 171548 378500
tri 171548 378220 171828 378500 nw
tri 166452 375672 169000 378220 ne
tri 169000 375672 171548 378220 nw
tri 6699 326500 8286 327800 ne
rect 8286 326500 71000 327800
tri 115796 326500 118172 328876 ne
rect 118172 328500 121452 328876
tri 121452 328500 121828 328876 sw
rect 118172 326500 119000 328500
tri 118172 325672 119000 326500 ne
tri 119000 325672 121828 328500 nw
rect 142000 326500 171000 330500
tri 731 315574 907 315750 se
rect 907 315574 5493 315750
tri 5493 315574 5669 315750 sw
tri 376 315219 731 315574 se
rect 731 315493 5669 315574
tri 5669 315493 5750 315574 sw
rect 731 315219 5750 315493
tri 200 315043 376 315219 se
rect 376 315043 5750 315219
tri 5750 315043 6200 315493 sw
rect 200 310457 6200 315043
tri 200 310281 376 310457 ne
rect 376 310281 6200 310457
tri 376 309750 907 310281 ne
rect 907 310007 6200 310281
tri 6200 310007 8348 312401 sw
rect 907 309750 8348 310007
tri 3205 306914 5750 309750 ne
rect 5750 307490 8348 309750
tri 8348 307490 10607 310007 sw
rect 5750 306915 10607 307490
tri 10607 306915 11123 307490 sw
rect 5750 306914 11123 306915
tri 5750 303250 9037 306914 ne
rect 9037 305500 11123 306914
tri 11123 305500 12393 306914 sw
rect 9037 303250 94828 305500
tri 94828 303250 97078 305500 sw
tri 9037 302672 9555 303250 ne
rect 9555 302672 97078 303250
tri 97078 302672 97656 303250 sw
tri 9555 301500 10607 302672 ne
rect 10607 301500 97656 302672
tri 97656 301500 98828 302672 sw
tri 93172 295844 98828 301500 ne
tri 98828 295844 104484 301500 sw
tri 98828 295250 99422 295844 ne
rect 99422 295250 104484 295844
tri 735 295078 907 295250 se
rect 907 295078 5493 295250
tri 5493 295078 5665 295250 sw
tri 99422 295078 99594 295250 ne
rect 99594 295078 104484 295250
tri 372 294715 735 295078 se
rect 735 294805 5665 295078
tri 5665 294805 5938 295078 sw
tri 99594 294805 99867 295078 ne
rect 99867 294805 104484 295078
rect 735 294715 5938 294805
tri 200 294543 372 294715 se
rect 372 294543 5938 294715
tri 5938 294543 6200 294805 sw
rect 200 289957 6200 294543
tri 99867 292026 102646 294805 ne
rect 102646 292026 104484 294805
tri 200 289785 372 289957 ne
rect 372 289785 6200 289957
tri 372 289250 907 289785 ne
rect 907 289696 6200 289785
tri 6200 289696 8454 292026 sw
tri 102646 290188 104484 292026 ne
tri 104484 290188 110140 295844 sw
rect 907 289250 8454 289696
tri 104484 289695 104977 290188 ne
rect 104977 289695 110140 290188
tri 3319 286543 5938 289250 ne
rect 5938 286543 8454 289250
tri 8454 286543 11504 289695 sw
tri 104977 286543 108129 289695 ne
rect 108129 286543 110140 289695
tri 5938 280789 11504 286543 ne
tri 11504 282253 15652 286543 sw
tri 108129 284532 110140 286543 ne
tri 110140 284532 115796 290188 sw
tri 110140 282253 112419 284532 ne
rect 112419 282253 115796 284532
rect 11504 280789 15652 282253
tri 15652 280789 17068 282253 sw
tri 112419 280789 113883 282253 ne
rect 113883 281328 115796 282253
tri 115796 281328 119000 284532 sw
rect 113883 280789 119000 281328
tri 11504 276500 15652 280789 ne
rect 15652 280500 17068 280789
tri 17068 280500 17348 280789 sw
tri 113883 280500 114172 280789 ne
rect 114172 280500 119000 280789
rect 15652 276500 71000 280500
tri 114172 278876 115796 280500 ne
rect 115796 278876 119000 280500
tri 119000 278876 121452 281328 sw
tri 115796 276500 118172 278876 ne
rect 118172 278500 121452 278876
tri 121452 278500 121828 278876 sw
rect 118172 276500 119000 278500
tri 118172 275672 119000 276500 ne
tri 119000 275672 121828 278500 nw
tri 735 274578 907 274750 se
rect 907 274578 5493 274750
tri 5493 274578 5665 274750 sw
tri 372 274215 735 274578 se
rect 735 274215 5665 274578
tri 200 274043 372 274215 se
rect 372 274190 5665 274215
tri 5665 274190 6053 274578 sw
rect 372 274043 6053 274190
tri 6053 274043 6200 274190 sw
rect 200 269457 6200 274043
tri 200 269285 372 269457 ne
rect 372 269310 6200 269457
tri 6200 269310 8501 271592 sw
rect 372 269285 8501 269310
tri 372 268750 907 269285 ne
rect 907 268750 8501 269285
tri 3385 266250 5907 268750 ne
rect 5907 268000 8501 268750
tri 8501 268000 9823 269310 sw
rect 5907 266250 44828 268000
tri 44828 266250 46578 268000 sw
tri 5907 266106 6053 266250 ne
rect 6053 266106 46578 266250
tri 46578 266106 46722 266250 sw
tri 6053 264000 8177 266106 ne
rect 8177 264000 46722 266106
tri 46722 264000 48828 266106 sw
tri 43172 260250 46922 264000 ne
rect 46922 260250 48828 264000
tri 48828 260250 52578 264000 sw
tri 46922 258344 48828 260250 ne
rect 48828 258344 52578 260250
tri 52578 258344 54484 260250 sw
tri 48828 254250 52922 258344 ne
rect 52922 255500 54484 258344
tri 54484 255500 57328 258344 sw
rect 52922 254250 94828 255500
tri 732 254075 907 254250 se
rect 907 254075 5493 254250
tri 5493 254075 5668 254250 sw
tri 52922 254075 53097 254250 ne
rect 53097 254075 94828 254250
tri 375 253718 732 254075 se
rect 732 253718 5668 254075
tri 200 253543 375 253718 se
rect 375 253543 5668 253718
tri 5668 253543 6200 254075 sw
rect 200 251232 6200 253543
tri 53097 252688 54484 254075 ne
rect 54484 252688 94828 254075
tri 94828 252688 97640 255500 sw
tri 54484 251500 55672 252688 ne
rect 55672 251500 97640 252688
tri 97640 251500 98828 252688 sw
tri 93172 251232 93440 251500 ne
rect 93440 251232 98828 251500
rect 200 251109 6201 251232
tri 6201 251109 6337 251232 sw
tri 93440 251109 93563 251232 ne
rect 93563 251109 98828 251232
rect 200 248957 6337 251109
tri 200 248782 375 248957 ne
rect 375 248782 6337 248957
tri 375 248250 907 248782 ne
rect 907 248250 6337 248782
tri 3533 245713 6337 248250 ne
tri 6337 248000 9771 251109 sw
tri 93563 248000 96672 251109 ne
rect 96672 248000 98828 251109
rect 6337 245713 52328 248000
tri 52328 245713 54615 248000 sw
tri 96672 245844 98828 248000 ne
tri 98828 245844 104484 251500 sw
tri 98828 245713 98959 245844 ne
rect 98959 245713 104484 245844
tri 6337 244750 7400 245713 ne
rect 7400 244750 54615 245713
tri 54615 244750 55578 245713 sw
tri 98959 244750 99922 245713 ne
rect 99922 244750 104484 245713
tri 104484 244750 105578 245844 sw
tri 7400 244000 8229 244750 ne
rect 8229 244000 55578 244750
tri 55578 244000 56328 244750 sw
tri 99922 244000 100672 244750 ne
rect 100672 244000 105578 244750
tri 50672 238750 55922 244000 ne
rect 55922 238750 56328 244000
tri 56328 238750 61578 244000 sw
tri 100672 240188 104484 244000 ne
rect 104484 240188 105578 244000
tri 105578 240188 110140 244750 sw
tri 104484 238750 105922 240188 ne
rect 105922 238750 110140 240188
tri 110140 238750 111578 240188 sw
tri 55922 238344 56328 238750 ne
rect 56328 238344 61578 238750
tri 61578 238344 61984 238750 sw
tri 105922 238344 106328 238750 ne
rect 106328 238344 111578 238750
tri 56328 233750 60922 238344 ne
rect 60922 233750 61984 238344
tri 735 233578 907 233750 se
rect 907 233578 5493 233750
tri 5493 233578 5665 233750 sw
tri 60922 233578 61094 233750 ne
rect 61094 233578 61984 233750
tri 372 233215 735 233578 se
rect 735 233215 5665 233578
tri 200 233043 372 233215 se
rect 372 233078 5665 233215
tri 5665 233078 6165 233578 sw
tri 61094 233078 61594 233578 ne
rect 61594 233078 61984 233578
rect 372 233043 6165 233078
tri 6165 233043 6200 233078 sw
rect 200 228457 6200 233043
tri 61594 232688 61984 233078 ne
tri 61984 232688 67640 238344 sw
tri 106328 234532 110140 238344 ne
rect 110140 234532 111578 238344
tri 111578 234532 115796 238750 sw
tri 110140 232688 111984 234532 ne
rect 111984 232688 115796 234532
tri 61984 230651 64021 232688 ne
rect 64021 230651 67640 232688
tri 200 228285 372 228457 ne
rect 372 228422 6200 228457
tri 6200 228422 8534 230651 sw
tri 64021 228422 66250 230651 ne
rect 66250 228500 67640 230651
tri 67640 228500 71828 232688 sw
tri 111984 228876 115796 232688 ne
tri 115796 231328 119000 234532 sw
rect 115796 228876 119000 231328
tri 119000 228876 121452 231328 sw
rect 66250 228422 70360 228500
rect 372 228285 8534 228422
tri 372 227750 907 228285 ne
rect 907 227750 8534 228285
tri 3445 225153 6165 227750 ne
rect 6165 225153 8534 227750
tri 8534 225153 11958 228422 sw
tri 66250 227032 67640 228422 ne
rect 67640 227032 70360 228422
tri 70360 227032 71828 228500 nw
tri 115796 227032 117640 228876 ne
rect 117640 228500 121452 228876
tri 121452 228500 121828 228876 sw
rect 117640 227032 119000 228500
tri 67640 225672 69000 227032 ne
tri 69000 225672 70360 227032 nw
tri 117640 225672 119000 227032 ne
tri 119000 225672 121828 228500 nw
tri 6165 223250 8157 225153 ne
rect 8157 223250 11958 225153
tri 11958 223250 13950 225153 sw
tri 8157 219621 11958 223250 ne
rect 11958 219621 13950 223250
tri 13950 219621 17751 223250 sw
rect 142000 220172 146000 326500
rect 187000 309250 191000 397750
tri 191000 397672 191078 397750 nw
tri 202844 397672 202922 397750 se
rect 202922 397672 206078 397750
tri 200422 395250 202844 397672 se
rect 202844 395250 206078 397672
tri 206078 395250 210672 399844 nw
tri 236860 399188 237516 399844 se
rect 237516 399188 242516 399844
tri 242516 399188 243172 399844 nw
tri 235697 398025 236860 399188 se
rect 236860 398025 241353 399188
tri 241353 398025 242516 399188 nw
tri 250697 398025 252516 399844 se
rect 252516 398025 380481 399844
tri 380481 398025 382169 399844 sw
tri 232922 395250 235697 398025 se
rect 235697 395250 238578 398025
tri 238578 395250 241353 398025 nw
tri 247922 395250 250697 398025 se
rect 250697 396500 382169 398025
rect 250697 395250 253240 396500
tri 199360 394188 200422 395250 se
rect 200422 394188 205016 395250
tri 205016 394188 206078 395250 nw
tri 232584 394912 232922 395250 se
rect 232922 394912 238240 395250
tri 238240 394912 238578 395250 nw
tri 247584 394912 247922 395250 se
rect 247922 394912 253240 395250
tri 253240 394912 254828 396500 nw
tri 378127 394912 379600 396500 ne
rect 379600 395251 382169 396500
tri 382169 395251 384743 398025 sw
rect 379600 395250 384743 395251
rect 379600 394912 387093 395250
tri 232516 394844 232584 394912 se
rect 232584 394844 238172 394912
tri 238172 394844 238240 394912 nw
tri 247516 394844 247584 394912 se
rect 247584 394844 253172 394912
tri 253172 394844 253240 394912 nw
tri 379600 394844 379663 394912 ne
rect 379663 394844 387093 394912
tri 231860 394188 232516 394844 se
rect 232516 394188 237516 394844
tri 237516 394188 238172 394844 nw
tri 246860 394188 247516 394844 se
rect 247516 394188 247656 394844
tri 197000 391828 199360 394188 se
rect 199360 391828 202656 394188
tri 202656 391828 205016 394188 nw
tri 231204 393532 231860 394188 se
rect 231860 393532 236860 394188
tri 236860 393532 237516 394188 nw
tri 229500 391828 231204 393532 se
rect 231204 391828 235156 393532
tri 235156 391828 236860 393532 nw
tri 244500 391828 246860 394188 se
rect 246860 391828 247656 394188
rect 197000 317776 201000 391828
tri 201000 390172 202656 391828 nw
tri 227844 390172 229500 391828 se
rect 229500 390172 233500 391828
tri 233500 390172 235156 391828 nw
tri 242844 390172 244500 391828 se
rect 244500 390172 247656 391828
tri 225548 387876 227844 390172 se
rect 227844 387876 231204 390172
tri 231204 387876 233500 390172 nw
tri 242000 389328 242844 390172 se
rect 242844 389328 247656 390172
tri 247656 389328 253172 394844 nw
tri 379663 392541 381800 394844 ne
rect 381800 394717 387093 394844
tri 387093 394717 387626 395250 sw
rect 381800 394543 387626 394717
tri 387626 394543 387800 394717 sw
rect 381800 389957 387800 394543
tri 381800 389588 382169 389957 ne
rect 382169 389783 387626 389957
tri 387626 389783 387800 389957 nw
rect 382169 389588 387267 389783
tri 382169 389424 382333 389588 ne
rect 382333 389424 387267 389588
tri 387267 389424 387626 389783 nw
rect 242000 389250 247578 389328
tri 247578 389250 247656 389328 nw
tri 382333 389250 382507 389424 ne
rect 382507 389250 387093 389424
tri 387093 389250 387267 389424 nw
tri 219892 382220 225548 387876 se
tri 225548 382220 231204 387876 nw
tri 216172 378500 219892 382220 se
rect 219892 378500 221828 382220
tri 221828 378500 225548 382220 nw
tri 216172 375672 219000 378500 ne
tri 219000 375672 221828 378500 nw
tri 216172 328500 219000 331328 se
tri 219000 330750 219578 331328 sw
rect 219000 328500 219578 330750
tri 216172 327608 217064 328500 ne
rect 217064 327608 219578 328500
tri 219578 327608 222720 330750 sw
tri 217064 325672 219000 327608 ne
rect 219000 325672 222720 327608
tri 219000 321952 222720 325672 ne
tri 222720 324750 225578 327608 sw
rect 222720 321952 225578 324750
tri 225578 321952 228376 324750 sw
tri 222720 319224 225448 321952 ne
rect 225448 319224 228376 321952
tri 228376 319224 231104 321952 sw
tri 201000 317776 202207 319224 sw
tri 225448 317776 226896 319224 ne
rect 226896 317776 231104 319224
tri 231104 317776 232552 319224 sw
tri 197000 311528 202207 317776 ne
tri 202207 311528 207414 317776 sw
tri 226896 316296 228376 317776 ne
rect 228376 316296 232552 317776
tri 232552 316296 234032 317776 sw
tri 228376 311528 233144 316296 ne
rect 233144 314328 234032 316296
tri 234032 314328 236000 316296 sw
rect 233144 313984 236000 314328
tri 236000 313984 236344 314328 sw
tri 241656 313984 242000 314328 se
rect 242000 313984 246000 389250
tri 246000 387672 247578 389250 nw
tri 266172 378500 269000 381328 se
tri 266172 378124 266548 378500 ne
rect 266548 378124 269000 378500
tri 269000 378124 272204 381328 sw
rect 317000 378124 377289 380500
tri 377289 378124 379833 380500 sw
tri 266548 375672 269000 378124 ne
rect 269000 375672 272204 378124
tri 269000 372468 272204 375672 ne
tri 272204 373750 276578 378124 sw
rect 317000 376500 379833 378124
tri 375711 376320 375903 376500 ne
rect 375903 376320 379833 376500
tri 379833 376320 381765 378124 sw
tri 375903 375027 377289 376320 ne
rect 377289 375027 381765 376320
tri 377289 373750 378656 375027 ne
rect 378656 373750 381765 375027
tri 381765 373750 384517 376320 sw
rect 272204 372468 276578 373750
tri 276578 372468 277860 373750 sw
tri 378656 372468 380029 373750 ne
rect 380029 373216 387093 373750
tri 387093 373216 387627 373750 sw
rect 380029 373043 387627 373216
tri 387627 373043 387800 373216 sw
rect 380029 372468 387800 373043
tri 272204 366812 277860 372468 ne
tri 277860 367750 282578 372468 sw
tri 380029 370847 381765 372468 ne
rect 381765 370847 387800 372468
tri 381765 370814 381800 370847 ne
rect 381800 368457 387800 370847
tri 381800 367923 382334 368457 ne
rect 382334 368284 387627 368457
tri 387627 368284 387800 368457 nw
rect 382334 367923 387266 368284
tri 387266 367923 387627 368284 nw
tri 382334 367750 382507 367923 ne
rect 382507 367750 387093 367923
tri 387093 367750 387266 367923 nw
rect 277860 366812 282578 367750
tri 282578 366812 283516 367750 sw
tri 277860 361156 283516 366812 ne
tri 283516 361156 289172 366812 sw
tri 283516 355500 289172 361156 ne
tri 289172 355500 294828 361156 sw
tri 289172 355418 289254 355500 ne
rect 289254 355418 382479 355500
tri 382479 355418 382542 355500 sw
tri 289254 352250 292422 355418 ne
rect 292422 352250 382542 355418
tri 382542 352250 385002 355418 sw
tri 292422 351500 293172 352250 ne
rect 293172 351737 387093 352250
tri 387093 351737 387606 352250 sw
rect 293172 351543 387606 351737
tri 387606 351543 387800 351737 sw
rect 293172 351500 387800 351543
tri 380521 349852 381800 351500 ne
rect 381800 346957 387800 351500
tri 381800 346250 382507 346957 ne
rect 382507 346763 387606 346957
tri 387606 346763 387800 346957 nw
rect 382507 346444 387287 346763
tri 387287 346444 387606 346763 nw
rect 382507 346250 387093 346444
tri 387093 346250 387287 346444 nw
tri 266172 328500 269000 331328 se
tri 269000 330750 269578 331328 sw
rect 269000 328500 269578 330750
tri 266172 328124 266548 328500 ne
rect 266548 328124 269578 328500
tri 269578 328124 272204 330750 sw
tri 382257 330500 382507 330750 se
rect 382507 330500 387093 330750
tri 387093 330500 387343 330750 sw
rect 317000 330482 381724 330500
tri 381724 330482 381800 330500 sw
tri 382239 330482 382257 330500 se
rect 382257 330482 387343 330500
rect 317000 330405 381803 330482
tri 381803 330405 382135 330482 sw
tri 382162 330405 382239 330482 se
rect 382239 330405 387343 330482
rect 317000 330400 382139 330405
tri 382139 330400 382156 330405 sw
tri 382157 330400 382162 330405 se
rect 382162 330400 387343 330405
rect 317000 330043 387343 330400
tri 387343 330043 387800 330500 sw
tri 266548 325672 269000 328124 ne
rect 269000 325672 272204 328124
tri 269000 322468 272204 325672 ne
tri 272204 324750 275578 328124 sw
rect 317000 326500 387800 330043
tri 381276 326380 381800 326500 ne
rect 381800 325457 387800 326500
tri 381800 325356 381901 325457 ne
rect 381901 325356 387699 325457
tri 387699 325356 387800 325457 nw
tri 381901 324750 382507 325356 ne
rect 382507 324750 387093 325356
tri 387093 324750 387699 325356 nw
rect 272204 322468 275578 324750
tri 275578 322468 277860 324750 sw
tri 272204 316812 277860 322468 ne
tri 277860 316812 283516 322468 sw
rect 233144 311528 236344 313984
tri 236344 311528 238800 313984 sw
tri 239200 311528 241656 313984 se
rect 241656 312672 246000 313984
rect 241656 311528 242578 312672
tri 202207 309328 204040 311528 ne
rect 204040 309328 207414 311528
tri 191000 309250 191078 309328 sw
tri 204040 309250 204105 309328 ne
rect 204105 309250 207414 309328
tri 207414 309250 209312 311528 sw
tri 233144 310640 234032 311528 ne
rect 234032 311328 238800 311528
tri 238800 311328 239000 311528 sw
tri 239000 311328 239200 311528 se
rect 239200 311328 242578 311528
rect 234032 310640 242578 311328
tri 234032 309250 235422 310640 ne
rect 235422 309250 242578 310640
tri 242578 309250 246000 312672 nw
tri 277860 311156 283516 316812 ne
tri 283516 311156 289172 316812 sw
tri 283516 309250 285422 311156 ne
rect 285422 309250 289172 311156
tri 289172 309250 291078 311156 sw
rect 187000 308328 191078 309250
tri 191078 308328 192000 309250 sw
tri 204105 308329 204873 309250 ne
rect 204873 308328 209312 309250
rect 187000 307672 192000 308328
tri 192000 307672 192656 308328 sw
tri 204873 307672 205420 308328 ne
rect 205420 307672 209312 308328
tri 187000 303250 191422 307672 ne
rect 191422 304328 192656 307672
tri 192656 304328 196000 307672 sw
tri 205420 305280 207414 307672 ne
rect 207414 305500 209312 307672
tri 209312 305500 212437 309250 sw
tri 235422 308672 236000 309250 ne
rect 236000 308672 242000 309250
tri 242000 308672 242578 309250 nw
tri 285422 308672 286000 309250 ne
rect 286000 308729 291078 309250
tri 291078 308729 291599 309250 sw
tri 381986 308729 382507 309250 se
rect 382507 308729 387093 309250
tri 387093 308729 387614 309250 sw
rect 286000 308672 291599 308729
tri 291599 308672 291656 308729 sw
tri 236000 308500 236172 308672 ne
rect 236172 308500 241828 308672
tri 241828 308500 242000 308672 nw
tri 236172 305672 239000 308500 ne
rect 239000 308328 241828 308500
tri 241828 308328 242000 308500 sw
tri 286000 308328 286344 308672 ne
rect 286344 308328 291656 308672
tri 291656 308328 292000 308672 sw
tri 381800 308543 381986 308729 se
rect 381986 308543 387614 308729
tri 387614 308543 387800 308729 sw
rect 239000 305672 242000 308328
tri 242000 305672 244656 308328 sw
tri 286344 305672 289000 308328 ne
rect 289000 305672 292000 308328
tri 292000 305672 294656 308328 sw
tri 239000 305500 239172 305672 ne
rect 239172 305500 244656 305672
tri 244656 305500 244828 305672 sw
tri 289000 305500 289172 305672 ne
rect 289172 305500 294656 305672
tri 294656 305500 294828 305672 sw
rect 381800 305500 387800 308543
rect 207414 305280 227328 305500
tri 227328 305280 227548 305500 sw
tri 239172 305280 239392 305500 ne
rect 239392 305280 244828 305500
tri 244828 305280 245048 305500 sw
tri 289172 305280 289392 305500 ne
rect 289392 305280 387800 305500
rect 191422 303250 196000 304328
tri 207414 303250 209105 305280 ne
rect 209105 303250 227548 305280
tri 227548 303250 229578 305280 sw
tri 239392 304984 239688 305280 ne
rect 239688 304984 245048 305280
tri 245048 304984 245344 305280 sw
tri 289392 304984 289688 305280 ne
rect 289688 304984 387800 305280
tri 239688 303250 241422 304984 ne
rect 241422 303250 245344 304984
tri 245344 303250 247078 304984 sw
tri 289688 303250 291422 304984 ne
rect 291422 303957 387800 304984
rect 291422 303436 387279 303957
tri 387279 303436 387800 303957 nw
rect 291422 303250 387093 303436
tri 387093 303250 387279 303436 nw
tri 191422 302672 192000 303250 ne
rect 192000 285500 196000 303250
tri 209105 301500 210563 303250 ne
rect 210563 301500 229578 303250
tri 229578 301500 231328 303250 sw
tri 241422 301500 243172 303250 ne
rect 243172 301500 247078 303250
tri 247078 301500 248828 303250 sw
tri 291422 301500 293172 303250 ne
rect 293172 301500 385501 303250
tri 385501 301500 386010 303250 nw
tri 225672 295844 231328 301500 ne
tri 231328 295844 236984 301500 sw
tri 243172 299328 245344 301500 ne
rect 245344 299328 248828 301500
tri 248828 299328 251000 301500 sw
tri 245344 297672 247000 299328 ne
tri 231328 290188 236984 295844 ne
tri 236984 291828 241000 295844 sw
rect 236984 290188 241000 291828
tri 236984 290172 237000 290188 ne
tri 188454 284532 189422 285500 se
rect 189422 284532 196000 285500
tri 185422 281500 188454 284532 se
rect 188454 281500 196000 284532
tri 185250 281328 185422 281500 se
rect 185422 281328 190906 281500
tri 190906 281328 191078 281500 nw
tri 184422 280500 185250 281328 se
rect 185250 280500 188454 281328
rect 167000 278876 188454 280500
tri 188454 278876 190906 281328 nw
rect 167000 276500 186078 278876
tri 186078 276500 188454 278876 nw
rect 192000 275500 196000 281500
tri 196922 275500 201922 280500 se
rect 201922 276500 221000 280500
rect 201922 275500 202578 276500
tri 202578 275500 203578 276500 nw
rect 192000 271500 198578 275500
tri 198578 271500 202578 275500 nw
rect 192000 235500 196000 271500
rect 237000 258328 241000 290188
rect 247000 267672 251000 299328
tri 382333 287576 382507 287750 se
rect 382507 287576 387093 287750
tri 387093 287576 387267 287750 sw
tri 381800 287043 382333 287576 se
rect 382333 287217 387267 287576
tri 387267 287217 387626 287576 sw
rect 382333 287043 387626 287217
tri 387626 287043 387800 287217 sw
tri 379288 281750 381800 284457 se
rect 381800 282457 387800 287043
rect 381800 282283 387626 282457
tri 387626 282283 387800 282457 nw
rect 381800 281750 387093 282283
tri 387093 281750 387626 282283 nw
tri 379238 281696 379288 281750 se
rect 379288 281696 384694 281750
tri 384694 281696 384744 281750 nw
tri 378896 281328 379238 281696 se
rect 379238 281328 383584 281696
tri 266172 278500 269000 281328 se
tri 266172 277468 267204 278500 ne
rect 267204 277468 269000 278500
tri 269000 277468 272860 281328 sw
tri 378128 280500 378896 281328 se
rect 378896 280500 383584 281328
tri 383584 280500 384694 281696 nw
rect 317000 277468 380770 280500
tri 380770 277468 383584 280500 nw
tri 267204 275672 269000 277468 ne
rect 269000 275672 272860 277468
tri 269000 271812 272860 275672 ne
tri 272860 271812 278516 277468 sw
rect 317000 276500 379872 277468
tri 379872 276500 380770 277468 nw
tri 247000 266812 247860 267672 ne
rect 247860 266812 251000 267672
tri 251000 266812 253516 269328 sw
tri 247860 263672 251000 266812 ne
rect 251000 266156 253516 266812
tri 253516 266156 254172 266812 sw
tri 272860 266156 278516 271812 ne
tri 278516 266250 284078 271812 sw
rect 278516 266156 284078 266250
tri 284078 266156 284172 266250 sw
rect 251000 263672 254172 266156
tri 251000 261156 253516 263672 ne
rect 253516 261156 254172 263672
tri 254172 261156 259172 266156 sw
tri 253516 259328 255344 261156 ne
rect 255344 260500 259172 261156
tri 259172 260500 259828 261156 sw
tri 278516 260500 284172 266156 ne
tri 284172 266034 284294 266156 sw
tri 382291 266034 382507 266250 se
rect 382507 266034 387093 266250
tri 387093 266034 387309 266250 sw
rect 284172 262437 284294 266034
tri 284294 262437 287891 266034 sw
tri 381800 265543 382291 266034 se
rect 382291 265759 387309 266034
tri 387309 265759 387584 266034 sw
rect 382291 265543 387584 265759
tri 387584 265543 387800 265759 sw
rect 284172 260500 287891 262437
tri 287891 260500 289828 262437 sw
tri 380454 260500 381800 262437 se
rect 381800 260957 387800 265543
rect 381800 260741 387584 260957
tri 387584 260741 387800 260957 nw
rect 381800 260500 387343 260741
tri 387343 260500 387584 260741 nw
rect 255344 260250 259828 260500
tri 259828 260250 260078 260500 sw
tri 284172 260250 284422 260500 ne
rect 284422 260250 387093 260500
tri 387093 260250 387343 260500 nw
rect 255344 259328 260078 260250
tri 260078 259328 261000 260250 sw
tri 284422 259328 285344 260250 ne
rect 285344 259328 382546 260250
tri 241000 258328 242000 259328 sw
tri 255344 258328 256344 259328 ne
rect 256344 258328 261000 259328
tri 261000 258328 262000 259328 sw
tri 285344 258328 286344 259328 ne
rect 286344 258328 382546 259328
rect 237000 257672 242000 258328
tri 242000 257672 242656 258328 sw
tri 256344 257672 257000 258328 ne
rect 257000 257672 262000 258328
tri 262000 257672 262656 258328 sw
tri 286344 257672 287000 258328 ne
rect 287000 257672 382546 258328
tri 237000 252672 242000 257672 ne
rect 242000 254328 242656 257672
tri 242656 254328 246000 257672 sw
tri 257000 255500 259172 257672 ne
rect 259172 256500 262656 257672
tri 262656 256500 263828 257672 sw
tri 287000 256500 288172 257672 ne
rect 288172 256500 382546 257672
tri 382546 256500 385151 260250 nw
rect 259172 255500 263828 256500
tri 263828 255500 264828 256500 sw
tri 188454 234532 189422 235500 se
rect 189422 234532 196000 235500
tri 185422 231500 188454 234532 se
rect 188454 231500 196000 234532
tri 185250 231328 185422 231500 se
rect 185422 231328 190906 231500
tri 190906 231328 191078 231500 nw
tri 184422 230500 185250 231328 se
rect 185250 230500 188454 231328
rect 167000 228876 188454 230500
tri 188454 228876 190906 231328 nw
rect 167000 226500 186078 228876
tri 186078 226500 188454 228876 nw
rect 192000 225500 196000 231500
rect 242000 235172 246000 254328
tri 259172 251500 263172 255500 ne
rect 263172 251500 282328 255500
tri 280672 250500 281672 251500 ne
rect 281672 250500 282328 251500
tri 282328 250500 287328 255500 sw
tri 281672 249844 282328 250500 ne
rect 282328 249844 379918 250500
tri 282328 247674 284498 249844 ne
rect 284498 247674 379918 249844
tri 379918 247674 382346 250500 sw
tri 284498 246500 285672 247674 ne
rect 285672 246500 382346 247674
tri 378082 244589 379723 246500 ne
rect 379723 244750 382346 246500
tri 382346 244750 384858 247674 sw
rect 379723 244589 387093 244750
tri 379723 242172 381800 244589 ne
rect 381800 244223 387093 244589
tri 387093 244223 387620 244750 sw
rect 381800 244043 387620 244223
tri 387620 244043 387800 244223 sw
rect 381800 239457 387800 244043
tri 381800 238930 382327 239457 ne
rect 382327 239277 387620 239457
tri 387620 239277 387800 239457 nw
rect 382327 238930 387273 239277
tri 387273 238930 387620 239277 nw
tri 382327 238750 382507 238930 ne
rect 382507 238750 387093 238930
tri 387093 238750 387273 238930 nw
tri 246000 235172 247656 236828 sw
tri 242000 231328 245844 235172 ne
rect 245844 231328 247656 235172
tri 247656 231328 251500 235172 sw
tri 245844 230500 246672 231328 ne
rect 246672 230500 251500 231328
tri 251500 230500 252328 231328 sw
tri 268172 230500 269000 231328 se
tri 269000 230500 269828 231328 sw
tri 200298 228876 201922 230500 se
rect 201922 228876 221000 230500
tri 246672 229516 247656 230500 ne
rect 247656 229516 271000 230500
tri 197922 226500 200298 228876 se
rect 200298 226500 221000 228876
tri 247656 228124 249048 229516 ne
rect 249048 228124 271000 229516
rect 317000 229328 377325 230500
tri 377325 229328 378503 230500 sw
tri 271000 228124 272204 229328 sw
rect 317000 228124 378503 229328
tri 378503 228124 379714 229328 sw
tri 249048 226500 250672 228124 ne
rect 250672 226500 272204 228124
tri 272204 226500 273828 228124 sw
rect 317000 226500 379714 228124
tri 379714 226500 381348 228124 sw
tri 197094 225672 197922 226500 se
rect 197922 225672 202578 226500
tri 196922 225500 197094 225672 se
rect 197094 225500 202578 225672
tri 202578 225500 203578 226500 nw
tri 268172 225672 269000 226500 ne
rect 269000 225672 273828 226500
tri 269000 225500 269172 225672 ne
rect 269172 225500 273828 225672
tri 273828 225500 274828 226500 sw
tri 375675 225898 376280 226500 ne
rect 376280 225898 381348 226500
tri 381348 225898 381954 226500 sw
tri 376280 225500 376681 225898 ne
rect 376681 225500 381954 225898
tri 381954 225500 382354 225898 sw
rect 192000 225153 202231 225500
tri 202231 225153 202578 225500 nw
tri 269172 225153 269519 225500 ne
rect 269519 225153 274828 225500
tri 274828 225153 275175 225500 sw
tri 376681 225153 377030 225500 ne
rect 377030 225153 382354 225500
tri 382354 225153 382703 225500 sw
rect 192000 223250 200328 225153
tri 200328 223250 202231 225153 nw
tri 269519 223250 271422 225153 ne
rect 271422 223250 275175 225153
tri 275175 223250 277078 225153 sw
tri 377030 224860 377325 225153 ne
rect 377325 224860 382703 225153
tri 377325 223250 378944 224860 ne
rect 378944 223250 382703 224860
tri 382703 223250 384618 225153 sw
tri 142000 219621 142551 220172 ne
rect 142551 219621 146000 220172
tri 146000 219621 148207 221828 sw
rect 192000 221500 198578 223250
tri 198578 221500 200328 223250 nw
tri 271422 222468 272204 223250 ne
rect 272204 222468 277078 223250
tri 277078 222468 277860 223250 sw
tri 378944 222697 379501 223250 ne
rect 379501 222715 387093 223250
tri 387093 222715 387628 223250 sw
rect 379501 222697 387628 222715
tri 379501 222468 379731 222697 ne
rect 379731 222543 387628 222697
tri 387628 222543 387800 222715 sw
rect 379731 222468 387800 222543
tri 272204 221500 273172 222468 ne
rect 273172 221500 277860 222468
tri 277860 221500 278828 222468 sw
tri 379731 221500 380705 222468 ne
rect 380705 221500 387800 222468
tri 11958 217250 14440 219621 ne
rect 14440 217250 17751 219621
tri 17751 217250 20233 219621 sw
tri 142551 217250 144922 219621 ne
rect 144922 217250 148207 219621
tri 148207 217250 150578 219621 sw
tri 14440 214089 17751 217250 ne
rect 17751 214089 20233 217250
tri 20233 214089 23544 217250 sw
tri 144922 216812 145360 217250 ne
rect 145360 216812 150578 217250
tri 150578 216812 151016 217250 sw
tri 145360 216172 146000 216812 ne
rect 146000 216172 151016 216812
tri 146000 214089 148083 216172 ne
rect 148083 214089 151016 216172
tri 151016 214089 153739 216812 sw
tri 17751 213250 18629 214089 ne
rect 18629 213250 23544 214089
tri 733 213076 907 213250 se
rect 907 213076 5493 213250
tri 5493 213076 5667 213250 sw
tri 18629 213076 18811 213250 ne
rect 18811 213076 23544 213250
tri 374 212717 733 213076 se
rect 733 212935 5667 213076
tri 5667 212935 5808 213076 sw
tri 18811 212935 18959 213076 ne
rect 18959 212935 23544 213076
rect 733 212717 5808 212935
tri 200 212543 374 212717 se
rect 374 212543 5808 212717
tri 5808 212543 6200 212935 sw
rect 200 207957 6200 212543
tri 18959 209942 22093 212935 ne
rect 22093 210500 23544 212935
tri 23544 210500 27302 214089 sw
tri 148083 211156 151016 214089 ne
rect 151016 211156 153739 214089
tri 153739 211156 156672 214089 sw
tri 151016 210500 151672 211156 ne
rect 151672 210500 156672 211156
tri 156672 210500 157328 211156 sw
rect 22093 209942 102328 210500
tri 200 207783 374 207957 ne
rect 374 207783 6200 207957
tri 374 207250 907 207783 ne
rect 907 207565 6200 207783
tri 6200 207565 8385 209942 sw
tri 22093 208557 23544 209942 ne
rect 23544 208557 102328 209942
tri 102328 208557 104271 210500 sw
tri 151672 208557 153615 210500 ne
rect 153615 208557 157328 210500
tri 157328 208557 159271 210500 sw
tri 23544 207565 24582 208557 ne
rect 24582 207565 104271 208557
rect 907 207250 8385 207565
tri 3241 204458 5808 207250 ne
rect 5808 204458 8385 207250
tri 8385 204458 11241 207565 sw
tri 24582 206500 25698 207565 ne
rect 25698 207156 104271 207565
tri 104271 207156 105672 208557 sw
tri 153615 207156 155016 208557 ne
rect 155016 207156 159271 208557
tri 159271 207156 160672 208557 sw
rect 25698 206500 105672 207156
tri 105672 206500 106328 207156 sw
tri 155016 206500 155672 207156 ne
rect 155672 206500 160672 207156
tri 160672 206500 161328 207156 sw
tri 100672 204458 102714 206500 ne
rect 102714 205500 106328 206500
tri 106328 205500 107328 206500 sw
tri 155672 205500 156672 206500 ne
rect 156672 205500 161328 206500
tri 161328 205500 162328 206500 sw
rect 102714 204458 144828 205500
tri 5808 201750 8297 204458 ne
rect 8297 201750 11241 204458
tri 11241 201750 13729 204458 sw
tri 102714 201750 105422 204458 ne
rect 105422 201750 144828 204458
tri 144828 201750 148578 205500 sw
tri 156672 201750 160422 205500 ne
rect 160422 201750 174828 205500
tri 174828 201750 178578 205500 sw
rect 192000 203328 196000 221500
tri 273172 216812 277860 221500 ne
rect 277860 217250 278828 221500
tri 278828 217250 283078 221500 sw
tri 380705 220412 381800 221500 ne
rect 381800 217957 387800 221500
tri 381800 217803 381954 217957 ne
rect 381954 217803 387628 217957
tri 381954 217422 382335 217803 ne
rect 382335 217785 387628 217803
tri 387628 217785 387800 217957 nw
rect 382335 217422 387265 217785
tri 387265 217422 387628 217785 nw
tri 382335 217250 382507 217422 ne
rect 382507 217250 387093 217422
tri 387093 217250 387265 217422 nw
rect 277860 216812 283078 217250
tri 283078 216812 283516 217250 sw
tri 277860 211156 283516 216812 ne
tri 283516 211156 289172 216812 sw
tri 283516 205500 289172 211156 ne
tri 289172 205500 294828 211156 sw
tri 289172 204328 290344 205500 ne
rect 290344 204328 379714 205500
tri 379714 204328 381144 205500 sw
tri 196000 203328 197000 204328 sw
tri 290344 204200 290472 204328 ne
rect 290472 204200 381144 204328
tri 381144 204200 381301 204328 sw
tri 290472 203328 291344 204200 ne
rect 291344 203328 381301 204200
tri 381301 203328 382365 204200 sw
rect 192000 202672 197000 203328
tri 197000 202672 197656 203328 sw
tri 291344 202672 292000 203328 ne
rect 292000 202672 382365 203328
tri 382365 202672 383167 203328 sw
tri 192000 201750 192922 202672 ne
rect 192922 201750 197656 202672
tri 197656 201750 198578 202672 sw
tri 292000 201750 292922 202672 ne
rect 292922 201750 383167 202672
tri 383167 201750 384293 202672 sw
tri 8297 198547 11241 201750 ne
rect 11241 200500 13729 201750
tri 13729 200500 14878 201750 sw
tri 105422 201500 105672 201750 ne
rect 105672 201500 148578 201750
tri 148578 201500 148828 201750 sw
tri 160422 201500 160672 201750 ne
rect 160672 201500 178578 201750
tri 178578 201500 178828 201750 sw
tri 192922 201500 193172 201750 ne
rect 193172 201500 198578 201750
tri 143172 200500 144172 201500 ne
rect 144172 200500 148828 201500
rect 11241 198547 99828 200500
tri 99828 198547 101781 200500 sw
tri 144172 198547 146125 200500 ne
rect 146125 198547 148828 200500
tri 11241 196500 13122 198547 ne
rect 13122 196500 101781 198547
tri 101781 196500 103828 198547 sw
tri 146125 196500 148172 198547 ne
rect 148172 196500 148828 198547
tri 98172 195750 98922 196500 ne
rect 98922 195750 103828 196500
tri 103828 195750 104578 196500 sw
tri 148172 195844 148828 196500 ne
tri 148828 195844 154484 201500 sw
tri 173172 200640 174032 201500 ne
rect 174032 200640 178828 201500
tri 178828 200640 179688 201500 sw
tri 174032 199844 174828 200640 ne
rect 174828 199844 179688 200640
tri 174828 195844 178828 199844 ne
rect 178828 197672 179688 199844
tri 179688 197672 182656 200640 sw
tri 193172 197672 197000 201500 ne
rect 197000 199328 198578 201500
tri 198578 199328 201000 201750 sw
tri 292922 201500 293172 201750 ne
rect 293172 201500 387093 201750
rect 178828 195844 182656 197672
tri 182656 195844 184484 197672 sw
tri 148828 195750 148922 195844 ne
rect 148922 195750 154484 195844
tri 154484 195750 154578 195844 sw
tri 178828 195750 178922 195844 ne
rect 178922 195750 184484 195844
tri 184484 195750 184578 195844 sw
tri 98922 192750 101922 195750 ne
rect 101922 192750 104578 195750
tri 735 192578 907 192750 se
rect 907 192578 5493 192750
tri 5493 192578 5665 192750 sw
tri 101922 192578 102094 192750 ne
rect 102094 192578 104578 192750
tri 372 192215 735 192578 se
rect 735 192326 5665 192578
tri 5665 192326 5917 192578 sw
tri 102094 192326 102346 192578 ne
rect 102346 192326 104578 192578
rect 735 192215 5917 192326
tri 200 192043 372 192215 se
rect 372 192043 5917 192215
tri 5917 192043 6200 192326 sw
rect 200 187457 6200 192043
tri 102346 190844 103828 192326 ne
rect 103828 190844 104578 192326
tri 104578 190844 109484 195750 sw
tri 148922 190844 153828 195750 ne
rect 153828 190844 154578 195750
tri 103828 189513 105159 190844 ne
rect 105159 189513 109484 190844
tri 200 187285 372 187457 ne
rect 372 187285 6200 187457
tri 372 186750 907 187285 ne
rect 907 187174 6200 187285
tri 6200 187174 8445 189513 sw
tri 105159 187174 107498 189513 ne
rect 107498 187174 109484 189513
rect 907 186750 8445 187174
tri 3308 184033 5917 186750 ne
rect 5917 184033 8445 186750
tri 8445 184033 11461 187174 sw
tri 107498 185188 109484 187174 ne
tri 109484 185188 115140 190844 sw
tri 153828 190188 154484 190844 ne
rect 154484 190188 154578 190844
tri 154578 190188 160140 195750 sw
tri 178922 194984 179688 195750 ne
rect 179688 194984 184578 195750
tri 184578 194984 185344 195750 sw
tri 179688 190188 184484 194984 ne
rect 184484 190188 185344 194984
tri 185344 190188 190140 194984 sw
tri 154484 185188 159484 190188 ne
rect 159484 185188 160140 190188
tri 109484 184033 110639 185188 ne
rect 110639 184033 115140 185188
tri 5917 180250 9548 184033 ne
rect 9548 180500 11461 184033
tri 11461 180500 14852 184033 sw
tri 110639 180500 114172 184033 ne
rect 114172 181328 115140 184033
tri 115140 181328 119000 185188 sw
tri 159484 184532 160140 185188 ne
tri 160140 184532 165796 190188 sw
tri 184484 189328 185344 190188 ne
rect 185344 189328 190140 190188
tri 190140 189328 191000 190188 sw
tri 185344 187672 187000 189328 ne
tri 160140 181328 163344 184532 ne
rect 163344 181328 165796 184532
tri 165796 181328 169000 184532 sw
rect 114172 180500 119000 181328
rect 9548 180250 71000 180500
tri 114172 180250 114422 180500 ne
rect 114422 180250 119000 180500
tri 119000 180250 120078 181328 sw
tri 163344 180250 164422 181328 ne
rect 164422 180250 169000 181328
tri 169000 180250 170078 181328 sw
tri 9548 178258 11461 180250 ne
rect 11461 178258 71000 180250
tri 114422 179532 115140 180250 ne
rect 115140 179532 120078 180250
tri 120078 179532 120796 180250 sw
tri 164422 179532 165140 180250 ne
rect 165140 179532 170078 180250
tri 11461 176500 13148 178258 ne
rect 13148 176500 71000 178258
tri 115140 176500 118172 179532 ne
rect 118172 178500 120796 179532
tri 120796 178500 121828 179532 sw
tri 165140 178876 165796 179532 ne
rect 165796 178876 170078 179532
tri 170078 178876 171452 180250 sw
rect 118172 176500 119000 178500
tri 118172 175672 119000 176500 ne
tri 119000 175672 121828 178500 nw
tri 165796 175672 169000 178876 ne
rect 169000 178500 171452 178876
tri 171452 178500 171828 178876 sw
tri 169000 175672 171828 178500 nw
tri 735 172078 907 172250 se
rect 907 172078 5493 172250
tri 5493 172078 5665 172250 sw
tri 372 171715 735 172078 se
rect 735 171715 5665 172078
tri 200 171543 372 171715 se
rect 372 171701 5665 171715
tri 5665 171701 6042 172078 sw
rect 372 171543 6042 171701
tri 6042 171543 6200 171701 sw
rect 200 166957 6200 171543
tri 200 166785 372 166957 ne
rect 372 166799 6200 166957
tri 6200 166799 8497 169085 sw
rect 372 166785 8497 166799
tri 372 166250 907 166785 ne
rect 907 166250 8497 166785
tri 3379 163600 6042 166250 ne
rect 6042 163600 8497 166250
tri 8497 163600 11712 166799 sw
tri 6042 158750 10914 163600 ne
rect 10914 160500 11712 163600
tri 11712 160500 14826 163600 sw
rect 10914 158750 139828 160500
tri 139828 158750 141578 160500 sw
tri 10914 157956 11712 158750 ne
rect 11712 157956 141578 158750
tri 141578 157956 142372 158750 sw
tri 11712 156500 13174 157956 ne
rect 13174 156500 142372 157956
tri 142372 156500 143828 157956 sw
tri 138172 152750 141922 156500 ne
rect 141922 152750 143828 156500
tri 143828 152750 147578 156500 sw
tri 141922 151750 142922 152750 ne
rect 142922 151750 147578 152750
tri 200 151043 907 151750 se
rect 907 151043 5493 151750
tri 5493 151043 6200 151750 sw
rect 200 150622 6200 151043
tri 142922 150844 143828 151750 ne
rect 143828 150844 147578 151750
tri 147578 150844 149484 152750 sw
tri 143828 150622 144050 150844 ne
rect 144050 150622 149484 150844
rect 200 150500 6210 150622
tri 6210 150500 9043 150622 sw
tri 144050 150500 144172 150622 ne
rect 144172 150500 149484 150622
rect 200 146838 99828 150500
tri 99828 146838 103490 150500 sw
tri 144172 146838 147834 150500 ne
rect 147834 146838 149484 150500
rect 200 146618 103490 146838
rect 200 146457 6200 146618
tri 6219 146500 8957 146618 ne
rect 8957 146500 103490 146618
tri 103490 146500 103828 146838 sw
tri 147834 146500 148172 146838 ne
rect 148172 146500 149484 146838
tri 200 145750 907 146457 ne
rect 907 145750 5493 146457
tri 5493 145750 6200 146457 nw
tri 98172 145750 98922 146500 ne
rect 98922 145750 103828 146500
tri 98922 140844 103828 145750 ne
tri 103828 140844 109484 146500 sw
tri 148172 145188 149484 146500 ne
tri 149484 145188 155140 150844 sw
tri 149484 140844 153828 145188 ne
rect 153828 140844 155140 145188
tri 103828 137250 107422 140844 ne
rect 107422 137250 109484 140844
tri 109484 137250 113078 140844 sw
tri 153828 139532 155140 140844 ne
tri 155140 139532 160796 145188 sw
tri 155140 137250 157422 139532 ne
rect 157422 137250 160796 139532
tri 160796 137250 163078 139532 sw
tri 107422 135188 109484 137250 ne
rect 109484 135188 113078 137250
tri 113078 135188 115140 137250 sw
tri 157422 135188 159484 137250 ne
rect 159484 135188 163078 137250
tri 109484 131250 113422 135188 ne
rect 113422 131328 115140 135188
tri 115140 131328 119000 135188 sw
tri 159484 133876 160796 135188 ne
rect 160796 133876 163078 135188
tri 163078 133876 166452 137250 sw
tri 160796 131328 163344 133876 ne
rect 163344 131328 166452 133876
rect 113422 131250 119000 131328
tri 119000 131250 119078 131328 sw
tri 163344 131250 163422 131328 ne
rect 163422 131250 166452 131328
tri 166452 131250 169078 133876 sw
tri 200 130543 907 131250 se
rect 907 130543 5493 131250
tri 5493 130543 6200 131250 sw
rect 200 130381 6200 130543
tri 113422 130500 114172 131250 ne
rect 114172 130500 119078 131250
tri 6200 130381 8957 130500 se
rect 8957 130381 71000 130500
rect 200 126500 71000 130381
tri 114172 129532 115140 130500 ne
rect 115140 129532 119078 130500
tri 119078 129532 120796 131250 sw
tri 163422 129532 165140 131250 ne
rect 165140 129532 169078 131250
tri 115140 126500 118172 129532 ne
rect 118172 128500 120796 129532
tri 120796 128500 121828 129532 sw
rect 118172 126500 119000 128500
rect 200 126378 6210 126500
tri 6210 126378 9043 126500 nw
tri 118172 126378 118294 126500 ne
rect 118294 126378 119000 126500
rect 200 125957 6200 126378
tri 200 125250 907 125957 ne
rect 907 125250 5493 125957
tri 5493 125250 6200 125957 nw
tri 118294 125672 119000 126378 ne
tri 119000 125672 121828 128500 nw
tri 165140 128220 166452 129532 ne
rect 166452 128500 169078 129532
tri 169078 128500 171828 131250 sw
rect 166452 128220 171548 128500
tri 171548 128220 171828 128500 nw
tri 166452 125672 169000 128220 ne
tri 169000 125672 171548 128220 nw
tri 185344 120172 187000 121828 se
rect 187000 120172 191000 189328
tri 182984 117812 185344 120172 se
rect 185344 117812 188640 120172
tri 188640 117812 191000 120172 nw
rect 197000 155500 201000 199328
tri 378286 199030 381301 201500 ne
rect 381301 201228 387093 201500
tri 387093 201228 387615 201750 sw
rect 381301 201043 387615 201228
tri 387615 201043 387800 201228 sw
rect 381301 199030 387800 201043
tri 381301 198621 381800 199030 ne
rect 381800 196457 387800 199030
tri 381800 195935 382322 196457 ne
rect 382322 196272 387615 196457
tri 387615 196272 387800 196457 nw
rect 382322 195935 387278 196272
tri 387278 195935 387615 196272 nw
tri 382322 195750 382507 195935 ne
rect 382507 195750 387093 195935
tri 387093 195750 387278 195935 nw
tri 217922 180250 219000 181328 se
tri 219000 180250 220078 181328 sw
tri 267922 180250 269000 181328 se
tri 269000 180250 270078 181328 sw
rect 317000 180250 385095 180500
tri 385095 180250 385255 180500 sw
tri 216548 178876 217922 180250 se
rect 217922 178876 220078 180250
tri 220078 178876 221452 180250 sw
tri 266548 178876 267922 180250 se
rect 267922 178876 270078 180250
tri 270078 178876 271452 180250 sw
rect 317000 179780 387093 180250
tri 387093 179780 387563 180250 sw
rect 317000 179543 387563 179780
tri 387563 179543 387800 179780 sw
tri 216172 178500 216548 178876 se
rect 216548 178500 221452 178876
tri 216172 177608 217064 178500 ne
rect 217064 177608 221452 178500
tri 221452 177608 222720 178876 sw
tri 266172 178500 266548 178876 se
tri 266172 178124 266548 178500 ne
rect 266548 178124 271452 178876
tri 271452 178124 272204 178876 sw
tri 266548 177608 267064 178124 ne
rect 267064 177608 272204 178124
tri 272204 177608 272720 178124 sw
tri 217064 175672 219000 177608 ne
rect 219000 175672 222720 177608
tri 222720 175672 224656 177608 sw
tri 267064 175672 269000 177608 ne
rect 269000 175672 272720 177608
tri 272720 175672 274656 177608 sw
rect 317000 176500 387800 179543
tri 219000 172250 222422 175672 ne
rect 222422 174250 224656 175672
tri 224656 174250 226078 175672 sw
tri 269000 174250 270422 175672 ne
rect 270422 174250 274656 175672
tri 274656 174250 276078 175672 sw
rect 381800 174957 387800 176500
tri 381800 174250 382507 174957 ne
rect 382507 174720 387563 174957
tri 387563 174720 387800 174957 nw
rect 382507 174487 387330 174720
tri 387330 174487 387563 174720 nw
rect 382507 174250 387093 174487
tri 387093 174250 387330 174487 nw
rect 222422 172250 226078 174250
tri 226078 172250 228078 174250 sw
tri 270422 172468 272204 174250 ne
rect 272204 172468 276078 174250
tri 276078 172468 277860 174250 sw
tri 272204 172250 272422 172468 ne
rect 272422 172250 277860 172468
tri 277860 172250 278078 172468 sw
tri 222422 172078 222594 172250 ne
rect 222594 172078 228078 172250
tri 228078 172078 228250 172250 sw
tri 272422 172078 272594 172250 ne
rect 272594 172078 278078 172250
tri 278078 172078 278250 172250 sw
tri 222594 171952 222720 172078 ne
rect 222720 171952 228250 172078
tri 228250 171952 228376 172078 sw
tri 272594 171952 272720 172078 ne
rect 272720 171952 278250 172078
tri 278250 171952 278376 172078 sw
tri 222720 171701 222971 171952 ne
rect 222971 171701 228376 171952
tri 228376 171701 228627 171952 sw
tri 272720 171701 272971 171952 ne
rect 272971 171701 278376 171952
tri 278376 171701 278627 171952 sw
tri 222971 169085 225587 171701 ne
rect 225587 169085 228627 171701
tri 228627 169085 231243 171701 sw
tri 272971 169085 275587 171701 ne
rect 275587 169085 278627 171701
tri 278627 169085 281243 171701 sw
tri 225587 166799 227873 169085 ne
rect 227873 166799 231243 169085
tri 231243 166799 233529 169085 sw
tri 275587 166812 277860 169085 ne
rect 277860 166812 281243 169085
tri 281243 166812 283516 169085 sw
tri 277860 166799 277873 166812 ne
rect 277873 166799 283516 166812
tri 283516 166799 283529 166812 sw
tri 227873 166296 228376 166799 ne
rect 228376 166296 233529 166799
tri 233529 166296 234032 166799 sw
tri 277873 166296 278376 166799 ne
rect 278376 166296 283529 166799
tri 283529 166296 284032 166799 sw
tri 228376 163600 231072 166296 ne
rect 231072 163600 234032 166296
tri 234032 163600 236728 166296 sw
tri 278376 163600 281072 166296 ne
rect 281072 163600 284032 166296
tri 284032 163600 286728 166296 sw
tri 231072 160640 234032 163600 ne
rect 234032 160640 236728 163600
tri 236728 160640 239688 163600 sw
tri 281072 161156 283516 163600 ne
rect 283516 161156 286728 163600
tri 286728 161156 289172 163600 sw
tri 283516 160640 284032 161156 ne
rect 284032 160640 289172 161156
tri 289172 160640 289688 161156 sw
tri 234032 160500 234172 160640 ne
rect 234172 160500 239688 160640
tri 239688 160500 239828 160640 sw
tri 284032 160500 284172 160640 ne
rect 284172 160500 289688 160640
tri 289688 160500 289828 160640 sw
tri 234172 158750 235922 160500 ne
rect 235922 158750 239828 160500
tri 239828 158750 241578 160500 sw
tri 284172 158750 285922 160500 ne
rect 285922 158750 289828 160500
tri 289828 158750 291578 160500 sw
tri 235922 157956 236716 158750 ne
rect 236716 157956 241578 158750
tri 241578 157956 242372 158750 sw
tri 285922 157956 286716 158750 ne
rect 286716 157956 291578 158750
tri 291578 157956 292372 158750 sw
tri 381800 158043 382507 158750 se
rect 382507 158304 387093 158750
tri 387093 158304 387539 158750 sw
rect 382507 158043 387539 158304
tri 387539 158043 387800 158304 sw
tri 236716 156500 238172 157956 ne
rect 238172 156500 242372 157956
tri 242372 156500 243828 157956 sw
tri 286716 156500 288172 157956 ne
rect 288172 156500 292372 157956
tri 292372 156500 293828 157956 sw
rect 197000 154984 227328 155500
tri 227328 154984 227844 155500 sw
tri 238172 154984 239688 156500 ne
rect 239688 154984 243828 156500
tri 243828 154984 245344 156500 sw
tri 288172 155500 289172 156500 ne
rect 289172 155500 293828 156500
tri 293828 155500 294828 156500 sw
rect 381800 155500 387800 158043
tri 289172 154984 289688 155500 ne
rect 289688 154984 387800 155500
rect 197000 153140 227844 154984
tri 227844 153140 229688 154984 sw
rect 197000 152750 229688 153140
tri 229688 152750 230078 153140 sw
tri 239688 152750 241922 154984 ne
rect 241922 152750 245344 154984
tri 245344 152750 247578 154984 sw
tri 289688 152750 291922 154984 ne
rect 291922 153457 387800 154984
rect 291922 153011 387354 153457
tri 387354 153011 387800 153457 nw
rect 291922 152750 387093 153011
tri 387093 152750 387354 153011 nw
rect 197000 151500 230078 152750
tri 177328 112156 182984 117812 se
tri 182984 112156 188640 117812 nw
tri 175922 110750 177328 112156 se
rect 177328 111828 182656 112156
tri 182656 111828 182984 112156 nw
rect 177328 110750 181578 111828
tri 181578 110750 182656 111828 nw
tri 195922 110750 197000 111828 se
rect 197000 110750 201000 151500
tri 225672 150844 226328 151500 ne
rect 226328 150844 230078 151500
tri 230078 150844 231984 152750 sw
tri 241922 150844 243828 152750 ne
rect 243828 150844 247578 152750
tri 247578 150844 249484 152750 sw
tri 291922 151500 293172 152750 ne
rect 293172 152749 385856 152750
rect 293172 151500 385412 152749
tri 385412 151500 385856 152749 nw
tri 226328 147484 229688 150844 ne
rect 229688 149328 231984 150844
tri 231984 149328 233500 150844 sw
tri 243828 149328 245344 150844 ne
rect 245344 149328 249484 150844
tri 249484 149328 251000 150844 sw
rect 229688 147672 233500 149328
tri 233500 147672 235156 149328 sw
tri 245344 147672 247000 149328 ne
rect 229688 147484 235156 147672
tri 235156 147484 235344 147672 sw
tri 229688 145188 231984 147484 ne
rect 231984 145188 235344 147484
tri 235344 145188 237640 147484 sw
tri 231984 141828 235344 145188 ne
rect 235344 141828 237640 145188
tri 237640 141828 241000 145188 sw
tri 235344 140172 237000 141828 ne
tri 215922 110750 217000 111828 se
rect 217000 110750 221000 130500
tri 713 110556 907 110750 se
rect 907 110556 5493 110750
tri 394 110237 713 110556 se
rect 713 110237 5493 110556
tri 200 110043 394 110237 se
rect 394 110043 5493 110237
tri 5493 110043 6200 110750 sw
tri 175672 110500 175922 110750 se
rect 175922 110500 181000 110750
rect 200 105500 6200 110043
tri 147319 107147 150672 110500 se
rect 150672 110172 181000 110500
tri 181000 110172 181578 110750 nw
tri 195344 110172 195922 110750 se
rect 195922 110172 201000 110750
tri 215344 110172 215922 110750 se
rect 215922 110172 221000 110750
rect 150672 107147 177975 110172
tri 177975 107147 181000 110172 nw
tri 192319 107147 195344 110172 se
rect 195344 107147 197975 110172
tri 197975 107147 201000 110172 nw
tri 212319 107147 215344 110172 se
rect 215344 109750 220578 110172
tri 220578 109750 221000 110172 nw
rect 215344 107147 217975 109750
tri 217975 107147 220578 109750 nw
tri 6200 105500 7479 107147 sw
tri 146672 106500 147319 107147 se
rect 147319 107140 177968 107147
tri 177968 107140 177975 107147 nw
tri 192312 107140 192319 107147 se
rect 192319 107140 197968 107147
tri 197968 107140 197975 107147 nw
tri 212312 107140 212319 107147 se
rect 212319 107140 217968 107147
tri 217968 107140 217975 107147 nw
rect 147319 106500 177328 107140
tri 177328 106500 177968 107140 nw
tri 146656 106484 146672 106500 se
rect 146672 106484 152312 106500
tri 152312 106484 152328 106500 nw
tri 145672 105500 146656 106484 se
rect 146656 106172 152000 106484
tri 152000 106172 152312 106484 nw
tri 191344 106172 192312 107140 se
rect 192312 106172 197000 107140
tri 197000 106172 197968 107140 nw
rect 146656 105500 151328 106172
tri 151328 105500 152000 106172 nw
tri 190672 105500 191344 106172 se
rect 191344 105500 196328 106172
tri 196328 105500 197000 106172 nw
tri 210672 105500 212312 107140 se
rect 212312 105500 216328 107140
tri 216328 105500 217968 107140 nw
rect 200 105457 94828 105500
tri 200 105263 394 105457 ne
rect 394 105263 94828 105457
tri 394 104750 907 105263 ne
rect 907 104750 94828 105263
tri 94828 104750 95578 105500 sw
tri 144922 104750 145672 105500 se
rect 145672 104750 150578 105500
tri 150578 104750 151328 105500 nw
tri 189922 104750 190672 105500 se
rect 190672 104750 195578 105500
tri 195578 104750 196328 105500 nw
tri 209922 104750 210672 105500 se
rect 210672 104750 215578 105500
tri 215578 104750 216328 105500 nw
tri 2997 101582 5458 104750 ne
rect 5458 101582 95578 104750
tri 95578 101582 98746 104750 sw
tri 141754 101582 144922 104750 se
rect 144922 101582 147410 104750
tri 147410 101582 150578 104750 nw
tri 186754 101582 189922 104750 se
rect 189922 101582 192410 104750
tri 192410 101582 195578 104750 nw
tri 206754 101582 209922 104750 se
rect 209922 101582 212410 104750
tri 212410 101582 215578 104750 nw
tri 5458 101500 5521 101582 ne
rect 5521 101500 98746 101582
tri 98746 101500 98828 101582 sw
tri 141672 101500 141754 101582 se
rect 141754 101500 147328 101582
tri 147328 101500 147410 101582 nw
tri 186672 101500 186754 101582 se
rect 186754 101500 192328 101582
tri 192328 101500 192410 101582 nw
tri 206672 101500 206754 101582 se
rect 206754 101500 212328 101582
tri 212328 101500 212410 101582 nw
tri 93172 95844 98828 101500 ne
tri 98828 95844 104484 101500 sw
tri 141000 100828 141672 101500 se
rect 141672 101484 147312 101500
tri 147312 101484 147328 101500 nw
tri 186656 101484 186672 101500 se
rect 186672 101484 192312 101500
tri 192312 101484 192328 101500 nw
tri 206656 101484 206672 101500 se
rect 206672 101484 212312 101500
tri 212312 101484 212328 101500 nw
rect 141672 100828 146656 101484
tri 146656 100828 147312 101484 nw
tri 137000 96828 141000 100828 se
rect 141000 100516 146344 100828
tri 146344 100516 146656 100828 nw
tri 185688 100516 186656 101484 se
rect 186656 100516 191344 101484
tri 191344 100516 192312 101484 nw
rect 141000 100500 146328 100516
tri 146328 100500 146344 100516 nw
tri 185672 100500 185688 100516 se
rect 185688 100500 186672 100516
rect 141000 96828 142328 100500
rect 137000 96500 142328 96828
tri 142328 96500 146328 100500 nw
tri 151672 96500 155672 100500 se
rect 155672 97796 177328 100500
tri 177328 97796 180032 100500 sw
tri 182968 97796 185672 100500 se
rect 185672 97796 186672 100500
rect 155672 96500 180032 97796
tri 180032 96500 181328 97796 sw
tri 181672 96500 182968 97796 se
rect 182968 96500 186672 97796
rect 137000 95844 141672 96500
tri 141672 95844 142328 96500 nw
tri 151016 95844 151672 96500 se
rect 151672 95844 156672 96500
tri 156672 95844 157328 96500 nw
tri 175672 95844 176328 96500 ne
rect 176328 96328 181328 96500
tri 181328 96328 181500 96500 sw
tri 181500 96328 181672 96500 se
rect 181672 96328 186672 96500
rect 176328 95844 186672 96328
tri 186672 95844 191344 100516 nw
tri 201016 95844 206656 101484 se
rect 206656 95844 206672 101484
tri 206672 95844 212312 101484 nw
tri 98828 94250 100422 95844 ne
rect 100422 94250 104484 95844
tri 104484 94250 106078 95844 sw
rect 137000 95828 141656 95844
tri 141656 95828 141672 95844 nw
tri 151000 95828 151016 95844 se
rect 151016 95828 156656 95844
tri 156656 95828 156672 95844 nw
tri 176328 95828 176344 95844 ne
rect 176344 95828 186656 95844
tri 186656 95828 186672 95844 nw
tri 201000 95828 201016 95844 se
rect 201016 95828 206656 95844
tri 206656 95828 206672 95844 nw
tri 100422 90250 104422 94250 ne
rect 104422 90250 106078 94250
tri 734 90077 907 90250 se
rect 907 90077 5493 90250
tri 5493 90077 5666 90250 sw
tri 104422 90188 104484 90250 ne
rect 104484 90188 106078 90250
tri 106078 90188 110140 94250 sw
tri 104484 90077 104595 90188 ne
rect 104595 90077 110140 90188
tri 373 89716 734 90077 se
rect 734 89857 5666 90077
tri 5666 89857 5886 90077 sw
tri 104595 89857 104815 90077 ne
rect 104815 89857 110140 90077
rect 734 89716 5886 89857
tri 200 89543 373 89716 se
rect 373 89543 5886 89716
tri 5886 89543 6200 89857 sw
rect 200 84957 6200 89543
tri 104815 88250 106422 89857 ne
rect 106422 88250 110140 89857
tri 110140 88250 112078 90188 sw
tri 106422 86993 107679 88250 ne
rect 107679 86993 112078 88250
tri 200 84784 373 84957 ne
rect 373 84784 6200 84957
tri 373 84250 907 84784 ne
rect 907 84643 6200 84784
tri 6200 84643 8429 86993 sw
tri 107679 84643 110029 86993 ne
rect 110029 84643 112078 86993
rect 907 84250 8429 84643
tri 3289 81513 5886 84250 ne
rect 5886 82313 8429 84250
tri 8429 82313 10640 84643 sw
tri 110029 84532 110140 84643 ne
rect 110140 84532 112078 84643
tri 112078 84532 115796 88250 sw
tri 110140 82313 112359 84532 ne
rect 112359 82313 115796 84532
rect 5886 81514 10640 82313
tri 10640 81514 11398 82313 sw
rect 5886 81513 11398 81514
tri 112359 81513 113159 82313 ne
rect 113159 81513 115796 82313
tri 5886 76500 10640 81513 ne
rect 10640 80500 11398 81513
tri 11398 80500 12360 81513 sw
tri 113159 80500 114172 81513 ne
rect 114172 81328 115796 81513
tri 115796 81328 119000 84532 sw
rect 114172 80500 119000 81328
rect 10640 76500 71000 80500
tri 114172 78876 115796 80500 ne
rect 115796 78876 119000 80500
tri 119000 78876 121452 81328 sw
tri 115796 76500 118172 78876 ne
rect 118172 78500 121452 78876
tri 121452 78500 121828 78876 sw
rect 118172 76500 119000 78500
tri 118172 75672 119000 76500 ne
tri 119000 75672 121828 78500 nw
tri 135344 70172 137000 71828 se
rect 137000 70172 141000 95828
tri 141000 95172 141656 95828 nw
tri 149422 94250 151000 95828 se
rect 151000 94250 155078 95828
tri 155078 94250 156656 95828 nw
tri 176344 94250 177922 95828 ne
rect 177922 94860 185688 95828
tri 185688 94860 186656 95828 nw
rect 177922 94250 185078 94860
tri 185078 94250 185688 94860 nw
tri 199422 94250 201000 95828 se
rect 201000 94250 205078 95828
tri 205078 94250 206656 95828 nw
tri 134922 69750 135344 70172 se
rect 135344 69750 140578 70172
tri 140578 69750 141000 70172 nw
tri 147000 91828 149422 94250 se
rect 149422 91828 151016 94250
rect 147000 90188 151016 91828
tri 151016 90188 155078 94250 nw
tri 177922 93500 178672 94250 ne
rect 178672 93500 184328 94250
tri 184328 93500 185078 94250 nw
tri 178672 90844 181328 93500 ne
rect 181328 92750 184328 93500
tri 184328 92750 185078 93500 sw
rect 181328 92140 185078 92750
tri 185078 92140 185688 92750 sw
rect 181328 90844 185688 92140
tri 185688 90844 186984 92140 sw
tri 197000 91828 199422 94250 se
rect 199422 94078 204906 94250
tri 204906 94078 205078 94250 nw
rect 199422 91828 201973 94078
rect 197000 91145 201973 91828
tri 201973 91145 204906 94078 nw
tri 181328 90672 181500 90844 ne
rect 181500 90672 186984 90844
tri 181500 90188 181984 90672 ne
rect 181984 90188 186984 90672
tri 735 69578 907 69750 se
rect 907 69578 5493 69750
tri 5493 69578 5665 69750 sw
tri 372 69215 735 69578 se
rect 735 69215 5665 69578
tri 200 69043 372 69215 se
rect 372 69204 5665 69215
tri 5665 69204 6039 69578 sw
rect 372 69043 6039 69204
tri 6039 69043 6200 69204 sw
rect 200 64457 6200 69043
tri 132984 67812 134922 69750 se
rect 134922 67812 138640 69750
tri 138640 67812 140578 69750 nw
tri 200 64285 372 64457 ne
rect 372 64296 6200 64457
tri 6200 64296 8497 66584 sw
tri 129468 64296 132984 67812 se
rect 132984 66828 137656 67812
tri 137656 66828 138640 67812 nw
rect 132984 65172 136000 66828
tri 136000 65172 137656 66828 nw
tri 145344 65172 147000 66828 se
rect 147000 65172 151000 90188
tri 151000 90172 151016 90188 nw
tri 181984 90172 182000 90188 ne
rect 182000 90172 186984 90188
tri 182000 88250 183922 90172 ne
rect 183922 88250 186984 90172
tri 183922 85188 186984 88250 ne
tri 186984 86828 191000 90844 sw
rect 186984 85188 191000 86828
tri 186984 85172 187000 85188 ne
tri 166548 78876 169000 81328 se
tri 169000 78876 171452 81328 sw
tri 166172 78500 166548 78876 se
rect 166548 78500 171452 78876
tri 171452 78500 171828 78876 sw
tri 164156 76484 166172 78500 se
rect 166172 76484 169812 78500
tri 169812 76484 171828 78500 nw
tri 163344 75672 164156 76484 se
rect 164156 75672 169000 76484
tri 169000 75672 169812 76484 nw
tri 158500 70828 163344 75672 se
rect 163344 72750 166078 75672
tri 166078 72750 169000 75672 nw
rect 163344 70828 164156 72750
tri 164156 70828 166078 72750 nw
tri 157422 69750 158500 70828 se
rect 158500 69750 163078 70828
tri 163078 69750 164156 70828 nw
rect 132984 64296 135124 65172
tri 135124 64296 136000 65172 nw
rect 372 64285 8497 64296
tri 372 63750 907 64285 ne
rect 907 63750 8497 64285
tri 3378 63468 3661 63750 ne
rect 3661 63468 8497 63750
tri 3661 61100 6039 63468 ne
rect 6039 62156 8497 63468
tri 8497 62156 10645 64296 sw
tri 127328 62156 129468 64296 se
rect 129468 63750 134578 64296
tri 134578 63750 135124 64296 nw
tri 143922 63750 145344 65172 se
rect 145344 63750 149578 65172
tri 149578 63750 151000 65172 nw
tri 154500 66828 157422 69750 se
rect 157422 66828 160078 69750
rect 154500 66750 160078 66828
tri 160078 66750 163078 69750 nw
tri 186922 66750 187000 66828 se
rect 187000 66750 191000 85188
rect 129468 63468 134296 63750
tri 134296 63468 134578 63750 nw
tri 143640 63468 143922 63750 se
rect 143922 63468 149296 63750
tri 149296 63468 149578 63750 nw
rect 129468 62156 132984 63468
tri 132984 62156 134296 63468 nw
tri 142328 62156 143640 63468 se
rect 143640 62156 147656 63468
rect 6039 61100 10645 62156
tri 10645 61100 11706 62156 sw
tri 126272 61100 127328 62156 se
rect 127328 61100 131928 62156
tri 131928 61100 132984 62156 nw
tri 6039 57812 9339 61100 ne
rect 9339 60500 11706 61100
tri 11706 60500 12308 61100 sw
tri 125672 60500 126272 61100 se
rect 126272 60500 128640 61100
rect 9339 57812 12308 60500
tri 9339 55454 11706 57812 ne
rect 11706 56500 12308 57812
tri 12308 56500 16322 60500 sw
tri 89172 56500 93172 60500 se
rect 93172 57812 128640 60500
tri 128640 57812 131928 61100 nw
tri 137984 57812 142328 62156 se
rect 142328 61828 147656 62156
tri 147656 61828 149296 63468 nw
rect 142328 60172 146000 61828
tri 146000 60172 147656 61828 nw
tri 152844 60172 154500 61828 se
rect 154500 60172 158500 66750
tri 158500 65172 160078 66750 nw
tri 185344 65172 186922 66750 se
rect 186922 65172 191000 66750
tri 181344 61172 185344 65172 se
rect 185344 61172 187000 65172
tri 187000 61172 191000 65172 nw
rect 197000 90188 201016 91145
tri 201016 90188 201973 91145 nw
rect 142328 59640 145468 60172
tri 145468 59640 146000 60172 nw
tri 152312 59640 152844 60172 se
rect 152844 59640 157968 60172
tri 157968 59640 158500 60172 nw
tri 179812 59640 181344 61172 se
rect 142328 57812 143640 59640
tri 143640 57812 145468 59640 nw
tri 150484 57812 152312 59640 se
rect 152312 57812 153828 59640
rect 93172 56500 127328 57812
tri 127328 56500 128640 57812 nw
tri 136672 56500 137984 57812 se
rect 137984 56500 139812 57812
rect 11706 55500 16322 56500
tri 16322 55500 17326 56500 sw
tri 88172 55500 89172 56500 se
rect 89172 55500 93782 56500
rect 11706 55454 93782 55500
tri 93782 55454 94828 56500 nw
tri 11706 52156 15015 55454 ne
rect 15015 52156 90484 55454
tri 90484 52156 93782 55454 nw
tri 132328 52156 136672 56500 se
rect 136672 53984 139812 56500
tri 139812 53984 143640 57812 nw
tri 146656 53984 150484 57812 se
rect 150484 55500 153828 57812
tri 153828 55500 157968 59640 nw
tri 175688 55516 179812 59640 se
rect 179812 55516 181344 59640
tri 181344 55516 187000 61172 nw
tri 175672 55500 175688 55516 se
rect 175688 55500 181328 55516
tri 181328 55500 181344 55516 nw
rect 150484 53984 152312 55500
tri 152312 53984 153828 55500 nw
tri 161656 53984 163172 55500 se
rect 163172 53984 177328 55500
rect 136672 52156 137984 53984
tri 137984 52156 139812 53984 nw
tri 144828 52156 146656 53984 se
rect 146656 52156 149578 53984
tri 15015 51500 15674 52156 ne
rect 15674 51500 89828 52156
tri 89828 51500 90484 52156 nw
tri 130672 50500 132328 52156 se
rect 132328 50500 135078 52156
tri 99422 49250 100672 50500 se
rect 100672 49250 135078 50500
tri 135078 49250 137984 52156 nw
tri 141922 49250 144828 52156 se
rect 144828 51250 149578 52156
tri 149578 51250 152312 53984 nw
tri 158922 51250 161656 53984 se
rect 161656 51500 177328 53984
tri 177328 51500 181328 55500 nw
rect 161656 51250 163172 51500
rect 144828 49250 147578 51250
tri 147578 49250 149578 51250 nw
tri 157516 49844 158922 51250 se
rect 158922 49844 163172 51250
tri 163172 49844 164828 51500 nw
tri 156922 49250 157516 49844 se
tri 735 49078 907 49250 se
rect 907 49078 5493 49250
tri 5493 49078 5665 49250 sw
tri 99250 49078 99422 49250 se
rect 99422 49078 134906 49250
tri 134906 49078 135078 49250 nw
tri 141750 49078 141922 49250 se
rect 141922 49078 147406 49250
tri 147406 49078 147578 49250 nw
tri 156750 49078 156922 49250 se
rect 156922 49078 157516 49250
tri 372 48715 735 49078 se
rect 735 48715 5665 49078
tri 200 48543 372 48715 se
rect 372 48625 5665 48715
tri 5665 48625 6118 49078 sw
tri 98797 48625 99250 49078 se
rect 99250 48625 134453 49078
tri 134453 48625 134906 49078 nw
tri 141297 48625 141750 49078 se
rect 141750 48625 146953 49078
tri 146953 48625 147406 49078 nw
tri 156297 48625 156750 49078 se
rect 156750 48625 157516 49078
rect 372 48543 6118 48625
tri 6118 48543 6200 48625 sw
rect 200 45250 6200 48543
tri 96672 46500 98797 48625 se
rect 98797 48328 134156 48625
tri 134156 48328 134453 48625 nw
tri 141000 48328 141297 48625 se
rect 141297 48328 146656 48625
tri 146656 48328 146953 48625 nw
tri 156000 48328 156297 48625 se
rect 156297 48328 157516 48625
rect 98797 46500 132328 48328
tri 132328 46500 134156 48328 nw
tri 96299 46127 96672 46500 se
rect 96672 46127 101955 46500
tri 101955 46127 102328 46500 nw
tri 138799 46127 141000 48328 se
rect 141000 46127 144455 48328
tri 144455 46127 146656 48328 nw
tri 153799 46127 156000 48328 se
rect 156000 46127 157516 48328
tri 6200 45250 7104 46127 sw
tri 96000 45828 96299 46127 se
rect 96299 45828 101656 46127
tri 101656 45828 101955 46127 nw
tri 95422 45250 96000 45828 se
rect 96000 45250 101078 45828
tri 101078 45250 101656 45828 nw
tri 137922 45250 138799 46127 se
rect 138799 45250 143578 46127
tri 143578 45250 144455 46127 nw
tri 152922 45250 153799 46127 se
rect 153799 45250 157516 46127
rect 200 43957 7104 45250
tri 200 43785 372 43957 ne
rect 372 43875 7104 43957
tri 7104 43875 8522 45250 sw
tri 94047 43875 95422 45250 se
rect 95422 43875 99703 45250
tri 99703 43875 101078 45250 nw
tri 137000 44328 137922 45250 se
rect 137922 44328 142203 45250
rect 137000 43875 142203 44328
tri 142203 43875 143578 45250 nw
tri 151860 44188 152922 45250 se
rect 152922 44188 157516 45250
tri 157516 44188 163172 49844 nw
tri 151547 43875 151860 44188 se
rect 151860 43875 152656 44188
rect 372 43785 8522 43875
tri 372 43250 907 43785 ne
rect 907 43250 8522 43785
tri 3420 40634 6118 43250 ne
rect 6118 40634 8522 43250
tri 8522 40634 11864 43875 sw
tri 92000 41828 94047 43875 se
rect 94047 41828 96462 43875
rect 92000 40634 96462 41828
tri 96462 40634 99703 43875 nw
tri 6118 35061 11864 40634 ne
tri 11864 35061 17610 40634 sw
tri 11864 29487 17610 35061 ne
tri 17610 30500 22311 35061 sw
rect 17610 29487 71000 30500
tri 17610 26500 20689 29487 ne
rect 20689 26500 71000 29487
tri 91672 26500 92000 26828 se
rect 92000 26500 96000 40634
tri 96000 40172 96462 40634 nw
tri 118172 30500 119000 31328 se
tri 119000 30500 119828 31328 sw
tri 116172 28500 118172 30500 se
rect 118172 28500 119828 30500
tri 119828 28500 121828 30500 sw
tri 114172 26500 116172 28500 se
rect 116172 26500 119828 28500
tri 119828 26500 121828 28500 nw
tri 90344 25172 91672 26500 se
rect 91672 25172 96000 26500
tri 88640 23468 90344 25172 se
rect 90344 23468 94296 25172
tri 94296 23468 96000 25172 nw
tri 111140 23468 114172 26500 se
rect 114172 23468 116796 26500
tri 116796 23468 119828 26500 nw
tri 82984 17812 88640 23468 se
tri 88640 17812 94296 23468 nw
tri 105484 17812 111140 23468 se
tri 111140 17812 116796 23468 nw
tri 135484 17812 137000 19328 se
rect 137000 17812 141000 43875
tri 141000 42672 142203 43875 nw
tri 150344 42672 151547 43875 se
rect 151547 42672 152656 43875
tri 77328 12156 82984 17812 se
tri 82984 12156 88640 17812 nw
tri 99828 12156 105484 17812 se
tri 105484 12156 111140 17812 nw
tri 135344 17672 135484 17812 se
rect 135484 17672 141000 17812
tri 129828 12156 135344 17672 se
rect 135344 12156 135484 17672
tri 135484 12156 141000 17672 nw
tri 147000 39328 150344 42672 se
rect 150344 39328 152656 42672
tri 152656 39328 157516 44188 nw
tri 144841 12156 147000 14326 se
rect 147000 12674 151000 39328
tri 151000 37672 152656 39328 nw
tri 195344 32672 197000 34328 se
rect 197000 32672 201000 90188
tri 201000 90172 201016 90188 nw
rect 217000 60172 221000 80500
rect 237000 66156 241000 141828
rect 247000 67672 251000 149328
tri 382335 137078 382507 137250 se
rect 382507 137078 387093 137250
tri 387093 137078 387265 137250 sw
tri 381800 136543 382335 137078 se
rect 382335 136715 387265 137078
tri 387265 136715 387628 137078 sw
rect 382335 136543 387628 136715
tri 387628 136543 387800 136715 sw
tri 381583 133876 381800 134091 se
rect 381800 133876 387800 136543
tri 379132 131446 381583 133876 se
rect 381583 131957 387800 133876
rect 381583 131785 387628 131957
tri 387628 131785 387800 131957 nw
rect 381583 131446 387289 131785
tri 387289 131446 387628 131785 nw
tri 379013 131328 379132 131446 se
rect 379132 131328 387093 131446
tri 268922 131250 269000 131328 se
tri 269000 131250 269078 131328 sw
tri 378934 131250 379013 131328 se
rect 379013 131250 387093 131328
tri 387093 131250 387289 131446 nw
tri 268172 130500 268922 131250 se
rect 268922 130500 269078 131250
tri 269078 130500 269828 131250 sw
tri 378177 130500 378934 131250 se
rect 378934 130500 383858 131250
tri 383858 130500 384614 131250 nw
tri 266172 128500 268172 130500 se
rect 268172 128500 269828 130500
tri 266172 128124 266548 128500 ne
rect 266548 128124 269828 128500
tri 269828 128124 272204 130500 sw
rect 317000 128124 381461 130500
tri 381461 128124 383858 130500 nw
tri 266548 125672 269000 128124 ne
rect 269000 125672 272204 128124
tri 269000 122468 272204 125672 ne
tri 272204 122468 277860 128124 sw
rect 317000 126500 379823 128124
tri 379823 126500 381461 128124 nw
tri 272204 116812 277860 122468 ne
tri 277860 116812 283516 122468 sw
tri 277860 111156 283516 116812 ne
tri 283516 115750 284578 116812 sw
rect 283516 115574 284578 115750
tri 284578 115574 284754 115750 sw
tri 382331 115574 382507 115750 se
rect 382507 115574 387093 115750
tri 387093 115574 387269 115750 sw
rect 283516 112401 284754 115574
tri 284754 112401 287927 115574 sw
tri 381800 115043 382331 115574 se
rect 382331 115219 387269 115574
tri 387269 115219 387624 115574 sw
rect 382331 115043 387624 115219
tri 387624 115043 387800 115219 sw
rect 283516 111156 287927 112401
tri 287927 111156 289172 112401 sw
tri 283516 109750 284922 111156 ne
rect 284922 109750 289172 111156
tri 289172 109750 290578 111156 sw
tri 379421 109750 381800 112401 se
rect 381800 110457 387800 115043
rect 381800 110281 387624 110457
tri 387624 110281 387800 110457 nw
rect 381800 109750 387093 110281
tri 387093 109750 387624 110281 nw
tri 284922 107147 287525 109750 ne
rect 287525 109584 290578 109750
tri 290578 109584 290744 109750 sw
tri 379272 109584 379421 109750 se
rect 379421 109584 384647 109750
tri 384647 109584 384796 109750 nw
rect 287525 107147 290744 109584
tri 290744 107147 293181 109584 sw
tri 377085 107147 379272 109584 se
rect 379272 107147 380982 109584
tri 287525 107140 287532 107147 ne
rect 287532 107140 293181 107147
tri 293181 107140 293188 107147 sw
tri 377079 107140 377085 107147 se
rect 377085 107140 380982 107147
tri 287532 105500 289172 107140 ne
rect 289172 105500 293188 107140
tri 293188 105500 294828 107140 sw
tri 375607 105500 377079 107140 se
rect 377079 105500 380982 107140
tri 380982 105500 384647 109584 nw
tri 289172 104750 289922 105500 ne
rect 289922 104750 377393 105500
tri 289922 101582 293090 104750 ne
rect 293090 101582 377393 104750
tri 293090 101500 293172 101582 ne
rect 293172 101500 377393 101582
tri 377393 101500 380982 105500 nw
tri 382335 94078 382507 94250 se
rect 382507 94078 387093 94250
tri 387093 94078 387265 94250 sw
tri 381800 93543 382335 94078 se
rect 382335 93715 387265 94078
tri 387265 93715 387628 94078 sw
rect 382335 93543 387628 93715
tri 387628 93543 387800 93715 sw
tri 380802 90188 381800 91145 se
rect 381800 90188 387800 93543
tri 379079 88536 380802 90188 se
rect 380802 88957 387800 90188
rect 380802 88785 387628 88957
tri 387628 88785 387800 88957 nw
rect 380802 88536 387379 88785
tri 387379 88536 387628 88785 nw
tri 378781 88250 379079 88536 se
rect 379079 88250 387093 88536
tri 387093 88250 387379 88536 nw
tri 374902 84532 378781 88250 se
rect 378781 84532 379079 88250
tri 373298 82994 374902 84532 se
rect 374902 82994 379079 84532
tri 379079 82994 384562 88250 nw
tri 371560 81328 373298 82994 se
rect 373298 81328 376477 82994
tri 370696 80500 371560 81328 se
rect 371560 80500 376477 81328
tri 376477 80500 379079 82994 nw
rect 267000 77468 287328 80500
tri 287328 77468 290360 80500 sw
rect 317000 77468 373314 80500
tri 373314 77468 376477 80500 nw
rect 267000 76500 290360 77468
tri 285672 71812 290360 76500 ne
tri 290360 72750 295078 77468 sw
rect 317000 76500 372304 77468
tri 372304 76500 373314 77468 nw
rect 290360 72578 295078 72750
tri 295078 72578 295250 72750 sw
tri 382335 72578 382507 72750 se
rect 382507 72578 387093 72750
tri 387093 72578 387265 72750 sw
rect 290360 71812 295250 72578
tri 295250 71812 296016 72578 sw
tri 381800 72043 382335 72578 se
rect 382335 72215 387265 72578
tri 387265 72215 387628 72578 sw
rect 382335 72043 387628 72215
tri 387628 72043 387800 72215 sw
tri 241000 66156 241672 66828 sw
tri 247000 66156 248516 67672 ne
rect 248516 66156 251000 67672
tri 251000 66156 254172 69328 sw
tri 290360 66156 296016 71812 ne
tri 296016 69513 298315 71812 sw
rect 296016 66801 298315 69513
tri 298315 66801 301027 69513 sw
tri 379197 66801 381800 69513 se
rect 381800 67457 387800 72043
rect 381800 67285 387628 67457
tri 387628 67285 387800 67457 nw
rect 381800 66801 387144 67285
tri 387144 66801 387628 67285 nw
rect 296016 66750 301027 66801
tri 301027 66750 301078 66801 sw
tri 379148 66750 379197 66801 se
rect 379197 66750 387093 66801
tri 387093 66750 387144 66801 nw
rect 296016 66156 301078 66750
tri 301078 66156 301672 66750 sw
rect 237000 65172 241672 66156
tri 237000 61828 240344 65172 ne
rect 240344 63672 241672 65172
tri 241672 63672 244156 66156 sw
tri 248516 63672 251000 66156 ne
rect 251000 63672 254172 66156
rect 240344 61828 244156 63672
tri 244156 61828 246000 63672 sw
tri 251000 61828 252844 63672 ne
rect 252844 61828 254172 63672
tri 254172 61828 258500 66156 sw
tri 296016 61828 300344 66156 ne
rect 300344 61828 301672 66156
tri 301672 61828 306000 66156 sw
tri 374424 61828 379148 66750 se
rect 379148 61828 379197 66750
tri 217000 59640 217532 60172 ne
rect 217532 59640 221000 60172
tri 221000 59640 223188 61828 sw
tri 240344 61812 240360 61828 ne
rect 240360 61812 246000 61828
tri 246000 61812 246016 61828 sw
tri 240360 61172 241000 61812 ne
rect 241000 61172 246016 61812
tri 241000 59640 242532 61172 ne
rect 242532 60500 246016 61172
tri 246016 60500 247328 61812 sw
tri 252844 60500 254172 61828 ne
rect 254172 60500 258500 61828
tri 258500 60500 259828 61828 sw
tri 300344 60500 301672 61828 ne
rect 301672 61025 306000 61828
tri 306000 61025 306803 61828 sw
tri 373653 61025 374424 61828 se
rect 374424 61025 379197 61828
tri 379197 61025 384693 66750 nw
rect 301672 60500 306803 61025
tri 306803 60500 307328 61025 sw
tri 373148 60500 373653 61025 se
rect 373653 60500 378693 61025
tri 378693 60500 379197 61025 nw
rect 242532 59640 247328 60500
tri 247328 59640 248188 60500 sw
tri 254172 59640 255032 60500 ne
rect 255032 59640 289828 60500
tri 289828 59640 290688 60500 sw
tri 301672 59640 302532 60500 ne
rect 302532 59640 374852 60500
tri 217532 59452 217720 59640 ne
rect 217720 59452 223188 59640
tri 223188 59452 223376 59640 sw
tri 242532 59452 242720 59640 ne
rect 242720 59452 248188 59640
tri 248188 59452 248376 59640 sw
tri 255032 59452 255220 59640 ne
rect 255220 59452 290688 59640
tri 290688 59452 290876 59640 sw
tri 302532 59452 302720 59640 ne
rect 302720 59452 374852 59640
tri 217720 56172 221000 59452 ne
rect 221000 56172 223376 59452
tri 221000 53984 223188 56172 ne
rect 223188 53984 223376 56172
tri 223376 53984 228844 59452 sw
tri 242720 56156 246016 59452 ne
rect 246016 56500 248376 59452
tri 248376 56500 251328 59452 sw
tri 255220 56500 258172 59452 ne
rect 258172 56500 290876 59452
tri 290876 56500 293828 59452 sw
tri 302720 56500 305672 59452 ne
rect 305672 56500 374852 59452
tri 374852 56500 378693 60500 nw
rect 246016 56156 251328 56500
tri 251328 56156 251672 56500 sw
tri 288172 56156 288516 56500 ne
rect 288516 56156 293828 56500
tri 293828 56156 294172 56500 sw
tri 246016 53984 248188 56156 ne
rect 248188 54844 251672 56156
tri 251672 54844 252984 56156 sw
tri 288516 54844 289828 56156 ne
rect 289828 54844 294172 56156
rect 248188 53984 252984 54844
tri 252984 53984 253844 54844 sw
tri 289828 53984 290688 54844 ne
rect 290688 53984 294172 54844
tri 294172 53984 296344 56156 sw
tri 223188 53796 223376 53984 ne
rect 223376 53796 228844 53984
tri 228844 53796 229032 53984 sw
tri 248188 53796 248376 53984 ne
rect 248376 53796 253844 53984
tri 253844 53796 254032 53984 sw
tri 290688 53796 290876 53984 ne
rect 290876 53796 296344 53984
tri 296344 53796 296532 53984 sw
tri 223376 51250 225922 53796 ne
rect 225922 51250 229032 53796
tri 229032 51250 231578 53796 sw
tri 248376 51250 250922 53796 ne
rect 250922 51250 254032 53796
tri 254032 51250 256578 53796 sw
tri 290876 51250 293422 53796 ne
rect 293422 51250 296532 53796
tri 296532 51250 299078 53796 sw
tri 225922 49250 227922 51250 ne
rect 227922 49250 231578 51250
tri 231578 49250 233578 51250 sw
tri 250922 50500 251672 51250 ne
rect 251672 50500 256578 51250
tri 256578 50500 257328 51250 sw
tri 293422 50500 294172 51250 ne
rect 294172 50500 299078 51250
tri 299078 50500 299828 51250 sw
tri 381800 50543 382507 51250 se
rect 382507 50543 387093 51250
tri 387093 50543 387800 51250 sw
tri 251672 49250 252922 50500 ne
rect 252922 50162 284828 50500
tri 284828 50162 285166 50500 sw
tri 294172 50162 294510 50500 ne
rect 294510 50381 379043 50500
tri 379043 50381 381800 50500 sw
rect 381800 50381 387800 50543
rect 294510 50162 387800 50381
rect 252922 49250 285166 50162
tri 285166 49250 286078 50162 sw
tri 294510 49250 295422 50162 ne
rect 295422 49250 387800 50162
tri 227922 49078 228094 49250 ne
rect 228094 49078 233578 49250
tri 233578 49078 233750 49250 sw
tri 252922 49078 253094 49250 ne
rect 253094 49078 286078 49250
tri 286078 49078 286250 49250 sw
tri 295422 49078 295594 49250 ne
rect 295594 49078 387800 49250
tri 228094 48625 228547 49078 ne
rect 228547 48625 233750 49078
tri 233750 48625 234203 49078 sw
tri 253094 48625 253547 49078 ne
rect 253547 48625 286250 49078
tri 286250 48625 286703 49078 sw
tri 295594 48625 296047 49078 ne
rect 296047 48625 387800 49078
tri 228547 48328 228844 48625 ne
rect 228844 48328 234203 48625
tri 234203 48328 234500 48625 sw
tri 253547 48328 253844 48625 ne
rect 253844 48328 286703 48625
tri 286703 48328 287000 48625 sw
tri 296047 48328 296344 48625 ne
rect 296344 48328 387800 48625
tri 228844 48140 229032 48328 ne
rect 229032 48140 234500 48328
tri 234500 48140 234688 48328 sw
tri 253844 48140 254032 48328 ne
rect 254032 48140 287000 48328
tri 287000 48140 287188 48328 sw
tri 296344 48140 296532 48328 ne
rect 296532 48140 387800 48328
tri 229032 46127 231045 48140 ne
rect 231045 46127 234688 48140
tri 234688 46127 236701 48140 sw
tri 254032 46500 255672 48140 ne
rect 255672 46500 287188 48140
tri 287188 46500 288828 48140 sw
tri 296532 46500 298172 48140 ne
rect 298172 46500 387800 48140
tri 283172 46127 283545 46500 ne
rect 283545 46377 288828 46500
tri 288828 46377 288951 46500 sw
tri 378957 46377 381800 46500 ne
rect 283545 46127 288951 46377
tri 288951 46127 289201 46377 sw
tri 231045 45250 231922 46127 ne
rect 231922 45250 236701 46127
tri 236701 45250 237578 46127 sw
tri 283545 45250 284422 46127 ne
rect 284422 45250 289201 46127
tri 289201 45250 290078 46127 sw
rect 381800 45957 387800 46500
tri 381800 45250 382507 45957 ne
rect 382507 45250 387093 45957
tri 387093 45250 387800 45957 nw
tri 231922 43875 233297 45250 ne
rect 233297 43875 237578 45250
tri 237578 43875 238953 45250 sw
tri 284422 44984 284688 45250 ne
rect 284688 44984 290078 45250
tri 290078 44984 290344 45250 sw
tri 284688 44844 284828 44984 ne
rect 284828 44844 290344 44984
tri 284828 43875 285797 44844 ne
rect 285797 43875 290344 44844
tri 290344 43875 291453 44984 sw
tri 233297 42672 234500 43875 ne
rect 234500 42672 238953 43875
tri 238953 42672 240156 43875 sw
tri 285797 42672 287000 43875 ne
rect 287000 42672 291453 43875
tri 291453 42672 292656 43875 sw
tri 234500 42484 234688 42672 ne
rect 234688 42484 240156 42672
tri 240156 42484 240344 42672 sw
tri 287000 42484 287188 42672 ne
rect 287188 42484 292656 42672
tri 292656 42484 292844 42672 sw
tri 234688 36828 240344 42484 ne
tri 240344 36828 246000 42484 sw
tri 287188 39328 290344 42484 ne
rect 290344 39328 292844 42484
tri 292844 39328 296000 42484 sw
tri 290344 37672 292000 39328 ne
tri 240344 35172 242000 36828 ne
tri 193172 30500 195344 32672 se
rect 195344 30500 198828 32672
tri 198828 30500 201000 32672 nw
tri 75672 10500 77328 12156 se
rect 77328 10500 81328 12156
tri 81328 10500 82984 12156 nw
tri 98172 10500 99828 12156 se
tri 56703 6500 60666 10500 se
rect 60666 6500 77328 10500
tri 77328 6500 81328 10500 nw
tri 84203 6500 88166 10500 se
rect 88166 6500 99828 10500
tri 99828 6500 105484 12156 nw
tri 128172 10500 129828 12156 se
rect 129828 10500 130146 12156
tri 111703 6500 115666 10500 se
rect 115666 6818 130146 10500
tri 130146 6818 135484 12156 nw
tri 141357 8654 144841 12156 se
rect 144841 8654 147000 12156
tri 147000 8654 151000 12674 nw
tri 139530 6818 141357 8654 se
rect 141357 6818 145172 8654
tri 145172 6818 147000 8654 nw
rect 115666 6500 129828 6818
tri 129828 6500 130146 6818 nw
tri 139213 6500 139530 6818 se
rect 139530 6500 144856 6818
tri 144856 6500 145172 6818 nw
tri 166688 6500 167000 6818 se
rect 167000 6500 171000 30500
tri 56406 6200 56703 6500 se
rect 56703 6200 62037 6500
tri 62037 6200 62334 6500 nw
tri 83906 6200 84203 6500 se
rect 84203 6200 89537 6500
tri 89537 6200 89834 6500 nw
tri 111406 6200 111703 6500 se
rect 111703 6200 117037 6500
tri 117037 6200 117334 6500 nw
tri 138915 6200 139213 6500 se
rect 139213 6200 144557 6500
tri 144557 6200 144856 6500 nw
tri 166393 6200 166688 6500 se
rect 166688 6200 171000 6500
tri 192000 29328 193172 30500 se
rect 193172 29328 196000 30500
rect 192000 6200 196000 29328
tri 196000 27672 198828 30500 nw
rect 217000 6200 221000 30500
rect 242000 9038 246000 36828
rect 267000 10214 271000 30500
rect 292000 12704 296000 39328
tri 318172 30500 319000 31328 se
tri 319000 30500 319828 31328 sw
tri 316172 28500 318172 30500 se
rect 318172 28500 319828 30500
tri 316172 28140 316532 28500 ne
rect 316532 28140 319828 28500
tri 319828 28140 322188 30500 sw
tri 316532 25672 319000 28140 ne
rect 319000 25672 322188 28140
tri 319000 22484 322188 25672 ne
tri 322188 22484 327844 28140 sw
tri 322188 16828 327844 22484 ne
tri 327844 16828 333500 22484 sw
tri 327844 15172 329500 16828 ne
tri 292000 11786 292868 12704 ne
rect 292868 11786 296000 12704
tri 296000 11786 298375 14296 sw
tri 246000 9038 246203 9265 sw
rect 242000 8972 246203 9038
tri 246203 8972 246262 9038 sw
tri 267000 8972 268154 10214 ne
rect 268154 8972 271000 10214
tri 271000 8972 273615 11786 sw
tri 292868 8972 295532 11786 ne
rect 295532 8972 298375 11786
tri 298375 8972 301038 11786 sw
rect 242000 7735 246262 8972
tri 242000 6705 242923 7735 ne
rect 242923 6704 246262 7735
tri 246262 6704 248294 8972 sw
tri 268154 6704 270262 8972 ne
rect 270262 6704 273615 8972
tri 273615 6704 275723 8972 sw
tri 295532 8940 295562 8972 ne
rect 295562 8940 301038 8972
tri 301038 8940 301069 8972 sw
tri 295562 8478 296000 8940 ne
rect 296000 8478 301069 8940
tri 296000 6704 297678 8478 ne
rect 297678 6704 301069 8478
tri 301069 6704 303185 8940 sw
tri 221000 6200 221405 6704 sw
tri 242923 6200 243375 6704 ne
rect 243375 6200 248294 6704
tri 248294 6200 248746 6704 sw
tri 270262 6200 270731 6704 ne
rect 270731 6200 275723 6704
tri 275723 6200 276192 6704 sw
tri 297678 6200 298155 6704 ne
rect 298155 6200 303185 6704
tri 303185 6200 303663 6704 sw
rect 329500 6200 333500 16828
tri 53813 6056 53957 6200 se
rect 53957 6056 61894 6200
tri 61894 6056 62037 6200 nw
tri 81313 6056 81457 6200 se
rect 81457 6056 89394 6200
tri 89394 6056 89537 6200 nw
tri 108813 6056 108957 6200 se
rect 108957 6056 116894 6200
tri 116894 6056 117037 6200 nw
tri 53422 5665 53813 6056 se
rect 53813 5665 61507 6056
tri 61507 5665 61894 6056 nw
tri 80922 5665 81313 6056 se
rect 81313 5665 86750 6056
tri 53250 5493 53422 5665 se
rect 53422 5493 59250 5665
rect 53250 907 59250 5493
tri 59250 3387 61507 5665 nw
tri 80750 5493 80922 5665 se
rect 80922 5493 86750 5665
tri 53250 735 53422 907 ne
rect 53422 735 58715 907
tri 53422 372 53785 735 ne
rect 53785 372 58715 735
tri 58715 372 59250 907 nw
rect 80750 907 86750 5493
tri 86750 3387 89394 6056 nw
tri 108422 5665 108813 6056 se
rect 108813 5665 114250 6056
tri 108250 5493 108422 5665 se
rect 108422 5493 114250 5665
tri 80750 735 80922 907 ne
rect 80922 735 86215 907
tri 80922 372 81285 735 ne
rect 81285 372 86215 735
tri 86215 372 86750 907 nw
rect 108250 907 114250 5493
tri 114250 3387 116894 6056 nw
tri 135922 5665 136457 6200 se
rect 136457 5886 144245 6200
tri 144245 5886 144557 6200 nw
rect 136457 5679 144039 5886
tri 144039 5679 144245 5886 nw
rect 136457 5665 141750 5679
tri 135750 5493 135922 5665 se
rect 135922 5493 141750 5665
tri 108250 735 108422 907 ne
rect 108422 735 113715 907
tri 108422 372 108785 735 ne
rect 108785 372 113715 735
tri 113715 372 114250 907 nw
rect 135750 907 141750 5493
tri 141750 3380 144039 5679 nw
tri 163250 5493 163957 6200 se
rect 163957 5493 171000 6200
rect 163250 5182 171000 5493
tri 135750 735 135922 907 ne
rect 135922 735 141564 907
tri 135922 372 136285 735 ne
rect 136285 721 141564 735
tri 141564 721 141750 907 nw
rect 163250 907 169250 5182
tri 169250 3401 171000 5182 nw
tri 190750 5493 191457 6200 se
rect 191457 5493 196043 6200
tri 196043 5493 196750 6200 sw
tri 163250 735 163422 907 ne
rect 163422 735 168715 907
rect 136285 372 141215 721
tri 141215 372 141564 721 nw
tri 163422 372 163785 735 ne
rect 163785 372 168715 735
tri 168715 372 169250 907 nw
rect 190750 907 196750 5493
rect 217000 5681 223543 6200
tri 223543 5681 224062 6200 sw
tri 243375 5946 243603 6200 ne
rect 243603 5946 251043 6200
tri 243603 5681 243840 5946 ne
rect 243840 5681 251043 5946
rect 217000 5493 224062 5681
tri 224062 5493 224250 5681 sw
rect 217000 5296 224250 5493
tri 217000 3740 218250 5296 ne
tri 190750 724 190933 907 ne
rect 190933 724 196043 907
tri 190933 383 191274 724 ne
rect 191274 383 196043 724
tri 53785 200 53957 372 ne
rect 53957 200 58543 372
tri 58543 200 58715 372 nw
tri 81285 200 81457 372 ne
rect 81457 200 86043 372
tri 86043 200 86215 372 nw
tri 108785 200 108957 372 ne
rect 108957 200 113543 372
tri 113543 200 113715 372 nw
tri 136285 200 136457 372 ne
rect 136457 200 141043 372
tri 141043 200 141215 372 nw
tri 163785 200 163957 372 ne
rect 163957 200 168543 372
tri 168543 200 168715 372 nw
tri 191274 200 191457 383 ne
rect 191457 200 196043 383
tri 196043 200 196750 907 nw
rect 218250 907 224250 5296
tri 243840 3550 245750 5681 ne
rect 245750 5669 251043 5681
tri 251043 5669 251574 6200 sw
tri 270731 5911 271000 6200 ne
rect 271000 5911 278543 6200
tri 271000 5858 271049 5911 ne
rect 271049 5858 278543 5911
rect 245750 5493 251574 5669
tri 251574 5493 251750 5669 sw
tri 218250 388 218769 907 ne
rect 218769 719 224062 907
tri 224062 719 224250 907 nw
rect 245750 907 251750 5493
tri 271049 3489 273250 5858 ne
rect 273250 5666 278543 5858
tri 278543 5666 279077 6200 sw
tri 298155 5812 298523 6200 ne
rect 298523 5812 306043 6200
tri 298523 5666 298661 5812 ne
rect 298661 5666 306043 5812
tri 306043 5666 306577 6200 sw
rect 273250 5493 279077 5666
tri 279077 5493 279250 5666 sw
rect 218769 388 223731 719
tri 223731 388 224062 719 nw
tri 245750 454 246203 907 ne
rect 246203 731 251574 907
tri 251574 731 251750 907 nw
rect 273250 907 279250 5493
tri 298661 3459 300750 5666 ne
rect 300750 5493 306577 5666
tri 306577 5493 306750 5666 sw
rect 246203 454 251219 731
tri 218769 200 218957 388 ne
rect 218957 200 223543 388
tri 223543 200 223731 388 nw
tri 246203 376 246281 454 ne
rect 246281 376 251219 454
tri 251219 376 251574 731 nw
tri 273250 542 273615 907 ne
rect 273615 734 279077 907
tri 279077 734 279250 907 nw
rect 300750 907 306750 5493
rect 273615 542 278716 734
tri 246281 200 246457 376 ne
rect 246457 200 251043 376
tri 251043 200 251219 376 nw
tri 273615 373 273784 542 ne
rect 273784 373 278716 542
tri 278716 373 279077 734 nw
tri 300750 588 301069 907 ne
rect 301069 734 306577 907
tri 306577 734 306750 907 nw
tri 328250 5493 328957 6200 se
rect 328957 5493 333543 6200
tri 333543 5493 334250 6200 sw
rect 328250 907 334250 5493
rect 301069 588 306216 734
tri 301069 373 301284 588 ne
rect 301284 373 306216 588
tri 306216 373 306577 734 nw
tri 273784 200 273957 373 ne
rect 273957 200 278543 373
tri 278543 200 278716 373 nw
tri 301284 200 301457 373 ne
rect 301457 200 306043 373
tri 306043 200 306216 373 nw
tri 328250 200 328957 907 ne
rect 328957 200 333543 907
tri 333543 200 334250 907 nw
use bump_bond0  bump_bond0_0
timestamp 1679504633
transform -1 0 69000 0 -1 28500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_1
timestamp 1679504633
transform 0 1 169000 -1 0 28500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_2
timestamp 1679504633
transform 0 1 219000 -1 0 28500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_3
timestamp 1679504633
transform 0 1 269000 -1 0 28500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_4
timestamp 1679504633
transform -1 0 69000 0 -1 78500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_5
timestamp 1679504633
transform 0 1 219000 -1 0 78500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_6
timestamp 1679504633
transform 1 0 269000 0 1 78500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_7
timestamp 1679504633
transform 1 0 319000 0 1 78500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_8
timestamp 1679504633
transform -1 0 69000 0 -1 128500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_9
timestamp 1679504633
transform 0 1 219000 -1 0 128500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_10
timestamp 1679504633
transform 1 0 319000 0 1 128500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_11
timestamp 1679504633
transform -1 0 69000 0 -1 178500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_12
timestamp 1679504633
transform 1 0 319000 0 1 178500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_13
timestamp 1679504633
transform 1 0 169000 0 1 228500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_14
timestamp 1679504633
transform -1 0 219000 0 -1 228500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_15
timestamp 1679504633
transform 1 0 319000 0 1 228500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_16
timestamp 1679504633
transform -1 0 69000 0 -1 278500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_17
timestamp 1679504633
transform 1 0 169000 0 1 278500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_18
timestamp 1679504633
transform -1 0 219000 0 -1 278500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_19
timestamp 1679504633
transform 1 0 319000 0 1 278500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_20
timestamp 1679504633
transform -1 0 69000 0 -1 328500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_21
timestamp 1679504633
transform -1 0 169000 0 -1 328500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_22
timestamp 1679504633
transform 1 0 319000 0 1 328500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_23
timestamp 1679504633
transform -1 0 69000 0 -1 378500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_24
timestamp 1679504633
transform -1 0 119000 0 -1 378500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_25
timestamp 1679504633
transform 1 0 319000 0 1 378500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_26
timestamp 1679504633
transform -1 0 69000 0 -1 428500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_27
timestamp 1679504633
transform 0 -1 119000 1 0 478500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_28
timestamp 1679504633
transform 0 -1 169000 1 0 478500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_29
timestamp 1679504633
transform 0 -1 219000 1 0 478500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_30
timestamp 1679504633
transform 0 -1 269000 1 0 478500
box -13449 -13449 19092 13449
use bump_bond0  bump_bond0_31
timestamp 1679504633
transform -1 0 269000 0 -1 228500
box -13449 -13449 19092 13449
use bump_bond45  bump_bond45_0
timestamp 1679504633
transform -1 0 119000 0 -1 28500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_1
timestamp 1679504633
transform 0 1 319000 -1 0 28500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_2
timestamp 1679504633
transform 0 -1 119000 1 0 78500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_3
timestamp 1679504633
transform -1 0 169000 0 -1 78500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_4
timestamp 1679504633
transform 0 -1 119000 1 0 128500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_5
timestamp 1679504633
transform 0 -1 169000 1 0 128500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_6
timestamp 1679504633
transform 0 1 269000 -1 0 128500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_7
timestamp 1679504633
transform 0 -1 119000 1 0 178500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_8
timestamp 1679504633
transform 0 -1 169000 1 0 178500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_9
timestamp 1679504633
transform 0 1 219000 -1 0 178500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_10
timestamp 1679504633
transform 0 1 269000 -1 0 178500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_11
timestamp 1679504633
transform 0 -1 69000 1 0 228500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_12
timestamp 1679504633
transform 0 -1 119000 1 0 228500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_13
timestamp 1679504633
transform 0 1 269000 -1 0 228500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_14
timestamp 1679504633
transform 0 -1 119000 1 0 278500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_15
timestamp 1679504633
transform 0 1 269000 -1 0 278500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_16
timestamp 1679504633
transform 0 -1 119000 1 0 328500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_17
timestamp 1679504633
transform 0 1 219000 -1 0 328500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_18
timestamp 1679504633
transform 0 1 269000 -1 0 328500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_19
timestamp 1679504633
transform 0 -1 169000 1 0 378500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_20
timestamp 1679504633
transform 1 0 219000 0 1 378500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_21
timestamp 1679504633
transform 0 1 269000 -1 0 378500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_22
timestamp 1679504633
transform 0 -1 119000 1 0 428500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_23
timestamp 1679504633
transform 0 -1 169000 1 0 428500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_24
timestamp 1679504633
transform 1 0 219000 0 1 428500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_25
timestamp 1679504633
transform 1 0 269000 0 1 428500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_26
timestamp 1679504633
transform 1 0 319000 0 1 428500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_27
timestamp 1679504633
transform 0 -1 69000 1 0 478500
box -13500 -13500 13500 13500
use bump_bond45  bump_bond45_28
timestamp 1679504633
transform 1 0 319000 0 1 478500
box -13500 -13500 13500 13500
<< end >>
