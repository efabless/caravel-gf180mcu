magic
tech gf180mcuC
magscale 1 10
timestamp 1655304105
<< metal1 >>
rect -41 -212 -29 -160
rect 85 -212 97 -160
<< via1 >>
rect -29 -212 85 -160
<< metal2 >>
rect -43 -160 99 -158
rect -43 -212 -29 -160
rect 85 -212 99 -160
rect -43 -214 99 -212
<< end >>
