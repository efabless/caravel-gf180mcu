magic
tech gf180mcuC
magscale 1 10
timestamp 1655473121
<< obsm1 >>
rect 336 724 5696 33962
<< metal2 >>
rect 2212 33962 2268 35200
rect 2660 33124 2716 35200
rect 3108 32564 3164 35200
rect 3556 34468 3612 35200
rect 4900 34944 6100 35000
rect 5348 33488 6100 33544
rect 5460 31926 6100 31982
rect 5796 30470 6100 30526
rect 5796 28906 6100 28962
rect 5796 27450 6100 27506
rect 5796 25886 6100 25942
rect 5796 24430 6100 24486
rect 5516 22866 6100 22922
rect 5796 21410 6100 21466
rect -100 14252 100 14328
rect -100 13731 100 13807
rect -100 13502 100 13578
rect -100 13360 100 13436
rect -100 12858 100 12934
rect -100 12647 100 12723
rect -100 1190 100 1266
rect -100 1044 100 1120
rect -100 898 100 974
rect -100 752 100 828
rect 2212 -200 2268 2604
rect 2660 -200 2716 1372
rect 3108 -200 3164 3388
rect 3556 -200 3612 588
<< obsm2 >>
rect 84 33902 2152 34944
rect 2328 33902 2600 34944
rect 84 33064 2600 33902
rect 2776 33064 3048 34944
rect 84 32504 3048 33064
rect 3224 34408 3496 34944
rect 3672 34884 4840 34944
rect 3672 34408 5964 34884
rect 3224 33604 5964 34408
rect 3224 33428 5288 33604
rect 3224 32504 5964 33428
rect 84 32042 5964 32504
rect 84 31866 5400 32042
rect 84 30586 5964 31866
rect 84 30410 5736 30586
rect 84 29022 5964 30410
rect 84 28846 5736 29022
rect 84 27566 5964 28846
rect 84 27390 5736 27566
rect 84 26002 5964 27390
rect 84 25826 5736 26002
rect 84 24546 5964 25826
rect 84 24370 5736 24546
rect 84 22982 5964 24370
rect 84 22806 5456 22982
rect 84 21526 5964 22806
rect 84 21350 5736 21526
rect 84 14388 5964 21350
rect 160 14192 5964 14388
rect 84 13867 5964 14192
rect 160 13671 5964 13867
rect 84 13638 5964 13671
rect 160 13300 5964 13638
rect 84 12994 5964 13300
rect 160 12798 5964 12994
rect 84 12783 5964 12798
rect 160 12587 5964 12783
rect 84 3448 5964 12587
rect 84 2664 3048 3448
rect 84 1326 2152 2664
rect 160 692 2152 1326
rect 84 532 2152 692
rect 2328 1432 3048 2664
rect 2328 532 2600 1432
rect 2776 532 3048 1432
rect 3224 648 5964 3448
rect 3224 532 3496 648
rect 3672 532 5964 648
<< metal3 >>
rect 5068 18900 6000 18956
rect 5404 18452 6000 18508
rect 5800 18004 6000 18060
rect 3836 17556 6000 17612
rect 4844 17108 6000 17164
rect 4788 16660 6000 16716
rect 5292 16212 6000 16268
rect 4844 15764 6000 15820
<< obsm3 >>
rect 74 19016 5974 33740
rect 74 18840 5008 19016
rect 74 18568 5974 18840
rect 74 18392 5344 18568
rect 74 18120 5974 18392
rect 74 17944 5740 18120
rect 74 17672 5974 17944
rect 74 17496 3776 17672
rect 74 17224 5974 17496
rect 74 17048 4784 17224
rect 74 16776 5974 17048
rect 74 16600 4728 16776
rect 74 16328 5974 16600
rect 74 16152 5232 16328
rect 74 15880 5974 16152
rect 74 15704 4784 15880
rect 74 756 5974 15704
<< metal4 >>
rect 376 724 696 33772
rect 1376 724 1696 33772
rect 2376 724 2696 33772
rect 3376 724 3696 33772
rect 4376 724 4696 33772
rect 5376 724 5696 33772
<< obsm4 >>
rect 196 2762 316 32182
rect 756 2762 1316 32182
rect 1756 2762 2316 32182
rect 2756 2762 3316 32182
rect 3756 2762 4316 32182
rect 4756 2762 5316 32182
rect 5756 2762 5964 32182
<< metal5 >>
rect 276 32424 5696 32744
rect 276 28924 5660 29244
rect 276 25424 5696 25744
rect 276 21924 5660 22244
rect 276 18424 5696 18744
rect 276 14924 5660 15244
rect 276 11424 5696 11744
rect 276 7924 5660 8244
rect 276 4424 5696 4744
rect 276 924 5660 1244
<< labels >>
rlabel metal4 s 376 724 696 33772 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 2376 724 2696 33772 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 4376 724 4696 33772 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 276 924 5660 1244 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 276 7924 5660 8244 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 276 14924 5660 15244 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 276 21924 5660 22244 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 276 28924 5660 29244 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 1376 724 1696 33772 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 3376 724 3696 33772 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 5376 724 5696 33772 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 276 4424 5696 4744 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 276 11424 5696 11744 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 276 18424 5696 18744 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 276 25424 5696 25744 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 276 32424 5696 32744 6 VSS
port 2 nsew ground bidirectional
rlabel metal2 s 4900 34944 6100 35000 6 gpio_defaults[0]
port 3 nsew signal input
rlabel metal2 s 5348 33488 6100 33544 6 gpio_defaults[1]
port 4 nsew signal input
rlabel metal2 s 5460 31926 6100 31982 6 gpio_defaults[2]
port 5 nsew signal input
rlabel metal2 s 5796 30470 6100 30526 6 gpio_defaults[3]
port 6 nsew signal input
rlabel metal2 s 5796 28906 6100 28962 6 gpio_defaults[4]
port 7 nsew signal input
rlabel metal2 s 5796 27450 6100 27506 6 gpio_defaults[5]
port 8 nsew signal input
rlabel metal2 s 5796 25886 6100 25942 6 gpio_defaults[6]
port 9 nsew signal input
rlabel metal2 s 5796 24430 6100 24486 6 gpio_defaults[7]
port 10 nsew signal input
rlabel metal2 s 5516 22866 6100 22922 6 gpio_defaults[8]
port 11 nsew signal input
rlabel metal2 s 5796 21410 6100 21466 6 gpio_defaults[9]
port 12 nsew signal input
rlabel metal3 s 4844 15764 6000 15820 6 mgmt_gpio_in
port 13 nsew signal output
rlabel metal3 s 3836 17556 6000 17612 6 mgmt_gpio_oeb
port 14 nsew signal input
rlabel metal3 s 5404 18452 6000 18508 6 mgmt_gpio_out
port 15 nsew signal input
rlabel metal3 s 4788 16660 6000 16716 6 one
port 16 nsew signal output
rlabel metal2 s -100 13502 100 13578 4 pad_gpio_drive_sel[0]
port 17 nsew signal output
rlabel metal2 s -100 13360 100 13436 4 pad_gpio_drive_sel[1]
port 18 nsew signal output
rlabel metal2 s -100 752 100 828 4 pad_gpio_in
port 19 nsew signal input
rlabel metal2 s -100 12647 100 12723 4 pad_gpio_inen
port 20 nsew signal output
rlabel metal2 s -100 1044 100 1120 4 pad_gpio_out
port 21 nsew signal output
rlabel metal2 s -100 898 100 974 4 pad_gpio_outen
port 22 nsew signal output
rlabel metal2 s -100 12858 100 12934 4 pad_gpio_pulldown_sel
port 23 nsew signal output
rlabel metal2 s -100 13731 100 13807 4 pad_gpio_pullup_sel
port 24 nsew signal output
rlabel metal2 s -100 14252 100 14328 4 pad_gpio_schmitt_sel
port 25 nsew signal output
rlabel metal2 s -100 1190 100 1266 4 pad_gpio_slew_sel
port 26 nsew signal output
rlabel metal2 s 2212 33962 2268 35200 6 resetn
port 27 nsew signal input
rlabel metal2 s 2212 -200 2268 2604 6 resetn_out
port 28 nsew signal output
rlabel metal2 s 3108 32564 3164 35200 6 serial_clock
port 29 nsew signal input
rlabel metal2 s 3108 -200 3164 3388 6 serial_clock_out
port 30 nsew signal output
rlabel metal2 s 3556 34468 3612 35200 6 serial_data_in
port 31 nsew signal input
rlabel metal2 s 2660 -200 2716 1372 6 serial_data_out
port 32 nsew signal output
rlabel metal2 s 2660 33124 2716 35200 6 serial_load
port 33 nsew signal input
rlabel metal2 s 3556 -200 3612 588 6 serial_load_out
port 34 nsew signal output
rlabel metal3 s 5292 16212 6000 16268 6 user_gpio_in
port 35 nsew signal output
rlabel metal3 s 5800 18004 6000 18060 6 user_gpio_oeb
port 36 nsew signal input
rlabel metal3 s 5068 18900 6000 18956 6 user_gpio_out
port 37 nsew signal input
rlabel metal3 s 4844 17108 6000 17164 6 zero
port 38 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 6000 35000
string GDS_END 346608
string GDS_FILE ../gds/gpio_control_block.gds.gz
string GDS_START 79228
string LEFclass BLOCK
string LEFview TRUE
<< end >>
