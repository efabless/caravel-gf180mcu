magic
tech gf180mcuD
magscale 1 10
timestamp 1655307388
<< error_p >>
rect -58 -655 -47 -609
<< nwell >>
rect -378 -886 368 886
<< mvpmos >>
rect -60 -576 50 624
<< mvpdiff >>
rect -148 611 -60 624
rect -148 -563 -135 611
rect -89 -563 -60 611
rect -148 -576 -60 -563
rect 50 611 138 624
rect 50 -563 79 611
rect 125 -563 138 611
rect 50 -576 138 -563
<< mvpdiffc >>
rect -135 -563 -89 611
rect 79 -563 125 611
<< mvnsubdiff >>
rect -292 787 282 800
rect -292 741 -176 787
rect 166 741 282 787
rect -292 728 282 741
rect -292 684 -220 728
rect -292 -684 -279 684
rect -233 -684 -220 684
rect 210 684 282 728
rect -292 -728 -220 -684
rect 210 -684 223 684
rect 269 -684 282 684
rect 210 -728 282 -684
rect -292 -800 282 -728
<< mvnsubdiffcont >>
rect -176 741 166 787
rect -279 -684 -233 684
rect 223 -684 269 684
<< polysilicon >>
rect -60 624 50 668
rect -60 -609 50 -576
rect -60 -655 -47 -609
rect 37 -655 50 -609
rect -60 -668 50 -655
<< polycontact >>
rect -47 -655 37 -609
<< metal1 >>
rect -279 741 -176 787
rect 166 741 269 787
rect -279 684 -233 741
rect 223 684 269 741
rect -135 611 -89 622
rect -135 -574 -89 -563
rect 79 611 125 622
rect 79 -574 125 -563
rect -58 -655 -47 -609
rect 37 -655 48 -609
rect -279 -741 -233 -684
rect 223 -741 269 -684
rect -279 -787 269 -741
<< properties >>
string FIXED_BBOX -246 -764 246 764
string gencell pmos_6p0
string library gf180mcu
string parameters w 6.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.5 wmin 0.3 full_metal 1 compatible {pmos_3p3 pmos_6p0}
<< end >>
