magic
tech micross
timestamp 1679504633
<< rdl >>
tri -2344 13295 0 13500 se
rect 0 13295 13500 13500
tri -4617 12686 -2344 13295 se
rect -2344 12686 13500 13295
tri -6750 11691 -4617 12686 se
rect -4617 11691 13500 12686
tri -8678 10342 -6750 11691 se
rect -6750 10342 13500 11691
tri -10342 8678 -8678 10342 se
rect -8678 8678 13500 10342
tri -11691 6750 -10342 8678 se
rect -10342 6750 13500 8678
tri -12686 4617 -11691 6750 se
rect -11691 4617 13500 6750
tri -13295 2344 -12686 4617 se
rect -12686 2344 13500 4617
tri -13500 0 -13295 2344 se
rect -13295 0 13500 2344
tri -13500 -2344 -13295 0 ne
rect -13295 -2344 13295 0
tri 13295 -2344 13500 0 nw
tri -13295 -4617 -12686 -2344 ne
rect -12686 -4617 12686 -2344
tri 12686 -4617 13295 -2344 nw
tri -12686 -6750 -11691 -4617 ne
rect -11691 -6750 11691 -4617
tri 11691 -6750 12686 -4617 nw
tri -11691 -8678 -10342 -6750 ne
rect -10342 -8678 10342 -6750
tri 10342 -8678 11691 -6750 nw
tri -10342 -10342 -8678 -8678 ne
rect -8678 -10342 8678 -8678
tri 8678 -10342 10342 -8678 nw
tri -8678 -11691 -6750 -10342 ne
rect -6750 -11691 6750 -10342
tri 6750 -11691 8678 -10342 nw
tri -6750 -12686 -4617 -11691 ne
rect -4617 -12686 4617 -11691
tri 4617 -12686 6750 -11691 nw
tri -4617 -13295 -2344 -12686 ne
rect -2344 -13295 2344 -12686
tri 2344 -13295 4617 -12686 nw
tri -2344 -13500 0 -13295 ne
tri 0 -13500 2344 -13295 nw
<< pi2 >>
tri -1910 10833 0 11000 se
tri 0 10833 1910 11000 sw
tri -3762 10337 -1910 10833 se
rect -1910 10337 1910 10833
tri 1910 10337 3762 10833 sw
tri -5500 9526 -3762 10337 se
rect -3762 9526 3762 10337
tri 3762 9526 5500 10337 sw
tri -7071 8426 -5500 9526 se
rect -5500 8426 5500 9526
tri 5500 8426 7071 9526 sw
tri -8426 7071 -7071 8426 se
rect -7071 7071 7071 8426
tri 7071 7071 8426 8426 sw
tri -9526 5500 -8426 7071 se
rect -8426 5500 8426 7071
tri 8426 5500 9526 7071 sw
tri -10337 3762 -9526 5500 se
rect -9526 3762 9526 5500
tri 9526 3762 10337 5500 sw
tri -10833 1910 -10337 3762 se
rect -10337 1910 10337 3762
tri 10337 1910 10833 3762 sw
tri -11000 0 -10833 1910 se
tri -11000 -1910 -10833 0 ne
rect -10833 -1910 10833 1910
tri 10833 0 11000 1910 sw
tri 10833 -1910 11000 0 nw
tri -10833 -3762 -10337 -1910 ne
rect -10337 -3762 10337 -1910
tri 10337 -3762 10833 -1910 nw
tri -10337 -5500 -9526 -3762 ne
rect -9526 -5500 9526 -3762
tri 9526 -5500 10337 -3762 nw
tri -9526 -7071 -8426 -5500 ne
rect -8426 -7071 8426 -5500
tri 8426 -7071 9526 -5500 nw
tri -8426 -8426 -7071 -7071 ne
rect -7071 -8426 7071 -7071
tri 7071 -8426 8426 -7071 nw
tri -7071 -9526 -5500 -8426 ne
rect -5500 -9526 5500 -8426
tri 5500 -9526 7071 -8426 nw
tri -5500 -10337 -3762 -9526 ne
rect -3762 -10337 3762 -9526
tri 3762 -10337 5500 -9526 nw
tri -3762 -10833 -1910 -10337 ne
rect -1910 -10833 1910 -10337
tri 1910 -10833 3762 -10337 nw
tri -1910 -11000 0 -10833 ne
tri 0 -11000 1910 -10833 nw
<< ubm >>
tri -2171 12310 0 12500 se
tri 0 12310 2171 12500 sw
tri -4275 11746 -2171 12310 se
rect -2171 11746 2171 12310
tri 2171 11746 4275 12310 sw
tri -6250 10825 -4275 11746 se
rect -4275 10825 4275 11746
tri 4275 10825 6250 11746 sw
tri -8035 9576 -6250 10825 se
rect -6250 9576 6250 10825
tri 6250 9576 8035 10825 sw
tri -9576 8035 -8035 9576 se
rect -8035 8035 8035 9576
tri 8035 8035 9576 9576 sw
tri -10825 6250 -9576 8035 se
rect -9576 6250 9576 8035
tri 9576 6250 10825 8035 sw
tri -11746 4275 -10825 6250 se
rect -10825 4275 10825 6250
tri 10825 4275 11746 6250 sw
tri -12310 2171 -11746 4275 se
rect -11746 2171 11746 4275
tri 11746 2171 12310 4275 sw
tri -12500 0 -12310 2171 se
tri -12500 -2171 -12310 0 ne
rect -12310 -2171 12310 2171
tri 12310 0 12500 2171 sw
tri 12310 -2171 12500 0 nw
tri -12310 -4275 -11746 -2171 ne
rect -11746 -4275 11746 -2171
tri 11746 -4275 12310 -2171 nw
tri -11746 -6250 -10825 -4275 ne
rect -10825 -6250 10825 -4275
tri 10825 -6250 11746 -4275 nw
tri -10825 -8035 -9576 -6250 ne
rect -9576 -8035 9576 -6250
tri 9576 -8035 10825 -6250 nw
tri -9576 -9576 -8035 -8035 ne
rect -8035 -9576 8035 -8035
tri 8035 -9576 9576 -8035 nw
tri -8035 -10825 -6250 -9576 ne
rect -6250 -10825 6250 -9576
tri 6250 -10825 8035 -9576 nw
tri -6250 -11746 -4275 -10825 ne
rect -4275 -11746 4275 -10825
tri 4275 -11746 6250 -10825 nw
tri -4275 -12310 -2171 -11746 ne
rect -2171 -12310 2171 -11746
tri 2171 -12310 4275 -11746 nw
tri -2171 -12500 0 -12310 ne
tri 0 -12500 2171 -12310 nw
<< properties >>
string FIXED_BBOX -13500 -13500 13500 13500
<< end >>
