magic
tech gf180mcuD
magscale 6 5
timestamp 1654634570
<< metal5 >>
rect 0 648 324 756
rect 0 540 108 648
rect 0 432 324 540
rect 0 108 108 432
rect 216 108 324 432
rect 0 0 324 108
<< properties >>
string FIXED_BBOX 0 0 432 756
<< end >>
