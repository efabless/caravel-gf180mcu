magic
tech gf180mcuD
magscale 1 10
timestamp 1655304105
<< metal1 >>
rect 265 1350 1460 1650
rect 266 392 466 540
rect 602 496 765 1350
rect 979 1273 1031 1290
rect 979 687 1031 699
rect 811 622 1045 627
rect 811 570 824 622
rect 1028 570 1045 622
rect 811 567 1045 570
rect 1258 393 1458 538
rect 266 340 545 392
rect 749 340 761 392
rect 1023 341 1035 393
rect 1239 341 1458 393
rect 1258 338 1458 341
rect 529 -1050 692 253
rect 750 154 1051 160
rect 750 102 808 154
rect 1012 102 1051 154
rect 750 99 1051 102
rect 874 -158 926 -146
rect 874 -745 926 -732
rect 1110 -1050 1273 257
rect 265 -1350 1460 -1050
<< via1 >>
rect 979 699 1031 1273
rect 824 570 1028 622
rect 545 340 749 392
rect 1035 341 1239 393
rect 808 102 1012 154
rect 874 -732 926 -158
<< metal2 >>
rect 977 1273 1033 1292
rect 977 699 979 1273
rect 1031 740 1033 1273
rect 1031 699 1162 740
rect 977 683 1162 699
rect 807 622 1045 624
rect 807 570 824 622
rect 1028 570 1045 622
rect 807 568 1045 570
rect 856 394 962 568
rect 1105 396 1162 683
rect 533 392 962 394
rect 533 340 545 392
rect 749 340 962 392
rect 533 338 962 340
rect 1021 393 1254 396
rect 1021 341 1035 393
rect 1239 341 1254 393
rect 1021 338 1254 341
rect 856 156 962 338
rect 796 154 1024 156
rect 796 102 808 154
rect 1012 102 1024 154
rect 796 100 1024 102
rect 1105 29 1162 338
rect 871 -28 1162 29
rect 871 -156 928 -28
rect 872 -158 928 -156
rect 872 -732 874 -158
rect 926 -732 928 -158
rect 872 -747 928 -732
use pmos_6p0_MUW2NR  XM0 primitives
timestamp 1655304105
transform 1 0 900 0 1 -424
box -480 -786 480 786
use nmos_6p0_BUMBJU  XM1 primitives
timestamp 1655304105
transform 1 0 880 0 1 962
box -334 -532 334 532
<< labels >>
flabel metal1 1258 338 1458 538 0 FreeSans 1280 0 0 0 Vout
port 3 nsew
flabel metal1 266 340 466 540 0 FreeSans 1280 0 0 0 Vin
port 2 nsew
flabel metal1 780 1419 980 1619 0 FreeSans 1280 0 0 0 VSS
port 1 nsew
flabel metal1 758 -1302 958 -1102 0 FreeSans 1280 0 0 0 VDD
port 0 nsew
<< end >>
