magic
tech gf180mcuC
magscale 1 10
timestamp 1670265380
<< obsm1 >>
rect 1120 1508 14878 11820
<< metal2 >>
rect 0 13200 112 14000
rect 1344 13200 1456 14000
rect 2688 13200 2800 14000
rect 4032 13200 4144 14000
rect 5376 13200 5488 14000
rect 6720 13200 6832 14000
rect 8064 13200 8176 14000
rect 9408 13200 9520 14000
rect 10752 13200 10864 14000
rect 12096 13200 12208 14000
rect 13440 13200 13552 14000
rect 14784 13200 14896 14000
rect 0 0 112 800
rect 1344 0 1456 800
rect 2688 0 2800 800
rect 4032 0 4144 800
rect 5376 0 5488 800
rect 6720 0 6832 800
rect 8064 0 8176 800
rect 9408 0 9520 800
rect 10752 0 10864 800
rect 12096 0 12208 800
rect 13440 0 13552 800
rect 14784 0 14896 800
<< obsm2 >>
rect 172 13140 1284 13300
rect 1516 13140 2628 13300
rect 2860 13140 3972 13300
rect 4204 13140 5316 13300
rect 5548 13140 6660 13300
rect 6892 13140 8004 13300
rect 8236 13140 9348 13300
rect 9580 13140 10692 13300
rect 10924 13140 12036 13300
rect 12268 13140 13380 13300
rect 13612 13140 14724 13300
rect 28 860 14868 13140
rect 172 690 1284 860
rect 1516 690 2628 860
rect 2860 690 3972 860
rect 4204 690 5316 860
rect 5548 690 6660 860
rect 6892 690 8004 860
rect 8236 690 9348 860
rect 9580 690 10692 860
rect 10924 690 12036 860
rect 12268 690 13380 860
rect 13612 690 14724 860
<< metal3 >>
rect 0 12768 800 12880
rect 14200 12768 15000 12880
rect 0 11424 800 11536
rect 14200 11424 15000 11536
rect 0 10080 800 10192
rect 14200 10080 15000 10192
rect 0 8736 800 8848
rect 14200 8736 15000 8848
rect 0 7392 800 7504
rect 14200 7392 15000 7504
rect 0 6048 800 6160
rect 14200 6048 15000 6160
rect 0 4704 800 4816
rect 14200 4704 15000 4816
rect 0 3360 800 3472
rect 14200 3360 15000 3472
rect 0 2016 800 2128
rect 14200 2016 15000 2128
rect 0 672 800 784
rect 14200 672 15000 784
<< obsm3 >>
rect 860 12708 14140 12852
rect 18 11596 14206 12708
rect 860 11364 14140 11596
rect 18 10252 14206 11364
rect 860 10020 14140 10252
rect 18 8908 14206 10020
rect 860 8676 14140 8908
rect 18 7564 14206 8676
rect 860 7332 14140 7564
rect 18 6220 14206 7332
rect 860 5988 14140 6220
rect 18 4876 14206 5988
rect 860 4644 14140 4876
rect 18 3532 14206 4644
rect 860 3300 14140 3532
rect 18 2188 14206 3300
rect 860 1956 14140 2188
rect 18 844 14206 1956
rect 860 700 14140 844
<< metal4 >>
rect 4224 1508 4544 11820
rect 5819 1508 6139 11820
rect 7414 1508 7734 11820
rect 9009 1508 9329 11820
rect 10604 1508 10924 11820
rect 12199 1508 12519 11820
<< metal5 >>
rect 1060 6096 13836 6416
rect 1060 4738 13836 5058
<< labels >>
rlabel metal4 s 4224 1508 4544 11820 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 7414 1508 7734 11820 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 10604 1508 10924 11820 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 1060 4738 13836 5058 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 5819 1508 6139 11820 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 9009 1508 9329 11820 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 12199 1508 12519 11820 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 1060 6096 13836 6416 6 VSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 4704 800 4816 6 spare_xfq[0]
port 3 nsew signal output
rlabel metal2 s 13440 0 13552 800 6 spare_xfq[1]
port 4 nsew signal output
rlabel metal2 s 6720 13200 6832 14000 6 spare_xi[0]
port 5 nsew signal output
rlabel metal2 s 5376 0 5488 800 6 spare_xi[1]
port 6 nsew signal output
rlabel metal3 s 14200 2016 15000 2128 6 spare_xi[2]
port 7 nsew signal output
rlabel metal3 s 0 10080 800 10192 6 spare_xi[3]
port 8 nsew signal output
rlabel metal3 s 14200 672 15000 784 6 spare_xib
port 9 nsew signal output
rlabel metal2 s 14784 0 14896 800 6 spare_xmx[0]
port 10 nsew signal output
rlabel metal3 s 14200 10080 15000 10192 6 spare_xmx[1]
port 11 nsew signal output
rlabel metal2 s 0 13200 112 14000 6 spare_xna[0]
port 12 nsew signal output
rlabel metal2 s 8064 0 8176 800 6 spare_xna[1]
port 13 nsew signal output
rlabel metal3 s 0 3360 800 3472 6 spare_xno[0]
port 14 nsew signal output
rlabel metal2 s 10752 0 10864 800 6 spare_xno[1]
port 15 nsew signal output
rlabel metal3 s 14200 11424 15000 11536 6 spare_xz[0]
port 16 nsew signal output
rlabel metal3 s 0 7392 800 7504 6 spare_xz[10]
port 17 nsew signal output
rlabel metal2 s 2688 0 2800 800 6 spare_xz[11]
port 18 nsew signal output
rlabel metal2 s 13440 13200 13552 14000 6 spare_xz[12]
port 19 nsew signal output
rlabel metal2 s 9408 13200 9520 14000 6 spare_xz[13]
port 20 nsew signal output
rlabel metal3 s 14200 7392 15000 7504 6 spare_xz[14]
port 21 nsew signal output
rlabel metal2 s 12096 13200 12208 14000 6 spare_xz[15]
port 22 nsew signal output
rlabel metal3 s 0 2016 800 2128 6 spare_xz[16]
port 23 nsew signal output
rlabel metal3 s 14200 12768 15000 12880 6 spare_xz[17]
port 24 nsew signal output
rlabel metal2 s 2688 13200 2800 14000 6 spare_xz[18]
port 25 nsew signal output
rlabel metal2 s 0 0 112 800 6 spare_xz[19]
port 26 nsew signal output
rlabel metal2 s 8064 13200 8176 14000 6 spare_xz[1]
port 27 nsew signal output
rlabel metal3 s 14200 8736 15000 8848 6 spare_xz[20]
port 28 nsew signal output
rlabel metal2 s 1344 13200 1456 14000 6 spare_xz[21]
port 29 nsew signal output
rlabel metal3 s 0 672 800 784 6 spare_xz[22]
port 30 nsew signal output
rlabel metal2 s 12096 0 12208 800 6 spare_xz[23]
port 31 nsew signal output
rlabel metal2 s 10752 13200 10864 14000 6 spare_xz[24]
port 32 nsew signal output
rlabel metal3 s 14200 3360 15000 3472 6 spare_xz[25]
port 33 nsew signal output
rlabel metal2 s 1344 0 1456 800 6 spare_xz[26]
port 34 nsew signal output
rlabel metal2 s 4032 0 4144 800 6 spare_xz[27]
port 35 nsew signal output
rlabel metal3 s 0 11424 800 11536 6 spare_xz[28]
port 36 nsew signal output
rlabel metal3 s 14200 4704 15000 4816 6 spare_xz[29]
port 37 nsew signal output
rlabel metal2 s 6720 0 6832 800 6 spare_xz[2]
port 38 nsew signal output
rlabel metal3 s 0 8736 800 8848 6 spare_xz[30]
port 39 nsew signal output
rlabel metal2 s 14784 13200 14896 14000 6 spare_xz[3]
port 40 nsew signal output
rlabel metal2 s 4032 13200 4144 14000 6 spare_xz[4]
port 41 nsew signal output
rlabel metal2 s 5376 13200 5488 14000 6 spare_xz[5]
port 42 nsew signal output
rlabel metal2 s 9408 0 9520 800 6 spare_xz[6]
port 43 nsew signal output
rlabel metal3 s 0 6048 800 6160 6 spare_xz[7]
port 44 nsew signal output
rlabel metal3 s 0 12768 800 12880 6 spare_xz[8]
port 45 nsew signal output
rlabel metal3 s 14200 6048 15000 6160 6 spare_xz[9]
port 46 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 15000 14000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 190582
string GDS_FILE /home/hosni/GF180/PnR_2/caravel-gf180mcu/openlane/spare_logic_block/runs/RUN_2022.12.05_18.35.53/results/signoff/spare_logic_block.magic.gds
string GDS_START 83874
<< end >>

