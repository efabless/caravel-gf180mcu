VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO housekeeping
  CLASS BLOCK ;
  FOREIGN housekeeping ;
  ORIGIN 0.000 0.000 ;
  SIZE 620.000 BY 780.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT -0.880 8.080 0.720 768.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.880 8.080 620.800 9.680 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.880 766.480 620.800 768.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 619.200 8.080 620.800 768.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 22.240 4.780 23.840 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.040 4.780 100.640 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 4.780 177.440 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 4.780 254.240 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 4.780 331.040 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 4.780 407.840 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 4.780 484.640 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 4.780 561.440 771.380 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 21.290 624.100 22.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 81.290 624.100 82.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 141.290 624.100 142.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 201.290 624.100 202.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 261.290 624.100 262.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 321.290 624.100 322.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 381.290 624.100 382.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 441.290 624.100 442.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 501.290 624.100 502.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 561.290 624.100 562.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 621.290 624.100 622.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 681.290 624.100 682.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 741.290 624.100 742.890 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT -4.180 4.780 -2.580 771.380 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 4.780 624.100 6.380 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 769.780 624.100 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 622.500 4.780 624.100 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 25.540 4.780 27.140 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 102.340 4.780 103.940 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 179.140 4.780 180.740 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 255.940 4.780 257.540 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 332.740 4.780 334.340 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 409.540 4.780 411.140 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 486.340 4.780 487.940 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 563.140 4.780 564.740 771.380 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 51.290 624.100 52.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 111.290 624.100 112.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 171.290 624.100 172.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 231.290 624.100 232.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 291.290 624.100 292.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 351.290 624.100 352.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 411.290 624.100 412.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 471.290 624.100 472.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 531.290 624.100 532.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 591.290 624.100 592.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 651.290 624.100 652.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 711.290 624.100 712.890 ;
    END
  END VSS
  PIN debug_in
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 22.960 4.000 23.520 ;
    END
  END debug_in
  PIN debug_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 29.120 4.000 29.680 ;
    END
  END debug_mode
  PIN debug_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 35.280 4.000 35.840 ;
    END
  END debug_oeb
  PIN debug_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 41.440 4.000 42.000 ;
    END
  END debug_out
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.760 4.000 54.320 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.920 4.000 60.480 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 66.080 4.000 66.640 ;
    END
  END irq[2]
  PIN mask_rev_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 393.680 0.000 394.240 4.000 ;
    END
  END mask_rev_in[0]
  PIN mask_rev_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 460.880 0.000 461.440 4.000 ;
    END
  END mask_rev_in[10]
  PIN mask_rev_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 467.600 0.000 468.160 4.000 ;
    END
  END mask_rev_in[11]
  PIN mask_rev_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 474.320 0.000 474.880 4.000 ;
    END
  END mask_rev_in[12]
  PIN mask_rev_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 481.040 0.000 481.600 4.000 ;
    END
  END mask_rev_in[13]
  PIN mask_rev_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 487.760 0.000 488.320 4.000 ;
    END
  END mask_rev_in[14]
  PIN mask_rev_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 494.480 0.000 495.040 4.000 ;
    END
  END mask_rev_in[15]
  PIN mask_rev_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 501.200 0.000 501.760 4.000 ;
    END
  END mask_rev_in[16]
  PIN mask_rev_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 507.920 0.000 508.480 4.000 ;
    END
  END mask_rev_in[17]
  PIN mask_rev_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 514.640 0.000 515.200 4.000 ;
    END
  END mask_rev_in[18]
  PIN mask_rev_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 521.360 0.000 521.920 4.000 ;
    END
  END mask_rev_in[19]
  PIN mask_rev_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 400.400 0.000 400.960 4.000 ;
    END
  END mask_rev_in[1]
  PIN mask_rev_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 528.080 0.000 528.640 4.000 ;
    END
  END mask_rev_in[20]
  PIN mask_rev_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 534.800 0.000 535.360 4.000 ;
    END
  END mask_rev_in[21]
  PIN mask_rev_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 541.520 0.000 542.080 4.000 ;
    END
  END mask_rev_in[22]
  PIN mask_rev_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 548.240 0.000 548.800 4.000 ;
    END
  END mask_rev_in[23]
  PIN mask_rev_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 554.960 0.000 555.520 4.000 ;
    END
  END mask_rev_in[24]
  PIN mask_rev_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 561.680 0.000 562.240 4.000 ;
    END
  END mask_rev_in[25]
  PIN mask_rev_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 568.400 0.000 568.960 4.000 ;
    END
  END mask_rev_in[26]
  PIN mask_rev_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 575.120 0.000 575.680 4.000 ;
    END
  END mask_rev_in[27]
  PIN mask_rev_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 581.840 0.000 582.400 4.000 ;
    END
  END mask_rev_in[28]
  PIN mask_rev_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 588.560 0.000 589.120 4.000 ;
    END
  END mask_rev_in[29]
  PIN mask_rev_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 407.120 0.000 407.680 4.000 ;
    END
  END mask_rev_in[2]
  PIN mask_rev_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 595.280 0.000 595.840 4.000 ;
    END
  END mask_rev_in[30]
  PIN mask_rev_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 602.000 0.000 602.560 4.000 ;
    END
  END mask_rev_in[31]
  PIN mask_rev_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.840 0.000 414.400 4.000 ;
    END
  END mask_rev_in[3]
  PIN mask_rev_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 420.560 0.000 421.120 4.000 ;
    END
  END mask_rev_in[4]
  PIN mask_rev_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 427.280 0.000 427.840 4.000 ;
    END
  END mask_rev_in[5]
  PIN mask_rev_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 434.000 0.000 434.560 4.000 ;
    END
  END mask_rev_in[6]
  PIN mask_rev_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 440.720 0.000 441.280 4.000 ;
    END
  END mask_rev_in[7]
  PIN mask_rev_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 447.440 0.000 448.000 4.000 ;
    END
  END mask_rev_in[8]
  PIN mask_rev_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 454.160 0.000 454.720 4.000 ;
    END
  END mask_rev_in[9]
  PIN mgmt_gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 72.240 620.000 72.800 ;
    END
  END mgmt_gpio_in[0]
  PIN mgmt_gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 425.040 620.000 425.600 ;
    END
  END mgmt_gpio_in[10]
  PIN mgmt_gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 460.320 620.000 460.880 ;
    END
  END mgmt_gpio_in[11]
  PIN mgmt_gpio_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 495.600 620.000 496.160 ;
    END
  END mgmt_gpio_in[12]
  PIN mgmt_gpio_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 530.880 620.000 531.440 ;
    END
  END mgmt_gpio_in[13]
  PIN mgmt_gpio_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 566.160 620.000 566.720 ;
    END
  END mgmt_gpio_in[14]
  PIN mgmt_gpio_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 601.440 620.000 602.000 ;
    END
  END mgmt_gpio_in[15]
  PIN mgmt_gpio_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 636.720 620.000 637.280 ;
    END
  END mgmt_gpio_in[16]
  PIN mgmt_gpio_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 672.000 620.000 672.560 ;
    END
  END mgmt_gpio_in[17]
  PIN mgmt_gpio_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 707.280 620.000 707.840 ;
    END
  END mgmt_gpio_in[18]
  PIN mgmt_gpio_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 742.560 620.000 743.120 ;
    END
  END mgmt_gpio_in[19]
  PIN mgmt_gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 107.520 620.000 108.080 ;
    END
  END mgmt_gpio_in[1]
  PIN mgmt_gpio_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 429.520 4.000 430.080 ;
    END
  END mgmt_gpio_in[20]
  PIN mgmt_gpio_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 448.000 4.000 448.560 ;
    END
  END mgmt_gpio_in[21]
  PIN mgmt_gpio_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 466.480 4.000 467.040 ;
    END
  END mgmt_gpio_in[22]
  PIN mgmt_gpio_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 484.960 4.000 485.520 ;
    END
  END mgmt_gpio_in[23]
  PIN mgmt_gpio_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 503.440 4.000 504.000 ;
    END
  END mgmt_gpio_in[24]
  PIN mgmt_gpio_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 521.920 4.000 522.480 ;
    END
  END mgmt_gpio_in[25]
  PIN mgmt_gpio_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 540.400 4.000 540.960 ;
    END
  END mgmt_gpio_in[26]
  PIN mgmt_gpio_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 558.880 4.000 559.440 ;
    END
  END mgmt_gpio_in[27]
  PIN mgmt_gpio_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 577.360 4.000 577.920 ;
    END
  END mgmt_gpio_in[28]
  PIN mgmt_gpio_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 595.840 4.000 596.400 ;
    END
  END mgmt_gpio_in[29]
  PIN mgmt_gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 142.800 620.000 143.360 ;
    END
  END mgmt_gpio_in[2]
  PIN mgmt_gpio_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 614.320 4.000 614.880 ;
    END
  END mgmt_gpio_in[30]
  PIN mgmt_gpio_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 632.800 4.000 633.360 ;
    END
  END mgmt_gpio_in[31]
  PIN mgmt_gpio_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 651.280 4.000 651.840 ;
    END
  END mgmt_gpio_in[32]
  PIN mgmt_gpio_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 669.760 4.000 670.320 ;
    END
  END mgmt_gpio_in[33]
  PIN mgmt_gpio_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 688.240 4.000 688.800 ;
    END
  END mgmt_gpio_in[34]
  PIN mgmt_gpio_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 706.720 4.000 707.280 ;
    END
  END mgmt_gpio_in[35]
  PIN mgmt_gpio_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 725.200 4.000 725.760 ;
    END
  END mgmt_gpio_in[36]
  PIN mgmt_gpio_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 743.680 4.000 744.240 ;
    END
  END mgmt_gpio_in[37]
  PIN mgmt_gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 178.080 620.000 178.640 ;
    END
  END mgmt_gpio_in[3]
  PIN mgmt_gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 213.360 620.000 213.920 ;
    END
  END mgmt_gpio_in[4]
  PIN mgmt_gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 248.640 620.000 249.200 ;
    END
  END mgmt_gpio_in[5]
  PIN mgmt_gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 283.920 620.000 284.480 ;
    END
  END mgmt_gpio_in[6]
  PIN mgmt_gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 319.200 620.000 319.760 ;
    END
  END mgmt_gpio_in[7]
  PIN mgmt_gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 354.480 620.000 355.040 ;
    END
  END mgmt_gpio_in[8]
  PIN mgmt_gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 389.760 620.000 390.320 ;
    END
  END mgmt_gpio_in[9]
  PIN mgmt_gpio_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 84.000 620.000 84.560 ;
    END
  END mgmt_gpio_oeb[0]
  PIN mgmt_gpio_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 436.800 620.000 437.360 ;
    END
  END mgmt_gpio_oeb[10]
  PIN mgmt_gpio_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 472.080 620.000 472.640 ;
    END
  END mgmt_gpio_oeb[11]
  PIN mgmt_gpio_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 507.360 620.000 507.920 ;
    END
  END mgmt_gpio_oeb[12]
  PIN mgmt_gpio_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 542.640 620.000 543.200 ;
    END
  END mgmt_gpio_oeb[13]
  PIN mgmt_gpio_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 577.920 620.000 578.480 ;
    END
  END mgmt_gpio_oeb[14]
  PIN mgmt_gpio_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 613.200 620.000 613.760 ;
    END
  END mgmt_gpio_oeb[15]
  PIN mgmt_gpio_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 648.480 620.000 649.040 ;
    END
  END mgmt_gpio_oeb[16]
  PIN mgmt_gpio_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 683.760 620.000 684.320 ;
    END
  END mgmt_gpio_oeb[17]
  PIN mgmt_gpio_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 719.040 620.000 719.600 ;
    END
  END mgmt_gpio_oeb[18]
  PIN mgmt_gpio_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 754.320 620.000 754.880 ;
    END
  END mgmt_gpio_oeb[19]
  PIN mgmt_gpio_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 119.280 620.000 119.840 ;
    END
  END mgmt_gpio_oeb[1]
  PIN mgmt_gpio_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 435.680 4.000 436.240 ;
    END
  END mgmt_gpio_oeb[20]
  PIN mgmt_gpio_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 454.160 4.000 454.720 ;
    END
  END mgmt_gpio_oeb[21]
  PIN mgmt_gpio_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 472.640 4.000 473.200 ;
    END
  END mgmt_gpio_oeb[22]
  PIN mgmt_gpio_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 491.120 4.000 491.680 ;
    END
  END mgmt_gpio_oeb[23]
  PIN mgmt_gpio_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 509.600 4.000 510.160 ;
    END
  END mgmt_gpio_oeb[24]
  PIN mgmt_gpio_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 528.080 4.000 528.640 ;
    END
  END mgmt_gpio_oeb[25]
  PIN mgmt_gpio_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 546.560 4.000 547.120 ;
    END
  END mgmt_gpio_oeb[26]
  PIN mgmt_gpio_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 565.040 4.000 565.600 ;
    END
  END mgmt_gpio_oeb[27]
  PIN mgmt_gpio_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 583.520 4.000 584.080 ;
    END
  END mgmt_gpio_oeb[28]
  PIN mgmt_gpio_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 602.000 4.000 602.560 ;
    END
  END mgmt_gpio_oeb[29]
  PIN mgmt_gpio_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 154.560 620.000 155.120 ;
    END
  END mgmt_gpio_oeb[2]
  PIN mgmt_gpio_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 620.480 4.000 621.040 ;
    END
  END mgmt_gpio_oeb[30]
  PIN mgmt_gpio_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 638.960 4.000 639.520 ;
    END
  END mgmt_gpio_oeb[31]
  PIN mgmt_gpio_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 657.440 4.000 658.000 ;
    END
  END mgmt_gpio_oeb[32]
  PIN mgmt_gpio_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 675.920 4.000 676.480 ;
    END
  END mgmt_gpio_oeb[33]
  PIN mgmt_gpio_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 694.400 4.000 694.960 ;
    END
  END mgmt_gpio_oeb[34]
  PIN mgmt_gpio_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 712.880 4.000 713.440 ;
    END
  END mgmt_gpio_oeb[35]
  PIN mgmt_gpio_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 731.360 4.000 731.920 ;
    END
  END mgmt_gpio_oeb[36]
  PIN mgmt_gpio_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 749.840 4.000 750.400 ;
    END
  END mgmt_gpio_oeb[37]
  PIN mgmt_gpio_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 189.840 620.000 190.400 ;
    END
  END mgmt_gpio_oeb[3]
  PIN mgmt_gpio_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 225.120 620.000 225.680 ;
    END
  END mgmt_gpio_oeb[4]
  PIN mgmt_gpio_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 260.400 620.000 260.960 ;
    END
  END mgmt_gpio_oeb[5]
  PIN mgmt_gpio_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 295.680 620.000 296.240 ;
    END
  END mgmt_gpio_oeb[6]
  PIN mgmt_gpio_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 330.960 620.000 331.520 ;
    END
  END mgmt_gpio_oeb[7]
  PIN mgmt_gpio_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 366.240 620.000 366.800 ;
    END
  END mgmt_gpio_oeb[8]
  PIN mgmt_gpio_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 401.520 620.000 402.080 ;
    END
  END mgmt_gpio_oeb[9]
  PIN mgmt_gpio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 95.760 620.000 96.320 ;
    END
  END mgmt_gpio_out[0]
  PIN mgmt_gpio_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 448.560 620.000 449.120 ;
    END
  END mgmt_gpio_out[10]
  PIN mgmt_gpio_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 483.840 620.000 484.400 ;
    END
  END mgmt_gpio_out[11]
  PIN mgmt_gpio_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 519.120 620.000 519.680 ;
    END
  END mgmt_gpio_out[12]
  PIN mgmt_gpio_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 554.400 620.000 554.960 ;
    END
  END mgmt_gpio_out[13]
  PIN mgmt_gpio_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 589.680 620.000 590.240 ;
    END
  END mgmt_gpio_out[14]
  PIN mgmt_gpio_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 624.960 620.000 625.520 ;
    END
  END mgmt_gpio_out[15]
  PIN mgmt_gpio_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 660.240 620.000 660.800 ;
    END
  END mgmt_gpio_out[16]
  PIN mgmt_gpio_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 695.520 620.000 696.080 ;
    END
  END mgmt_gpio_out[17]
  PIN mgmt_gpio_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 730.800 620.000 731.360 ;
    END
  END mgmt_gpio_out[18]
  PIN mgmt_gpio_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 766.080 620.000 766.640 ;
    END
  END mgmt_gpio_out[19]
  PIN mgmt_gpio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 131.040 620.000 131.600 ;
    END
  END mgmt_gpio_out[1]
  PIN mgmt_gpio_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 441.840 4.000 442.400 ;
    END
  END mgmt_gpio_out[20]
  PIN mgmt_gpio_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 460.320 4.000 460.880 ;
    END
  END mgmt_gpio_out[21]
  PIN mgmt_gpio_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 478.800 4.000 479.360 ;
    END
  END mgmt_gpio_out[22]
  PIN mgmt_gpio_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 497.280 4.000 497.840 ;
    END
  END mgmt_gpio_out[23]
  PIN mgmt_gpio_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 515.760 4.000 516.320 ;
    END
  END mgmt_gpio_out[24]
  PIN mgmt_gpio_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 534.240 4.000 534.800 ;
    END
  END mgmt_gpio_out[25]
  PIN mgmt_gpio_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 552.720 4.000 553.280 ;
    END
  END mgmt_gpio_out[26]
  PIN mgmt_gpio_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 571.200 4.000 571.760 ;
    END
  END mgmt_gpio_out[27]
  PIN mgmt_gpio_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 589.680 4.000 590.240 ;
    END
  END mgmt_gpio_out[28]
  PIN mgmt_gpio_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 608.160 4.000 608.720 ;
    END
  END mgmt_gpio_out[29]
  PIN mgmt_gpio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 166.320 620.000 166.880 ;
    END
  END mgmt_gpio_out[2]
  PIN mgmt_gpio_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 626.640 4.000 627.200 ;
    END
  END mgmt_gpio_out[30]
  PIN mgmt_gpio_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 645.120 4.000 645.680 ;
    END
  END mgmt_gpio_out[31]
  PIN mgmt_gpio_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 663.600 4.000 664.160 ;
    END
  END mgmt_gpio_out[32]
  PIN mgmt_gpio_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 682.080 4.000 682.640 ;
    END
  END mgmt_gpio_out[33]
  PIN mgmt_gpio_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 700.560 4.000 701.120 ;
    END
  END mgmt_gpio_out[34]
  PIN mgmt_gpio_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 719.040 4.000 719.600 ;
    END
  END mgmt_gpio_out[35]
  PIN mgmt_gpio_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 737.520 4.000 738.080 ;
    END
  END mgmt_gpio_out[36]
  PIN mgmt_gpio_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 756.000 4.000 756.560 ;
    END
  END mgmt_gpio_out[37]
  PIN mgmt_gpio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 201.600 620.000 202.160 ;
    END
  END mgmt_gpio_out[3]
  PIN mgmt_gpio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 236.880 620.000 237.440 ;
    END
  END mgmt_gpio_out[4]
  PIN mgmt_gpio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 272.160 620.000 272.720 ;
    END
  END mgmt_gpio_out[5]
  PIN mgmt_gpio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 307.440 620.000 308.000 ;
    END
  END mgmt_gpio_out[6]
  PIN mgmt_gpio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 342.720 620.000 343.280 ;
    END
  END mgmt_gpio_out[7]
  PIN mgmt_gpio_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 378.000 620.000 378.560 ;
    END
  END mgmt_gpio_out[8]
  PIN mgmt_gpio_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 413.280 620.000 413.840 ;
    END
  END mgmt_gpio_out[9]
  PIN pad_flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 17.360 0.000 17.920 4.000 ;
    END
  END pad_flash_clk
  PIN pad_flash_clk_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 24.080 0.000 24.640 4.000 ;
    END
  END pad_flash_clk_oe
  PIN pad_flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.800 0.000 31.360 4.000 ;
    END
  END pad_flash_csb
  PIN pad_flash_csb_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 37.520 0.000 38.080 4.000 ;
    END
  END pad_flash_csb_oe
  PIN pad_flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 44.240 0.000 44.800 4.000 ;
    END
  END pad_flash_io0_di
  PIN pad_flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.960 0.000 51.520 4.000 ;
    END
  END pad_flash_io0_do
  PIN pad_flash_io0_ie
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.680 0.000 58.240 4.000 ;
    END
  END pad_flash_io0_ie
  PIN pad_flash_io0_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 64.400 0.000 64.960 4.000 ;
    END
  END pad_flash_io0_oe
  PIN pad_flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 71.120 0.000 71.680 4.000 ;
    END
  END pad_flash_io1_di
  PIN pad_flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.840 0.000 78.400 4.000 ;
    END
  END pad_flash_io1_do
  PIN pad_flash_io1_ie
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.560 0.000 85.120 4.000 ;
    END
  END pad_flash_io1_ie
  PIN pad_flash_io1_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 91.280 0.000 91.840 4.000 ;
    END
  END pad_flash_io1_oe
  PIN pll90_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.640 0.000 179.200 4.000 ;
    END
  END pll90_sel[0]
  PIN pll90_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 185.360 0.000 185.920 4.000 ;
    END
  END pll90_sel[1]
  PIN pll90_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 192.080 0.000 192.640 4.000 ;
    END
  END pll90_sel[2]
  PIN pll_bypass
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 373.520 0.000 374.080 4.000 ;
    END
  END pll_bypass
  PIN pll_dco_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 118.160 0.000 118.720 4.000 ;
    END
  END pll_dco_ena
  PIN pll_div[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.880 0.000 125.440 4.000 ;
    END
  END pll_div[0]
  PIN pll_div[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.600 0.000 132.160 4.000 ;
    END
  END pll_div[1]
  PIN pll_div[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 138.320 0.000 138.880 4.000 ;
    END
  END pll_div[2]
  PIN pll_div[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 145.040 0.000 145.600 4.000 ;
    END
  END pll_div[3]
  PIN pll_div[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.760 0.000 152.320 4.000 ;
    END
  END pll_div[4]
  PIN pll_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 111.440 0.000 112.000 4.000 ;
    END
  END pll_ena
  PIN pll_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 158.480 0.000 159.040 4.000 ;
    END
  END pll_sel[0]
  PIN pll_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 165.200 0.000 165.760 4.000 ;
    END
  END pll_sel[1]
  PIN pll_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.920 0.000 172.480 4.000 ;
    END
  END pll_sel[2]
  PIN pll_trim[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 198.800 0.000 199.360 4.000 ;
    END
  END pll_trim[0]
  PIN pll_trim[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 266.000 0.000 266.560 4.000 ;
    END
  END pll_trim[10]
  PIN pll_trim[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.720 0.000 273.280 4.000 ;
    END
  END pll_trim[11]
  PIN pll_trim[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 279.440 0.000 280.000 4.000 ;
    END
  END pll_trim[12]
  PIN pll_trim[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 286.160 0.000 286.720 4.000 ;
    END
  END pll_trim[13]
  PIN pll_trim[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.880 0.000 293.440 4.000 ;
    END
  END pll_trim[14]
  PIN pll_trim[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.600 0.000 300.160 4.000 ;
    END
  END pll_trim[15]
  PIN pll_trim[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 306.320 0.000 306.880 4.000 ;
    END
  END pll_trim[16]
  PIN pll_trim[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 313.040 0.000 313.600 4.000 ;
    END
  END pll_trim[17]
  PIN pll_trim[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 319.760 0.000 320.320 4.000 ;
    END
  END pll_trim[18]
  PIN pll_trim[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 326.480 0.000 327.040 4.000 ;
    END
  END pll_trim[19]
  PIN pll_trim[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 205.520 0.000 206.080 4.000 ;
    END
  END pll_trim[1]
  PIN pll_trim[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 333.200 0.000 333.760 4.000 ;
    END
  END pll_trim[20]
  PIN pll_trim[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 339.920 0.000 340.480 4.000 ;
    END
  END pll_trim[21]
  PIN pll_trim[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 346.640 0.000 347.200 4.000 ;
    END
  END pll_trim[22]
  PIN pll_trim[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 353.360 0.000 353.920 4.000 ;
    END
  END pll_trim[23]
  PIN pll_trim[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 360.080 0.000 360.640 4.000 ;
    END
  END pll_trim[24]
  PIN pll_trim[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.800 0.000 367.360 4.000 ;
    END
  END pll_trim[25]
  PIN pll_trim[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 212.240 0.000 212.800 4.000 ;
    END
  END pll_trim[2]
  PIN pll_trim[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.960 0.000 219.520 4.000 ;
    END
  END pll_trim[3]
  PIN pll_trim[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.680 0.000 226.240 4.000 ;
    END
  END pll_trim[4]
  PIN pll_trim[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 232.400 0.000 232.960 4.000 ;
    END
  END pll_trim[5]
  PIN pll_trim[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 239.120 0.000 239.680 4.000 ;
    END
  END pll_trim[6]
  PIN pll_trim[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.840 0.000 246.400 4.000 ;
    END
  END pll_trim[7]
  PIN pll_trim[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.560 0.000 253.120 4.000 ;
    END
  END pll_trim[8]
  PIN pll_trim[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 259.280 0.000 259.840 4.000 ;
    END
  END pll_trim[9]
  PIN porb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 98.000 0.000 98.560 4.000 ;
    END
  END porb
  PIN pwr_ctrl_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 608.720 0.000 609.280 4.000 ;
    END
  END pwr_ctrl_out
  PIN qspi_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 115.360 4.000 115.920 ;
    END
  END qspi_enabled
  PIN reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.720 0.000 105.280 4.000 ;
    END
  END reset
  PIN ser_rx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 109.200 4.000 109.760 ;
    END
  END ser_rx
  PIN ser_tx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 103.040 4.000 103.600 ;
    END
  END ser_tx
  PIN serial_clock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 13.440 620.000 14.000 ;
    END
  END serial_clock
  PIN serial_data_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 48.720 620.000 49.280 ;
    END
  END serial_data_1
  PIN serial_data_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 60.480 620.000 61.040 ;
    END
  END serial_data_2
  PIN serial_load
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 36.960 620.000 37.520 ;
    END
  END serial_load
  PIN serial_resetn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 25.200 620.000 25.760 ;
    END
  END serial_resetn
  PIN spi_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.720 4.000 91.280 ;
    END
  END spi_csb
  PIN spi_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END spi_enabled
  PIN spi_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.560 4.000 85.120 ;
    END
  END spi_sck
  PIN spi_sdi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 96.880 4.000 97.440 ;
    END
  END spi_sdi
  PIN spi_sdo
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 78.400 4.000 78.960 ;
    END
  END spi_sdo
  PIN spi_sdoenb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 72.240 4.000 72.800 ;
    END
  END spi_sdoenb
  PIN spimemio_flash_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 343.280 4.000 343.840 ;
    END
  END spimemio_flash_clk
  PIN spimemio_flash_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 349.440 4.000 350.000 ;
    END
  END spimemio_flash_csb
  PIN spimemio_flash_io0_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 355.600 4.000 356.160 ;
    END
  END spimemio_flash_io0_di
  PIN spimemio_flash_io0_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 361.760 4.000 362.320 ;
    END
  END spimemio_flash_io0_do
  PIN spimemio_flash_io0_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 367.920 4.000 368.480 ;
    END
  END spimemio_flash_io0_oeb
  PIN spimemio_flash_io1_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 374.080 4.000 374.640 ;
    END
  END spimemio_flash_io1_di
  PIN spimemio_flash_io1_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 380.240 4.000 380.800 ;
    END
  END spimemio_flash_io1_do
  PIN spimemio_flash_io1_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 386.400 4.000 386.960 ;
    END
  END spimemio_flash_io1_oeb
  PIN spimemio_flash_io2_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 392.560 4.000 393.120 ;
    END
  END spimemio_flash_io2_di
  PIN spimemio_flash_io2_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 398.720 4.000 399.280 ;
    END
  END spimemio_flash_io2_do
  PIN spimemio_flash_io2_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 404.880 4.000 405.440 ;
    END
  END spimemio_flash_io2_oeb
  PIN spimemio_flash_io3_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 411.040 4.000 411.600 ;
    END
  END spimemio_flash_io3_di
  PIN spimemio_flash_io3_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 417.200 4.000 417.760 ;
    END
  END spimemio_flash_io3_do
  PIN spimemio_flash_io3_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 423.360 4.000 423.920 ;
    END
  END spimemio_flash_io3_oeb
  PIN trap
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 47.600 4.000 48.160 ;
    END
  END trap
  PIN uart_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 121.520 4.000 122.080 ;
    END
  END uart_enabled
  PIN user_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.640 0.000 11.200 4.000 ;
    END
  END user_clock
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 133.840 4.000 134.400 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.600 776.000 20.160 780.000 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.600 776.000 104.160 780.000 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 776.000 112.560 780.000 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.400 776.000 120.960 780.000 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 776.000 129.360 780.000 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.200 776.000 137.760 780.000 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 776.000 146.160 780.000 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.000 776.000 154.560 780.000 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 776.000 162.960 780.000 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 170.800 776.000 171.360 780.000 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 776.000 179.760 780.000 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 776.000 28.560 780.000 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.600 776.000 188.160 780.000 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 776.000 196.560 780.000 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.400 776.000 204.960 780.000 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 776.000 213.360 780.000 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.200 776.000 221.760 780.000 ;
    END
  END wb_adr_i[24]
  PIN wb_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 776.000 230.160 780.000 ;
    END
  END wb_adr_i[25]
  PIN wb_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.000 776.000 238.560 780.000 ;
    END
  END wb_adr_i[26]
  PIN wb_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 246.400 776.000 246.960 780.000 ;
    END
  END wb_adr_i[27]
  PIN wb_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 254.800 776.000 255.360 780.000 ;
    END
  END wb_adr_i[28]
  PIN wb_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 776.000 263.760 780.000 ;
    END
  END wb_adr_i[29]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.400 776.000 36.960 780.000 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 271.600 776.000 272.160 780.000 ;
    END
  END wb_adr_i[30]
  PIN wb_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 776.000 280.560 780.000 ;
    END
  END wb_adr_i[31]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 776.000 45.360 780.000 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.200 776.000 53.760 780.000 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 776.000 62.160 780.000 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.000 776.000 70.560 780.000 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 776.000 78.960 780.000 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.800 776.000 87.360 780.000 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 776.000 95.760 780.000 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 380.240 0.000 380.800 4.000 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 599.200 776.000 599.760 780.000 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.400 776.000 288.960 780.000 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.400 776.000 372.960 780.000 ;
    END
  END wb_dat_i[10]
  PIN wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 380.800 776.000 381.360 780.000 ;
    END
  END wb_dat_i[11]
  PIN wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 389.200 776.000 389.760 780.000 ;
    END
  END wb_dat_i[12]
  PIN wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 397.600 776.000 398.160 780.000 ;
    END
  END wb_dat_i[13]
  PIN wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.000 776.000 406.560 780.000 ;
    END
  END wb_dat_i[14]
  PIN wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 776.000 414.960 780.000 ;
    END
  END wb_dat_i[15]
  PIN wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 422.800 776.000 423.360 780.000 ;
    END
  END wb_dat_i[16]
  PIN wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 431.200 776.000 431.760 780.000 ;
    END
  END wb_dat_i[17]
  PIN wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 439.600 776.000 440.160 780.000 ;
    END
  END wb_dat_i[18]
  PIN wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 448.000 776.000 448.560 780.000 ;
    END
  END wb_dat_i[19]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 776.000 297.360 780.000 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.400 776.000 456.960 780.000 ;
    END
  END wb_dat_i[20]
  PIN wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 464.800 776.000 465.360 780.000 ;
    END
  END wb_dat_i[21]
  PIN wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.200 776.000 473.760 780.000 ;
    END
  END wb_dat_i[22]
  PIN wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 481.600 776.000 482.160 780.000 ;
    END
  END wb_dat_i[23]
  PIN wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 490.000 776.000 490.560 780.000 ;
    END
  END wb_dat_i[24]
  PIN wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 498.400 776.000 498.960 780.000 ;
    END
  END wb_dat_i[25]
  PIN wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 506.800 776.000 507.360 780.000 ;
    END
  END wb_dat_i[26]
  PIN wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 515.200 776.000 515.760 780.000 ;
    END
  END wb_dat_i[27]
  PIN wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 523.600 776.000 524.160 780.000 ;
    END
  END wb_dat_i[28]
  PIN wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 532.000 776.000 532.560 780.000 ;
    END
  END wb_dat_i[29]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 305.200 776.000 305.760 780.000 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 540.400 776.000 540.960 780.000 ;
    END
  END wb_dat_i[30]
  PIN wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 548.800 776.000 549.360 780.000 ;
    END
  END wb_dat_i[31]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 313.600 776.000 314.160 780.000 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.000 776.000 322.560 780.000 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 330.400 776.000 330.960 780.000 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 338.800 776.000 339.360 780.000 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 347.200 776.000 347.760 780.000 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 355.600 776.000 356.160 780.000 ;
    END
  END wb_dat_i[8]
  PIN wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 364.000 776.000 364.560 780.000 ;
    END
  END wb_dat_i[9]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 146.160 4.000 146.720 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.760 4.000 208.320 ;
    END
  END wb_dat_o[10]
  PIN wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 213.920 4.000 214.480 ;
    END
  END wb_dat_o[11]
  PIN wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 220.080 4.000 220.640 ;
    END
  END wb_dat_o[12]
  PIN wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 226.240 4.000 226.800 ;
    END
  END wb_dat_o[13]
  PIN wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 232.400 4.000 232.960 ;
    END
  END wb_dat_o[14]
  PIN wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 238.560 4.000 239.120 ;
    END
  END wb_dat_o[15]
  PIN wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 244.720 4.000 245.280 ;
    END
  END wb_dat_o[16]
  PIN wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 250.880 4.000 251.440 ;
    END
  END wb_dat_o[17]
  PIN wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 257.040 4.000 257.600 ;
    END
  END wb_dat_o[18]
  PIN wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 263.200 4.000 263.760 ;
    END
  END wb_dat_o[19]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 152.320 4.000 152.880 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 269.360 4.000 269.920 ;
    END
  END wb_dat_o[20]
  PIN wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 275.520 4.000 276.080 ;
    END
  END wb_dat_o[21]
  PIN wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 281.680 4.000 282.240 ;
    END
  END wb_dat_o[22]
  PIN wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 287.840 4.000 288.400 ;
    END
  END wb_dat_o[23]
  PIN wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.000 4.000 294.560 ;
    END
  END wb_dat_o[24]
  PIN wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 300.160 4.000 300.720 ;
    END
  END wb_dat_o[25]
  PIN wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 306.320 4.000 306.880 ;
    END
  END wb_dat_o[26]
  PIN wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 312.480 4.000 313.040 ;
    END
  END wb_dat_o[27]
  PIN wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.640 4.000 319.200 ;
    END
  END wb_dat_o[28]
  PIN wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 324.800 4.000 325.360 ;
    END
  END wb_dat_o[29]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 158.480 4.000 159.040 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 330.960 4.000 331.520 ;
    END
  END wb_dat_o[30]
  PIN wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 337.120 4.000 337.680 ;
    END
  END wb_dat_o[31]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 4.000 165.200 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 170.800 4.000 171.360 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 176.960 4.000 177.520 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 183.120 4.000 183.680 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 189.280 4.000 189.840 ;
    END
  END wb_dat_o[7]
  PIN wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 195.440 4.000 196.000 ;
    END
  END wb_dat_o[8]
  PIN wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END wb_dat_o[9]
  PIN wb_rstn_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.960 0.000 387.520 4.000 ;
    END
  END wb_rstn_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 557.200 776.000 557.760 780.000 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 565.600 776.000 566.160 780.000 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 574.000 776.000 574.560 780.000 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 582.400 776.000 582.960 780.000 ;
    END
  END wb_sel_i[3]
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 140.000 4.000 140.560 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 590.800 776.000 591.360 780.000 ;
    END
  END wb_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 613.200 762.010 ;
      LAYER Metal2 ;
        RECT 4.060 775.700 19.300 776.580 ;
        RECT 20.460 775.700 27.700 776.580 ;
        RECT 28.860 775.700 36.100 776.580 ;
        RECT 37.260 775.700 44.500 776.580 ;
        RECT 45.660 775.700 52.900 776.580 ;
        RECT 54.060 775.700 61.300 776.580 ;
        RECT 62.460 775.700 69.700 776.580 ;
        RECT 70.860 775.700 78.100 776.580 ;
        RECT 79.260 775.700 86.500 776.580 ;
        RECT 87.660 775.700 94.900 776.580 ;
        RECT 96.060 775.700 103.300 776.580 ;
        RECT 104.460 775.700 111.700 776.580 ;
        RECT 112.860 775.700 120.100 776.580 ;
        RECT 121.260 775.700 128.500 776.580 ;
        RECT 129.660 775.700 136.900 776.580 ;
        RECT 138.060 775.700 145.300 776.580 ;
        RECT 146.460 775.700 153.700 776.580 ;
        RECT 154.860 775.700 162.100 776.580 ;
        RECT 163.260 775.700 170.500 776.580 ;
        RECT 171.660 775.700 178.900 776.580 ;
        RECT 180.060 775.700 187.300 776.580 ;
        RECT 188.460 775.700 195.700 776.580 ;
        RECT 196.860 775.700 204.100 776.580 ;
        RECT 205.260 775.700 212.500 776.580 ;
        RECT 213.660 775.700 220.900 776.580 ;
        RECT 222.060 775.700 229.300 776.580 ;
        RECT 230.460 775.700 237.700 776.580 ;
        RECT 238.860 775.700 246.100 776.580 ;
        RECT 247.260 775.700 254.500 776.580 ;
        RECT 255.660 775.700 262.900 776.580 ;
        RECT 264.060 775.700 271.300 776.580 ;
        RECT 272.460 775.700 279.700 776.580 ;
        RECT 280.860 775.700 288.100 776.580 ;
        RECT 289.260 775.700 296.500 776.580 ;
        RECT 297.660 775.700 304.900 776.580 ;
        RECT 306.060 775.700 313.300 776.580 ;
        RECT 314.460 775.700 321.700 776.580 ;
        RECT 322.860 775.700 330.100 776.580 ;
        RECT 331.260 775.700 338.500 776.580 ;
        RECT 339.660 775.700 346.900 776.580 ;
        RECT 348.060 775.700 355.300 776.580 ;
        RECT 356.460 775.700 363.700 776.580 ;
        RECT 364.860 775.700 372.100 776.580 ;
        RECT 373.260 775.700 380.500 776.580 ;
        RECT 381.660 775.700 388.900 776.580 ;
        RECT 390.060 775.700 397.300 776.580 ;
        RECT 398.460 775.700 405.700 776.580 ;
        RECT 406.860 775.700 414.100 776.580 ;
        RECT 415.260 775.700 422.500 776.580 ;
        RECT 423.660 775.700 430.900 776.580 ;
        RECT 432.060 775.700 439.300 776.580 ;
        RECT 440.460 775.700 447.700 776.580 ;
        RECT 448.860 775.700 456.100 776.580 ;
        RECT 457.260 775.700 464.500 776.580 ;
        RECT 465.660 775.700 472.900 776.580 ;
        RECT 474.060 775.700 481.300 776.580 ;
        RECT 482.460 775.700 489.700 776.580 ;
        RECT 490.860 775.700 498.100 776.580 ;
        RECT 499.260 775.700 506.500 776.580 ;
        RECT 507.660 775.700 514.900 776.580 ;
        RECT 516.060 775.700 523.300 776.580 ;
        RECT 524.460 775.700 531.700 776.580 ;
        RECT 532.860 775.700 540.100 776.580 ;
        RECT 541.260 775.700 548.500 776.580 ;
        RECT 549.660 775.700 556.900 776.580 ;
        RECT 558.060 775.700 565.300 776.580 ;
        RECT 566.460 775.700 573.700 776.580 ;
        RECT 574.860 775.700 582.100 776.580 ;
        RECT 583.260 775.700 590.500 776.580 ;
        RECT 591.660 775.700 598.900 776.580 ;
        RECT 600.060 775.700 617.540 776.580 ;
        RECT 4.060 4.300 617.540 775.700 ;
        RECT 4.060 0.090 10.340 4.300 ;
        RECT 11.500 0.090 17.060 4.300 ;
        RECT 18.220 0.090 23.780 4.300 ;
        RECT 24.940 0.090 30.500 4.300 ;
        RECT 31.660 0.090 37.220 4.300 ;
        RECT 38.380 0.090 43.940 4.300 ;
        RECT 45.100 0.090 50.660 4.300 ;
        RECT 51.820 0.090 57.380 4.300 ;
        RECT 58.540 0.090 64.100 4.300 ;
        RECT 65.260 0.090 70.820 4.300 ;
        RECT 71.980 0.090 77.540 4.300 ;
        RECT 78.700 0.090 84.260 4.300 ;
        RECT 85.420 0.090 90.980 4.300 ;
        RECT 92.140 0.090 97.700 4.300 ;
        RECT 98.860 0.090 104.420 4.300 ;
        RECT 105.580 0.090 111.140 4.300 ;
        RECT 112.300 0.090 117.860 4.300 ;
        RECT 119.020 0.090 124.580 4.300 ;
        RECT 125.740 0.090 131.300 4.300 ;
        RECT 132.460 0.090 138.020 4.300 ;
        RECT 139.180 0.090 144.740 4.300 ;
        RECT 145.900 0.090 151.460 4.300 ;
        RECT 152.620 0.090 158.180 4.300 ;
        RECT 159.340 0.090 164.900 4.300 ;
        RECT 166.060 0.090 171.620 4.300 ;
        RECT 172.780 0.090 178.340 4.300 ;
        RECT 179.500 0.090 185.060 4.300 ;
        RECT 186.220 0.090 191.780 4.300 ;
        RECT 192.940 0.090 198.500 4.300 ;
        RECT 199.660 0.090 205.220 4.300 ;
        RECT 206.380 0.090 211.940 4.300 ;
        RECT 213.100 0.090 218.660 4.300 ;
        RECT 219.820 0.090 225.380 4.300 ;
        RECT 226.540 0.090 232.100 4.300 ;
        RECT 233.260 0.090 238.820 4.300 ;
        RECT 239.980 0.090 245.540 4.300 ;
        RECT 246.700 0.090 252.260 4.300 ;
        RECT 253.420 0.090 258.980 4.300 ;
        RECT 260.140 0.090 265.700 4.300 ;
        RECT 266.860 0.090 272.420 4.300 ;
        RECT 273.580 0.090 279.140 4.300 ;
        RECT 280.300 0.090 285.860 4.300 ;
        RECT 287.020 0.090 292.580 4.300 ;
        RECT 293.740 0.090 299.300 4.300 ;
        RECT 300.460 0.090 306.020 4.300 ;
        RECT 307.180 0.090 312.740 4.300 ;
        RECT 313.900 0.090 319.460 4.300 ;
        RECT 320.620 0.090 326.180 4.300 ;
        RECT 327.340 0.090 332.900 4.300 ;
        RECT 334.060 0.090 339.620 4.300 ;
        RECT 340.780 0.090 346.340 4.300 ;
        RECT 347.500 0.090 353.060 4.300 ;
        RECT 354.220 0.090 359.780 4.300 ;
        RECT 360.940 0.090 366.500 4.300 ;
        RECT 367.660 0.090 373.220 4.300 ;
        RECT 374.380 0.090 379.940 4.300 ;
        RECT 381.100 0.090 386.660 4.300 ;
        RECT 387.820 0.090 393.380 4.300 ;
        RECT 394.540 0.090 400.100 4.300 ;
        RECT 401.260 0.090 406.820 4.300 ;
        RECT 407.980 0.090 413.540 4.300 ;
        RECT 414.700 0.090 420.260 4.300 ;
        RECT 421.420 0.090 426.980 4.300 ;
        RECT 428.140 0.090 433.700 4.300 ;
        RECT 434.860 0.090 440.420 4.300 ;
        RECT 441.580 0.090 447.140 4.300 ;
        RECT 448.300 0.090 453.860 4.300 ;
        RECT 455.020 0.090 460.580 4.300 ;
        RECT 461.740 0.090 467.300 4.300 ;
        RECT 468.460 0.090 474.020 4.300 ;
        RECT 475.180 0.090 480.740 4.300 ;
        RECT 481.900 0.090 487.460 4.300 ;
        RECT 488.620 0.090 494.180 4.300 ;
        RECT 495.340 0.090 500.900 4.300 ;
        RECT 502.060 0.090 507.620 4.300 ;
        RECT 508.780 0.090 514.340 4.300 ;
        RECT 515.500 0.090 521.060 4.300 ;
        RECT 522.220 0.090 527.780 4.300 ;
        RECT 528.940 0.090 534.500 4.300 ;
        RECT 535.660 0.090 541.220 4.300 ;
        RECT 542.380 0.090 547.940 4.300 ;
        RECT 549.100 0.090 554.660 4.300 ;
        RECT 555.820 0.090 561.380 4.300 ;
        RECT 562.540 0.090 568.100 4.300 ;
        RECT 569.260 0.090 574.820 4.300 ;
        RECT 575.980 0.090 581.540 4.300 ;
        RECT 582.700 0.090 588.260 4.300 ;
        RECT 589.420 0.090 594.980 4.300 ;
        RECT 596.140 0.090 601.700 4.300 ;
        RECT 602.860 0.090 608.420 4.300 ;
        RECT 609.580 0.090 617.540 4.300 ;
      LAYER Metal3 ;
        RECT 1.210 765.780 615.700 766.500 ;
        RECT 1.210 756.860 617.590 765.780 ;
        RECT 4.300 755.700 617.590 756.860 ;
        RECT 1.210 755.180 617.590 755.700 ;
        RECT 1.210 754.020 615.700 755.180 ;
        RECT 1.210 750.700 617.590 754.020 ;
        RECT 4.300 749.540 617.590 750.700 ;
        RECT 1.210 744.540 617.590 749.540 ;
        RECT 4.300 743.420 617.590 744.540 ;
        RECT 4.300 743.380 615.700 743.420 ;
        RECT 1.210 742.260 615.700 743.380 ;
        RECT 1.210 738.380 617.590 742.260 ;
        RECT 4.300 737.220 617.590 738.380 ;
        RECT 1.210 732.220 617.590 737.220 ;
        RECT 4.300 731.660 617.590 732.220 ;
        RECT 4.300 731.060 615.700 731.660 ;
        RECT 1.210 730.500 615.700 731.060 ;
        RECT 1.210 726.060 617.590 730.500 ;
        RECT 4.300 724.900 617.590 726.060 ;
        RECT 1.210 719.900 617.590 724.900 ;
        RECT 4.300 718.740 615.700 719.900 ;
        RECT 1.210 713.740 617.590 718.740 ;
        RECT 4.300 712.580 617.590 713.740 ;
        RECT 1.210 708.140 617.590 712.580 ;
        RECT 1.210 707.580 615.700 708.140 ;
        RECT 4.300 706.980 615.700 707.580 ;
        RECT 4.300 706.420 617.590 706.980 ;
        RECT 1.210 701.420 617.590 706.420 ;
        RECT 4.300 700.260 617.590 701.420 ;
        RECT 1.210 696.380 617.590 700.260 ;
        RECT 1.210 695.260 615.700 696.380 ;
        RECT 4.300 695.220 615.700 695.260 ;
        RECT 4.300 694.100 617.590 695.220 ;
        RECT 1.210 689.100 617.590 694.100 ;
        RECT 4.300 687.940 617.590 689.100 ;
        RECT 1.210 684.620 617.590 687.940 ;
        RECT 1.210 683.460 615.700 684.620 ;
        RECT 1.210 682.940 617.590 683.460 ;
        RECT 4.300 681.780 617.590 682.940 ;
        RECT 1.210 676.780 617.590 681.780 ;
        RECT 4.300 675.620 617.590 676.780 ;
        RECT 1.210 672.860 617.590 675.620 ;
        RECT 1.210 671.700 615.700 672.860 ;
        RECT 1.210 670.620 617.590 671.700 ;
        RECT 4.300 669.460 617.590 670.620 ;
        RECT 1.210 664.460 617.590 669.460 ;
        RECT 4.300 663.300 617.590 664.460 ;
        RECT 1.210 661.100 617.590 663.300 ;
        RECT 1.210 659.940 615.700 661.100 ;
        RECT 1.210 658.300 617.590 659.940 ;
        RECT 4.300 657.140 617.590 658.300 ;
        RECT 1.210 652.140 617.590 657.140 ;
        RECT 4.300 650.980 617.590 652.140 ;
        RECT 1.210 649.340 617.590 650.980 ;
        RECT 1.210 648.180 615.700 649.340 ;
        RECT 1.210 645.980 617.590 648.180 ;
        RECT 4.300 644.820 617.590 645.980 ;
        RECT 1.210 639.820 617.590 644.820 ;
        RECT 4.300 638.660 617.590 639.820 ;
        RECT 1.210 637.580 617.590 638.660 ;
        RECT 1.210 636.420 615.700 637.580 ;
        RECT 1.210 633.660 617.590 636.420 ;
        RECT 4.300 632.500 617.590 633.660 ;
        RECT 1.210 627.500 617.590 632.500 ;
        RECT 4.300 626.340 617.590 627.500 ;
        RECT 1.210 625.820 617.590 626.340 ;
        RECT 1.210 624.660 615.700 625.820 ;
        RECT 1.210 621.340 617.590 624.660 ;
        RECT 4.300 620.180 617.590 621.340 ;
        RECT 1.210 615.180 617.590 620.180 ;
        RECT 4.300 614.060 617.590 615.180 ;
        RECT 4.300 614.020 615.700 614.060 ;
        RECT 1.210 612.900 615.700 614.020 ;
        RECT 1.210 609.020 617.590 612.900 ;
        RECT 4.300 607.860 617.590 609.020 ;
        RECT 1.210 602.860 617.590 607.860 ;
        RECT 4.300 602.300 617.590 602.860 ;
        RECT 4.300 601.700 615.700 602.300 ;
        RECT 1.210 601.140 615.700 601.700 ;
        RECT 1.210 596.700 617.590 601.140 ;
        RECT 4.300 595.540 617.590 596.700 ;
        RECT 1.210 590.540 617.590 595.540 ;
        RECT 4.300 589.380 615.700 590.540 ;
        RECT 1.210 584.380 617.590 589.380 ;
        RECT 4.300 583.220 617.590 584.380 ;
        RECT 1.210 578.780 617.590 583.220 ;
        RECT 1.210 578.220 615.700 578.780 ;
        RECT 4.300 577.620 615.700 578.220 ;
        RECT 4.300 577.060 617.590 577.620 ;
        RECT 1.210 572.060 617.590 577.060 ;
        RECT 4.300 570.900 617.590 572.060 ;
        RECT 1.210 567.020 617.590 570.900 ;
        RECT 1.210 565.900 615.700 567.020 ;
        RECT 4.300 565.860 615.700 565.900 ;
        RECT 4.300 564.740 617.590 565.860 ;
        RECT 1.210 559.740 617.590 564.740 ;
        RECT 4.300 558.580 617.590 559.740 ;
        RECT 1.210 555.260 617.590 558.580 ;
        RECT 1.210 554.100 615.700 555.260 ;
        RECT 1.210 553.580 617.590 554.100 ;
        RECT 4.300 552.420 617.590 553.580 ;
        RECT 1.210 547.420 617.590 552.420 ;
        RECT 4.300 546.260 617.590 547.420 ;
        RECT 1.210 543.500 617.590 546.260 ;
        RECT 1.210 542.340 615.700 543.500 ;
        RECT 1.210 541.260 617.590 542.340 ;
        RECT 4.300 540.100 617.590 541.260 ;
        RECT 1.210 535.100 617.590 540.100 ;
        RECT 4.300 533.940 617.590 535.100 ;
        RECT 1.210 531.740 617.590 533.940 ;
        RECT 1.210 530.580 615.700 531.740 ;
        RECT 1.210 528.940 617.590 530.580 ;
        RECT 4.300 527.780 617.590 528.940 ;
        RECT 1.210 522.780 617.590 527.780 ;
        RECT 4.300 521.620 617.590 522.780 ;
        RECT 1.210 519.980 617.590 521.620 ;
        RECT 1.210 518.820 615.700 519.980 ;
        RECT 1.210 516.620 617.590 518.820 ;
        RECT 4.300 515.460 617.590 516.620 ;
        RECT 1.210 510.460 617.590 515.460 ;
        RECT 4.300 509.300 617.590 510.460 ;
        RECT 1.210 508.220 617.590 509.300 ;
        RECT 1.210 507.060 615.700 508.220 ;
        RECT 1.210 504.300 617.590 507.060 ;
        RECT 4.300 503.140 617.590 504.300 ;
        RECT 1.210 498.140 617.590 503.140 ;
        RECT 4.300 496.980 617.590 498.140 ;
        RECT 1.210 496.460 617.590 496.980 ;
        RECT 1.210 495.300 615.700 496.460 ;
        RECT 1.210 491.980 617.590 495.300 ;
        RECT 4.300 490.820 617.590 491.980 ;
        RECT 1.210 485.820 617.590 490.820 ;
        RECT 4.300 484.700 617.590 485.820 ;
        RECT 4.300 484.660 615.700 484.700 ;
        RECT 1.210 483.540 615.700 484.660 ;
        RECT 1.210 479.660 617.590 483.540 ;
        RECT 4.300 478.500 617.590 479.660 ;
        RECT 1.210 473.500 617.590 478.500 ;
        RECT 4.300 472.940 617.590 473.500 ;
        RECT 4.300 472.340 615.700 472.940 ;
        RECT 1.210 471.780 615.700 472.340 ;
        RECT 1.210 467.340 617.590 471.780 ;
        RECT 4.300 466.180 617.590 467.340 ;
        RECT 1.210 461.180 617.590 466.180 ;
        RECT 4.300 460.020 615.700 461.180 ;
        RECT 1.210 455.020 617.590 460.020 ;
        RECT 4.300 453.860 617.590 455.020 ;
        RECT 1.210 449.420 617.590 453.860 ;
        RECT 1.210 448.860 615.700 449.420 ;
        RECT 4.300 448.260 615.700 448.860 ;
        RECT 4.300 447.700 617.590 448.260 ;
        RECT 1.210 442.700 617.590 447.700 ;
        RECT 4.300 441.540 617.590 442.700 ;
        RECT 1.210 437.660 617.590 441.540 ;
        RECT 1.210 436.540 615.700 437.660 ;
        RECT 4.300 436.500 615.700 436.540 ;
        RECT 4.300 435.380 617.590 436.500 ;
        RECT 1.210 430.380 617.590 435.380 ;
        RECT 4.300 429.220 617.590 430.380 ;
        RECT 1.210 425.900 617.590 429.220 ;
        RECT 1.210 424.740 615.700 425.900 ;
        RECT 1.210 424.220 617.590 424.740 ;
        RECT 4.300 423.060 617.590 424.220 ;
        RECT 1.210 418.060 617.590 423.060 ;
        RECT 4.300 416.900 617.590 418.060 ;
        RECT 1.210 414.140 617.590 416.900 ;
        RECT 1.210 412.980 615.700 414.140 ;
        RECT 1.210 411.900 617.590 412.980 ;
        RECT 4.300 410.740 617.590 411.900 ;
        RECT 1.210 405.740 617.590 410.740 ;
        RECT 4.300 404.580 617.590 405.740 ;
        RECT 1.210 402.380 617.590 404.580 ;
        RECT 1.210 401.220 615.700 402.380 ;
        RECT 1.210 399.580 617.590 401.220 ;
        RECT 4.300 398.420 617.590 399.580 ;
        RECT 1.210 393.420 617.590 398.420 ;
        RECT 4.300 392.260 617.590 393.420 ;
        RECT 1.210 390.620 617.590 392.260 ;
        RECT 1.210 389.460 615.700 390.620 ;
        RECT 1.210 387.260 617.590 389.460 ;
        RECT 4.300 386.100 617.590 387.260 ;
        RECT 1.210 381.100 617.590 386.100 ;
        RECT 4.300 379.940 617.590 381.100 ;
        RECT 1.210 378.860 617.590 379.940 ;
        RECT 1.210 377.700 615.700 378.860 ;
        RECT 1.210 374.940 617.590 377.700 ;
        RECT 4.300 373.780 617.590 374.940 ;
        RECT 1.210 368.780 617.590 373.780 ;
        RECT 4.300 367.620 617.590 368.780 ;
        RECT 1.210 367.100 617.590 367.620 ;
        RECT 1.210 365.940 615.700 367.100 ;
        RECT 1.210 362.620 617.590 365.940 ;
        RECT 4.300 361.460 617.590 362.620 ;
        RECT 1.210 356.460 617.590 361.460 ;
        RECT 4.300 355.340 617.590 356.460 ;
        RECT 4.300 355.300 615.700 355.340 ;
        RECT 1.210 354.180 615.700 355.300 ;
        RECT 1.210 350.300 617.590 354.180 ;
        RECT 4.300 349.140 617.590 350.300 ;
        RECT 1.210 344.140 617.590 349.140 ;
        RECT 4.300 343.580 617.590 344.140 ;
        RECT 4.300 342.980 615.700 343.580 ;
        RECT 1.210 342.420 615.700 342.980 ;
        RECT 1.210 337.980 617.590 342.420 ;
        RECT 4.300 336.820 617.590 337.980 ;
        RECT 1.210 331.820 617.590 336.820 ;
        RECT 4.300 330.660 615.700 331.820 ;
        RECT 1.210 325.660 617.590 330.660 ;
        RECT 4.300 324.500 617.590 325.660 ;
        RECT 1.210 320.060 617.590 324.500 ;
        RECT 1.210 319.500 615.700 320.060 ;
        RECT 4.300 318.900 615.700 319.500 ;
        RECT 4.300 318.340 617.590 318.900 ;
        RECT 1.210 313.340 617.590 318.340 ;
        RECT 4.300 312.180 617.590 313.340 ;
        RECT 1.210 308.300 617.590 312.180 ;
        RECT 1.210 307.180 615.700 308.300 ;
        RECT 4.300 307.140 615.700 307.180 ;
        RECT 4.300 306.020 617.590 307.140 ;
        RECT 1.210 301.020 617.590 306.020 ;
        RECT 4.300 299.860 617.590 301.020 ;
        RECT 1.210 296.540 617.590 299.860 ;
        RECT 1.210 295.380 615.700 296.540 ;
        RECT 1.210 294.860 617.590 295.380 ;
        RECT 4.300 293.700 617.590 294.860 ;
        RECT 1.210 288.700 617.590 293.700 ;
        RECT 4.300 287.540 617.590 288.700 ;
        RECT 1.210 284.780 617.590 287.540 ;
        RECT 1.210 283.620 615.700 284.780 ;
        RECT 1.210 282.540 617.590 283.620 ;
        RECT 4.300 281.380 617.590 282.540 ;
        RECT 1.210 276.380 617.590 281.380 ;
        RECT 4.300 275.220 617.590 276.380 ;
        RECT 1.210 273.020 617.590 275.220 ;
        RECT 1.210 271.860 615.700 273.020 ;
        RECT 1.210 270.220 617.590 271.860 ;
        RECT 4.300 269.060 617.590 270.220 ;
        RECT 1.210 264.060 617.590 269.060 ;
        RECT 4.300 262.900 617.590 264.060 ;
        RECT 1.210 261.260 617.590 262.900 ;
        RECT 1.210 260.100 615.700 261.260 ;
        RECT 1.210 257.900 617.590 260.100 ;
        RECT 4.300 256.740 617.590 257.900 ;
        RECT 1.210 251.740 617.590 256.740 ;
        RECT 4.300 250.580 617.590 251.740 ;
        RECT 1.210 249.500 617.590 250.580 ;
        RECT 1.210 248.340 615.700 249.500 ;
        RECT 1.210 245.580 617.590 248.340 ;
        RECT 4.300 244.420 617.590 245.580 ;
        RECT 1.210 239.420 617.590 244.420 ;
        RECT 4.300 238.260 617.590 239.420 ;
        RECT 1.210 237.740 617.590 238.260 ;
        RECT 1.210 236.580 615.700 237.740 ;
        RECT 1.210 233.260 617.590 236.580 ;
        RECT 4.300 232.100 617.590 233.260 ;
        RECT 1.210 227.100 617.590 232.100 ;
        RECT 4.300 225.980 617.590 227.100 ;
        RECT 4.300 225.940 615.700 225.980 ;
        RECT 1.210 224.820 615.700 225.940 ;
        RECT 1.210 220.940 617.590 224.820 ;
        RECT 4.300 219.780 617.590 220.940 ;
        RECT 1.210 214.780 617.590 219.780 ;
        RECT 4.300 214.220 617.590 214.780 ;
        RECT 4.300 213.620 615.700 214.220 ;
        RECT 1.210 213.060 615.700 213.620 ;
        RECT 1.210 208.620 617.590 213.060 ;
        RECT 4.300 207.460 617.590 208.620 ;
        RECT 1.210 202.460 617.590 207.460 ;
        RECT 4.300 201.300 615.700 202.460 ;
        RECT 1.210 196.300 617.590 201.300 ;
        RECT 4.300 195.140 617.590 196.300 ;
        RECT 1.210 190.700 617.590 195.140 ;
        RECT 1.210 190.140 615.700 190.700 ;
        RECT 4.300 189.540 615.700 190.140 ;
        RECT 4.300 188.980 617.590 189.540 ;
        RECT 1.210 183.980 617.590 188.980 ;
        RECT 4.300 182.820 617.590 183.980 ;
        RECT 1.210 178.940 617.590 182.820 ;
        RECT 1.210 177.820 615.700 178.940 ;
        RECT 4.300 177.780 615.700 177.820 ;
        RECT 4.300 176.660 617.590 177.780 ;
        RECT 1.210 171.660 617.590 176.660 ;
        RECT 4.300 170.500 617.590 171.660 ;
        RECT 1.210 167.180 617.590 170.500 ;
        RECT 1.210 166.020 615.700 167.180 ;
        RECT 1.210 165.500 617.590 166.020 ;
        RECT 4.300 164.340 617.590 165.500 ;
        RECT 1.210 159.340 617.590 164.340 ;
        RECT 4.300 158.180 617.590 159.340 ;
        RECT 1.210 155.420 617.590 158.180 ;
        RECT 1.210 154.260 615.700 155.420 ;
        RECT 1.210 153.180 617.590 154.260 ;
        RECT 4.300 152.020 617.590 153.180 ;
        RECT 1.210 147.020 617.590 152.020 ;
        RECT 4.300 145.860 617.590 147.020 ;
        RECT 1.210 143.660 617.590 145.860 ;
        RECT 1.210 142.500 615.700 143.660 ;
        RECT 1.210 140.860 617.590 142.500 ;
        RECT 4.300 139.700 617.590 140.860 ;
        RECT 1.210 134.700 617.590 139.700 ;
        RECT 4.300 133.540 617.590 134.700 ;
        RECT 1.210 131.900 617.590 133.540 ;
        RECT 1.210 130.740 615.700 131.900 ;
        RECT 1.210 128.540 617.590 130.740 ;
        RECT 4.300 127.380 617.590 128.540 ;
        RECT 1.210 122.380 617.590 127.380 ;
        RECT 4.300 121.220 617.590 122.380 ;
        RECT 1.210 120.140 617.590 121.220 ;
        RECT 1.210 118.980 615.700 120.140 ;
        RECT 1.210 116.220 617.590 118.980 ;
        RECT 4.300 115.060 617.590 116.220 ;
        RECT 1.210 110.060 617.590 115.060 ;
        RECT 4.300 108.900 617.590 110.060 ;
        RECT 1.210 108.380 617.590 108.900 ;
        RECT 1.210 107.220 615.700 108.380 ;
        RECT 1.210 103.900 617.590 107.220 ;
        RECT 4.300 102.740 617.590 103.900 ;
        RECT 1.210 97.740 617.590 102.740 ;
        RECT 4.300 96.620 617.590 97.740 ;
        RECT 4.300 96.580 615.700 96.620 ;
        RECT 1.210 95.460 615.700 96.580 ;
        RECT 1.210 91.580 617.590 95.460 ;
        RECT 4.300 90.420 617.590 91.580 ;
        RECT 1.210 85.420 617.590 90.420 ;
        RECT 4.300 84.860 617.590 85.420 ;
        RECT 4.300 84.260 615.700 84.860 ;
        RECT 1.210 83.700 615.700 84.260 ;
        RECT 1.210 79.260 617.590 83.700 ;
        RECT 4.300 78.100 617.590 79.260 ;
        RECT 1.210 73.100 617.590 78.100 ;
        RECT 4.300 71.940 615.700 73.100 ;
        RECT 1.210 66.940 617.590 71.940 ;
        RECT 4.300 65.780 617.590 66.940 ;
        RECT 1.210 61.340 617.590 65.780 ;
        RECT 1.210 60.780 615.700 61.340 ;
        RECT 4.300 60.180 615.700 60.780 ;
        RECT 4.300 59.620 617.590 60.180 ;
        RECT 1.210 54.620 617.590 59.620 ;
        RECT 4.300 53.460 617.590 54.620 ;
        RECT 1.210 49.580 617.590 53.460 ;
        RECT 1.210 48.460 615.700 49.580 ;
        RECT 4.300 48.420 615.700 48.460 ;
        RECT 4.300 47.300 617.590 48.420 ;
        RECT 1.210 42.300 617.590 47.300 ;
        RECT 4.300 41.140 617.590 42.300 ;
        RECT 1.210 37.820 617.590 41.140 ;
        RECT 1.210 36.660 615.700 37.820 ;
        RECT 1.210 36.140 617.590 36.660 ;
        RECT 4.300 34.980 617.590 36.140 ;
        RECT 1.210 29.980 617.590 34.980 ;
        RECT 4.300 28.820 617.590 29.980 ;
        RECT 1.210 26.060 617.590 28.820 ;
        RECT 1.210 24.900 615.700 26.060 ;
        RECT 1.210 23.820 617.590 24.900 ;
        RECT 4.300 22.660 617.590 23.820 ;
        RECT 1.210 14.300 617.590 22.660 ;
        RECT 1.210 13.140 615.700 14.300 ;
        RECT 1.210 0.140 617.590 13.140 ;
      LAYER Metal4 ;
        RECT 1.260 4.480 21.940 759.270 ;
        RECT 24.140 4.480 25.240 759.270 ;
        RECT 27.440 4.480 98.740 759.270 ;
        RECT 100.940 4.480 102.040 759.270 ;
        RECT 104.240 4.480 175.540 759.270 ;
        RECT 177.740 4.480 178.840 759.270 ;
        RECT 181.040 4.480 252.340 759.270 ;
        RECT 254.540 4.480 255.640 759.270 ;
        RECT 257.840 4.480 329.140 759.270 ;
        RECT 331.340 4.480 332.440 759.270 ;
        RECT 334.640 4.480 405.940 759.270 ;
        RECT 408.140 4.480 409.240 759.270 ;
        RECT 411.440 4.480 482.740 759.270 ;
        RECT 484.940 4.480 486.040 759.270 ;
        RECT 488.240 4.480 559.540 759.270 ;
        RECT 561.740 4.480 562.840 759.270 ;
        RECT 565.040 4.480 611.380 759.270 ;
        RECT 1.260 0.090 611.380 4.480 ;
      LAYER Metal5 ;
        RECT 1.180 593.390 611.460 618.180 ;
        RECT 1.180 563.390 611.460 590.790 ;
        RECT 1.180 533.390 611.460 560.790 ;
        RECT 1.180 503.390 611.460 530.790 ;
        RECT 1.180 473.390 611.460 500.790 ;
        RECT 1.180 443.390 611.460 470.790 ;
        RECT 1.180 413.390 611.460 440.790 ;
        RECT 1.180 383.390 611.460 410.790 ;
        RECT 1.180 353.390 611.460 380.790 ;
        RECT 1.180 323.390 611.460 350.790 ;
        RECT 1.180 293.390 611.460 320.790 ;
        RECT 1.180 263.390 611.460 290.790 ;
        RECT 1.180 233.390 611.460 260.790 ;
        RECT 1.180 203.390 611.460 230.790 ;
        RECT 1.180 173.390 611.460 200.790 ;
        RECT 1.180 143.390 611.460 170.790 ;
        RECT 1.180 113.390 611.460 140.790 ;
        RECT 1.180 83.390 611.460 110.790 ;
        RECT 1.180 53.390 611.460 80.790 ;
        RECT 1.180 23.390 611.460 50.790 ;
        RECT 1.180 10.180 611.460 20.790 ;
        RECT 1.180 6.880 611.460 7.580 ;
        RECT 1.180 1.180 611.460 4.280 ;
  END
END housekeeping
END LIBRARY

