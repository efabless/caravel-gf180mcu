magic
tech gf180mcuC
magscale 1 10
timestamp 1654631816
<< metal1 >>
rect 672 12570 34832 12604
rect 672 12518 4818 12570
rect 4870 12518 4922 12570
rect 4974 12518 5026 12570
rect 5078 12518 13370 12570
rect 13422 12518 13474 12570
rect 13526 12518 13578 12570
rect 13630 12518 21922 12570
rect 21974 12518 22026 12570
rect 22078 12518 22130 12570
rect 22182 12518 30474 12570
rect 30526 12518 30578 12570
rect 30630 12518 30682 12570
rect 30734 12518 34832 12570
rect 672 12484 34832 12518
rect 6918 12346 6970 12358
rect 6918 12282 6970 12294
rect 12406 12346 12458 12358
rect 12406 12282 12458 12294
rect 18342 12346 18394 12358
rect 18342 12282 18394 12294
rect 21422 12346 21474 12358
rect 21422 12282 21474 12294
rect 1822 12234 1874 12246
rect 1822 12170 1874 12182
rect 13358 12178 13410 12190
rect 2538 12070 2550 12122
rect 2602 12070 2614 12122
rect 9930 12114 9942 12166
rect 9994 12114 10006 12166
rect 10378 12114 10390 12166
rect 10442 12114 10454 12166
rect 19742 12178 19794 12190
rect 23370 12182 23382 12234
rect 23434 12182 23446 12234
rect 10826 12070 10838 12122
rect 10890 12070 10902 12122
rect 13358 12114 13410 12126
rect 13750 12122 13802 12134
rect 14746 12114 14758 12166
rect 14810 12114 14822 12166
rect 15306 12114 15318 12166
rect 15370 12114 15382 12166
rect 24154 12138 24166 12190
rect 24218 12138 24230 12190
rect 19742 12114 19794 12126
rect 20134 12122 20186 12134
rect 13750 12058 13802 12070
rect 14074 12024 14086 12076
rect 14138 12024 14150 12076
rect 18958 12066 19010 12078
rect 1934 12010 1986 12022
rect 1934 11946 1986 11958
rect 2158 12010 2210 12022
rect 10670 12010 10722 12022
rect 5002 11958 5014 12010
rect 5066 11958 5078 12010
rect 7578 11958 7590 12010
rect 7642 11958 7654 12010
rect 2158 11946 2210 11958
rect 10670 11946 10722 11958
rect 11006 12010 11058 12022
rect 11006 11946 11058 11958
rect 11398 12010 11450 12022
rect 11398 11946 11450 11958
rect 11734 12010 11786 12022
rect 11734 11946 11786 11958
rect 12070 12010 12122 12022
rect 12070 11946 12122 11958
rect 13022 12010 13074 12022
rect 13022 11946 13074 11958
rect 14590 12010 14642 12022
rect 20134 12058 20186 12070
rect 21086 12122 21138 12134
rect 17658 11958 17670 12010
rect 17722 11958 17734 12010
rect 18958 12002 19010 12014
rect 19406 12010 19458 12022
rect 20514 12014 20526 12066
rect 20578 12014 20590 12066
rect 21086 12058 21138 12070
rect 21814 12122 21866 12134
rect 24714 12114 24726 12166
rect 24778 12114 24790 12166
rect 25386 12114 25398 12166
rect 25450 12114 25462 12166
rect 28746 12126 28758 12178
rect 28810 12126 28822 12178
rect 30650 12114 30662 12166
rect 30714 12114 30726 12166
rect 31322 12114 31334 12166
rect 31386 12114 31398 12166
rect 21814 12058 21866 12070
rect 22138 12010 22150 12062
rect 22202 12010 22214 12062
rect 22654 12010 22706 12022
rect 14590 11946 14642 11958
rect 19406 11946 19458 11958
rect 27626 12004 27638 12056
rect 27690 12004 27702 12056
rect 28590 12010 28642 12022
rect 22654 11946 22706 11958
rect 29418 11958 29430 12010
rect 29482 11958 29494 12010
rect 33562 12004 33574 12056
rect 33626 12004 33638 12056
rect 34526 12010 34578 12022
rect 28590 11946 28642 11958
rect 34526 11946 34578 11958
rect 672 11786 34832 11820
rect 672 11734 9094 11786
rect 9146 11734 9198 11786
rect 9250 11734 9302 11786
rect 9354 11734 17646 11786
rect 17698 11734 17750 11786
rect 17802 11734 17854 11786
rect 17906 11734 26198 11786
rect 26250 11734 26302 11786
rect 26354 11734 26406 11786
rect 26458 11734 34832 11786
rect 672 11700 34832 11734
rect 2830 11562 2882 11574
rect 11174 11562 11226 11574
rect 2830 11498 2882 11510
rect 1374 11450 1426 11462
rect 1374 11386 1426 11398
rect 2606 11450 2658 11462
rect 2606 11386 2658 11398
rect 3278 11450 3330 11462
rect 3278 11386 3330 11398
rect 7142 11450 7194 11462
rect 8362 11458 8374 11510
rect 8426 11458 8438 11510
rect 11174 11498 11226 11510
rect 11790 11562 11842 11574
rect 11790 11498 11842 11510
rect 15990 11562 16042 11574
rect 7142 11386 7194 11398
rect 8710 11450 8762 11462
rect 12070 11450 12122 11462
rect 13794 11454 13806 11506
rect 13858 11454 13870 11506
rect 15990 11498 16042 11510
rect 16494 11562 16546 11574
rect 16494 11498 16546 11510
rect 17054 11562 17106 11574
rect 29934 11562 29986 11574
rect 17434 11510 17446 11562
rect 17498 11510 17510 11562
rect 17054 11498 17106 11510
rect 17894 11450 17946 11462
rect 8710 11386 8762 11398
rect 1710 11338 1762 11350
rect 2202 11330 2214 11382
rect 2266 11330 2278 11382
rect 3054 11338 3106 11350
rect 1710 11274 1762 11286
rect 3658 11330 3670 11382
rect 3722 11330 3734 11382
rect 4006 11338 4058 11350
rect 3054 11274 3106 11286
rect 4330 11330 4342 11382
rect 4394 11330 4406 11382
rect 4778 11330 4790 11382
rect 4842 11330 4854 11382
rect 9930 11360 9942 11412
rect 9994 11360 10006 11412
rect 9438 11338 9490 11350
rect 10490 11342 10502 11394
rect 10554 11342 10566 11394
rect 12070 11386 12122 11398
rect 16270 11394 16322 11406
rect 16874 11398 16886 11450
rect 16938 11398 16950 11450
rect 4006 11274 4058 11286
rect 11498 11330 11510 11382
rect 11562 11330 11574 11382
rect 12394 11330 12406 11382
rect 12458 11330 12470 11382
rect 13122 11342 13134 11394
rect 13186 11342 13198 11394
rect 17894 11386 17946 11398
rect 18790 11450 18842 11462
rect 18790 11386 18842 11398
rect 19294 11450 19346 11462
rect 19294 11386 19346 11398
rect 20022 11450 20074 11462
rect 20402 11454 20414 11506
rect 20466 11454 20478 11506
rect 29934 11498 29986 11510
rect 30270 11562 30322 11574
rect 30270 11498 30322 11510
rect 20022 11386 20074 11398
rect 21590 11450 21642 11462
rect 25118 11450 25170 11462
rect 21590 11386 21642 11398
rect 16270 11330 16322 11342
rect 20918 11338 20970 11350
rect 9438 11274 9490 11286
rect 1878 11226 1930 11238
rect 1878 11162 1930 11174
rect 7814 11226 7866 11238
rect 7814 11162 7866 11174
rect 9102 11226 9154 11238
rect 9102 11162 9154 11174
rect 10278 11226 10330 11238
rect 10602 11236 10614 11288
rect 10666 11236 10678 11288
rect 23930 11330 23942 11382
rect 23994 11330 24006 11382
rect 24490 11354 24502 11406
rect 24554 11354 24566 11406
rect 28970 11426 28982 11478
rect 29034 11426 29046 11478
rect 25118 11386 25170 11398
rect 26058 11354 26070 11406
rect 26122 11354 26134 11406
rect 26730 11354 26742 11406
rect 26794 11354 26806 11406
rect 33574 11394 33626 11406
rect 30046 11338 30098 11350
rect 30818 11342 30830 11394
rect 30882 11342 30894 11394
rect 20918 11274 20970 11286
rect 31210 11330 31222 11382
rect 31274 11330 31286 11382
rect 33574 11330 33626 11342
rect 30046 11274 30098 11286
rect 10278 11162 10330 11174
rect 10894 11226 10946 11238
rect 25006 11226 25058 11238
rect 16426 11174 16438 11226
rect 16490 11174 16502 11226
rect 18442 11174 18454 11226
rect 18506 11174 18518 11226
rect 10894 11162 10946 11174
rect 19630 11170 19682 11182
rect 25006 11162 25058 11174
rect 25342 11226 25394 11238
rect 25342 11162 25394 11174
rect 25678 11226 25730 11238
rect 25678 11162 25730 11174
rect 25790 11226 25842 11238
rect 34458 11174 34470 11226
rect 34522 11174 34534 11226
rect 25790 11162 25842 11174
rect 19630 11106 19682 11118
rect 672 11002 34832 11036
rect 672 10950 4818 11002
rect 4870 10950 4922 11002
rect 4974 10950 5026 11002
rect 5078 10950 13370 11002
rect 13422 10950 13474 11002
rect 13526 10950 13578 11002
rect 13630 10950 21922 11002
rect 21974 10950 22026 11002
rect 22078 10950 22130 11002
rect 22182 10950 30474 11002
rect 30526 10950 30578 11002
rect 30630 10950 30682 11002
rect 30734 10950 34832 11002
rect 672 10916 34832 10950
rect 9550 10778 9602 10790
rect 5854 10666 5906 10678
rect 1082 10566 1094 10618
rect 1146 10566 1158 10618
rect 3894 10610 3946 10622
rect 1586 10558 1598 10610
rect 1650 10558 1662 10610
rect 6414 10666 6466 10678
rect 8026 10670 8038 10722
rect 8090 10670 8102 10722
rect 9550 10714 9602 10726
rect 13806 10778 13858 10790
rect 13806 10714 13858 10726
rect 14422 10778 14474 10790
rect 14422 10714 14474 10726
rect 5854 10602 5906 10614
rect 5966 10610 6018 10622
rect 3894 10546 3946 10558
rect 5562 10546 5574 10598
rect 5626 10546 5638 10598
rect 5966 10546 6018 10558
rect 6246 10610 6298 10622
rect 8766 10666 8818 10678
rect 16314 10668 16326 10720
rect 16378 10668 16390 10720
rect 6414 10602 6466 10614
rect 6246 10546 6298 10558
rect 6906 10546 6918 10598
rect 6970 10546 6982 10598
rect 7242 10570 7254 10622
rect 7306 10570 7318 10622
rect 7758 10610 7810 10622
rect 7466 10546 7478 10598
rect 7530 10546 7542 10598
rect 17054 10666 17106 10678
rect 8766 10602 8818 10614
rect 9438 10610 9490 10622
rect 16102 10610 16154 10622
rect 7758 10546 7810 10558
rect 8990 10554 9042 10566
rect 9438 10546 9490 10558
rect 9930 10546 9942 10598
rect 9994 10546 10006 10598
rect 10602 10546 10614 10598
rect 10666 10546 10678 10598
rect 14970 10558 14982 10610
rect 15034 10558 15046 10610
rect 17054 10602 17106 10614
rect 17782 10666 17834 10678
rect 17782 10602 17834 10614
rect 19014 10666 19066 10678
rect 26014 10666 26066 10678
rect 19014 10602 19066 10614
rect 8990 10490 9042 10502
rect 12842 10474 12854 10526
rect 12906 10474 12918 10526
rect 14074 10502 14086 10554
rect 14138 10502 14150 10554
rect 14746 10502 14758 10554
rect 14810 10502 14822 10554
rect 16102 10546 16154 10558
rect 16762 10546 16774 10598
rect 16826 10546 16838 10598
rect 17434 10540 17446 10592
rect 17498 10540 17510 10592
rect 18330 10540 18342 10592
rect 18394 10540 18406 10592
rect 22026 10570 22038 10622
rect 22090 10570 22102 10622
rect 26014 10602 26066 10614
rect 26294 10666 26346 10678
rect 26294 10602 26346 10614
rect 34470 10666 34522 10678
rect 22586 10546 22598 10598
rect 22650 10546 22662 10598
rect 25722 10546 25734 10598
rect 25786 10546 25798 10598
rect 26966 10554 27018 10566
rect 29306 10546 29318 10598
rect 29370 10546 29382 10598
rect 29754 10546 29766 10598
rect 29818 10546 29830 10598
rect 30986 10546 30998 10598
rect 31050 10546 31062 10598
rect 31378 10558 31390 10610
rect 31442 10558 31454 10610
rect 34470 10602 34522 10614
rect 4790 10442 4842 10454
rect 4790 10378 4842 10390
rect 5070 10442 5122 10454
rect 5070 10378 5122 10390
rect 5182 10442 5234 10454
rect 18006 10442 18058 10454
rect 22822 10442 22874 10454
rect 24994 10446 25006 10498
rect 25058 10446 25070 10498
rect 26966 10490 27018 10502
rect 5182 10378 5234 10390
rect 5742 10386 5794 10398
rect 8094 10386 8146 10398
rect 5742 10322 5794 10334
rect 7242 10308 7254 10360
rect 7306 10308 7318 10360
rect 8094 10322 8146 10334
rect 8318 10386 8370 10398
rect 9146 10390 9158 10442
rect 9210 10390 9222 10442
rect 15754 10390 15766 10442
rect 15818 10390 15830 10442
rect 8318 10322 8370 10334
rect 16382 10386 16434 10398
rect 16382 10322 16434 10334
rect 16606 10386 16658 10398
rect 19674 10390 19686 10442
rect 19738 10390 19750 10442
rect 18006 10378 18058 10390
rect 22822 10378 22874 10390
rect 30158 10442 30210 10454
rect 30158 10378 30210 10390
rect 30270 10442 30322 10454
rect 33786 10390 33798 10442
rect 33850 10390 33862 10442
rect 30270 10378 30322 10390
rect 16606 10322 16658 10334
rect 672 10218 34832 10252
rect 672 10166 9094 10218
rect 9146 10166 9198 10218
rect 9250 10166 9302 10218
rect 9354 10166 17646 10218
rect 17698 10166 17750 10218
rect 17802 10166 17854 10218
rect 17906 10166 26198 10218
rect 26250 10166 26302 10218
rect 26354 10166 26406 10218
rect 26458 10166 34832 10218
rect 672 10132 34832 10166
rect 5406 10050 5458 10062
rect 7534 10050 7586 10062
rect 5406 9986 5458 9998
rect 7086 9994 7138 10006
rect 6234 9942 6246 9994
rect 6298 9942 6310 9994
rect 14522 10024 14534 10076
rect 14586 10024 14598 10076
rect 20682 10024 20694 10076
rect 20746 10024 20758 10076
rect 7534 9986 7586 9998
rect 7646 9994 7698 10006
rect 7086 9930 7138 9942
rect 7646 9930 7698 9942
rect 8542 9994 8594 10006
rect 8542 9930 8594 9942
rect 8878 9994 8930 10006
rect 10558 9994 10610 10006
rect 16102 9994 16154 10006
rect 19742 9994 19794 10006
rect 9762 9942 9774 9994
rect 9826 9942 9838 9994
rect 11162 9942 11174 9994
rect 11226 9942 11238 9994
rect 13514 9942 13526 9994
rect 13578 9942 13590 9994
rect 19450 9942 19462 9994
rect 19514 9942 19526 9994
rect 8878 9930 8930 9942
rect 10558 9930 10610 9942
rect 16102 9930 16154 9942
rect 19742 9930 19794 9942
rect 20078 9994 20130 10006
rect 22430 9994 22482 10006
rect 21690 9942 21702 9994
rect 21754 9942 21766 9994
rect 24378 9967 24390 10019
rect 24442 9967 24454 10019
rect 25946 9967 25958 10019
rect 26010 9967 26022 10019
rect 26518 9994 26570 10006
rect 20078 9930 20130 9942
rect 22430 9930 22482 9942
rect 26518 9930 26570 9942
rect 28534 9994 28586 10006
rect 28534 9930 28586 9942
rect 32958 9994 33010 10006
rect 32958 9930 33010 9942
rect 33182 9994 33234 10006
rect 33182 9930 33234 9942
rect 3894 9882 3946 9894
rect 5182 9882 5234 9894
rect 1082 9786 1094 9838
rect 1146 9786 1158 9838
rect 1530 9786 1542 9838
rect 1594 9786 1606 9838
rect 4778 9830 4790 9882
rect 4842 9830 4854 9882
rect 6638 9882 6690 9894
rect 3894 9818 3946 9830
rect 5182 9818 5234 9830
rect 6458 9790 6470 9842
rect 6522 9790 6534 9842
rect 6638 9818 6690 9830
rect 6974 9882 7026 9894
rect 6974 9818 7026 9830
rect 7758 9882 7810 9894
rect 10110 9882 10162 9894
rect 8698 9830 8710 9882
rect 8762 9830 8774 9882
rect 9202 9830 9214 9882
rect 9266 9830 9278 9882
rect 13694 9882 13746 9894
rect 17558 9882 17610 9894
rect 7758 9818 7810 9830
rect 4566 9770 4618 9782
rect 4566 9706 4618 9718
rect 5854 9770 5906 9782
rect 5854 9706 5906 9718
rect 7086 9770 7138 9782
rect 7914 9768 7926 9820
rect 7978 9768 7990 9820
rect 8250 9774 8262 9826
rect 8314 9774 8326 9826
rect 10110 9818 10162 9830
rect 10334 9826 10386 9838
rect 11454 9826 11506 9838
rect 10334 9762 10386 9774
rect 10714 9754 10726 9806
rect 10778 9754 10790 9806
rect 11230 9770 11282 9782
rect 7086 9706 7138 9718
rect 11454 9762 11506 9774
rect 11734 9823 11786 9835
rect 12170 9792 12182 9844
rect 12234 9792 12246 9844
rect 13246 9826 13298 9838
rect 11734 9759 11786 9771
rect 13694 9818 13746 9830
rect 14298 9786 14310 9838
rect 14362 9786 14374 9838
rect 13246 9762 13298 9774
rect 14634 9762 14646 9814
rect 14698 9762 14710 9814
rect 14858 9786 14870 9838
rect 14922 9786 14934 9838
rect 15474 9830 15486 9882
rect 15538 9830 15550 9882
rect 16370 9830 16382 9882
rect 16434 9830 16446 9882
rect 17558 9818 17610 9830
rect 17838 9882 17890 9894
rect 17838 9818 17890 9830
rect 18062 9882 18114 9894
rect 20974 9882 21026 9894
rect 18442 9830 18454 9882
rect 18506 9830 18518 9882
rect 19898 9830 19910 9882
rect 19962 9830 19974 9882
rect 18062 9818 18114 9830
rect 16942 9770 16994 9782
rect 11230 9706 11282 9718
rect 16942 9706 16994 9718
rect 17166 9770 17218 9782
rect 18778 9774 18790 9826
rect 18842 9774 18854 9826
rect 20974 9818 21026 9830
rect 21366 9882 21418 9894
rect 27918 9882 27970 9894
rect 21366 9818 21418 9830
rect 22206 9826 22258 9838
rect 22810 9830 22822 9882
rect 22874 9830 22886 9882
rect 20346 9762 20358 9814
rect 20410 9762 20422 9814
rect 20682 9762 20694 9814
rect 20746 9762 20758 9814
rect 22206 9762 22258 9774
rect 22990 9770 23042 9782
rect 23706 9774 23718 9826
rect 23770 9774 23782 9826
rect 25274 9774 25286 9826
rect 25338 9774 25350 9826
rect 26394 9803 26406 9855
rect 26458 9803 26470 9855
rect 27022 9826 27074 9838
rect 26574 9770 26626 9782
rect 17166 9706 17218 9718
rect 23482 9718 23494 9770
rect 23546 9718 23558 9770
rect 25050 9718 25062 9770
rect 25114 9718 25126 9770
rect 27694 9826 27746 9838
rect 27022 9762 27074 9774
rect 27470 9770 27522 9782
rect 22990 9706 23042 9718
rect 26574 9706 26626 9718
rect 27918 9818 27970 9830
rect 28198 9882 28250 9894
rect 33686 9882 33738 9894
rect 28198 9818 28250 9830
rect 29430 9826 29482 9838
rect 27694 9762 27746 9774
rect 33686 9818 33738 9830
rect 29430 9762 29482 9774
rect 31770 9762 31782 9814
rect 31834 9762 31846 9814
rect 32330 9766 32342 9818
rect 32394 9766 32406 9818
rect 27470 9706 27522 9718
rect 6078 9658 6130 9670
rect 5114 9606 5126 9658
rect 5178 9606 5190 9658
rect 6078 9594 6130 9606
rect 9438 9658 9490 9670
rect 12518 9658 12570 9670
rect 10042 9606 10054 9658
rect 10106 9606 10118 9658
rect 9438 9594 9490 9606
rect 12518 9594 12570 9606
rect 13134 9658 13186 9670
rect 13134 9594 13186 9606
rect 13918 9658 13970 9670
rect 15710 9658 15762 9670
rect 15250 9606 15262 9658
rect 15314 9606 15326 9658
rect 13918 9594 13970 9606
rect 15710 9594 15762 9606
rect 16718 9658 16770 9670
rect 32566 9658 32618 9670
rect 17770 9606 17782 9658
rect 17834 9606 17846 9658
rect 22362 9606 22374 9658
rect 22426 9606 22438 9658
rect 16718 9594 16770 9606
rect 26798 9602 26850 9614
rect 27962 9606 27974 9658
rect 28026 9606 28038 9658
rect 32566 9594 32618 9606
rect 34470 9658 34522 9670
rect 34470 9594 34522 9606
rect 26798 9538 26850 9550
rect 672 9434 34832 9468
rect 672 9382 4818 9434
rect 4870 9382 4922 9434
rect 4974 9382 5026 9434
rect 5078 9382 13370 9434
rect 13422 9382 13474 9434
rect 13526 9382 13578 9434
rect 13630 9382 21922 9434
rect 21974 9382 22026 9434
rect 22078 9382 22130 9434
rect 22182 9382 30474 9434
rect 30526 9382 30578 9434
rect 30630 9382 30682 9434
rect 30734 9382 34832 9434
rect 672 9348 34832 9382
rect 18286 9266 18338 9278
rect 5854 9210 5906 9222
rect 3994 9158 4006 9210
rect 4058 9158 4070 9210
rect 5854 9146 5906 9158
rect 6190 9210 6242 9222
rect 6190 9146 6242 9158
rect 7254 9210 7306 9222
rect 7254 9146 7306 9158
rect 7478 9210 7530 9222
rect 7478 9146 7530 9158
rect 7702 9210 7754 9222
rect 11566 9210 11618 9222
rect 10546 9158 10558 9210
rect 10610 9158 10622 9210
rect 12238 9210 12290 9222
rect 7702 9146 7754 9158
rect 1486 9098 1538 9110
rect 1486 9034 1538 9046
rect 1710 9098 1762 9110
rect 1710 9034 1762 9046
rect 1934 9098 1986 9110
rect 4846 9098 4898 9110
rect 1934 9034 1986 9046
rect 2494 9042 2546 9054
rect 2650 9046 2662 9098
rect 2714 9046 2726 9098
rect 3782 9042 3834 9054
rect 2494 8978 2546 8990
rect 3322 8972 3334 9024
rect 3386 8972 3398 9024
rect 6526 9098 6578 9110
rect 4846 9034 4898 9046
rect 3782 8978 3834 8990
rect 4958 8986 5010 8998
rect 5114 8996 5126 9048
rect 5178 8996 5190 9048
rect 5338 8990 5350 9042
rect 5402 8990 5414 9042
rect 6526 9034 6578 9046
rect 6974 9098 7026 9110
rect 9034 9102 9046 9154
rect 9098 9102 9110 9154
rect 11274 9096 11286 9148
rect 11338 9096 11350 9148
rect 11566 9146 11618 9158
rect 11946 9108 11958 9160
rect 12010 9108 12022 9160
rect 12238 9146 12290 9158
rect 12910 9210 12962 9222
rect 12910 9146 12962 9158
rect 13134 9210 13186 9222
rect 13134 9146 13186 9158
rect 15094 9210 15146 9222
rect 17098 9158 17110 9210
rect 17162 9158 17174 9210
rect 18286 9202 18338 9214
rect 20974 9266 21026 9278
rect 20974 9202 21026 9214
rect 22094 9210 22146 9222
rect 15094 9146 15146 9158
rect 18062 9154 18114 9166
rect 12686 9098 12738 9110
rect 6974 9034 7026 9046
rect 9662 9042 9714 9054
rect 19898 9102 19910 9154
rect 19962 9102 19974 9154
rect 21354 9112 21366 9164
rect 21418 9112 21430 9164
rect 22094 9146 22146 9158
rect 22430 9210 22482 9222
rect 22430 9146 22482 9158
rect 26630 9210 26682 9222
rect 26630 9146 26682 9158
rect 26854 9210 26906 9222
rect 26854 9146 26906 9158
rect 30886 9210 30938 9222
rect 30886 9146 30938 9158
rect 18062 9090 18114 9102
rect 2650 8912 2662 8964
rect 2714 8912 2726 8964
rect 4398 8930 4450 8942
rect 1374 8874 1426 8886
rect 1374 8810 1426 8822
rect 2270 8874 2322 8886
rect 2270 8810 2322 8822
rect 2998 8874 3050 8886
rect 2998 8810 3050 8822
rect 3950 8874 4002 8886
rect 5898 8982 5910 9034
rect 5962 8982 5974 9034
rect 10154 8990 10166 9042
rect 10218 8990 10230 9042
rect 8586 8934 8598 8986
rect 8650 8934 8662 8986
rect 9662 8978 9714 8990
rect 10490 8984 10502 9036
rect 10554 8984 10566 9036
rect 11162 8990 11174 9042
rect 11226 8990 11238 9042
rect 12686 9034 12738 9046
rect 12014 8986 12066 8998
rect 13738 8978 13750 9030
rect 13802 8978 13814 9030
rect 14074 8978 14086 9030
rect 14138 8978 14150 9030
rect 14298 9002 14310 9054
rect 14362 9002 14374 9054
rect 15418 9002 15430 9054
rect 15482 9002 15494 9054
rect 16090 9002 16102 9054
rect 16154 9002 16166 9054
rect 16314 9002 16326 9054
rect 16378 9002 16390 9054
rect 17782 9042 17834 9054
rect 16650 8978 16662 9030
rect 16714 8978 16726 9030
rect 16942 8986 16994 8998
rect 4958 8922 5010 8934
rect 12014 8922 12066 8934
rect 16942 8922 16994 8934
rect 17166 8986 17218 8998
rect 17166 8922 17218 8934
rect 17446 8986 17498 8998
rect 19562 8990 19574 9042
rect 19626 8990 19638 9042
rect 17782 8978 17834 8990
rect 20738 8934 20750 8986
rect 20802 8934 20814 8986
rect 21242 8970 21254 9022
rect 21306 8970 21318 9022
rect 21422 8986 21474 8998
rect 22138 8982 22150 9034
rect 22202 8982 22214 9034
rect 23034 9002 23046 9054
rect 23098 9002 23110 9054
rect 23594 8978 23606 9030
rect 23658 8978 23670 9030
rect 25958 8986 26010 8998
rect 17446 8922 17498 8934
rect 21422 8922 21474 8934
rect 29866 8978 29878 9030
rect 29930 8978 29942 9030
rect 30314 9002 30326 9054
rect 30378 9002 30390 9054
rect 33954 8990 33966 9042
rect 34018 8990 34030 9042
rect 34346 9002 34358 9054
rect 34410 9002 34422 9054
rect 25958 8922 26010 8934
rect 4398 8866 4450 8878
rect 8038 8874 8090 8886
rect 3950 8810 4002 8822
rect 4174 8818 4226 8830
rect 4174 8754 4226 8766
rect 4734 8818 4786 8830
rect 8038 8810 8090 8822
rect 8206 8874 8258 8886
rect 8206 8810 8258 8822
rect 8430 8874 8482 8886
rect 8430 8810 8482 8822
rect 8766 8874 8818 8886
rect 8766 8810 8818 8822
rect 9102 8874 9154 8886
rect 9102 8810 9154 8822
rect 9326 8874 9378 8886
rect 9326 8810 9378 8822
rect 9774 8874 9826 8886
rect 13526 8874 13578 8886
rect 9774 8810 9826 8822
rect 10670 8818 10722 8830
rect 4734 8754 4786 8766
rect 10670 8754 10722 8766
rect 10894 8818 10946 8830
rect 13526 8810 13578 8822
rect 14702 8874 14754 8886
rect 14702 8810 14754 8822
rect 15766 8874 15818 8886
rect 18846 8874 18898 8886
rect 21646 8874 21698 8886
rect 18330 8822 18342 8874
rect 18394 8822 18406 8874
rect 20234 8822 20246 8874
rect 20298 8822 20310 8874
rect 15766 8810 15818 8822
rect 10894 8754 10946 8766
rect 13962 8740 13974 8792
rect 14026 8740 14038 8792
rect 16426 8766 16438 8818
rect 16490 8766 16502 8818
rect 18846 8810 18898 8822
rect 21646 8810 21698 8822
rect 22654 8874 22706 8886
rect 27514 8822 27526 8874
rect 27578 8822 27590 8874
rect 31546 8822 31558 8874
rect 31610 8822 31622 8874
rect 22654 8810 22706 8822
rect 672 8650 34832 8684
rect 672 8598 9094 8650
rect 9146 8598 9198 8650
rect 9250 8598 9302 8650
rect 9354 8598 17646 8650
rect 17698 8598 17750 8650
rect 17802 8598 17854 8650
rect 17906 8598 26198 8650
rect 26250 8598 26302 8650
rect 26354 8598 26406 8650
rect 26458 8598 34832 8650
rect 672 8564 34832 8598
rect 14030 8482 14082 8494
rect 31782 8482 31834 8494
rect 10782 8426 10834 8438
rect 1642 8374 1654 8426
rect 1706 8374 1718 8426
rect 5406 8370 5458 8382
rect 14030 8418 14082 8430
rect 19910 8426 19962 8438
rect 21018 8430 21030 8482
rect 21082 8430 21094 8482
rect 10782 8362 10834 8374
rect 19910 8362 19962 8374
rect 24502 8426 24554 8438
rect 25386 8430 25398 8482
rect 25450 8430 25462 8482
rect 26394 8374 26406 8426
rect 26458 8374 26470 8426
rect 30202 8374 30214 8426
rect 30266 8374 30278 8426
rect 31782 8418 31834 8430
rect 34022 8426 34074 8438
rect 24502 8362 24554 8374
rect 34022 8362 34074 8374
rect 5406 8306 5458 8318
rect 6862 8314 6914 8326
rect 3994 8218 4006 8270
rect 4058 8218 4070 8270
rect 7466 8284 7478 8336
rect 7530 8284 7542 8336
rect 8026 8284 8038 8336
rect 8090 8284 8102 8336
rect 8430 8314 8482 8326
rect 6862 8250 6914 8262
rect 7310 8258 7362 8270
rect 982 8202 1034 8214
rect 4554 8194 4566 8246
rect 4618 8194 4630 8246
rect 6010 8194 6022 8246
rect 6074 8194 6086 8246
rect 6302 8202 6354 8214
rect 982 8138 1034 8150
rect 6302 8138 6354 8150
rect 6526 8202 6578 8214
rect 6526 8138 6578 8150
rect 6974 8202 7026 8214
rect 7310 8194 7362 8206
rect 7870 8258 7922 8270
rect 9214 8314 9266 8326
rect 8430 8250 8482 8262
rect 8698 8206 8710 8258
rect 8762 8206 8774 8258
rect 9034 8212 9046 8264
rect 9098 8212 9110 8264
rect 9998 8314 10050 8326
rect 11342 8314 11394 8326
rect 11902 8314 11954 8326
rect 9214 8250 9266 8262
rect 9438 8258 9490 8270
rect 7466 8150 7478 8202
rect 7530 8150 7542 8202
rect 7870 8194 7922 8206
rect 8026 8150 8038 8202
rect 8090 8150 8102 8202
rect 9438 8194 9490 8206
rect 9774 8258 9826 8270
rect 10938 8262 10950 8314
rect 11002 8262 11014 8314
rect 9998 8250 10050 8262
rect 11118 8258 11170 8270
rect 10210 8206 10222 8258
rect 10274 8206 10286 8258
rect 10378 8206 10390 8258
rect 10442 8206 10454 8258
rect 11722 8262 11734 8314
rect 11786 8262 11798 8314
rect 12394 8284 12406 8336
rect 12458 8284 12470 8336
rect 13022 8314 13074 8326
rect 13806 8314 13858 8326
rect 11342 8250 11394 8262
rect 11902 8250 11954 8262
rect 12238 8258 12290 8270
rect 9774 8194 9826 8206
rect 11118 8194 11170 8206
rect 13346 8262 13358 8314
rect 13410 8262 13422 8314
rect 13022 8250 13074 8262
rect 13806 8250 13858 8262
rect 14478 8314 14530 8326
rect 15150 8314 15202 8326
rect 21198 8314 21250 8326
rect 14478 8250 14530 8262
rect 14926 8258 14978 8270
rect 12238 8194 12290 8206
rect 12394 8150 12406 8202
rect 12458 8150 12470 8202
rect 13626 8186 13638 8238
rect 13690 8186 13702 8238
rect 13918 8202 13970 8214
rect 15530 8262 15542 8314
rect 15594 8262 15606 8314
rect 15150 8250 15202 8262
rect 14926 8194 14978 8206
rect 15822 8202 15874 8214
rect 6974 8138 7026 8150
rect 13918 8138 13970 8150
rect 16090 8198 16102 8250
rect 16154 8198 16166 8250
rect 16594 8206 16606 8258
rect 16658 8206 16670 8258
rect 18890 8194 18902 8246
rect 18954 8194 18966 8246
rect 20078 8202 20130 8214
rect 15822 8138 15874 8150
rect 20570 8194 20582 8246
rect 20634 8194 20646 8246
rect 20906 8218 20918 8270
rect 20970 8218 20982 8270
rect 26798 8314 26850 8326
rect 21198 8250 21250 8262
rect 20750 8202 20802 8214
rect 20078 8138 20130 8150
rect 21578 8194 21590 8246
rect 21642 8194 21654 8246
rect 25050 8218 25062 8270
rect 25114 8218 25126 8270
rect 33350 8314 33402 8326
rect 26798 8250 26850 8262
rect 25274 8194 25286 8246
rect 25338 8194 25350 8246
rect 25610 8194 25622 8246
rect 25674 8194 25686 8246
rect 26618 8194 26630 8246
rect 26682 8194 26694 8246
rect 27022 8202 27074 8214
rect 20750 8138 20802 8150
rect 27290 8194 27302 8246
rect 27354 8194 27366 8246
rect 27850 8218 27862 8270
rect 27914 8218 27926 8270
rect 31434 8206 31446 8258
rect 31498 8206 31510 8258
rect 32554 8224 32566 8276
rect 32618 8224 32630 8276
rect 33350 8250 33402 8262
rect 32902 8202 32954 8214
rect 31210 8150 31222 8202
rect 31274 8150 31286 8202
rect 5686 8090 5738 8102
rect 4778 8038 4790 8090
rect 4842 8038 4854 8090
rect 5182 8034 5234 8046
rect 9090 8038 9102 8090
rect 9154 8038 9166 8090
rect 10042 8084 10054 8136
rect 10106 8084 10118 8136
rect 11790 8090 11842 8102
rect 5686 8026 5738 8038
rect 11790 8026 11842 8038
rect 14590 8090 14642 8102
rect 22306 8094 22318 8146
rect 22370 8094 22382 8146
rect 27022 8138 27074 8150
rect 32902 8138 32954 8150
rect 33070 8202 33122 8214
rect 33674 8194 33686 8246
rect 33738 8194 33750 8246
rect 34346 8194 34358 8246
rect 34410 8194 34422 8246
rect 33070 8138 33122 8150
rect 26014 8090 26066 8102
rect 15082 8038 15094 8090
rect 15146 8038 15158 8090
rect 14590 8026 14642 8038
rect 26014 8026 26066 8038
rect 26238 8090 26290 8102
rect 26238 8026 26290 8038
rect 30886 8090 30938 8102
rect 30886 8026 30938 8038
rect 5182 7970 5234 7982
rect 672 7866 34832 7900
rect 672 7814 4818 7866
rect 4870 7814 4922 7866
rect 4974 7814 5026 7866
rect 5078 7814 13370 7866
rect 13422 7814 13474 7866
rect 13526 7814 13578 7866
rect 13630 7814 21922 7866
rect 21974 7814 22026 7866
rect 22078 7814 22130 7866
rect 22182 7814 30474 7866
rect 30526 7814 30578 7866
rect 30630 7814 30682 7866
rect 30734 7814 34832 7866
rect 672 7780 34832 7814
rect 7870 7698 7922 7710
rect 6134 7642 6186 7654
rect 6134 7578 6186 7590
rect 7534 7642 7586 7654
rect 7870 7634 7922 7646
rect 10334 7642 10386 7654
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 7534 7578 7586 7590
rect 10334 7578 10386 7590
rect 11342 7642 11394 7654
rect 11342 7578 11394 7590
rect 11454 7642 11506 7654
rect 11454 7578 11506 7590
rect 11846 7642 11898 7654
rect 11846 7578 11898 7590
rect 18510 7642 18562 7654
rect 9438 7530 9490 7542
rect 13582 7530 13634 7542
rect 14186 7534 14198 7586
rect 14250 7534 14262 7586
rect 18510 7578 18562 7590
rect 29990 7642 30042 7654
rect 2650 7410 2662 7462
rect 2714 7410 2726 7462
rect 3098 7434 3110 7486
rect 3162 7434 3174 7486
rect 9438 7466 9490 7478
rect 8262 7418 8314 7430
rect 9662 7418 9714 7430
rect 8262 7354 8314 7366
rect 8586 7320 8598 7372
rect 8650 7320 8662 7372
rect 9662 7354 9714 7366
rect 9998 7418 10050 7430
rect 10378 7422 10390 7474
rect 10442 7422 10454 7474
rect 10938 7434 10950 7486
rect 11002 7434 11014 7486
rect 12618 7478 12630 7530
rect 12682 7478 12694 7530
rect 22710 7530 22762 7542
rect 27794 7534 27806 7586
rect 27858 7534 27870 7586
rect 29990 7578 30042 7590
rect 30886 7642 30938 7654
rect 30886 7578 30938 7590
rect 9998 7354 10050 7366
rect 12238 7418 12290 7430
rect 12842 7422 12854 7474
rect 12906 7422 12918 7474
rect 13582 7466 13634 7478
rect 12238 7354 12290 7366
rect 13918 7418 13970 7430
rect 14354 7422 14366 7474
rect 14418 7422 14430 7474
rect 14634 7410 14646 7462
rect 14698 7410 14710 7462
rect 15306 7434 15318 7486
rect 15370 7434 15382 7486
rect 18834 7422 18846 7474
rect 18898 7422 18910 7474
rect 19506 7422 19518 7474
rect 19570 7422 19582 7474
rect 22710 7466 22762 7478
rect 21690 7410 21702 7462
rect 21754 7410 21766 7462
rect 23034 7409 23046 7461
rect 23098 7409 23110 7461
rect 23482 7410 23494 7462
rect 23546 7410 23558 7462
rect 25722 7434 25734 7486
rect 25786 7434 25798 7486
rect 27066 7410 27078 7462
rect 27130 7410 27142 7462
rect 30270 7418 30322 7430
rect 13918 7354 13970 7366
rect 17546 7338 17558 7390
rect 17610 7338 17622 7390
rect 33898 7410 33910 7462
rect 33962 7410 33974 7462
rect 34458 7410 34470 7462
rect 34522 7410 34534 7462
rect 30270 7354 30322 7366
rect 6414 7306 6466 7318
rect 5450 7254 5462 7306
rect 5514 7254 5526 7306
rect 6414 7242 6466 7254
rect 6862 7306 6914 7318
rect 6862 7242 6914 7254
rect 7086 7306 7138 7318
rect 7086 7242 7138 7254
rect 10614 7306 10666 7318
rect 26742 7306 26794 7318
rect 10614 7242 10666 7254
rect 14142 7250 14194 7262
rect 26742 7242 26794 7254
rect 30382 7306 30434 7318
rect 31546 7254 31558 7306
rect 31610 7254 31622 7306
rect 30382 7242 30434 7254
rect 14142 7186 14194 7198
rect 672 7082 34832 7116
rect 672 7030 9094 7082
rect 9146 7030 9198 7082
rect 9250 7030 9302 7082
rect 9354 7030 17646 7082
rect 17698 7030 17750 7082
rect 17802 7030 17854 7082
rect 17906 7030 26198 7082
rect 26250 7030 26302 7082
rect 26354 7030 26406 7082
rect 26458 7030 34832 7082
rect 672 6996 34832 7030
rect 3502 6858 3554 6870
rect 3502 6794 3554 6806
rect 4174 6858 4226 6870
rect 4174 6794 4226 6806
rect 12238 6858 12290 6870
rect 12238 6794 12290 6806
rect 13246 6858 13298 6870
rect 13246 6794 13298 6806
rect 13582 6858 13634 6870
rect 13582 6794 13634 6806
rect 14870 6858 14922 6870
rect 16202 6862 16214 6914
rect 16266 6862 16278 6914
rect 14870 6794 14922 6806
rect 18846 6858 18898 6870
rect 18846 6794 18898 6806
rect 19294 6858 19346 6870
rect 19294 6794 19346 6806
rect 20526 6858 20578 6870
rect 20906 6831 20918 6883
rect 20970 6831 20982 6883
rect 23930 6831 23942 6883
rect 23994 6831 24006 6883
rect 32958 6858 33010 6870
rect 25610 6806 25622 6858
rect 25674 6806 25686 6858
rect 20526 6794 20578 6806
rect 32958 6794 33010 6806
rect 7354 6722 7366 6774
rect 7418 6722 7430 6774
rect 11398 6746 11450 6758
rect 13806 6746 13858 6758
rect 2090 6626 2102 6678
rect 2154 6626 2166 6678
rect 4554 6650 4566 6702
rect 4618 6650 4630 6702
rect 13066 6694 13078 6746
rect 13130 6694 13142 6746
rect 3278 6634 3330 6646
rect 3278 6570 3330 6582
rect 3726 6634 3778 6646
rect 3726 6570 3778 6582
rect 3950 6634 4002 6646
rect 5170 6638 5182 6690
rect 5234 6638 5246 6690
rect 11398 6682 11450 6694
rect 13806 6682 13858 6694
rect 14086 6746 14138 6758
rect 20134 6746 20186 6758
rect 15474 6694 15486 6746
rect 15538 6694 15550 6746
rect 15698 6694 15710 6746
rect 15762 6694 15774 6746
rect 14086 6682 14138 6694
rect 3950 6570 4002 6582
rect 8318 6634 8370 6646
rect 8474 6626 8486 6678
rect 8538 6626 8550 6678
rect 9034 6626 9046 6678
rect 9098 6626 9110 6678
rect 12574 6634 12626 6646
rect 8318 6570 8370 6582
rect 12574 6570 12626 6582
rect 14366 6634 14418 6646
rect 14366 6570 14418 6582
rect 14590 6634 14642 6646
rect 14590 6570 14642 6582
rect 15262 6634 15314 6646
rect 15978 6626 15990 6678
rect 16042 6626 16054 6678
rect 16314 6626 16326 6678
rect 16378 6626 16390 6678
rect 16538 6626 16550 6678
rect 16602 6626 16614 6678
rect 17210 6656 17222 6708
rect 17274 6656 17286 6708
rect 20134 6682 20186 6694
rect 16886 6634 16938 6646
rect 15262 6570 15314 6582
rect 16886 6570 16938 6582
rect 17502 6634 17554 6646
rect 17502 6570 17554 6582
rect 17726 6634 17778 6646
rect 17726 6570 17778 6582
rect 18398 6634 18450 6646
rect 18398 6570 18450 6582
rect 18622 6634 18674 6646
rect 18622 6570 18674 6582
rect 19406 6634 19458 6646
rect 19406 6570 19458 6582
rect 19742 6634 19794 6646
rect 21354 6638 21366 6690
rect 21418 6638 21430 6690
rect 22094 6634 22146 6646
rect 21802 6582 21814 6634
rect 21866 6582 21878 6634
rect 22474 6626 22486 6678
rect 22538 6626 22550 6678
rect 22822 6634 22874 6646
rect 23370 6638 23382 6690
rect 23434 6638 23446 6690
rect 24334 6634 24386 6646
rect 19742 6570 19794 6582
rect 22094 6570 22146 6582
rect 23146 6582 23158 6634
rect 23210 6582 23222 6634
rect 27962 6626 27974 6678
rect 28026 6626 28038 6678
rect 28410 6626 28422 6678
rect 28474 6626 28486 6678
rect 29866 6650 29878 6702
rect 29930 6650 29942 6702
rect 32106 6626 32118 6678
rect 32170 6626 32182 6678
rect 32554 6630 32566 6682
rect 32618 6630 32630 6682
rect 33350 6634 33402 6646
rect 22822 6570 22874 6582
rect 24334 6570 24386 6582
rect 33350 6570 33402 6582
rect 33518 6634 33570 6646
rect 33518 6570 33570 6582
rect 33742 6634 33794 6646
rect 34346 6626 34358 6678
rect 34410 6626 34422 6678
rect 33742 6570 33794 6582
rect 1766 6522 1818 6534
rect 1766 6458 1818 6470
rect 12070 6522 12122 6534
rect 12070 6458 12122 6470
rect 13134 6522 13186 6534
rect 18062 6522 18114 6534
rect 13738 6470 13750 6522
rect 13802 6470 13814 6522
rect 13134 6458 13186 6470
rect 18062 6458 18114 6470
rect 18174 6522 18226 6534
rect 18174 6458 18226 6470
rect 19854 6522 19906 6534
rect 19854 6458 19906 6470
rect 24950 6522 25002 6534
rect 34022 6522 34074 6534
rect 28858 6470 28870 6522
rect 28922 6470 28934 6522
rect 24950 6458 25002 6470
rect 34022 6458 34074 6470
rect 672 6298 34832 6332
rect 672 6246 4818 6298
rect 4870 6246 4922 6298
rect 4974 6246 5026 6298
rect 5078 6246 13370 6298
rect 13422 6246 13474 6298
rect 13526 6246 13578 6298
rect 13630 6246 21922 6298
rect 21974 6246 22026 6298
rect 22078 6246 22130 6298
rect 22182 6246 30474 6298
rect 30526 6246 30578 6298
rect 30630 6246 30682 6298
rect 30734 6246 34832 6298
rect 672 6212 34832 6246
rect 24558 6130 24610 6142
rect 7758 6074 7810 6086
rect 6234 5966 6246 6018
rect 6298 5966 6310 6018
rect 7758 6010 7810 6022
rect 13414 6074 13466 6086
rect 13962 6022 13974 6074
rect 14026 6022 14038 6074
rect 18442 6022 18454 6074
rect 18506 6022 18518 6074
rect 24558 6066 24610 6078
rect 24782 6130 24834 6142
rect 24782 6066 24834 6078
rect 25006 6130 25058 6142
rect 25006 6066 25058 6078
rect 30886 6074 30938 6086
rect 29642 6022 29654 6074
rect 29706 6022 29718 6074
rect 8698 5961 8710 6013
rect 8762 5961 8774 6013
rect 13414 6010 13466 6022
rect 30886 6010 30938 6022
rect 1082 5841 1094 5893
rect 1146 5841 1158 5893
rect 1698 5854 1710 5906
rect 1762 5854 1774 5906
rect 3882 5842 3894 5894
rect 3946 5842 3958 5894
rect 6458 5866 6470 5918
rect 6522 5866 6534 5918
rect 7130 5866 7142 5918
rect 7194 5866 7206 5918
rect 6190 5850 6242 5862
rect 6190 5786 6242 5798
rect 6974 5850 7026 5862
rect 6974 5786 7026 5798
rect 7534 5850 7586 5862
rect 8250 5854 8262 5906
rect 8314 5854 8326 5906
rect 8586 5860 8598 5912
rect 8650 5860 8662 5912
rect 9930 5866 9942 5918
rect 9994 5866 10006 5918
rect 14030 5906 14082 5918
rect 7534 5786 7586 5798
rect 9214 5850 9266 5862
rect 10434 5854 10446 5906
rect 10498 5854 10510 5906
rect 12742 5850 12794 5862
rect 9370 5798 9382 5850
rect 9434 5798 9446 5850
rect 14634 5862 14646 5914
rect 14698 5862 14710 5914
rect 14030 5842 14082 5854
rect 14410 5798 14422 5850
rect 14474 5798 14486 5850
rect 15194 5842 15206 5894
rect 15258 5842 15270 5894
rect 17434 5866 17446 5918
rect 17498 5866 17510 5918
rect 23818 5910 23830 5962
rect 23882 5910 23894 5962
rect 18846 5850 18898 5862
rect 9214 5786 9266 5798
rect 12742 5786 12794 5798
rect 18846 5786 18898 5798
rect 19182 5850 19234 5862
rect 19450 5846 19462 5898
rect 19514 5846 19526 5898
rect 19898 5842 19910 5894
rect 19962 5842 19974 5894
rect 22822 5850 22874 5862
rect 23370 5854 23382 5906
rect 23434 5854 23446 5906
rect 25162 5875 25174 5927
rect 25226 5875 25238 5927
rect 25834 5862 25846 5914
rect 25898 5862 25910 5914
rect 19182 5786 19234 5798
rect 26394 5842 26406 5894
rect 26458 5842 26470 5894
rect 28634 5866 28646 5918
rect 28698 5866 28710 5918
rect 33954 5854 33966 5906
rect 34018 5854 34030 5906
rect 34346 5842 34358 5894
rect 34410 5842 34422 5894
rect 4902 5738 4954 5750
rect 4902 5674 4954 5686
rect 5182 5738 5234 5750
rect 5182 5674 5234 5686
rect 5574 5738 5626 5750
rect 8766 5738 8818 5750
rect 5574 5674 5626 5686
rect 5966 5682 6018 5694
rect 7354 5686 7366 5738
rect 7418 5686 7430 5738
rect 9550 5738 9602 5750
rect 8766 5674 8818 5686
rect 8990 5682 9042 5694
rect 5966 5618 6018 5630
rect 19294 5738 19346 5750
rect 20626 5742 20638 5794
rect 20690 5742 20702 5794
rect 22822 5786 22874 5798
rect 9550 5674 9602 5686
rect 13806 5682 13858 5694
rect 8990 5618 9042 5630
rect 24614 5738 24666 5750
rect 19294 5674 19346 5686
rect 23718 5678 23770 5690
rect 13806 5618 13858 5630
rect 24614 5674 24666 5686
rect 25454 5738 25506 5750
rect 25454 5674 25506 5686
rect 29878 5738 29930 5750
rect 29878 5674 29930 5686
rect 30214 5738 30266 5750
rect 31546 5686 31558 5738
rect 31610 5686 31622 5738
rect 30214 5674 30266 5686
rect 23718 5614 23770 5626
rect 672 5514 34832 5548
rect 672 5462 9094 5514
rect 9146 5462 9198 5514
rect 9250 5462 9302 5514
rect 9354 5462 17646 5514
rect 17698 5462 17750 5514
rect 17802 5462 17854 5514
rect 17906 5462 26198 5514
rect 26250 5462 26302 5514
rect 26354 5462 26406 5514
rect 26458 5462 34832 5514
rect 672 5428 34832 5462
rect 6078 5346 6130 5358
rect 4846 5290 4898 5302
rect 3882 5238 3894 5290
rect 3946 5238 3958 5290
rect 6078 5282 6130 5294
rect 6862 5346 6914 5358
rect 6862 5282 6914 5294
rect 7870 5346 7922 5358
rect 10110 5346 10162 5358
rect 7870 5282 7922 5294
rect 9886 5290 9938 5302
rect 4846 5226 4898 5238
rect 8318 5234 8370 5246
rect 5182 5178 5234 5190
rect 5182 5114 5234 5126
rect 5854 5178 5906 5190
rect 5854 5114 5906 5126
rect 7086 5178 7138 5190
rect 19518 5346 19570 5358
rect 10110 5282 10162 5294
rect 10894 5290 10946 5302
rect 9886 5226 9938 5238
rect 10894 5226 10946 5238
rect 12182 5290 12234 5302
rect 18666 5263 18678 5315
rect 18730 5263 18742 5315
rect 19518 5282 19570 5294
rect 19742 5346 19794 5358
rect 25498 5320 25510 5372
rect 25562 5320 25574 5372
rect 19742 5282 19794 5294
rect 23830 5290 23882 5302
rect 12182 5226 12234 5238
rect 8318 5170 8370 5182
rect 8654 5178 8706 5190
rect 9998 5178 10050 5190
rect 16594 5182 16606 5234
rect 16658 5182 16670 5234
rect 23830 5226 23882 5238
rect 26966 5290 27018 5302
rect 33462 5290 33514 5302
rect 29306 5238 29318 5290
rect 29370 5238 29382 5290
rect 26966 5226 27018 5238
rect 33462 5226 33514 5238
rect 34078 5290 34130 5302
rect 34078 5226 34130 5238
rect 34302 5290 34354 5302
rect 34302 5226 34354 5238
rect 27862 5178 27914 5190
rect 7086 5114 7138 5126
rect 7366 5122 7418 5134
rect 1082 5058 1094 5110
rect 1146 5058 1158 5110
rect 1530 5058 1542 5110
rect 1594 5058 1606 5110
rect 5450 5062 5462 5114
rect 5514 5062 5526 5114
rect 6346 5058 6358 5110
rect 6410 5058 6422 5110
rect 6682 5058 6694 5110
rect 6746 5058 6758 5110
rect 7366 5058 7418 5070
rect 7702 5122 7754 5134
rect 7702 5058 7754 5070
rect 8094 5122 8146 5134
rect 8654 5114 8706 5126
rect 8878 5122 8930 5134
rect 9258 5126 9270 5178
rect 9322 5126 9334 5178
rect 11050 5126 11062 5178
rect 11114 5126 11126 5178
rect 8094 5058 8146 5070
rect 8766 5066 8818 5078
rect 4566 4954 4618 4966
rect 5338 4964 5350 5016
rect 5402 4964 5414 5016
rect 9998 5114 10050 5126
rect 11230 5122 11282 5134
rect 8878 5058 8930 5070
rect 9550 5066 9602 5078
rect 5786 4958 5798 5010
rect 5850 4958 5862 5010
rect 8766 5002 8818 5014
rect 10266 5064 10278 5116
rect 10330 5064 10342 5116
rect 10490 5070 10502 5122
rect 10554 5070 10566 5122
rect 12282 5099 12294 5151
rect 12346 5099 12358 5151
rect 13066 5088 13078 5140
rect 13130 5088 13142 5140
rect 13626 5082 13638 5134
rect 13690 5082 13702 5134
rect 11230 5058 11282 5070
rect 12126 5066 12178 5078
rect 9550 5002 9602 5014
rect 11678 5010 11730 5022
rect 7130 4946 7142 4998
rect 7194 4946 7206 4998
rect 14298 5058 14310 5110
rect 14362 5058 14374 5110
rect 17994 5070 18006 5122
rect 18058 5070 18070 5122
rect 17770 5014 17782 5066
rect 17834 5014 17846 5066
rect 19338 5050 19350 5102
rect 19402 5050 19414 5102
rect 19630 5066 19682 5078
rect 12126 5002 12178 5014
rect 19630 5002 19682 5014
rect 20078 5066 20130 5078
rect 20402 5070 20414 5122
rect 20466 5070 20478 5122
rect 23706 5099 23718 5151
rect 23770 5099 23782 5151
rect 25162 5082 25174 5134
rect 25226 5082 25238 5134
rect 25386 5082 25398 5134
rect 25450 5082 25462 5134
rect 25722 5082 25734 5134
rect 25786 5082 25798 5134
rect 26058 5126 26070 5178
rect 26122 5126 26134 5178
rect 27862 5114 27914 5126
rect 28142 5178 28194 5190
rect 32566 5178 32618 5190
rect 28142 5114 28194 5126
rect 28366 5122 28418 5134
rect 26630 5066 26682 5078
rect 20078 5002 20130 5014
rect 23886 5010 23938 5022
rect 7802 4902 7814 4954
rect 7866 4902 7878 4954
rect 11678 4946 11730 4958
rect 11902 4954 11954 4966
rect 4566 4890 4618 4902
rect 11902 4890 11954 4902
rect 13414 4954 13466 4966
rect 13414 4890 13466 4902
rect 17502 4954 17554 4966
rect 17502 4890 17554 4902
rect 19070 4954 19122 4966
rect 21186 4958 21198 5010
rect 21250 4958 21262 5010
rect 28366 5058 28418 5070
rect 28758 5122 28810 5134
rect 29754 5082 29766 5134
rect 29818 5082 29830 5134
rect 32566 5114 32618 5126
rect 28758 5058 28810 5070
rect 30202 5058 30214 5110
rect 30266 5058 30278 5110
rect 33786 5058 33798 5110
rect 33850 5058 33862 5110
rect 26630 5002 26682 5014
rect 23258 4902 23270 4954
rect 23322 4902 23334 4954
rect 23886 4946 23938 4958
rect 24110 4954 24162 4966
rect 19070 4890 19122 4902
rect 24110 4890 24162 4902
rect 24334 4954 24386 4966
rect 24334 4890 24386 4902
rect 26406 4954 26458 4966
rect 26406 4890 26458 4902
rect 27358 4954 27410 4966
rect 27358 4890 27410 4902
rect 27470 4954 27522 4966
rect 29038 4954 29090 4966
rect 28074 4902 28086 4954
rect 28138 4902 28150 4954
rect 27470 4890 27522 4902
rect 29038 4890 29090 4902
rect 29262 4954 29314 4966
rect 29262 4890 29314 4902
rect 33238 4954 33290 4966
rect 33238 4890 33290 4902
rect 672 4730 34832 4764
rect 672 4678 4818 4730
rect 4870 4678 4922 4730
rect 4974 4678 5026 4730
rect 5078 4678 13370 4730
rect 13422 4678 13474 4730
rect 13526 4678 13578 4730
rect 13630 4678 21922 4730
rect 21974 4678 22026 4730
rect 22078 4678 22130 4730
rect 22182 4678 30474 4730
rect 30526 4678 30578 4730
rect 30630 4678 30682 4730
rect 30734 4678 34832 4730
rect 672 4644 34832 4678
rect 4790 4506 4842 4518
rect 10222 4506 10274 4518
rect 6066 4454 6078 4506
rect 6130 4454 6142 4506
rect 7354 4454 7366 4506
rect 7418 4454 7430 4506
rect 4790 4442 4842 4454
rect 9930 4404 9942 4456
rect 9994 4404 10006 4456
rect 10222 4442 10274 4454
rect 11174 4506 11226 4518
rect 11174 4442 11226 4454
rect 13022 4506 13074 4518
rect 16102 4506 16154 4518
rect 13458 4454 13470 4506
rect 13522 4454 13534 4506
rect 13738 4454 13750 4506
rect 13802 4454 13814 4506
rect 15418 4454 15430 4506
rect 15482 4454 15494 4506
rect 12170 4398 12182 4450
rect 12234 4398 12246 4450
rect 13022 4442 13074 4454
rect 16102 4442 16154 4454
rect 18286 4506 18338 4518
rect 26518 4506 26570 4518
rect 19786 4454 19798 4506
rect 19850 4454 19862 4506
rect 20682 4454 20694 4506
rect 20746 4454 20758 4506
rect 22698 4454 22710 4506
rect 22762 4454 22774 4506
rect 1194 4274 1206 4326
rect 1258 4274 1270 4326
rect 1754 4298 1766 4350
rect 1818 4298 1830 4350
rect 5226 4342 5238 4394
rect 5290 4342 5302 4394
rect 17994 4392 18006 4444
rect 18058 4392 18070 4444
rect 18286 4442 18338 4454
rect 26518 4442 26570 4454
rect 27918 4506 27970 4518
rect 27918 4442 27970 4454
rect 30886 4506 30938 4518
rect 18846 4394 18898 4406
rect 7310 4338 7362 4350
rect 4118 4282 4170 4294
rect 5674 4286 5686 4338
rect 5738 4286 5750 4338
rect 6010 4286 6022 4338
rect 6074 4286 6086 4338
rect 4118 4218 4170 4230
rect 5226 4208 5238 4260
rect 5290 4208 5302 4260
rect 6906 4230 6918 4282
rect 6970 4230 6982 4282
rect 7310 4274 7362 4286
rect 7982 4282 8034 4294
rect 8250 4280 8262 4332
rect 8314 4280 8326 4332
rect 8586 4286 8598 4338
rect 8650 4286 8662 4338
rect 8990 4282 9042 4294
rect 7982 4218 8034 4230
rect 9258 4274 9270 4326
rect 9322 4274 9334 4326
rect 9482 4298 9494 4350
rect 9546 4298 9558 4350
rect 12462 4338 12514 4350
rect 15262 4338 15314 4350
rect 13850 4286 13862 4338
rect 13914 4286 13926 4338
rect 11498 4230 11510 4282
rect 11562 4230 11574 4282
rect 12462 4274 12514 4286
rect 14646 4282 14698 4294
rect 13234 4230 13246 4282
rect 13298 4230 13310 4282
rect 17322 4298 17334 4350
rect 17386 4298 17398 4350
rect 15262 4274 15314 4286
rect 16718 4282 16770 4294
rect 17882 4286 17894 4338
rect 17946 4286 17958 4338
rect 18846 4330 18898 4342
rect 21086 4394 21138 4406
rect 29754 4398 29766 4450
rect 29818 4398 29830 4450
rect 30886 4442 30938 4454
rect 24322 4342 24334 4394
rect 24386 4342 24398 4394
rect 21086 4330 21138 4342
rect 29094 4338 29146 4350
rect 15866 4230 15878 4282
rect 15930 4230 15942 4282
rect 8990 4218 9042 4230
rect 5070 4170 5122 4182
rect 7534 4170 7586 4182
rect 5070 4106 5122 4118
rect 6190 4114 6242 4126
rect 6190 4050 6242 4062
rect 6414 4114 6466 4126
rect 9998 4170 10050 4182
rect 7534 4106 7586 4118
rect 7870 4114 7922 4126
rect 6414 4050 6466 4062
rect 7870 4050 7922 4062
rect 8094 4114 8146 4126
rect 9146 4062 9158 4114
rect 9210 4062 9222 4114
rect 9998 4106 10050 4118
rect 10502 4170 10554 4182
rect 10502 4106 10554 4118
rect 10894 4170 10946 4182
rect 10894 4106 10946 4118
rect 11902 4170 11954 4182
rect 11902 4106 11954 4118
rect 12126 4170 12178 4182
rect 12126 4106 12178 4118
rect 12630 4170 12682 4182
rect 14410 4174 14422 4226
rect 14474 4174 14486 4226
rect 14646 4218 14698 4230
rect 16718 4218 16770 4230
rect 19182 4282 19234 4294
rect 19182 4218 19234 4230
rect 19462 4282 19514 4294
rect 21690 4268 21702 4320
rect 21754 4268 21766 4320
rect 22038 4282 22090 4294
rect 19462 4218 19514 4230
rect 21310 4226 21362 4238
rect 16494 4170 16546 4182
rect 12630 4106 12682 4118
rect 15486 4114 15538 4126
rect 16494 4106 16546 4118
rect 16942 4170 16994 4182
rect 16942 4106 16994 4118
rect 17670 4170 17722 4182
rect 17670 4106 17722 4118
rect 20190 4170 20242 4182
rect 20190 4106 20242 4118
rect 20414 4170 20466 4182
rect 22038 4218 22090 4230
rect 22430 4282 22482 4294
rect 23034 4230 23046 4282
rect 23098 4230 23110 4282
rect 23594 4274 23606 4326
rect 23658 4274 23670 4326
rect 27526 4282 27578 4294
rect 28410 4230 28422 4282
rect 28474 4230 28486 4282
rect 29094 4274 29146 4286
rect 30314 4272 30326 4324
rect 30378 4272 30390 4324
rect 33898 4298 33910 4350
rect 33962 4298 33974 4350
rect 34458 4298 34470 4350
rect 34522 4298 34534 4350
rect 22430 4218 22482 4230
rect 27526 4218 27578 4230
rect 21310 4162 21362 4174
rect 23214 4170 23266 4182
rect 20414 4106 20466 4118
rect 22654 4114 22706 4126
rect 8094 4050 8146 4062
rect 15486 4050 15538 4062
rect 23214 4106 23266 4118
rect 26686 4170 26738 4182
rect 27134 4170 27186 4182
rect 26686 4106 26738 4118
rect 27022 4114 27074 4126
rect 22654 4050 22706 4062
rect 28030 4170 28082 4182
rect 29822 4170 29874 4182
rect 27134 4106 27186 4118
rect 27246 4114 27298 4126
rect 27022 4050 27074 4062
rect 29418 4118 29430 4170
rect 29482 4118 29494 4170
rect 28030 4106 28082 4118
rect 29822 4106 29874 4118
rect 30046 4114 30098 4126
rect 31546 4118 31558 4170
rect 31610 4118 31622 4170
rect 27246 4050 27298 4062
rect 30046 4050 30098 4062
rect 672 3946 34832 3980
rect 672 3894 9094 3946
rect 9146 3894 9198 3946
rect 9250 3894 9302 3946
rect 9354 3894 17646 3946
rect 17698 3894 17750 3946
rect 17802 3894 17854 3946
rect 17906 3894 26198 3946
rect 26250 3894 26302 3946
rect 26354 3894 26406 3946
rect 26458 3894 34832 3946
rect 672 3860 34832 3894
rect 9550 3778 9602 3790
rect 2158 3722 2210 3734
rect 2158 3658 2210 3670
rect 3726 3722 3778 3734
rect 3726 3658 3778 3670
rect 4062 3722 4114 3734
rect 4062 3658 4114 3670
rect 4174 3722 4226 3734
rect 4174 3658 4226 3670
rect 4566 3722 4618 3734
rect 4566 3658 4618 3670
rect 4902 3722 4954 3734
rect 4902 3658 4954 3670
rect 6470 3722 6522 3734
rect 7242 3726 7254 3778
rect 7306 3726 7318 3778
rect 6470 3658 6522 3670
rect 8094 3722 8146 3734
rect 14926 3778 14978 3790
rect 9550 3714 9602 3726
rect 9774 3722 9826 3734
rect 8094 3658 8146 3670
rect 9774 3658 9826 3670
rect 10110 3722 10162 3734
rect 10110 3658 10162 3670
rect 11286 3722 11338 3734
rect 11286 3658 11338 3670
rect 12350 3722 12402 3734
rect 12350 3658 12402 3670
rect 12910 3722 12962 3734
rect 12910 3658 12962 3670
rect 13134 3722 13186 3734
rect 14926 3714 14978 3726
rect 16382 3722 16434 3734
rect 13134 3658 13186 3670
rect 16382 3658 16434 3670
rect 16662 3722 16714 3734
rect 22934 3722 22986 3734
rect 20234 3670 20246 3722
rect 20298 3670 20310 3722
rect 23482 3695 23494 3747
rect 23546 3695 23558 3747
rect 25006 3722 25058 3734
rect 16662 3658 16714 3670
rect 22934 3658 22986 3670
rect 25006 3658 25058 3670
rect 25398 3722 25450 3734
rect 25398 3658 25450 3670
rect 25622 3722 25674 3734
rect 25622 3658 25674 3670
rect 25958 3722 26010 3734
rect 29754 3726 29766 3778
rect 29818 3726 29830 3778
rect 34246 3722 34298 3734
rect 27402 3670 27414 3722
rect 27466 3670 27478 3722
rect 25958 3658 26010 3670
rect 28254 3666 28306 3678
rect 28970 3670 28982 3722
rect 29034 3670 29046 3722
rect 8206 3610 8258 3622
rect 2874 3490 2886 3542
rect 2938 3490 2950 3542
rect 3502 3498 3554 3510
rect 5450 3490 5462 3542
rect 5514 3490 5526 3542
rect 6862 3498 6914 3510
rect 3502 3434 3554 3446
rect 5854 3442 5906 3454
rect 1766 3386 1818 3398
rect 1766 3322 1818 3334
rect 2550 3386 2602 3398
rect 2550 3322 2602 3334
rect 5126 3386 5178 3398
rect 7018 3490 7030 3542
rect 7082 3490 7094 3542
rect 7354 3490 7366 3542
rect 7418 3490 7430 3542
rect 7578 3514 7590 3566
rect 7642 3514 7654 3566
rect 7982 3554 8034 3566
rect 9326 3610 9378 3622
rect 10446 3610 10498 3622
rect 13526 3610 13578 3622
rect 8206 3546 8258 3558
rect 8362 3508 8374 3560
rect 8426 3508 8438 3560
rect 8698 3502 8710 3554
rect 8762 3502 8774 3554
rect 9034 3516 9046 3568
rect 9098 3516 9110 3568
rect 9930 3558 9942 3610
rect 9994 3558 10006 3610
rect 11778 3558 11790 3610
rect 11842 3558 11854 3610
rect 9326 3546 9378 3558
rect 10446 3546 10498 3558
rect 10826 3502 10838 3554
rect 10890 3502 10902 3554
rect 12058 3514 12070 3566
rect 12122 3514 12134 3566
rect 13526 3546 13578 3558
rect 13806 3610 13858 3622
rect 15150 3610 15202 3622
rect 27022 3610 27074 3622
rect 13806 3546 13858 3558
rect 14030 3554 14082 3566
rect 7982 3490 8034 3502
rect 11118 3498 11170 3510
rect 6862 3434 6914 3446
rect 9482 3390 9494 3442
rect 9546 3390 9558 3442
rect 10714 3396 10726 3448
rect 10778 3396 10790 3448
rect 11118 3434 11170 3446
rect 11342 3498 11394 3510
rect 11342 3434 11394 3446
rect 11566 3498 11618 3510
rect 14410 3502 14422 3554
rect 14474 3502 14486 3554
rect 14030 3490 14082 3502
rect 14746 3496 14758 3548
rect 14810 3496 14822 3548
rect 15150 3546 15202 3558
rect 15038 3498 15090 3510
rect 11566 3434 11618 3446
rect 15038 3434 15090 3446
rect 15710 3498 15762 3510
rect 16986 3490 16998 3542
rect 17050 3490 17062 3542
rect 17322 3514 17334 3566
rect 17386 3514 17398 3566
rect 21970 3558 21982 3610
rect 22034 3558 22046 3610
rect 17938 3502 17950 3554
rect 18002 3502 18014 3554
rect 22586 3520 22598 3572
rect 22650 3520 22662 3572
rect 26394 3558 26406 3610
rect 26458 3558 26470 3610
rect 21310 3498 21362 3510
rect 15710 3434 15762 3446
rect 21310 3434 21362 3446
rect 22206 3498 22258 3510
rect 24042 3502 24054 3554
rect 24106 3502 24118 3554
rect 27022 3546 27074 3558
rect 27246 3610 27298 3622
rect 34246 3658 34298 3670
rect 28254 3602 28306 3614
rect 29374 3610 29426 3622
rect 27246 3546 27298 3558
rect 28522 3514 28534 3566
rect 28586 3514 28598 3566
rect 34414 3610 34466 3622
rect 29374 3546 29426 3558
rect 26742 3498 26794 3510
rect 24266 3446 24278 3498
rect 24330 3446 24342 3498
rect 22206 3434 22258 3446
rect 26742 3434 26794 3446
rect 27582 3498 27634 3510
rect 27582 3434 27634 3446
rect 28702 3498 28754 3510
rect 28970 3490 28982 3542
rect 29034 3490 29046 3542
rect 29642 3514 29654 3566
rect 29706 3514 29718 3566
rect 29978 3490 29990 3542
rect 30042 3490 30054 3542
rect 30426 3515 30438 3567
rect 30490 3515 30502 3567
rect 30270 3498 30322 3510
rect 30930 3502 30942 3554
rect 30994 3502 31006 3554
rect 34414 3546 34466 3558
rect 28702 3434 28754 3446
rect 33226 3490 33238 3542
rect 33290 3490 33302 3542
rect 30270 3434 30322 3446
rect 5854 3378 5906 3390
rect 12462 3386 12514 3398
rect 20918 3386 20970 3398
rect 5126 3322 5178 3334
rect 6078 3330 6130 3342
rect 13850 3334 13862 3386
rect 13914 3334 13926 3386
rect 15474 3334 15486 3386
rect 15538 3334 15550 3386
rect 16034 3334 16046 3386
rect 16098 3334 16110 3386
rect 12462 3322 12514 3334
rect 20918 3322 20970 3334
rect 21198 3386 21250 3398
rect 27806 3386 27858 3398
rect 21634 3334 21646 3386
rect 21698 3334 21710 3386
rect 21198 3322 21250 3334
rect 27806 3322 27858 3334
rect 6078 3266 6130 3278
rect 672 3162 34832 3196
rect 672 3110 4818 3162
rect 4870 3110 4922 3162
rect 4974 3110 5026 3162
rect 5078 3110 13370 3162
rect 13422 3110 13474 3162
rect 13526 3110 13578 3162
rect 13630 3110 21922 3162
rect 21974 3110 22026 3162
rect 22078 3110 22130 3162
rect 22182 3110 30474 3162
rect 30526 3110 30578 3162
rect 30630 3110 30682 3162
rect 30734 3110 34832 3162
rect 672 3076 34832 3110
rect 26126 2994 26178 3006
rect 6078 2938 6130 2950
rect 6078 2874 6130 2886
rect 7086 2938 7138 2950
rect 6234 2824 6246 2876
rect 6298 2824 6310 2876
rect 7086 2874 7138 2886
rect 12742 2938 12794 2950
rect 12742 2874 12794 2886
rect 13358 2938 13410 2950
rect 24166 2938 24218 2950
rect 20122 2886 20134 2938
rect 20186 2886 20198 2938
rect 26126 2930 26178 2942
rect 26350 2938 26402 2950
rect 13358 2874 13410 2886
rect 24166 2874 24218 2886
rect 26350 2874 26402 2886
rect 29150 2938 29202 2950
rect 30326 2938 30378 2950
rect 29150 2874 29202 2886
rect 18510 2826 18562 2838
rect 2090 2726 2102 2778
rect 2154 2726 2166 2778
rect 7422 2770 7474 2782
rect 2594 2718 2606 2770
rect 2658 2718 2670 2770
rect 5854 2714 5906 2726
rect 6458 2718 6470 2770
rect 6522 2718 6534 2770
rect 8878 2770 8930 2782
rect 7422 2706 7474 2718
rect 7814 2714 7866 2726
rect 4834 2606 4846 2658
rect 4898 2606 4910 2658
rect 5854 2650 5906 2662
rect 8542 2714 8594 2726
rect 9258 2730 9270 2782
rect 9322 2730 9334 2782
rect 9762 2718 9774 2770
rect 9826 2718 9838 2770
rect 13178 2738 13190 2790
rect 13242 2738 13254 2790
rect 13582 2770 13634 2782
rect 14298 2730 14310 2782
rect 14362 2730 14374 2782
rect 14746 2726 14758 2778
rect 14810 2726 14822 2778
rect 24334 2826 24386 2838
rect 15362 2718 15374 2770
rect 15426 2718 15438 2770
rect 18510 2762 18562 2774
rect 19182 2770 19234 2782
rect 20570 2730 20582 2782
rect 20634 2730 20646 2782
rect 7814 2650 7866 2662
rect 8026 2616 8038 2668
rect 8090 2616 8102 2668
rect 8698 2662 8710 2714
rect 8762 2662 8774 2714
rect 8878 2706 8930 2718
rect 13582 2706 13634 2718
rect 8542 2650 8594 2662
rect 17546 2634 17558 2686
rect 17610 2634 17622 2686
rect 19002 2662 19014 2714
rect 19066 2662 19078 2714
rect 19182 2706 19234 2718
rect 20078 2714 20130 2726
rect 21074 2718 21086 2770
rect 21138 2718 21150 2770
rect 24334 2762 24386 2774
rect 25566 2826 25618 2838
rect 29306 2836 29318 2888
rect 29370 2836 29382 2888
rect 30326 2874 30378 2886
rect 34470 2938 34522 2950
rect 34470 2874 34522 2886
rect 25566 2762 25618 2774
rect 26630 2773 26682 2785
rect 27178 2774 27190 2826
rect 27242 2774 27254 2826
rect 19674 2662 19686 2714
rect 19738 2662 19750 2714
rect 20078 2650 20130 2662
rect 25678 2714 25730 2726
rect 26630 2709 26682 2721
rect 27402 2718 27414 2770
rect 27466 2718 27478 2770
rect 28186 2730 28198 2782
rect 28250 2730 28262 2782
rect 28522 2706 28534 2758
rect 28586 2706 28598 2758
rect 29418 2726 29430 2778
rect 29482 2726 29494 2778
rect 30874 2730 30886 2782
rect 30938 2730 30950 2782
rect 31434 2730 31446 2782
rect 31498 2730 31510 2782
rect 28814 2714 28866 2726
rect 25678 2650 25730 2662
rect 28814 2650 28866 2662
rect 29934 2714 29986 2726
rect 29934 2650 29986 2662
rect 33798 2714 33850 2726
rect 33798 2650 33850 2662
rect 13302 2602 13354 2614
rect 12058 2550 12070 2602
rect 12122 2550 12134 2602
rect 13302 2538 13354 2550
rect 13974 2602 14026 2614
rect 13974 2538 14026 2550
rect 18846 2602 18898 2614
rect 18846 2538 18898 2550
rect 19406 2602 19458 2614
rect 24558 2602 24610 2614
rect 19406 2538 19458 2550
rect 20302 2546 20354 2558
rect 23482 2550 23494 2602
rect 23546 2550 23558 2602
rect 24558 2538 24610 2550
rect 24894 2602 24946 2614
rect 24894 2538 24946 2550
rect 25118 2602 25170 2614
rect 25118 2538 25170 2550
rect 26406 2602 26458 2614
rect 26406 2538 26458 2550
rect 26910 2602 26962 2614
rect 26910 2538 26962 2550
rect 28410 2494 28422 2546
rect 28474 2494 28486 2546
rect 20302 2482 20354 2494
rect 672 2378 34832 2412
rect 672 2326 9094 2378
rect 9146 2326 9198 2378
rect 9250 2326 9302 2378
rect 9354 2326 17646 2378
rect 17698 2326 17750 2378
rect 17802 2326 17854 2378
rect 17906 2326 26198 2378
rect 26250 2326 26302 2378
rect 26354 2326 26406 2378
rect 26458 2326 34832 2378
rect 672 2292 34832 2326
rect 7422 2210 7474 2222
rect 4958 2154 5010 2166
rect 6906 2127 6918 2179
rect 6970 2127 6982 2179
rect 22206 2210 22258 2222
rect 7422 2146 7474 2158
rect 7534 2154 7586 2166
rect 4958 2090 5010 2102
rect 7534 2090 7586 2102
rect 8430 2154 8482 2166
rect 8430 2090 8482 2102
rect 9102 2154 9154 2166
rect 9102 2090 9154 2102
rect 9774 2154 9826 2166
rect 9774 2090 9826 2102
rect 10054 2154 10106 2166
rect 10054 2090 10106 2102
rect 10446 2154 10498 2166
rect 10446 2090 10498 2102
rect 11454 2154 11506 2166
rect 11454 2090 11506 2102
rect 11790 2154 11842 2166
rect 14254 2154 14306 2166
rect 13682 2102 13694 2154
rect 13746 2102 13758 2154
rect 11790 2090 11842 2102
rect 14254 2090 14306 2102
rect 14590 2154 14642 2166
rect 17726 2154 17778 2166
rect 15754 2102 15766 2154
rect 15818 2102 15830 2154
rect 14590 2090 14642 2102
rect 17726 2090 17778 2102
rect 18062 2154 18114 2166
rect 18062 2090 18114 2102
rect 18174 2154 18226 2166
rect 18174 2090 18226 2102
rect 18510 2154 18562 2166
rect 18510 2090 18562 2102
rect 18622 2154 18674 2166
rect 18622 2090 18674 2102
rect 19070 2154 19122 2166
rect 19070 2090 19122 2102
rect 19294 2154 19346 2166
rect 19294 2090 19346 2102
rect 19518 2154 19570 2166
rect 19518 2090 19570 2102
rect 19966 2154 20018 2166
rect 19966 2090 20018 2102
rect 20190 2154 20242 2166
rect 21646 2154 21698 2166
rect 20906 2102 20918 2154
rect 20970 2102 20982 2154
rect 22206 2146 22258 2158
rect 22430 2210 22482 2222
rect 22430 2146 22482 2158
rect 23102 2154 23154 2166
rect 20190 2090 20242 2102
rect 21646 2090 21698 2102
rect 23102 2090 23154 2102
rect 23550 2154 23602 2166
rect 23550 2090 23602 2102
rect 23774 2154 23826 2166
rect 23774 2090 23826 2102
rect 24334 2154 24386 2166
rect 24334 2090 24386 2102
rect 28814 2154 28866 2166
rect 28814 2090 28866 2102
rect 28926 2154 28978 2166
rect 28926 2090 28978 2102
rect 29598 2154 29650 2166
rect 29598 2090 29650 2102
rect 30438 2154 30490 2166
rect 30438 2090 30490 2102
rect 34470 2154 34522 2166
rect 34470 2090 34522 2102
rect 3894 2042 3946 2054
rect 1082 1946 1094 1998
rect 1146 1946 1158 1998
rect 1530 1946 1542 1998
rect 1594 1946 1606 1998
rect 3894 1978 3946 1990
rect 7646 2042 7698 2054
rect 4734 1930 4786 1942
rect 4734 1866 4786 1878
rect 5182 1930 5234 1942
rect 5182 1866 5234 1878
rect 5406 1930 5458 1942
rect 5406 1866 5458 1878
rect 5630 1930 5682 1942
rect 6234 1934 6246 1986
rect 6298 1934 6310 1986
rect 7646 1978 7698 1990
rect 7802 1963 7814 2015
rect 7866 1963 7878 2015
rect 8082 1990 8094 2042
rect 8146 1990 8158 2042
rect 8586 2012 8598 2064
rect 8650 2012 8662 2064
rect 8990 2042 9042 2054
rect 16158 2042 16210 2054
rect 11610 1990 11622 2042
rect 11674 1990 11686 2042
rect 13122 1990 13134 2042
rect 13186 1990 13198 2042
rect 8990 1978 9042 1990
rect 9326 1930 9378 1942
rect 6682 1878 6694 1930
rect 6746 1878 6758 1930
rect 8586 1878 8598 1930
rect 8650 1878 8662 1930
rect 5630 1866 5682 1878
rect 9326 1866 9378 1878
rect 9550 1930 9602 1942
rect 9550 1866 9602 1878
rect 10670 1930 10722 1942
rect 10670 1866 10722 1878
rect 11230 1930 11282 1942
rect 11230 1866 11282 1878
rect 12126 1930 12178 1942
rect 12506 1934 12518 1986
rect 12570 1934 12582 1986
rect 14074 1942 14086 1994
rect 14138 1942 14150 1994
rect 15978 1950 15990 2002
rect 16042 1950 16054 2002
rect 16158 1978 16210 1990
rect 17614 2042 17666 2054
rect 17614 1978 17666 1990
rect 20526 2042 20578 2054
rect 21310 2042 21362 2054
rect 20526 1978 20578 1990
rect 20682 1950 20694 2002
rect 20746 1950 20758 2002
rect 22810 1990 22822 2042
rect 22874 1990 22886 2042
rect 23258 2012 23270 2064
rect 23322 2012 23334 2064
rect 23998 2042 24050 2054
rect 27862 2042 27914 2054
rect 21310 1978 21362 1990
rect 23998 1978 24050 1990
rect 24938 1946 24950 1998
rect 25002 1946 25014 1998
rect 13358 1930 13410 1942
rect 12126 1866 12178 1878
rect 4566 1818 4618 1830
rect 12394 1828 12406 1880
rect 12458 1828 12470 1880
rect 13358 1866 13410 1878
rect 14366 1930 14418 1942
rect 14366 1866 14418 1878
rect 15598 1930 15650 1942
rect 15598 1866 15650 1878
rect 18846 1930 18898 1942
rect 18846 1866 18898 1878
rect 19742 1930 19794 1942
rect 19742 1866 19794 1878
rect 21870 1930 21922 1942
rect 25442 1934 25454 1986
rect 25506 1934 25518 1986
rect 27862 1978 27914 1990
rect 28534 1930 28586 1942
rect 23258 1878 23270 1930
rect 23322 1878 23334 1930
rect 21870 1866 21922 1878
rect 28534 1866 28586 1878
rect 29150 1930 29202 1942
rect 29150 1866 29202 1878
rect 29374 1930 29426 1942
rect 30090 1922 30102 1974
rect 30154 1922 30166 1974
rect 30818 1934 30830 1986
rect 30882 1934 30894 1986
rect 31266 1934 31278 1986
rect 31330 1934 31342 1986
rect 33450 1946 33462 1998
rect 33514 1946 33526 1998
rect 29374 1866 29426 1878
rect 4566 1754 4618 1766
rect 15374 1818 15426 1830
rect 15374 1754 15426 1766
rect 21086 1818 21138 1830
rect 22362 1766 22374 1818
rect 22426 1766 22438 1818
rect 21086 1754 21138 1766
rect 672 1594 34832 1628
rect 672 1542 4818 1594
rect 4870 1542 4922 1594
rect 4974 1542 5026 1594
rect 5078 1542 13370 1594
rect 13422 1542 13474 1594
rect 13526 1542 13578 1594
rect 13630 1542 21922 1594
rect 21974 1542 22026 1594
rect 22078 1542 22130 1594
rect 22182 1542 30474 1594
rect 30526 1542 30578 1594
rect 30630 1542 30682 1594
rect 30734 1542 34832 1594
rect 672 1508 34832 1542
rect 7982 1370 8034 1382
rect 7982 1306 8034 1318
rect 25398 1370 25450 1382
rect 25398 1306 25450 1318
rect 27470 1370 27522 1382
rect 31334 1370 31386 1382
rect 27470 1306 27522 1318
rect 4846 1258 4898 1270
rect 4846 1194 4898 1206
rect 12910 1258 12962 1270
rect 12910 1194 12962 1206
rect 13134 1258 13186 1270
rect 13134 1194 13186 1206
rect 17726 1258 17778 1270
rect 17726 1194 17778 1206
rect 18846 1258 18898 1270
rect 18846 1194 18898 1206
rect 19182 1258 19234 1270
rect 19182 1194 19234 1206
rect 19630 1258 19682 1270
rect 19630 1194 19682 1206
rect 19854 1258 19906 1270
rect 19854 1194 19906 1206
rect 20078 1258 20130 1270
rect 20078 1194 20130 1206
rect 20302 1258 20354 1270
rect 20302 1194 20354 1206
rect 20414 1258 20466 1270
rect 20414 1194 20466 1206
rect 20750 1258 20802 1270
rect 20750 1194 20802 1206
rect 20974 1258 21026 1270
rect 20974 1194 21026 1206
rect 21198 1258 21250 1270
rect 21198 1194 21250 1206
rect 21422 1258 21474 1270
rect 21422 1194 21474 1206
rect 21758 1258 21810 1270
rect 21758 1194 21810 1206
rect 22654 1258 22706 1270
rect 22654 1194 22706 1206
rect 22990 1258 23042 1270
rect 22990 1194 23042 1206
rect 23438 1258 23490 1270
rect 23438 1194 23490 1206
rect 23662 1258 23714 1270
rect 23662 1194 23714 1206
rect 24110 1258 24162 1270
rect 24110 1194 24162 1206
rect 24782 1258 24834 1270
rect 24782 1194 24834 1206
rect 25230 1258 25282 1270
rect 26014 1258 26066 1270
rect 25230 1194 25282 1206
rect 25722 1162 25734 1214
rect 25786 1162 25798 1214
rect 26014 1194 26066 1206
rect 26574 1258 26626 1270
rect 26574 1194 26626 1206
rect 26686 1258 26738 1270
rect 26686 1194 26738 1206
rect 26910 1258 26962 1270
rect 26910 1194 26962 1206
rect 27134 1258 27186 1270
rect 27626 1268 27638 1320
rect 27690 1268 27702 1320
rect 31334 1306 31386 1318
rect 32454 1370 32506 1382
rect 33518 1370 33570 1382
rect 32454 1306 32506 1318
rect 28142 1258 28194 1270
rect 27134 1194 27186 1206
rect 27738 1158 27750 1210
rect 27802 1158 27814 1210
rect 28142 1194 28194 1206
rect 28366 1258 28418 1270
rect 28366 1194 28418 1206
rect 28590 1258 28642 1270
rect 28590 1194 28642 1206
rect 28814 1258 28866 1270
rect 28814 1194 28866 1206
rect 28926 1258 28978 1270
rect 28926 1194 28978 1206
rect 29374 1258 29426 1270
rect 29374 1194 29426 1206
rect 29766 1258 29818 1270
rect 31502 1258 31554 1270
rect 33338 1268 33350 1320
rect 33402 1268 33414 1320
rect 33518 1306 33570 1318
rect 34022 1370 34074 1382
rect 34022 1306 34074 1318
rect 29766 1194 29818 1206
rect 7870 1146 7922 1158
rect 7870 1082 7922 1094
rect 19406 1146 19458 1158
rect 19406 1082 19458 1094
rect 22094 1146 22146 1158
rect 22094 1082 22146 1094
rect 26350 1146 26402 1158
rect 30090 1132 30102 1184
rect 30154 1132 30166 1184
rect 30986 1162 30998 1214
rect 31050 1162 31062 1214
rect 31502 1194 31554 1206
rect 31882 1132 31894 1184
rect 31946 1132 31958 1184
rect 32778 1162 32790 1214
rect 32842 1162 32854 1214
rect 32230 1146 32282 1158
rect 33114 1150 33126 1202
rect 33178 1150 33190 1202
rect 26350 1082 26402 1094
rect 32230 1082 32282 1094
rect 34414 1146 34466 1158
rect 34414 1082 34466 1094
rect 17502 1034 17554 1046
rect 17502 970 17554 982
rect 17950 1034 18002 1046
rect 17950 970 18002 982
rect 18174 1034 18226 1046
rect 18174 970 18226 982
rect 18398 1034 18450 1046
rect 18398 970 18450 982
rect 21646 1034 21698 1046
rect 21646 970 21698 982
rect 22318 1034 22370 1046
rect 22318 970 22370 982
rect 22542 1034 22594 1046
rect 22542 970 22594 982
rect 23102 1034 23154 1046
rect 23102 970 23154 982
rect 23774 1034 23826 1046
rect 23774 970 23826 982
rect 24222 1034 24274 1046
rect 24222 970 24274 982
rect 25006 1034 25058 1046
rect 25006 970 25058 982
rect 29486 1034 29538 1046
rect 29486 970 29538 982
rect 30718 1034 30770 1046
rect 30718 970 30770 982
rect 33854 1034 33906 1046
rect 33854 970 33906 982
rect 672 810 34832 844
rect 672 758 9094 810
rect 9146 758 9198 810
rect 9250 758 9302 810
rect 9354 758 17646 810
rect 17698 758 17750 810
rect 17802 758 17854 810
rect 17906 758 26198 810
rect 26250 758 26302 810
rect 26354 758 26406 810
rect 26458 758 34832 810
rect 672 724 34832 758
rect 20290 534 20302 586
rect 20354 583 20366 586
rect 21634 583 21646 586
rect 20354 537 21646 583
rect 20354 534 20366 537
rect 21634 534 21646 537
rect 21698 583 21710 586
rect 22530 583 22542 586
rect 21698 537 22542 583
rect 21698 534 21710 537
rect 22530 534 22542 537
rect 22594 534 22606 586
rect 20962 422 20974 474
rect 21026 471 21038 474
rect 22306 471 22318 474
rect 21026 425 22318 471
rect 21026 422 21038 425
rect 22306 422 22318 425
rect 22370 422 22382 474
<< via1 >>
rect 4818 12518 4870 12570
rect 4922 12518 4974 12570
rect 5026 12518 5078 12570
rect 13370 12518 13422 12570
rect 13474 12518 13526 12570
rect 13578 12518 13630 12570
rect 21922 12518 21974 12570
rect 22026 12518 22078 12570
rect 22130 12518 22182 12570
rect 30474 12518 30526 12570
rect 30578 12518 30630 12570
rect 30682 12518 30734 12570
rect 6918 12294 6970 12346
rect 12406 12294 12458 12346
rect 18342 12294 18394 12346
rect 21422 12294 21474 12346
rect 1822 12182 1874 12234
rect 2550 12070 2602 12122
rect 9942 12114 9994 12166
rect 10390 12114 10442 12166
rect 13358 12126 13410 12178
rect 23382 12182 23434 12234
rect 10838 12070 10890 12122
rect 13750 12070 13802 12122
rect 14758 12114 14810 12166
rect 15318 12114 15370 12166
rect 19742 12126 19794 12178
rect 24166 12138 24218 12190
rect 14086 12024 14138 12076
rect 1934 11958 1986 12010
rect 2158 11958 2210 12010
rect 5014 11958 5066 12010
rect 7590 11958 7642 12010
rect 10670 11958 10722 12010
rect 11006 11958 11058 12010
rect 11398 11958 11450 12010
rect 11734 11958 11786 12010
rect 12070 11958 12122 12010
rect 13022 11958 13074 12010
rect 18958 12014 19010 12066
rect 20134 12070 20186 12122
rect 21086 12070 21138 12122
rect 14590 11958 14642 12010
rect 17670 11958 17722 12010
rect 20526 12014 20578 12066
rect 21814 12070 21866 12122
rect 24726 12114 24778 12166
rect 25398 12114 25450 12166
rect 28758 12126 28810 12178
rect 30662 12114 30714 12166
rect 31334 12114 31386 12166
rect 22150 12010 22202 12062
rect 19406 11958 19458 12010
rect 22654 11958 22706 12010
rect 27638 12004 27690 12056
rect 28590 11958 28642 12010
rect 29430 11958 29482 12010
rect 33574 12004 33626 12056
rect 34526 11958 34578 12010
rect 9094 11734 9146 11786
rect 9198 11734 9250 11786
rect 9302 11734 9354 11786
rect 17646 11734 17698 11786
rect 17750 11734 17802 11786
rect 17854 11734 17906 11786
rect 26198 11734 26250 11786
rect 26302 11734 26354 11786
rect 26406 11734 26458 11786
rect 2830 11510 2882 11562
rect 11174 11510 11226 11562
rect 1374 11398 1426 11450
rect 2606 11398 2658 11450
rect 3278 11398 3330 11450
rect 8374 11458 8426 11510
rect 11790 11510 11842 11562
rect 15990 11510 16042 11562
rect 7142 11398 7194 11450
rect 8710 11398 8762 11450
rect 13806 11454 13858 11506
rect 16494 11510 16546 11562
rect 17054 11510 17106 11562
rect 17446 11510 17498 11562
rect 29934 11510 29986 11562
rect 1710 11286 1762 11338
rect 2214 11330 2266 11382
rect 3054 11286 3106 11338
rect 3670 11330 3722 11382
rect 4006 11286 4058 11338
rect 4342 11330 4394 11382
rect 4790 11330 4842 11382
rect 9942 11360 9994 11412
rect 12070 11398 12122 11450
rect 10502 11342 10554 11394
rect 16886 11398 16938 11450
rect 17894 11398 17946 11450
rect 9438 11286 9490 11338
rect 11510 11330 11562 11382
rect 12406 11330 12458 11382
rect 13134 11342 13186 11394
rect 16270 11342 16322 11394
rect 18790 11398 18842 11450
rect 19294 11398 19346 11450
rect 20414 11454 20466 11506
rect 30270 11510 30322 11562
rect 20022 11398 20074 11450
rect 21590 11398 21642 11450
rect 1878 11174 1930 11226
rect 7814 11174 7866 11226
rect 9102 11174 9154 11226
rect 10614 11236 10666 11288
rect 20918 11286 20970 11338
rect 23942 11330 23994 11382
rect 24502 11354 24554 11406
rect 25118 11398 25170 11450
rect 28982 11426 29034 11478
rect 26070 11354 26122 11406
rect 26742 11354 26794 11406
rect 30830 11342 30882 11394
rect 30046 11286 30098 11338
rect 31222 11330 31274 11382
rect 33574 11342 33626 11394
rect 10278 11174 10330 11226
rect 10894 11174 10946 11226
rect 16438 11174 16490 11226
rect 18454 11174 18506 11226
rect 19630 11118 19682 11170
rect 25006 11174 25058 11226
rect 25342 11174 25394 11226
rect 25678 11174 25730 11226
rect 25790 11174 25842 11226
rect 34470 11174 34522 11226
rect 4818 10950 4870 11002
rect 4922 10950 4974 11002
rect 5026 10950 5078 11002
rect 13370 10950 13422 11002
rect 13474 10950 13526 11002
rect 13578 10950 13630 11002
rect 21922 10950 21974 11002
rect 22026 10950 22078 11002
rect 22130 10950 22182 11002
rect 30474 10950 30526 11002
rect 30578 10950 30630 11002
rect 30682 10950 30734 11002
rect 9550 10726 9602 10778
rect 1094 10566 1146 10618
rect 1598 10558 1650 10610
rect 3894 10558 3946 10610
rect 5854 10614 5906 10666
rect 8038 10670 8090 10722
rect 13806 10726 13858 10778
rect 14422 10726 14474 10778
rect 5574 10546 5626 10598
rect 5966 10558 6018 10610
rect 6246 10558 6298 10610
rect 6414 10614 6466 10666
rect 16326 10668 16378 10720
rect 6918 10546 6970 10598
rect 7254 10570 7306 10622
rect 7478 10546 7530 10598
rect 7758 10558 7810 10610
rect 8766 10614 8818 10666
rect 8990 10502 9042 10554
rect 9438 10558 9490 10610
rect 9942 10546 9994 10598
rect 10614 10546 10666 10598
rect 14982 10558 15034 10610
rect 16102 10558 16154 10610
rect 17054 10614 17106 10666
rect 17782 10614 17834 10666
rect 19014 10614 19066 10666
rect 12854 10474 12906 10526
rect 14086 10502 14138 10554
rect 14758 10502 14810 10554
rect 16774 10546 16826 10598
rect 17446 10540 17498 10592
rect 18342 10540 18394 10592
rect 22038 10570 22090 10622
rect 26014 10614 26066 10666
rect 26294 10614 26346 10666
rect 34470 10614 34522 10666
rect 22598 10546 22650 10598
rect 25734 10546 25786 10598
rect 26966 10502 27018 10554
rect 29318 10546 29370 10598
rect 29766 10546 29818 10598
rect 30998 10546 31050 10598
rect 31390 10558 31442 10610
rect 4790 10390 4842 10442
rect 5070 10390 5122 10442
rect 25006 10446 25058 10498
rect 5182 10390 5234 10442
rect 5742 10334 5794 10386
rect 7254 10308 7306 10360
rect 8094 10334 8146 10386
rect 9158 10390 9210 10442
rect 15766 10390 15818 10442
rect 8318 10334 8370 10386
rect 16382 10334 16434 10386
rect 16606 10334 16658 10386
rect 18006 10390 18058 10442
rect 19686 10390 19738 10442
rect 22822 10390 22874 10442
rect 30158 10390 30210 10442
rect 30270 10390 30322 10442
rect 33798 10390 33850 10442
rect 9094 10166 9146 10218
rect 9198 10166 9250 10218
rect 9302 10166 9354 10218
rect 17646 10166 17698 10218
rect 17750 10166 17802 10218
rect 17854 10166 17906 10218
rect 26198 10166 26250 10218
rect 26302 10166 26354 10218
rect 26406 10166 26458 10218
rect 5406 9998 5458 10050
rect 6246 9942 6298 9994
rect 7086 9942 7138 9994
rect 7534 9998 7586 10050
rect 14534 10024 14586 10076
rect 20694 10024 20746 10076
rect 7646 9942 7698 9994
rect 8542 9942 8594 9994
rect 8878 9942 8930 9994
rect 9774 9942 9826 9994
rect 10558 9942 10610 9994
rect 11174 9942 11226 9994
rect 13526 9942 13578 9994
rect 16102 9942 16154 9994
rect 19462 9942 19514 9994
rect 19742 9942 19794 9994
rect 20078 9942 20130 9994
rect 21702 9942 21754 9994
rect 22430 9942 22482 9994
rect 24390 9967 24442 10019
rect 25958 9967 26010 10019
rect 26518 9942 26570 9994
rect 28534 9942 28586 9994
rect 32958 9942 33010 9994
rect 33182 9942 33234 9994
rect 1094 9786 1146 9838
rect 1542 9786 1594 9838
rect 3894 9830 3946 9882
rect 4790 9830 4842 9882
rect 5182 9830 5234 9882
rect 6470 9790 6522 9842
rect 6638 9830 6690 9882
rect 6974 9830 7026 9882
rect 7758 9830 7810 9882
rect 8710 9830 8762 9882
rect 9214 9830 9266 9882
rect 10110 9830 10162 9882
rect 4566 9718 4618 9770
rect 5854 9718 5906 9770
rect 7086 9718 7138 9770
rect 7926 9768 7978 9820
rect 8262 9774 8314 9826
rect 10334 9774 10386 9826
rect 10726 9754 10778 9806
rect 11230 9718 11282 9770
rect 11454 9774 11506 9826
rect 11734 9771 11786 9823
rect 12182 9792 12234 9844
rect 13246 9774 13298 9826
rect 13694 9830 13746 9882
rect 14310 9786 14362 9838
rect 14646 9762 14698 9814
rect 14870 9786 14922 9838
rect 15486 9830 15538 9882
rect 16382 9830 16434 9882
rect 17558 9830 17610 9882
rect 17838 9830 17890 9882
rect 18062 9830 18114 9882
rect 18454 9830 18506 9882
rect 19910 9830 19962 9882
rect 20974 9830 21026 9882
rect 16942 9718 16994 9770
rect 18790 9774 18842 9826
rect 21366 9830 21418 9882
rect 22822 9830 22874 9882
rect 17166 9718 17218 9770
rect 20358 9762 20410 9814
rect 20694 9762 20746 9814
rect 22206 9774 22258 9826
rect 23718 9774 23770 9826
rect 25286 9774 25338 9826
rect 26406 9803 26458 9855
rect 22990 9718 23042 9770
rect 23494 9718 23546 9770
rect 25062 9718 25114 9770
rect 26574 9718 26626 9770
rect 27022 9774 27074 9826
rect 27470 9718 27522 9770
rect 27694 9774 27746 9826
rect 27918 9830 27970 9882
rect 28198 9830 28250 9882
rect 29430 9774 29482 9826
rect 33686 9830 33738 9882
rect 31782 9762 31834 9814
rect 32342 9766 32394 9818
rect 5126 9606 5178 9658
rect 6078 9606 6130 9658
rect 9438 9606 9490 9658
rect 10054 9606 10106 9658
rect 12518 9606 12570 9658
rect 13134 9606 13186 9658
rect 13918 9606 13970 9658
rect 15262 9606 15314 9658
rect 15710 9606 15762 9658
rect 16718 9606 16770 9658
rect 17782 9606 17834 9658
rect 22374 9606 22426 9658
rect 27974 9606 28026 9658
rect 32566 9606 32618 9658
rect 26798 9550 26850 9602
rect 34470 9606 34522 9658
rect 4818 9382 4870 9434
rect 4922 9382 4974 9434
rect 5026 9382 5078 9434
rect 13370 9382 13422 9434
rect 13474 9382 13526 9434
rect 13578 9382 13630 9434
rect 21922 9382 21974 9434
rect 22026 9382 22078 9434
rect 22130 9382 22182 9434
rect 30474 9382 30526 9434
rect 30578 9382 30630 9434
rect 30682 9382 30734 9434
rect 4006 9158 4058 9210
rect 5854 9158 5906 9210
rect 6190 9158 6242 9210
rect 7254 9158 7306 9210
rect 7478 9158 7530 9210
rect 7702 9158 7754 9210
rect 10558 9158 10610 9210
rect 11566 9158 11618 9210
rect 1486 9046 1538 9098
rect 1710 9046 1762 9098
rect 1934 9046 1986 9098
rect 2662 9046 2714 9098
rect 2494 8990 2546 9042
rect 3334 8972 3386 9024
rect 3782 8990 3834 9042
rect 4846 9046 4898 9098
rect 5126 8996 5178 9048
rect 6526 9046 6578 9098
rect 5350 8990 5402 9042
rect 9046 9102 9098 9154
rect 6974 9046 7026 9098
rect 11286 9096 11338 9148
rect 11958 9108 12010 9160
rect 12238 9158 12290 9210
rect 12910 9158 12962 9210
rect 13134 9158 13186 9210
rect 18286 9214 18338 9266
rect 15094 9158 15146 9210
rect 17110 9158 17162 9210
rect 20974 9214 21026 9266
rect 12686 9046 12738 9098
rect 18062 9102 18114 9154
rect 19910 9102 19962 9154
rect 21366 9112 21418 9164
rect 22094 9158 22146 9210
rect 22430 9158 22482 9210
rect 26630 9158 26682 9210
rect 26854 9158 26906 9210
rect 30886 9158 30938 9210
rect 2662 8912 2714 8964
rect 1374 8822 1426 8874
rect 2270 8822 2322 8874
rect 2998 8822 3050 8874
rect 3950 8822 4002 8874
rect 4398 8878 4450 8930
rect 4958 8934 5010 8986
rect 5910 8982 5962 9034
rect 9662 8990 9714 9042
rect 10166 8990 10218 9042
rect 8598 8934 8650 8986
rect 10502 8984 10554 9036
rect 11174 8990 11226 9042
rect 12014 8934 12066 8986
rect 13750 8978 13802 9030
rect 14086 8978 14138 9030
rect 14310 9002 14362 9054
rect 15430 9002 15482 9054
rect 16102 9002 16154 9054
rect 16326 9002 16378 9054
rect 16662 8978 16714 9030
rect 16942 8934 16994 8986
rect 17166 8934 17218 8986
rect 17446 8934 17498 8986
rect 17782 8990 17834 9042
rect 19574 8990 19626 9042
rect 20750 8934 20802 8986
rect 21254 8970 21306 9022
rect 21422 8934 21474 8986
rect 22150 8982 22202 9034
rect 23046 9002 23098 9054
rect 23606 8978 23658 9030
rect 25958 8934 26010 8986
rect 29878 8978 29930 9030
rect 30326 9002 30378 9054
rect 33966 8990 34018 9042
rect 34358 9002 34410 9054
rect 4174 8766 4226 8818
rect 4734 8766 4786 8818
rect 8038 8822 8090 8874
rect 8206 8822 8258 8874
rect 8430 8822 8482 8874
rect 8766 8822 8818 8874
rect 9102 8822 9154 8874
rect 9326 8822 9378 8874
rect 9774 8822 9826 8874
rect 10670 8766 10722 8818
rect 10894 8766 10946 8818
rect 13526 8822 13578 8874
rect 14702 8822 14754 8874
rect 15766 8822 15818 8874
rect 18342 8822 18394 8874
rect 18846 8822 18898 8874
rect 20246 8822 20298 8874
rect 21646 8822 21698 8874
rect 13974 8740 14026 8792
rect 16438 8766 16490 8818
rect 22654 8822 22706 8874
rect 27526 8822 27578 8874
rect 31558 8822 31610 8874
rect 9094 8598 9146 8650
rect 9198 8598 9250 8650
rect 9302 8598 9354 8650
rect 17646 8598 17698 8650
rect 17750 8598 17802 8650
rect 17854 8598 17906 8650
rect 26198 8598 26250 8650
rect 26302 8598 26354 8650
rect 26406 8598 26458 8650
rect 1654 8374 1706 8426
rect 5406 8318 5458 8370
rect 10782 8374 10834 8426
rect 14030 8430 14082 8482
rect 21030 8430 21082 8482
rect 19910 8374 19962 8426
rect 25398 8430 25450 8482
rect 31782 8430 31834 8482
rect 24502 8374 24554 8426
rect 26406 8374 26458 8426
rect 30214 8374 30266 8426
rect 34022 8374 34074 8426
rect 4006 8218 4058 8270
rect 6862 8262 6914 8314
rect 7478 8284 7530 8336
rect 8038 8284 8090 8336
rect 982 8150 1034 8202
rect 4566 8194 4618 8246
rect 6022 8194 6074 8246
rect 6302 8150 6354 8202
rect 6526 8150 6578 8202
rect 6974 8150 7026 8202
rect 7310 8206 7362 8258
rect 7870 8206 7922 8258
rect 8430 8262 8482 8314
rect 8710 8206 8762 8258
rect 9046 8212 9098 8264
rect 9214 8262 9266 8314
rect 9438 8206 9490 8258
rect 7478 8150 7530 8202
rect 8038 8150 8090 8202
rect 9774 8206 9826 8258
rect 9998 8262 10050 8314
rect 10950 8262 11002 8314
rect 10222 8206 10274 8258
rect 10390 8206 10442 8258
rect 11118 8206 11170 8258
rect 11342 8262 11394 8314
rect 11734 8262 11786 8314
rect 11902 8262 11954 8314
rect 12406 8284 12458 8336
rect 12238 8206 12290 8258
rect 13022 8262 13074 8314
rect 13358 8262 13410 8314
rect 13806 8262 13858 8314
rect 14478 8262 14530 8314
rect 12406 8150 12458 8202
rect 13638 8186 13690 8238
rect 13918 8150 13970 8202
rect 14926 8206 14978 8258
rect 15150 8262 15202 8314
rect 15542 8262 15594 8314
rect 15822 8150 15874 8202
rect 16102 8198 16154 8250
rect 16606 8206 16658 8258
rect 18902 8194 18954 8246
rect 20078 8150 20130 8202
rect 20582 8194 20634 8246
rect 20918 8218 20970 8270
rect 21198 8262 21250 8314
rect 20750 8150 20802 8202
rect 21590 8194 21642 8246
rect 25062 8218 25114 8270
rect 26798 8262 26850 8314
rect 25286 8194 25338 8246
rect 25622 8194 25674 8246
rect 26630 8194 26682 8246
rect 27022 8150 27074 8202
rect 27302 8194 27354 8246
rect 27862 8218 27914 8270
rect 31446 8206 31498 8258
rect 32566 8224 32618 8276
rect 33350 8262 33402 8314
rect 31222 8150 31274 8202
rect 32902 8150 32954 8202
rect 4790 8038 4842 8090
rect 5182 7982 5234 8034
rect 5686 8038 5738 8090
rect 9102 8038 9154 8090
rect 10054 8084 10106 8136
rect 11790 8038 11842 8090
rect 22318 8094 22370 8146
rect 33070 8150 33122 8202
rect 33686 8194 33738 8246
rect 34358 8194 34410 8246
rect 14590 8038 14642 8090
rect 15094 8038 15146 8090
rect 26014 8038 26066 8090
rect 26238 8038 26290 8090
rect 30886 8038 30938 8090
rect 4818 7814 4870 7866
rect 4922 7814 4974 7866
rect 5026 7814 5078 7866
rect 13370 7814 13422 7866
rect 13474 7814 13526 7866
rect 13578 7814 13630 7866
rect 21922 7814 21974 7866
rect 22026 7814 22078 7866
rect 22130 7814 22182 7866
rect 30474 7814 30526 7866
rect 30578 7814 30630 7866
rect 30682 7814 30734 7866
rect 6134 7590 6186 7642
rect 7534 7590 7586 7642
rect 7870 7646 7922 7698
rect 9046 7590 9098 7642
rect 10334 7590 10386 7642
rect 11342 7590 11394 7642
rect 11454 7590 11506 7642
rect 11846 7590 11898 7642
rect 18510 7590 18562 7642
rect 14198 7534 14250 7586
rect 29990 7590 30042 7642
rect 2662 7410 2714 7462
rect 3110 7434 3162 7486
rect 9438 7478 9490 7530
rect 8262 7366 8314 7418
rect 8598 7320 8650 7372
rect 9662 7366 9714 7418
rect 10390 7422 10442 7474
rect 10950 7434 11002 7486
rect 12630 7478 12682 7530
rect 13582 7478 13634 7530
rect 27806 7534 27858 7586
rect 30886 7590 30938 7642
rect 9998 7366 10050 7418
rect 12854 7422 12906 7474
rect 12238 7366 12290 7418
rect 14366 7422 14418 7474
rect 13918 7366 13970 7418
rect 14646 7410 14698 7462
rect 15318 7434 15370 7486
rect 22710 7478 22762 7530
rect 18846 7422 18898 7474
rect 19518 7422 19570 7474
rect 21702 7410 21754 7462
rect 23046 7409 23098 7461
rect 23494 7410 23546 7462
rect 25734 7434 25786 7486
rect 27078 7410 27130 7462
rect 17558 7338 17610 7390
rect 30270 7366 30322 7418
rect 33910 7410 33962 7462
rect 34470 7410 34522 7462
rect 5462 7254 5514 7306
rect 6414 7254 6466 7306
rect 6862 7254 6914 7306
rect 7086 7254 7138 7306
rect 10614 7254 10666 7306
rect 14142 7198 14194 7250
rect 26742 7254 26794 7306
rect 30382 7254 30434 7306
rect 31558 7254 31610 7306
rect 9094 7030 9146 7082
rect 9198 7030 9250 7082
rect 9302 7030 9354 7082
rect 17646 7030 17698 7082
rect 17750 7030 17802 7082
rect 17854 7030 17906 7082
rect 26198 7030 26250 7082
rect 26302 7030 26354 7082
rect 26406 7030 26458 7082
rect 3502 6806 3554 6858
rect 4174 6806 4226 6858
rect 12238 6806 12290 6858
rect 13246 6806 13298 6858
rect 13582 6806 13634 6858
rect 16214 6862 16266 6914
rect 14870 6806 14922 6858
rect 18846 6806 18898 6858
rect 19294 6806 19346 6858
rect 20526 6806 20578 6858
rect 20918 6831 20970 6883
rect 23942 6831 23994 6883
rect 25622 6806 25674 6858
rect 32958 6806 33010 6858
rect 7366 6722 7418 6774
rect 2102 6626 2154 6678
rect 4566 6650 4618 6702
rect 11398 6694 11450 6746
rect 13078 6694 13130 6746
rect 13806 6694 13858 6746
rect 3278 6582 3330 6634
rect 3726 6582 3778 6634
rect 5182 6638 5234 6690
rect 14086 6694 14138 6746
rect 15486 6694 15538 6746
rect 15710 6694 15762 6746
rect 3950 6582 4002 6634
rect 8318 6582 8370 6634
rect 8486 6626 8538 6678
rect 9046 6626 9098 6678
rect 12574 6582 12626 6634
rect 14366 6582 14418 6634
rect 14590 6582 14642 6634
rect 15262 6582 15314 6634
rect 15990 6626 16042 6678
rect 16326 6626 16378 6678
rect 16550 6626 16602 6678
rect 17222 6656 17274 6708
rect 20134 6694 20186 6746
rect 16886 6582 16938 6634
rect 17502 6582 17554 6634
rect 17726 6582 17778 6634
rect 18398 6582 18450 6634
rect 18622 6582 18674 6634
rect 19406 6582 19458 6634
rect 21366 6638 21418 6690
rect 19742 6582 19794 6634
rect 21814 6582 21866 6634
rect 22094 6582 22146 6634
rect 22486 6626 22538 6678
rect 23382 6638 23434 6690
rect 22822 6582 22874 6634
rect 23158 6582 23210 6634
rect 24334 6582 24386 6634
rect 27974 6626 28026 6678
rect 28422 6626 28474 6678
rect 29878 6650 29930 6702
rect 32118 6626 32170 6678
rect 32566 6630 32618 6682
rect 33350 6582 33402 6634
rect 33518 6582 33570 6634
rect 33742 6582 33794 6634
rect 34358 6626 34410 6678
rect 1766 6470 1818 6522
rect 12070 6470 12122 6522
rect 13134 6470 13186 6522
rect 13750 6470 13802 6522
rect 18062 6470 18114 6522
rect 18174 6470 18226 6522
rect 19854 6470 19906 6522
rect 24950 6470 25002 6522
rect 28870 6470 28922 6522
rect 34022 6470 34074 6522
rect 4818 6246 4870 6298
rect 4922 6246 4974 6298
rect 5026 6246 5078 6298
rect 13370 6246 13422 6298
rect 13474 6246 13526 6298
rect 13578 6246 13630 6298
rect 21922 6246 21974 6298
rect 22026 6246 22078 6298
rect 22130 6246 22182 6298
rect 30474 6246 30526 6298
rect 30578 6246 30630 6298
rect 30682 6246 30734 6298
rect 7758 6022 7810 6074
rect 6246 5966 6298 6018
rect 24558 6078 24610 6130
rect 13414 6022 13466 6074
rect 13974 6022 14026 6074
rect 18454 6022 18506 6074
rect 24782 6078 24834 6130
rect 25006 6078 25058 6130
rect 29654 6022 29706 6074
rect 30886 6022 30938 6074
rect 8710 5961 8762 6013
rect 1094 5841 1146 5893
rect 1710 5854 1762 5906
rect 3894 5842 3946 5894
rect 6470 5866 6522 5918
rect 7142 5866 7194 5918
rect 6190 5798 6242 5850
rect 6974 5798 7026 5850
rect 8262 5854 8314 5906
rect 8598 5860 8650 5912
rect 9942 5866 9994 5918
rect 7534 5798 7586 5850
rect 10446 5854 10498 5906
rect 9214 5798 9266 5850
rect 9382 5798 9434 5850
rect 12742 5798 12794 5850
rect 14030 5854 14082 5906
rect 14646 5862 14698 5914
rect 14422 5798 14474 5850
rect 15206 5842 15258 5894
rect 17446 5866 17498 5918
rect 23830 5910 23882 5962
rect 18846 5798 18898 5850
rect 19182 5798 19234 5850
rect 19462 5846 19514 5898
rect 19910 5842 19962 5894
rect 23382 5854 23434 5906
rect 25174 5875 25226 5927
rect 25846 5862 25898 5914
rect 22822 5798 22874 5850
rect 26406 5842 26458 5894
rect 28646 5866 28698 5918
rect 33966 5854 34018 5906
rect 34358 5842 34410 5894
rect 4902 5686 4954 5738
rect 5182 5686 5234 5738
rect 5574 5686 5626 5738
rect 7366 5686 7418 5738
rect 8766 5686 8818 5738
rect 5966 5630 6018 5682
rect 8990 5630 9042 5682
rect 9550 5686 9602 5738
rect 20638 5742 20690 5794
rect 13806 5630 13858 5682
rect 19294 5686 19346 5738
rect 23718 5626 23770 5678
rect 24614 5686 24666 5738
rect 25454 5686 25506 5738
rect 29878 5686 29930 5738
rect 30214 5686 30266 5738
rect 31558 5686 31610 5738
rect 9094 5462 9146 5514
rect 9198 5462 9250 5514
rect 9302 5462 9354 5514
rect 17646 5462 17698 5514
rect 17750 5462 17802 5514
rect 17854 5462 17906 5514
rect 26198 5462 26250 5514
rect 26302 5462 26354 5514
rect 26406 5462 26458 5514
rect 3894 5238 3946 5290
rect 4846 5238 4898 5290
rect 6078 5294 6130 5346
rect 6862 5294 6914 5346
rect 7870 5294 7922 5346
rect 5182 5126 5234 5178
rect 5854 5126 5906 5178
rect 7086 5126 7138 5178
rect 8318 5182 8370 5234
rect 9886 5238 9938 5290
rect 10110 5294 10162 5346
rect 10894 5238 10946 5290
rect 12182 5238 12234 5290
rect 18678 5263 18730 5315
rect 19518 5294 19570 5346
rect 19742 5294 19794 5346
rect 25510 5320 25562 5372
rect 23830 5238 23882 5290
rect 16606 5182 16658 5234
rect 26966 5238 27018 5290
rect 29318 5238 29370 5290
rect 33462 5238 33514 5290
rect 34078 5238 34130 5290
rect 34302 5238 34354 5290
rect 1094 5058 1146 5110
rect 1542 5058 1594 5110
rect 5462 5062 5514 5114
rect 6358 5058 6410 5110
rect 6694 5058 6746 5110
rect 7366 5070 7418 5122
rect 7702 5070 7754 5122
rect 8094 5070 8146 5122
rect 8654 5126 8706 5178
rect 9270 5126 9322 5178
rect 9998 5126 10050 5178
rect 11062 5126 11114 5178
rect 5350 4964 5402 5016
rect 8766 5014 8818 5066
rect 8878 5070 8930 5122
rect 5798 4958 5850 5010
rect 9550 5014 9602 5066
rect 10278 5064 10330 5116
rect 10502 5070 10554 5122
rect 11230 5070 11282 5122
rect 12294 5099 12346 5151
rect 13078 5088 13130 5140
rect 13638 5082 13690 5134
rect 4566 4902 4618 4954
rect 7142 4946 7194 4998
rect 11678 4958 11730 5010
rect 12126 5014 12178 5066
rect 14310 5058 14362 5110
rect 18006 5070 18058 5122
rect 17782 5014 17834 5066
rect 19350 5050 19402 5102
rect 19630 5014 19682 5066
rect 20414 5070 20466 5122
rect 23718 5099 23770 5151
rect 25174 5082 25226 5134
rect 25398 5082 25450 5134
rect 25734 5082 25786 5134
rect 26070 5126 26122 5178
rect 27862 5126 27914 5178
rect 28142 5126 28194 5178
rect 20078 5014 20130 5066
rect 7814 4902 7866 4954
rect 11902 4902 11954 4954
rect 13414 4902 13466 4954
rect 17502 4902 17554 4954
rect 21198 4958 21250 5010
rect 23886 4958 23938 5010
rect 26630 5014 26682 5066
rect 28366 5070 28418 5122
rect 28758 5070 28810 5122
rect 29766 5082 29818 5134
rect 32566 5126 32618 5178
rect 30214 5058 30266 5110
rect 33798 5058 33850 5110
rect 19070 4902 19122 4954
rect 23270 4902 23322 4954
rect 24110 4902 24162 4954
rect 24334 4902 24386 4954
rect 26406 4902 26458 4954
rect 27358 4902 27410 4954
rect 27470 4902 27522 4954
rect 28086 4902 28138 4954
rect 29038 4902 29090 4954
rect 29262 4902 29314 4954
rect 33238 4902 33290 4954
rect 4818 4678 4870 4730
rect 4922 4678 4974 4730
rect 5026 4678 5078 4730
rect 13370 4678 13422 4730
rect 13474 4678 13526 4730
rect 13578 4678 13630 4730
rect 21922 4678 21974 4730
rect 22026 4678 22078 4730
rect 22130 4678 22182 4730
rect 30474 4678 30526 4730
rect 30578 4678 30630 4730
rect 30682 4678 30734 4730
rect 4790 4454 4842 4506
rect 6078 4454 6130 4506
rect 7366 4454 7418 4506
rect 9942 4404 9994 4456
rect 10222 4454 10274 4506
rect 11174 4454 11226 4506
rect 13022 4454 13074 4506
rect 13470 4454 13522 4506
rect 13750 4454 13802 4506
rect 15430 4454 15482 4506
rect 16102 4454 16154 4506
rect 12182 4398 12234 4450
rect 18286 4454 18338 4506
rect 19798 4454 19850 4506
rect 20694 4454 20746 4506
rect 22710 4454 22762 4506
rect 26518 4454 26570 4506
rect 1206 4274 1258 4326
rect 1766 4298 1818 4350
rect 5238 4342 5290 4394
rect 18006 4392 18058 4444
rect 27918 4454 27970 4506
rect 30886 4454 30938 4506
rect 5686 4286 5738 4338
rect 6022 4286 6074 4338
rect 7310 4286 7362 4338
rect 4118 4230 4170 4282
rect 5238 4208 5290 4260
rect 6918 4230 6970 4282
rect 7982 4230 8034 4282
rect 8262 4280 8314 4332
rect 8598 4286 8650 4338
rect 8990 4230 9042 4282
rect 9270 4274 9322 4326
rect 9494 4298 9546 4350
rect 12462 4286 12514 4338
rect 13862 4286 13914 4338
rect 11510 4230 11562 4282
rect 13246 4230 13298 4282
rect 14646 4230 14698 4282
rect 15262 4286 15314 4338
rect 17334 4298 17386 4350
rect 18846 4342 18898 4394
rect 17894 4286 17946 4338
rect 29766 4398 29818 4450
rect 21086 4342 21138 4394
rect 24334 4342 24386 4394
rect 15878 4230 15930 4282
rect 16718 4230 16770 4282
rect 5070 4118 5122 4170
rect 6190 4062 6242 4114
rect 6414 4062 6466 4114
rect 7534 4118 7586 4170
rect 7870 4062 7922 4114
rect 9998 4118 10050 4170
rect 8094 4062 8146 4114
rect 9158 4062 9210 4114
rect 10502 4118 10554 4170
rect 10894 4118 10946 4170
rect 11902 4118 11954 4170
rect 12126 4118 12178 4170
rect 14422 4174 14474 4226
rect 19182 4230 19234 4282
rect 19462 4230 19514 4282
rect 21702 4268 21754 4320
rect 12630 4118 12682 4170
rect 15486 4062 15538 4114
rect 16494 4118 16546 4170
rect 16942 4118 16994 4170
rect 17670 4118 17722 4170
rect 20190 4118 20242 4170
rect 20414 4118 20466 4170
rect 21310 4174 21362 4226
rect 22038 4230 22090 4282
rect 22430 4230 22482 4282
rect 23046 4230 23098 4282
rect 23606 4274 23658 4326
rect 29094 4286 29146 4338
rect 27526 4230 27578 4282
rect 28422 4230 28474 4282
rect 30326 4272 30378 4324
rect 33910 4298 33962 4350
rect 34470 4298 34522 4350
rect 22654 4062 22706 4114
rect 23214 4118 23266 4170
rect 26686 4118 26738 4170
rect 27022 4062 27074 4114
rect 27134 4118 27186 4170
rect 27246 4062 27298 4114
rect 28030 4118 28082 4170
rect 29430 4118 29482 4170
rect 29822 4118 29874 4170
rect 31558 4118 31610 4170
rect 30046 4062 30098 4114
rect 9094 3894 9146 3946
rect 9198 3894 9250 3946
rect 9302 3894 9354 3946
rect 17646 3894 17698 3946
rect 17750 3894 17802 3946
rect 17854 3894 17906 3946
rect 26198 3894 26250 3946
rect 26302 3894 26354 3946
rect 26406 3894 26458 3946
rect 2158 3670 2210 3722
rect 3726 3670 3778 3722
rect 4062 3670 4114 3722
rect 4174 3670 4226 3722
rect 4566 3670 4618 3722
rect 4902 3670 4954 3722
rect 7254 3726 7306 3778
rect 6470 3670 6522 3722
rect 8094 3670 8146 3722
rect 9550 3726 9602 3778
rect 9774 3670 9826 3722
rect 10110 3670 10162 3722
rect 11286 3670 11338 3722
rect 12350 3670 12402 3722
rect 12910 3670 12962 3722
rect 13134 3670 13186 3722
rect 14926 3726 14978 3778
rect 16382 3670 16434 3722
rect 16662 3670 16714 3722
rect 20246 3670 20298 3722
rect 22934 3670 22986 3722
rect 23494 3695 23546 3747
rect 25006 3670 25058 3722
rect 25398 3670 25450 3722
rect 25622 3670 25674 3722
rect 29766 3726 29818 3778
rect 25958 3670 26010 3722
rect 27414 3670 27466 3722
rect 28982 3670 29034 3722
rect 34246 3670 34298 3722
rect 2886 3490 2938 3542
rect 3502 3446 3554 3498
rect 5462 3490 5514 3542
rect 1766 3334 1818 3386
rect 2550 3334 2602 3386
rect 5126 3334 5178 3386
rect 5854 3390 5906 3442
rect 6862 3446 6914 3498
rect 7030 3490 7082 3542
rect 7366 3490 7418 3542
rect 7590 3514 7642 3566
rect 7982 3502 8034 3554
rect 8206 3558 8258 3610
rect 8374 3508 8426 3560
rect 8710 3502 8762 3554
rect 9046 3516 9098 3568
rect 9326 3558 9378 3610
rect 9942 3558 9994 3610
rect 10446 3558 10498 3610
rect 11790 3558 11842 3610
rect 10838 3502 10890 3554
rect 12070 3514 12122 3566
rect 13526 3558 13578 3610
rect 13806 3558 13858 3610
rect 15150 3558 15202 3610
rect 9494 3390 9546 3442
rect 10726 3396 10778 3448
rect 11118 3446 11170 3498
rect 11342 3446 11394 3498
rect 11566 3446 11618 3498
rect 14030 3502 14082 3554
rect 14422 3502 14474 3554
rect 14758 3496 14810 3548
rect 15038 3446 15090 3498
rect 15710 3446 15762 3498
rect 16998 3490 17050 3542
rect 17334 3514 17386 3566
rect 21982 3558 22034 3610
rect 17950 3502 18002 3554
rect 22598 3520 22650 3572
rect 26406 3558 26458 3610
rect 27022 3558 27074 3610
rect 21310 3446 21362 3498
rect 24054 3502 24106 3554
rect 27246 3558 27298 3610
rect 28254 3614 28306 3666
rect 28534 3514 28586 3566
rect 29374 3558 29426 3610
rect 22206 3446 22258 3498
rect 24278 3446 24330 3498
rect 26742 3446 26794 3498
rect 27582 3446 27634 3498
rect 28702 3446 28754 3498
rect 28982 3490 29034 3542
rect 29654 3514 29706 3566
rect 29990 3490 30042 3542
rect 30438 3515 30490 3567
rect 34414 3558 34466 3610
rect 30942 3502 30994 3554
rect 30270 3446 30322 3498
rect 33238 3490 33290 3542
rect 6078 3278 6130 3330
rect 12462 3334 12514 3386
rect 13862 3334 13914 3386
rect 15486 3334 15538 3386
rect 16046 3334 16098 3386
rect 20918 3334 20970 3386
rect 21198 3334 21250 3386
rect 21646 3334 21698 3386
rect 27806 3334 27858 3386
rect 4818 3110 4870 3162
rect 4922 3110 4974 3162
rect 5026 3110 5078 3162
rect 13370 3110 13422 3162
rect 13474 3110 13526 3162
rect 13578 3110 13630 3162
rect 21922 3110 21974 3162
rect 22026 3110 22078 3162
rect 22130 3110 22182 3162
rect 30474 3110 30526 3162
rect 30578 3110 30630 3162
rect 30682 3110 30734 3162
rect 6078 2886 6130 2938
rect 7086 2886 7138 2938
rect 6246 2824 6298 2876
rect 12742 2886 12794 2938
rect 13358 2886 13410 2938
rect 20134 2886 20186 2938
rect 24166 2886 24218 2938
rect 26126 2942 26178 2994
rect 26350 2886 26402 2938
rect 29150 2886 29202 2938
rect 2102 2726 2154 2778
rect 2606 2718 2658 2770
rect 6470 2718 6522 2770
rect 7422 2718 7474 2770
rect 5854 2662 5906 2714
rect 4846 2606 4898 2658
rect 7814 2662 7866 2714
rect 8878 2718 8930 2770
rect 9270 2730 9322 2782
rect 9774 2718 9826 2770
rect 13190 2738 13242 2790
rect 13582 2718 13634 2770
rect 14310 2730 14362 2782
rect 14758 2726 14810 2778
rect 18510 2774 18562 2826
rect 15374 2718 15426 2770
rect 19182 2718 19234 2770
rect 20582 2730 20634 2782
rect 24334 2774 24386 2826
rect 8038 2616 8090 2668
rect 8542 2662 8594 2714
rect 8710 2662 8762 2714
rect 17558 2634 17610 2686
rect 19014 2662 19066 2714
rect 21086 2718 21138 2770
rect 29318 2836 29370 2888
rect 30326 2886 30378 2938
rect 34470 2886 34522 2938
rect 25566 2774 25618 2826
rect 27190 2774 27242 2826
rect 19686 2662 19738 2714
rect 20078 2662 20130 2714
rect 25678 2662 25730 2714
rect 26630 2721 26682 2773
rect 27414 2718 27466 2770
rect 28198 2730 28250 2782
rect 28534 2706 28586 2758
rect 29430 2726 29482 2778
rect 30886 2730 30938 2782
rect 31446 2730 31498 2782
rect 28814 2662 28866 2714
rect 29934 2662 29986 2714
rect 33798 2662 33850 2714
rect 12070 2550 12122 2602
rect 13302 2550 13354 2602
rect 13974 2550 14026 2602
rect 18846 2550 18898 2602
rect 19406 2550 19458 2602
rect 23494 2550 23546 2602
rect 24558 2550 24610 2602
rect 20302 2494 20354 2546
rect 24894 2550 24946 2602
rect 25118 2550 25170 2602
rect 26406 2550 26458 2602
rect 26910 2550 26962 2602
rect 28422 2494 28474 2546
rect 9094 2326 9146 2378
rect 9198 2326 9250 2378
rect 9302 2326 9354 2378
rect 17646 2326 17698 2378
rect 17750 2326 17802 2378
rect 17854 2326 17906 2378
rect 26198 2326 26250 2378
rect 26302 2326 26354 2378
rect 26406 2326 26458 2378
rect 4958 2102 5010 2154
rect 6918 2127 6970 2179
rect 7422 2158 7474 2210
rect 7534 2102 7586 2154
rect 8430 2102 8482 2154
rect 9102 2102 9154 2154
rect 9774 2102 9826 2154
rect 10054 2102 10106 2154
rect 10446 2102 10498 2154
rect 11454 2102 11506 2154
rect 11790 2102 11842 2154
rect 13694 2102 13746 2154
rect 14254 2102 14306 2154
rect 14590 2102 14642 2154
rect 15766 2102 15818 2154
rect 17726 2102 17778 2154
rect 18062 2102 18114 2154
rect 18174 2102 18226 2154
rect 18510 2102 18562 2154
rect 18622 2102 18674 2154
rect 19070 2102 19122 2154
rect 19294 2102 19346 2154
rect 19518 2102 19570 2154
rect 19966 2102 20018 2154
rect 20190 2102 20242 2154
rect 20918 2102 20970 2154
rect 21646 2102 21698 2154
rect 22206 2158 22258 2210
rect 22430 2158 22482 2210
rect 23102 2102 23154 2154
rect 23550 2102 23602 2154
rect 23774 2102 23826 2154
rect 24334 2102 24386 2154
rect 28814 2102 28866 2154
rect 28926 2102 28978 2154
rect 29598 2102 29650 2154
rect 30438 2102 30490 2154
rect 34470 2102 34522 2154
rect 1094 1946 1146 1998
rect 1542 1946 1594 1998
rect 3894 1990 3946 2042
rect 7646 1990 7698 2042
rect 4734 1878 4786 1930
rect 5182 1878 5234 1930
rect 5406 1878 5458 1930
rect 6246 1934 6298 1986
rect 7814 1963 7866 2015
rect 8094 1990 8146 2042
rect 8598 2012 8650 2064
rect 8990 1990 9042 2042
rect 11622 1990 11674 2042
rect 13134 1990 13186 2042
rect 5630 1878 5682 1930
rect 6694 1878 6746 1930
rect 8598 1878 8650 1930
rect 9326 1878 9378 1930
rect 9550 1878 9602 1930
rect 10670 1878 10722 1930
rect 11230 1878 11282 1930
rect 12518 1934 12570 1986
rect 14086 1942 14138 1994
rect 15990 1950 16042 2002
rect 16158 1990 16210 2042
rect 17614 1990 17666 2042
rect 20526 1990 20578 2042
rect 20694 1950 20746 2002
rect 21310 1990 21362 2042
rect 22822 1990 22874 2042
rect 23270 2012 23322 2064
rect 23998 1990 24050 2042
rect 24950 1946 25002 1998
rect 27862 1990 27914 2042
rect 12126 1878 12178 1930
rect 12406 1828 12458 1880
rect 13358 1878 13410 1930
rect 14366 1878 14418 1930
rect 15598 1878 15650 1930
rect 18846 1878 18898 1930
rect 19742 1878 19794 1930
rect 25454 1934 25506 1986
rect 21870 1878 21922 1930
rect 23270 1878 23322 1930
rect 28534 1878 28586 1930
rect 29150 1878 29202 1930
rect 29374 1878 29426 1930
rect 30102 1922 30154 1974
rect 30830 1934 30882 1986
rect 31278 1934 31330 1986
rect 33462 1946 33514 1998
rect 4566 1766 4618 1818
rect 15374 1766 15426 1818
rect 21086 1766 21138 1818
rect 22374 1766 22426 1818
rect 4818 1542 4870 1594
rect 4922 1542 4974 1594
rect 5026 1542 5078 1594
rect 13370 1542 13422 1594
rect 13474 1542 13526 1594
rect 13578 1542 13630 1594
rect 21922 1542 21974 1594
rect 22026 1542 22078 1594
rect 22130 1542 22182 1594
rect 30474 1542 30526 1594
rect 30578 1542 30630 1594
rect 30682 1542 30734 1594
rect 7982 1318 8034 1370
rect 25398 1318 25450 1370
rect 27470 1318 27522 1370
rect 4846 1206 4898 1258
rect 12910 1206 12962 1258
rect 13134 1206 13186 1258
rect 17726 1206 17778 1258
rect 18846 1206 18898 1258
rect 19182 1206 19234 1258
rect 19630 1206 19682 1258
rect 19854 1206 19906 1258
rect 20078 1206 20130 1258
rect 20302 1206 20354 1258
rect 20414 1206 20466 1258
rect 20750 1206 20802 1258
rect 20974 1206 21026 1258
rect 21198 1206 21250 1258
rect 21422 1206 21474 1258
rect 21758 1206 21810 1258
rect 22654 1206 22706 1258
rect 22990 1206 23042 1258
rect 23438 1206 23490 1258
rect 23662 1206 23714 1258
rect 24110 1206 24162 1258
rect 24782 1206 24834 1258
rect 25230 1206 25282 1258
rect 25734 1162 25786 1214
rect 26014 1206 26066 1258
rect 26574 1206 26626 1258
rect 26686 1206 26738 1258
rect 26910 1206 26962 1258
rect 27638 1268 27690 1320
rect 31334 1318 31386 1370
rect 32454 1318 32506 1370
rect 27134 1206 27186 1258
rect 27750 1158 27802 1210
rect 28142 1206 28194 1258
rect 28366 1206 28418 1258
rect 28590 1206 28642 1258
rect 28814 1206 28866 1258
rect 28926 1206 28978 1258
rect 29374 1206 29426 1258
rect 29766 1206 29818 1258
rect 33350 1268 33402 1320
rect 33518 1318 33570 1370
rect 34022 1318 34074 1370
rect 7870 1094 7922 1146
rect 19406 1094 19458 1146
rect 22094 1094 22146 1146
rect 26350 1094 26402 1146
rect 30102 1132 30154 1184
rect 30998 1162 31050 1214
rect 31502 1206 31554 1258
rect 31894 1132 31946 1184
rect 32790 1162 32842 1214
rect 33126 1150 33178 1202
rect 32230 1094 32282 1146
rect 34414 1094 34466 1146
rect 17502 982 17554 1034
rect 17950 982 18002 1034
rect 18174 982 18226 1034
rect 18398 982 18450 1034
rect 21646 982 21698 1034
rect 22318 982 22370 1034
rect 22542 982 22594 1034
rect 23102 982 23154 1034
rect 23774 982 23826 1034
rect 24222 982 24274 1034
rect 25006 982 25058 1034
rect 29486 982 29538 1034
rect 30718 982 30770 1034
rect 33854 982 33906 1034
rect 9094 758 9146 810
rect 9198 758 9250 810
rect 9302 758 9354 810
rect 17646 758 17698 810
rect 17750 758 17802 810
rect 17854 758 17906 810
rect 26198 758 26250 810
rect 26302 758 26354 810
rect 26406 758 26458 810
rect 20302 534 20354 586
rect 21646 534 21698 586
rect 22542 534 22594 586
rect 20974 422 21026 474
rect 22318 422 22370 474
<< metal2 >>
rect 2520 13200 2632 14000
rect 7672 13200 7784 14000
rect 12824 13200 12936 14000
rect 17976 13200 18088 14000
rect 23128 13200 23240 14000
rect 28280 13200 28392 14000
rect 33432 13200 33544 14000
rect 1820 12236 1876 12246
rect 1820 12142 1876 12180
rect 2548 12236 2604 13200
rect 4816 12572 5080 12582
rect 4872 12516 4920 12572
rect 4976 12516 5024 12572
rect 4816 12506 5080 12516
rect 2548 12122 2604 12180
rect 2548 12070 2550 12122
rect 2602 12070 2604 12122
rect 2548 12058 2604 12070
rect 6916 12346 6972 12358
rect 6916 12294 6918 12346
rect 6970 12294 6972 12346
rect 1932 12012 1988 12022
rect 2156 12012 2212 12022
rect 1932 12010 2212 12012
rect 1932 11958 1934 12010
rect 1986 11958 2158 12010
rect 2210 11958 2212 12010
rect 1932 11956 2212 11958
rect 1932 11946 2044 11956
rect 1092 11452 1148 11462
rect 1092 10618 1148 11396
rect 1372 11452 1428 11462
rect 1372 11358 1428 11396
rect 1708 11338 1764 11350
rect 1708 11286 1710 11338
rect 1762 11286 1764 11338
rect 1708 10892 1764 11286
rect 1708 10826 1764 10836
rect 1876 11226 1932 11238
rect 1876 11174 1878 11226
rect 1930 11174 1932 11226
rect 1876 10668 1932 11174
rect 1092 10566 1094 10618
rect 1146 10566 1148 10618
rect 1092 9838 1148 10566
rect 1596 10612 1932 10668
rect 1596 10610 1652 10612
rect 1596 10558 1598 10610
rect 1650 10558 1652 10610
rect 1596 10546 1652 10558
rect 1092 9786 1094 9838
rect 1146 9786 1148 9838
rect 1092 9772 1148 9786
rect 1540 10444 1596 10454
rect 1540 9838 1596 10388
rect 1540 9786 1542 9838
rect 1594 9786 1596 9838
rect 1540 9774 1596 9786
rect 1092 9716 1484 9772
rect 1428 9110 1484 9716
rect 1988 9660 2044 11946
rect 2156 11676 2212 11956
rect 5012 12010 5068 12022
rect 5012 11958 5014 12010
rect 5066 11958 5068 12010
rect 2156 11610 2212 11620
rect 2828 11676 2884 11686
rect 2828 11562 2884 11620
rect 2828 11510 2830 11562
rect 2882 11510 2884 11562
rect 2828 11498 2884 11510
rect 3892 11676 3948 11686
rect 5012 11676 5068 11958
rect 2604 11452 2660 11462
rect 1708 9604 2044 9660
rect 2212 11382 2268 11394
rect 2212 11330 2214 11382
rect 2266 11330 2268 11382
rect 2604 11358 2660 11396
rect 3276 11452 3332 11462
rect 3276 11358 3332 11396
rect 3668 11382 3724 11394
rect 3052 11340 3108 11350
rect 2212 9660 2268 11330
rect 1316 9100 1372 9110
rect 1428 9098 1540 9110
rect 1708 9100 1764 9604
rect 2212 9594 2268 9604
rect 2996 11338 3108 11340
rect 2996 11286 3054 11338
rect 3106 11286 3108 11338
rect 2996 11274 3108 11286
rect 3668 11330 3670 11382
rect 3722 11330 3724 11382
rect 2492 9548 2548 9558
rect 1428 9046 1486 9098
rect 1538 9046 1540 9098
rect 1428 9044 1540 9046
rect 980 8988 1036 8998
rect 980 8202 1036 8932
rect 1316 8886 1372 9044
rect 1316 8874 1428 8886
rect 1316 8822 1374 8874
rect 1426 8822 1428 8874
rect 1316 8820 1428 8822
rect 1372 8810 1428 8820
rect 1484 8652 1540 9044
rect 1484 8586 1540 8596
rect 1652 9098 1764 9100
rect 1652 9046 1710 9098
rect 1762 9046 1764 9098
rect 1652 9034 1764 9046
rect 1932 9100 1988 9110
rect 1652 8426 1708 9034
rect 1932 9006 1988 9044
rect 2492 9100 2548 9492
rect 2996 9548 3052 11274
rect 3668 10332 3724 11330
rect 3668 10266 3724 10276
rect 3892 11228 3948 11620
rect 4900 11620 5068 11676
rect 4340 11452 4396 11462
rect 4340 11382 4396 11396
rect 4004 11340 4060 11350
rect 4004 11246 4060 11284
rect 4340 11330 4342 11382
rect 4394 11330 4396 11382
rect 3892 10610 3948 11172
rect 3892 10558 3894 10610
rect 3946 10558 3948 10610
rect 4340 10668 4396 11330
rect 4788 11382 4844 11394
rect 4788 11340 4790 11382
rect 4842 11340 4844 11382
rect 4788 11274 4844 11284
rect 4900 11228 4956 11620
rect 6916 11564 6972 12294
rect 6916 11498 6972 11508
rect 7588 12010 7644 12022
rect 7588 11958 7590 12010
rect 7642 11958 7644 12010
rect 4900 11162 4956 11172
rect 7140 11450 7196 11462
rect 7140 11398 7142 11450
rect 7194 11398 7196 11450
rect 7140 11228 7196 11398
rect 7140 11162 7196 11172
rect 7588 11228 7644 11958
rect 7700 11788 7756 13200
rect 12404 12348 12460 12358
rect 12404 12254 12460 12292
rect 12852 12348 12908 13200
rect 13368 12572 13632 12582
rect 13424 12516 13472 12572
rect 13528 12516 13576 12572
rect 13368 12506 13632 12516
rect 12852 12282 12908 12292
rect 13356 12236 13412 12256
rect 13356 12178 13412 12180
rect 9940 12166 9996 12178
rect 9940 12114 9942 12166
rect 9994 12114 9996 12166
rect 7700 11722 7756 11732
rect 9092 11788 9356 11798
rect 9148 11732 9196 11788
rect 9252 11732 9300 11788
rect 9092 11722 9356 11732
rect 9940 11788 9996 12114
rect 10388 12166 10444 12178
rect 10388 12124 10390 12166
rect 10442 12124 10444 12166
rect 10388 12058 10444 12068
rect 10836 12122 10892 12134
rect 10836 12070 10838 12122
rect 10890 12070 10892 12122
rect 10668 12012 10724 12022
rect 10668 12010 10780 12012
rect 10668 11958 10670 12010
rect 10722 11958 10780 12010
rect 10668 11946 10780 11958
rect 9940 11722 9996 11732
rect 10276 11676 10332 11686
rect 8372 11564 8428 11574
rect 8372 11458 8374 11508
rect 8426 11458 8428 11508
rect 9940 11564 9996 11574
rect 7588 11162 7644 11172
rect 7812 11228 7868 11238
rect 7812 11226 7980 11228
rect 7812 11174 7814 11226
rect 7866 11174 7980 11226
rect 7812 11172 7980 11174
rect 7812 11162 7868 11172
rect 4816 11004 5080 11014
rect 4872 10948 4920 11004
rect 4976 10948 5024 11004
rect 4816 10938 5080 10948
rect 7252 11004 7308 11014
rect 5964 10892 6020 10902
rect 4340 10602 4396 10612
rect 5460 10724 5740 10780
rect 2996 9482 3052 9492
rect 3892 9882 3948 10558
rect 4788 10442 4844 10454
rect 4788 10390 4790 10442
rect 4842 10390 4844 10442
rect 4788 10220 4844 10390
rect 5068 10444 5124 10454
rect 5068 10350 5124 10388
rect 5180 10442 5236 10454
rect 5180 10390 5182 10442
rect 5234 10390 5236 10442
rect 4788 10154 4844 10164
rect 5180 10108 5236 10390
rect 5460 10332 5516 10724
rect 5684 10668 5740 10724
rect 5852 10668 5908 10678
rect 5684 10666 5908 10668
rect 5684 10614 5854 10666
rect 5906 10614 5908 10666
rect 5684 10612 5908 10614
rect 5012 10052 5236 10108
rect 5404 10276 5516 10332
rect 5572 10598 5628 10610
rect 5852 10602 5908 10612
rect 5964 10610 6020 10836
rect 6412 10668 6468 10678
rect 5572 10546 5574 10598
rect 5626 10546 5628 10598
rect 5964 10558 5966 10610
rect 6018 10558 6020 10610
rect 5964 10546 6020 10558
rect 6244 10610 6300 10622
rect 6244 10558 6246 10610
rect 6298 10558 6300 10610
rect 6412 10574 6468 10612
rect 7252 10622 7308 10948
rect 6916 10598 6972 10610
rect 5012 9996 5068 10052
rect 5404 10050 5460 10276
rect 5404 9998 5406 10050
rect 5458 9998 5460 10050
rect 5404 9986 5460 9998
rect 5012 9930 5068 9940
rect 4788 9884 4844 9894
rect 3892 9830 3894 9882
rect 3946 9830 3948 9882
rect 3108 9324 3164 9334
rect 3892 9324 3948 9830
rect 4676 9882 4844 9884
rect 4676 9830 4790 9882
rect 4842 9830 4844 9882
rect 4676 9828 4844 9830
rect 4564 9772 4620 9782
rect 4564 9678 4620 9716
rect 2492 9042 2548 9044
rect 2492 8990 2494 9042
rect 2546 8990 2548 9042
rect 2660 9100 2716 9138
rect 2660 9034 2716 9044
rect 2492 8968 2548 8990
rect 2660 8964 2716 8976
rect 2660 8912 2662 8964
rect 2714 8912 2716 8964
rect 2268 8874 2324 8886
rect 2268 8822 2270 8874
rect 2322 8822 2324 8874
rect 2268 8764 2324 8822
rect 2660 8876 2716 8912
rect 2660 8810 2716 8820
rect 2996 8876 3052 8886
rect 2996 8782 3052 8820
rect 2268 8698 2324 8708
rect 1652 8374 1654 8426
rect 1706 8374 1708 8426
rect 1652 8362 1708 8374
rect 2660 8652 2716 8662
rect 980 8150 982 8202
rect 1034 8150 1036 8202
rect 980 8138 1036 8150
rect 2660 7462 2716 8596
rect 2660 7410 2662 7462
rect 2714 7410 2716 7462
rect 3108 7486 3164 9268
rect 3668 9268 3948 9324
rect 3332 9024 3388 9036
rect 3332 8988 3334 9024
rect 3386 8988 3388 9024
rect 3332 8922 3388 8932
rect 3108 7434 3110 7486
rect 3162 7434 3164 7486
rect 3108 7422 3164 7434
rect 2660 6860 2716 7410
rect 2660 6794 2716 6804
rect 3500 7196 3556 7206
rect 3500 6860 3556 7140
rect 3500 6728 3556 6804
rect 2100 6678 2156 6690
rect 1092 6636 1148 6646
rect 1092 5893 1148 6580
rect 2100 6626 2102 6678
rect 2154 6626 2156 6678
rect 3668 6646 3724 9268
rect 4004 9210 4060 9222
rect 4004 9158 4006 9210
rect 4058 9158 4060 9210
rect 3892 9100 3948 9110
rect 3780 9042 3836 9054
rect 3780 8990 3782 9042
rect 3834 8990 3836 9042
rect 3780 8092 3836 8990
rect 3892 8886 3948 9044
rect 4004 9056 4060 9158
rect 4676 9100 4732 9828
rect 4788 9818 4844 9828
rect 5180 9884 5236 9894
rect 5180 9882 5292 9884
rect 5180 9830 5182 9882
rect 5234 9830 5292 9882
rect 5180 9818 5292 9830
rect 5124 9660 5180 9670
rect 5124 9566 5180 9604
rect 5236 9548 5292 9818
rect 4816 9436 5080 9446
rect 4872 9380 4920 9436
rect 4976 9380 5024 9436
rect 4816 9370 5080 9380
rect 5124 9212 5180 9222
rect 4844 9100 4900 9110
rect 4676 9098 4900 9100
rect 4004 9000 4116 9056
rect 4676 9046 4846 9098
rect 4898 9046 4900 9098
rect 4676 9044 4900 9046
rect 4844 9034 4900 9044
rect 5124 9048 5180 9156
rect 3892 8874 4004 8886
rect 3892 8822 3950 8874
rect 4002 8822 4004 8874
rect 3892 8820 4004 8822
rect 3948 8810 4004 8820
rect 4060 8652 4116 9000
rect 4956 8988 5012 8998
rect 4396 8930 4452 8942
rect 4396 8878 4398 8930
rect 4450 8878 4452 8930
rect 5124 8996 5126 9048
rect 5178 8996 5180 9048
rect 5124 8984 5180 8996
rect 4956 8894 5012 8932
rect 4004 8596 4116 8652
rect 4172 8818 4228 8830
rect 4172 8766 4174 8818
rect 4226 8766 4228 8818
rect 4004 8270 4060 8596
rect 4004 8218 4006 8270
rect 4058 8218 4060 8270
rect 4172 8316 4228 8766
rect 4396 8764 4452 8878
rect 5236 8876 5292 9492
rect 5572 9212 5628 10546
rect 6132 10444 6188 10454
rect 5740 10386 5796 10398
rect 5740 10334 5742 10386
rect 5794 10334 5796 10386
rect 5740 9884 5796 10334
rect 6132 10230 6188 10388
rect 5348 9156 5628 9212
rect 5684 9828 5740 9884
rect 5684 9752 5796 9828
rect 6076 10220 6188 10230
rect 6132 10164 6188 10220
rect 5852 9772 5908 9782
rect 5684 9212 5740 9752
rect 5852 9678 5908 9716
rect 6076 9660 6132 10164
rect 6244 9994 6300 10558
rect 6916 10546 6918 10598
rect 6970 10546 6972 10598
rect 7252 10570 7254 10622
rect 7306 10570 7308 10622
rect 7756 10610 7812 10622
rect 7252 10558 7308 10570
rect 7476 10598 7532 10610
rect 6916 10108 6972 10546
rect 7476 10546 7478 10598
rect 7530 10546 7532 10598
rect 7756 10558 7758 10610
rect 7810 10558 7812 10610
rect 7756 10556 7812 10558
rect 7476 10444 7532 10546
rect 7476 10378 7532 10388
rect 7700 10500 7812 10556
rect 7252 10360 7308 10372
rect 7252 10308 7254 10360
rect 7306 10308 7308 10360
rect 7252 10220 7308 10308
rect 7252 10154 7308 10164
rect 7532 10220 7588 10230
rect 6916 10042 6972 10052
rect 7140 10108 7196 10118
rect 7140 10006 7196 10052
rect 6244 9942 6246 9994
rect 6298 9942 6300 9994
rect 6244 9930 6300 9942
rect 6468 9996 6524 10006
rect 6468 9842 6524 9940
rect 6468 9790 6470 9842
rect 6522 9790 6524 9842
rect 6636 9996 6692 10006
rect 6636 9882 6692 9940
rect 7084 9994 7196 10006
rect 7084 9942 7086 9994
rect 7138 9942 7196 9994
rect 7532 10050 7588 10164
rect 7700 10108 7756 10500
rect 7532 9998 7534 10050
rect 7586 9998 7588 10050
rect 7532 9986 7588 9998
rect 7644 10052 7756 10108
rect 7924 10108 7980 11172
rect 8372 11116 8428 11458
rect 8708 11452 8764 11462
rect 8708 11358 8764 11396
rect 9940 11412 9996 11508
rect 9940 11360 9942 11412
rect 9994 11360 9996 11412
rect 9436 11340 9492 11350
rect 9436 11246 9492 11284
rect 9100 11228 9156 11238
rect 9100 11134 9156 11172
rect 8372 11050 8428 11060
rect 9548 10780 9604 10790
rect 9940 10780 9996 11360
rect 8036 10722 8092 10734
rect 8036 10670 8038 10722
rect 8090 10670 8092 10722
rect 9548 10686 9604 10724
rect 9828 10724 9996 10780
rect 10276 11226 10332 11620
rect 10500 11564 10556 11574
rect 10500 11394 10556 11508
rect 10500 11342 10502 11394
rect 10554 11342 10556 11394
rect 10500 11330 10556 11342
rect 10612 11452 10668 11462
rect 10276 11174 10278 11226
rect 10330 11174 10332 11226
rect 10612 11288 10668 11396
rect 10612 11236 10614 11288
rect 10666 11236 10668 11288
rect 10612 11224 10668 11236
rect 8036 10556 8092 10670
rect 8764 10668 8820 10678
rect 8764 10574 8820 10612
rect 9436 10610 9492 10622
rect 8036 10490 8092 10500
rect 8988 10556 9044 10566
rect 9436 10558 9438 10610
rect 9490 10558 9492 10610
rect 9436 10556 9492 10558
rect 9828 10556 9884 10724
rect 9436 10500 9884 10556
rect 8988 10462 9044 10500
rect 9156 10444 9212 10454
rect 7644 9994 7700 10052
rect 7924 10042 7980 10052
rect 8092 10386 8148 10398
rect 8092 10334 8094 10386
rect 8146 10334 8148 10386
rect 7084 9940 7196 9942
rect 7644 9942 7646 9994
rect 7698 9942 7700 9994
rect 7084 9930 7140 9940
rect 7644 9930 7700 9942
rect 8092 9996 8148 10334
rect 8316 10386 8372 10398
rect 8316 10334 8318 10386
rect 8370 10334 8372 10386
rect 9156 10350 9212 10388
rect 8316 10220 8372 10334
rect 9092 10220 9356 10230
rect 8316 10164 8428 10220
rect 8092 9930 8148 9940
rect 6636 9830 6638 9882
rect 6690 9830 6692 9882
rect 6636 9818 6692 9830
rect 6972 9884 7028 9894
rect 6972 9790 7028 9828
rect 7756 9882 7812 9894
rect 7756 9830 7758 9882
rect 7810 9830 7812 9882
rect 6076 9658 6244 9660
rect 6076 9606 6078 9658
rect 6130 9606 6244 9658
rect 6076 9604 6244 9606
rect 6076 9594 6132 9604
rect 5852 9212 5908 9222
rect 5684 9210 5908 9212
rect 5684 9158 5854 9210
rect 5906 9158 5908 9210
rect 5684 9156 5908 9158
rect 5348 9042 5404 9156
rect 5348 8990 5350 9042
rect 5402 8990 5404 9042
rect 5348 8978 5404 8990
rect 5460 8988 5516 8998
rect 5460 8876 5516 8932
rect 4396 8698 4452 8708
rect 4732 8818 4788 8830
rect 4732 8766 4734 8818
rect 4786 8766 4788 8818
rect 5236 8810 5292 8820
rect 5404 8820 5516 8876
rect 4732 8652 4788 8766
rect 4732 8316 4788 8596
rect 5404 8370 5460 8820
rect 5404 8318 5406 8370
rect 5458 8318 5460 8370
rect 5572 8428 5628 9156
rect 5852 9146 5908 9156
rect 6188 9212 6244 9604
rect 6468 9436 6524 9790
rect 7084 9770 7140 9782
rect 7084 9718 7086 9770
rect 7138 9718 7140 9770
rect 7084 9660 7140 9718
rect 7476 9772 7532 9782
rect 7084 9604 7196 9660
rect 6468 9370 6524 9380
rect 6972 9436 7028 9446
rect 6188 9080 6244 9156
rect 6524 9100 6580 9110
rect 5908 9034 5964 9046
rect 5908 8988 5910 9034
rect 5962 8988 5964 9034
rect 6524 9006 6580 9044
rect 6972 9098 7028 9380
rect 6972 9046 6974 9098
rect 7026 9046 7028 9098
rect 6972 9034 7028 9046
rect 5908 8922 5964 8932
rect 6860 8988 6916 8998
rect 5572 8362 5628 8372
rect 4732 8260 5236 8316
rect 5404 8306 5460 8318
rect 6860 8314 6916 8932
rect 7140 8876 7196 9604
rect 7252 9212 7308 9222
rect 7252 9118 7308 9156
rect 7476 9210 7532 9716
rect 7756 9772 7812 9830
rect 7756 9706 7812 9716
rect 7924 9820 7980 9832
rect 7924 9768 7926 9820
rect 7978 9768 7980 9820
rect 7476 9158 7478 9210
rect 7530 9158 7532 9210
rect 7476 9146 7532 9158
rect 7700 9436 7756 9446
rect 7700 9210 7756 9380
rect 7700 9158 7702 9210
rect 7754 9158 7756 9210
rect 7700 9146 7756 9158
rect 7140 8810 7196 8820
rect 7924 8876 7980 9768
rect 8260 9826 8316 9838
rect 8260 9774 8262 9826
rect 8314 9774 8316 9826
rect 8260 9772 8316 9774
rect 8260 9706 8316 9716
rect 8372 9100 8428 10164
rect 9148 10164 9196 10220
rect 9252 10164 9300 10220
rect 9092 10154 9356 10164
rect 9828 10006 9884 10500
rect 9940 10598 9996 10610
rect 9940 10546 9942 10598
rect 9994 10546 9996 10598
rect 9940 10220 9996 10546
rect 9940 10154 9996 10164
rect 8484 9996 8596 10006
rect 8876 9996 8932 10006
rect 8540 9994 8596 9996
rect 8540 9942 8542 9994
rect 8594 9942 8596 9994
rect 8540 9940 8596 9942
rect 8484 9930 8596 9940
rect 8820 9940 8876 9996
rect 8820 9902 8932 9940
rect 9772 9994 9884 10006
rect 9772 9942 9774 9994
rect 9826 9942 9884 9994
rect 9772 9940 9884 9942
rect 10276 9996 10332 11174
rect 10724 10780 10780 11946
rect 10836 11564 10892 12070
rect 11844 12124 11900 12134
rect 10836 11498 10892 11508
rect 11004 12010 11060 12022
rect 11004 11958 11006 12010
rect 11058 11958 11060 12010
rect 11004 11676 11060 11958
rect 11396 12012 11452 12022
rect 11396 11918 11452 11956
rect 11732 12010 11788 12022
rect 11732 11958 11734 12010
rect 11786 11958 11788 12010
rect 11004 11452 11060 11620
rect 11172 11788 11228 11798
rect 11172 11562 11228 11732
rect 11732 11788 11788 11958
rect 11732 11722 11788 11732
rect 11844 11574 11900 12068
rect 13356 12126 13358 12178
rect 13410 12126 13412 12178
rect 14756 12166 14812 12178
rect 12068 12010 12124 12022
rect 12068 11958 12070 12010
rect 12122 11958 12124 12010
rect 12068 11676 12124 11958
rect 13020 12012 13076 12022
rect 13020 11918 13076 11956
rect 13188 12012 13244 12022
rect 12068 11610 12124 11620
rect 11172 11510 11174 11562
rect 11226 11510 11228 11562
rect 11172 11498 11228 11510
rect 11396 11564 11452 11574
rect 11004 11386 11060 11396
rect 10892 11228 10948 11238
rect 10892 11226 11004 11228
rect 10892 11174 10894 11226
rect 10946 11174 11004 11226
rect 10892 11162 11004 11174
rect 10724 10714 10780 10724
rect 10612 10598 10668 10610
rect 10612 10546 10614 10598
rect 10666 10546 10668 10598
rect 10612 10444 10668 10546
rect 10612 10378 10668 10388
rect 10948 10556 11004 11162
rect 9772 9930 9828 9940
rect 10276 9930 10332 9940
rect 10556 9996 10612 10006
rect 10948 9996 11004 10500
rect 11396 10108 11452 11508
rect 11788 11562 11900 11574
rect 11788 11510 11790 11562
rect 11842 11510 11900 11562
rect 11788 11508 11900 11510
rect 11956 11564 12012 11574
rect 11788 11498 11844 11508
rect 11956 11452 12012 11508
rect 12852 11564 12908 11574
rect 12068 11452 12124 11462
rect 11956 11450 12124 11452
rect 11956 11398 12070 11450
rect 12122 11398 12124 11450
rect 11956 11396 12124 11398
rect 11508 11382 11564 11394
rect 12068 11386 12124 11396
rect 11508 11340 11510 11382
rect 11562 11340 11564 11382
rect 11508 11274 11564 11284
rect 12404 11382 12460 11394
rect 12404 11330 12406 11382
rect 12458 11330 12460 11382
rect 12404 10780 12460 11330
rect 12404 10714 12460 10724
rect 12852 10526 12908 11508
rect 13188 11452 13244 11956
rect 13356 11900 13412 12126
rect 13748 12124 13804 12134
rect 13356 11834 13412 11844
rect 13636 12122 13804 12124
rect 13636 12070 13750 12122
rect 13802 12070 13804 12122
rect 13636 12068 13804 12070
rect 13636 11564 13692 12068
rect 13748 12058 13804 12068
rect 14084 12124 14140 12134
rect 14084 12024 14086 12068
rect 14138 12024 14140 12068
rect 14084 12012 14140 12024
rect 14756 12114 14758 12166
rect 14810 12114 14812 12166
rect 14588 12012 14644 12022
rect 14756 12012 14812 12114
rect 15316 12166 15372 12178
rect 15316 12124 15318 12166
rect 15370 12124 15372 12166
rect 15316 12058 15372 12068
rect 15988 12124 16044 12134
rect 14588 12010 14700 12012
rect 14588 11958 14590 12010
rect 14642 11958 14700 12010
rect 14588 11946 14700 11958
rect 14756 11946 14812 11956
rect 14420 11900 14476 11910
rect 13636 11498 13692 11508
rect 13804 11788 13860 11798
rect 13804 11506 13860 11732
rect 12852 10474 12854 10526
rect 12906 10474 12908 10526
rect 12852 10462 12908 10474
rect 12964 11396 13244 11452
rect 13804 11454 13806 11506
rect 13858 11454 13860 11506
rect 13804 11442 13860 11454
rect 13972 11564 14028 11574
rect 11396 10052 11508 10108
rect 11172 9996 11228 10006
rect 10556 9994 10892 9996
rect 10556 9942 10558 9994
rect 10610 9942 10892 9994
rect 10556 9940 10892 9942
rect 10948 9994 11228 9996
rect 10948 9942 11174 9994
rect 11226 9942 11228 9994
rect 10948 9940 11228 9942
rect 10556 9930 10612 9940
rect 8708 9882 8764 9894
rect 8708 9830 8710 9882
rect 8762 9830 8764 9882
rect 8708 9660 8764 9830
rect 8708 9594 8764 9604
rect 8820 9212 8876 9902
rect 9212 9884 9268 9894
rect 8820 9146 8876 9156
rect 9044 9324 9100 9334
rect 9044 9154 9100 9268
rect 8372 9034 8428 9044
rect 8596 9100 8652 9110
rect 9044 9102 9046 9154
rect 9098 9102 9100 9154
rect 9044 9090 9100 9102
rect 9212 9100 9268 9828
rect 10108 9884 10164 9894
rect 10108 9882 10220 9884
rect 10108 9830 10110 9882
rect 10162 9830 10220 9882
rect 10108 9818 10220 9830
rect 10164 9772 10220 9818
rect 9436 9658 9492 9670
rect 10052 9660 10108 9670
rect 9436 9606 9438 9658
rect 9490 9606 9492 9658
rect 9436 9548 9492 9606
rect 9436 9482 9492 9492
rect 9940 9658 10108 9660
rect 9940 9606 10054 9658
rect 10106 9606 10108 9658
rect 9940 9604 10108 9606
rect 8596 8986 8652 9044
rect 9940 9056 9996 9604
rect 10052 9594 10108 9604
rect 9212 9034 9268 9044
rect 9660 9042 9996 9056
rect 8596 8934 8598 8986
rect 8650 8934 8652 8986
rect 9660 8990 9662 9042
rect 9714 9000 9996 9042
rect 10164 9324 10220 9716
rect 10332 9826 10388 9838
rect 10332 9774 10334 9826
rect 10386 9774 10388 9826
rect 10332 9324 10388 9774
rect 10164 9042 10220 9268
rect 10276 9268 10388 9324
rect 10724 9806 10780 9818
rect 10724 9754 10726 9806
rect 10778 9754 10780 9806
rect 10276 9212 10332 9268
rect 10556 9212 10612 9222
rect 10276 9146 10332 9156
rect 10388 9210 10612 9212
rect 10388 9158 10558 9210
rect 10610 9158 10612 9210
rect 10388 9156 10612 9158
rect 9714 8990 9716 9000
rect 9660 8978 9716 8990
rect 10164 8990 10166 9042
rect 10218 8990 10220 9042
rect 10164 8978 10220 8990
rect 8596 8922 8652 8934
rect 7924 8810 7980 8820
rect 8036 8874 8092 8886
rect 8204 8876 8260 8886
rect 8428 8876 8484 8886
rect 8036 8822 8038 8874
rect 8090 8822 8092 8874
rect 8036 8764 8092 8822
rect 8036 8698 8092 8708
rect 8148 8874 8260 8876
rect 8148 8822 8206 8874
rect 8258 8822 8260 8874
rect 8148 8810 8260 8822
rect 8372 8874 8484 8876
rect 8372 8822 8430 8874
rect 8482 8822 8484 8874
rect 8372 8810 8484 8822
rect 8764 8876 8820 8886
rect 9100 8876 9156 8886
rect 8764 8874 8876 8876
rect 8764 8822 8766 8874
rect 8818 8822 8876 8874
rect 8764 8810 8876 8822
rect 8148 8540 8204 8810
rect 8372 8540 8428 8810
rect 7700 8484 8204 8540
rect 8260 8484 8428 8540
rect 7476 8372 7644 8428
rect 7476 8336 7532 8372
rect 4172 8250 4228 8260
rect 4004 8206 4060 8218
rect 4564 8246 4620 8258
rect 3780 8026 3836 8036
rect 4564 8194 4566 8246
rect 4618 8194 4620 8246
rect 4004 7532 4060 7542
rect 4004 6646 4060 7476
rect 4172 7196 4228 7206
rect 4172 6858 4228 7140
rect 4172 6806 4174 6858
rect 4226 6806 4228 6858
rect 4172 6794 4228 6806
rect 4564 7196 4620 8194
rect 4788 8092 4844 8130
rect 4788 8026 4844 8036
rect 5180 8034 5236 8260
rect 6860 8262 6862 8314
rect 6914 8262 6916 8314
rect 6020 8246 6076 8258
rect 6860 8250 6916 8262
rect 7028 8316 7084 8326
rect 7476 8284 7478 8336
rect 7530 8284 7532 8336
rect 7476 8272 7532 8284
rect 6020 8194 6022 8246
rect 6074 8194 6076 8246
rect 7028 8214 7084 8260
rect 5684 8092 5740 8102
rect 5180 7982 5182 8034
rect 5234 7982 5236 8034
rect 4816 7868 5080 7878
rect 4872 7812 4920 7868
rect 4976 7812 5024 7868
rect 4816 7802 5080 7812
rect 5180 7532 5236 7982
rect 5180 7466 5236 7476
rect 5572 8090 5740 8092
rect 5572 8038 5686 8090
rect 5738 8038 5740 8090
rect 5572 8036 5740 8038
rect 1764 6522 1820 6534
rect 1764 6470 1766 6522
rect 1818 6470 1820 6522
rect 1764 5918 1820 6470
rect 1092 5841 1094 5893
rect 1146 5841 1148 5893
rect 1708 5906 1820 5918
rect 1708 5854 1710 5906
rect 1762 5858 1820 5906
rect 1762 5854 1764 5858
rect 1708 5842 1764 5854
rect 1092 5110 1148 5841
rect 1092 5058 1094 5110
rect 1146 5058 1148 5110
rect 1092 4340 1148 5058
rect 1540 5110 1596 5122
rect 1540 5058 1542 5110
rect 1594 5058 1596 5110
rect 1092 4326 1260 4340
rect 1092 4284 1206 4326
rect 1204 4274 1206 4284
rect 1258 4274 1260 4326
rect 1092 3052 1148 3062
rect 1204 3052 1260 4274
rect 1540 3836 1596 5058
rect 2100 4844 2156 6626
rect 3276 6636 3332 6646
rect 3668 6636 3780 6646
rect 3668 6634 3836 6636
rect 3668 6582 3726 6634
rect 3778 6582 3836 6634
rect 3668 6580 3836 6582
rect 3276 6542 3332 6580
rect 3724 6570 3836 6580
rect 3948 6634 4060 6646
rect 4564 6702 4620 7140
rect 4564 6650 4566 6702
rect 4618 6650 4620 6702
rect 4564 6638 4620 6650
rect 4676 7308 4732 7318
rect 3948 6582 3950 6634
rect 4002 6582 4060 6634
rect 3948 6580 4060 6582
rect 3948 6570 4004 6580
rect 3780 5896 3836 6570
rect 3892 5896 3948 5906
rect 3780 5894 3948 5896
rect 3780 5842 3894 5894
rect 3946 5842 3948 5894
rect 3780 5840 3948 5842
rect 3892 5516 3948 5840
rect 4676 5516 4732 7252
rect 5460 7308 5516 7318
rect 5460 7214 5516 7252
rect 5572 6748 5628 8036
rect 5684 8026 5740 8036
rect 6020 7644 6076 8194
rect 6300 8204 6356 8214
rect 6524 8204 6580 8214
rect 6300 8202 6580 8204
rect 6300 8150 6302 8202
rect 6354 8150 6526 8202
rect 6578 8150 6580 8202
rect 6300 8148 6580 8150
rect 6300 8138 6412 8148
rect 6524 8138 6580 8148
rect 6972 8202 7084 8214
rect 6972 8150 6974 8202
rect 7026 8150 7084 8202
rect 6972 8138 7084 8150
rect 6020 7578 6076 7588
rect 6132 8092 6188 8102
rect 6132 7642 6188 8036
rect 6132 7590 6134 7642
rect 6186 7590 6188 7642
rect 6132 7578 6188 7590
rect 6356 7318 6412 8138
rect 7028 7318 7084 8138
rect 7308 8258 7364 8270
rect 7308 8206 7310 8258
rect 7362 8206 7364 8258
rect 7308 7756 7364 8206
rect 7476 8202 7532 8214
rect 7476 8150 7478 8202
rect 7530 8150 7532 8202
rect 7476 7868 7532 8150
rect 7588 7980 7644 8372
rect 7700 8316 7756 8484
rect 8036 8372 8204 8428
rect 8036 8336 8092 8372
rect 8036 8284 8038 8336
rect 8090 8284 8092 8336
rect 8036 8272 8092 8284
rect 7700 8250 7756 8260
rect 7868 8258 7924 8270
rect 7868 8206 7870 8258
rect 7922 8206 7924 8258
rect 7868 8204 7924 8206
rect 7868 8138 7924 8148
rect 8036 8204 8092 8214
rect 8036 8110 8092 8148
rect 7588 7924 8092 7980
rect 7476 7812 7756 7868
rect 7252 7700 7364 7756
rect 6356 7308 6468 7318
rect 6356 7252 6412 7308
rect 6412 7214 6468 7252
rect 6860 7306 6916 7318
rect 6860 7254 6862 7306
rect 6914 7254 6916 7306
rect 6860 7196 6916 7254
rect 7028 7308 7140 7318
rect 7028 7252 7084 7308
rect 6860 7130 6916 7140
rect 5180 6692 5628 6748
rect 7084 6748 7140 7252
rect 5180 6690 5236 6692
rect 5180 6638 5182 6690
rect 5234 6638 5236 6690
rect 7084 6682 7140 6692
rect 5180 6626 5236 6638
rect 4816 6300 5080 6310
rect 4872 6244 4920 6300
rect 4976 6244 5024 6300
rect 4816 6234 5080 6244
rect 7140 6188 7196 6198
rect 6244 6076 6300 6086
rect 6244 6018 6300 6020
rect 6244 5966 6246 6018
rect 6298 5966 6300 6018
rect 6244 5954 6300 5966
rect 6468 5964 6524 5974
rect 6468 5866 6470 5908
rect 6522 5866 6524 5908
rect 6188 5852 6244 5862
rect 6468 5854 6524 5866
rect 7140 5918 7196 6132
rect 7140 5866 7142 5918
rect 7194 5866 7196 5918
rect 6188 5758 6244 5796
rect 6972 5850 7028 5862
rect 7140 5854 7196 5866
rect 6972 5798 6974 5850
rect 7026 5798 7028 5850
rect 4900 5740 4956 5750
rect 5180 5740 5236 5750
rect 4900 5738 5236 5740
rect 4900 5686 4902 5738
rect 4954 5686 5182 5738
rect 5234 5686 5236 5738
rect 4900 5684 5236 5686
rect 4900 5674 4956 5684
rect 3892 5460 4900 5516
rect 3892 5290 3948 5460
rect 3892 5238 3894 5290
rect 3946 5238 3948 5290
rect 3892 5226 3948 5238
rect 2100 4778 2156 4788
rect 1764 4508 1820 4518
rect 1764 4350 1820 4452
rect 1764 4298 1766 4350
rect 1818 4298 1820 4350
rect 1764 4286 1820 4298
rect 1540 3770 1596 3780
rect 2212 4284 2268 4294
rect 4116 4284 4172 5460
rect 4844 5290 4900 5460
rect 4844 5238 4846 5290
rect 4898 5238 4900 5290
rect 4844 5226 4900 5238
rect 5180 5178 5236 5684
rect 5572 5740 5628 5750
rect 6972 5740 7028 5798
rect 5572 5646 5628 5684
rect 5964 5682 6020 5694
rect 5964 5630 5966 5682
rect 6018 5630 6020 5682
rect 5964 5404 6020 5630
rect 6692 5684 7028 5740
rect 6076 5404 6132 5414
rect 5964 5348 6076 5404
rect 6076 5346 6132 5348
rect 5572 5292 5628 5302
rect 6076 5294 6078 5346
rect 6130 5294 6132 5346
rect 6076 5282 6132 5294
rect 5180 5126 5182 5178
rect 5234 5126 5236 5178
rect 5180 5114 5236 5126
rect 5348 5180 5404 5190
rect 5348 5016 5404 5124
rect 2212 3734 2268 4228
rect 2156 3722 2268 3734
rect 2156 3670 2158 3722
rect 2210 3670 2268 3722
rect 2156 3668 2268 3670
rect 3724 4282 4172 4284
rect 3724 4230 4118 4282
rect 4170 4230 4172 4282
rect 3724 4228 4172 4230
rect 3724 3724 3780 4228
rect 4116 4218 4172 4228
rect 4564 4954 4620 4966
rect 4564 4902 4566 4954
rect 4618 4902 4620 4954
rect 4172 3948 4228 3958
rect 4060 3724 4116 3734
rect 3724 3722 3948 3724
rect 3724 3670 3726 3722
rect 3778 3670 3948 3722
rect 3724 3668 3948 3670
rect 2156 3658 2212 3668
rect 3724 3658 3780 3668
rect 2884 3542 2940 3554
rect 2884 3490 2886 3542
rect 2938 3490 2940 3542
rect 1764 3388 1820 3398
rect 1148 2996 1260 3052
rect 1540 3386 1820 3388
rect 1540 3334 1766 3386
rect 1818 3334 1820 3386
rect 1540 3332 1820 3334
rect 1092 1998 1148 2996
rect 1092 1946 1094 1998
rect 1146 1946 1148 1998
rect 1092 1934 1148 1946
rect 1540 1998 1596 3332
rect 1764 3322 1820 3332
rect 2548 3386 2604 3398
rect 2548 3334 2550 3386
rect 2602 3334 2604 3386
rect 2100 3052 2156 3062
rect 2100 2778 2156 2996
rect 2100 2726 2102 2778
rect 2154 2726 2156 2778
rect 2548 2828 2604 3334
rect 2884 2940 2940 3490
rect 3500 3498 3556 3510
rect 3500 3446 3502 3498
rect 3554 3446 3556 3498
rect 3500 3387 3556 3446
rect 3500 3331 3612 3387
rect 2884 2874 2940 2884
rect 3556 3052 3612 3331
rect 2548 2772 2660 2828
rect 2100 2714 2156 2726
rect 2604 2770 2660 2772
rect 2604 2718 2606 2770
rect 2658 2718 2660 2770
rect 2604 2706 2660 2718
rect 3556 2492 3612 2996
rect 3556 2426 3612 2436
rect 1540 1946 1542 1998
rect 1594 1946 1596 1998
rect 1540 1934 1596 1946
rect 3892 2042 3948 3668
rect 4060 3630 4116 3668
rect 4172 3722 4228 3892
rect 4172 3670 4174 3722
rect 4226 3670 4228 3722
rect 4172 3658 4228 3670
rect 4564 3724 4620 4902
rect 4676 4956 4732 4966
rect 5348 4964 5350 5016
rect 5402 4964 5404 5016
rect 5348 4952 5404 4964
rect 5460 5114 5516 5126
rect 5460 5062 5462 5114
rect 5514 5062 5516 5114
rect 5460 4956 5516 5062
rect 4676 4172 4732 4900
rect 5460 4890 5516 4900
rect 4816 4732 5080 4742
rect 5572 4732 5628 5236
rect 5852 5180 5908 5190
rect 5852 5178 5964 5180
rect 5852 5126 5854 5178
rect 5906 5126 5964 5178
rect 5852 5114 5964 5126
rect 4872 4676 4920 4732
rect 4976 4676 5024 4732
rect 4816 4666 5080 4676
rect 5236 4676 5628 4732
rect 5796 5010 5852 5022
rect 5796 4958 5798 5010
rect 5850 4958 5852 5010
rect 4788 4506 4844 4518
rect 4788 4454 4790 4506
rect 4842 4454 4844 4506
rect 4788 4396 4844 4454
rect 4788 4330 4844 4340
rect 5236 4394 5292 4676
rect 5796 4508 5852 4958
rect 5908 4508 5964 5114
rect 6356 5110 6412 5122
rect 6356 5068 6358 5110
rect 6410 5068 6412 5110
rect 6356 5002 6412 5012
rect 6692 5110 6748 5684
rect 7252 5628 7308 7700
rect 7532 7644 7588 7654
rect 7532 7550 7588 7588
rect 7364 6774 7420 6786
rect 7364 6748 7366 6774
rect 7418 6748 7420 6774
rect 7364 6682 7420 6692
rect 7700 6636 7756 7812
rect 7868 7756 7924 7766
rect 7868 7698 7924 7700
rect 7868 7646 7870 7698
rect 7922 7646 7924 7698
rect 7868 7634 7924 7646
rect 7700 6570 7756 6580
rect 8036 6188 8092 7924
rect 7756 6132 8092 6188
rect 7756 6076 7812 6132
rect 7700 6074 7812 6076
rect 7700 6022 7758 6074
rect 7810 6022 7812 6074
rect 7700 6010 7812 6022
rect 7532 5850 7588 5862
rect 7532 5798 7534 5850
rect 7586 5798 7588 5850
rect 6860 5572 7308 5628
rect 7364 5738 7420 5750
rect 7532 5740 7588 5798
rect 7364 5686 7366 5738
rect 7418 5686 7420 5738
rect 6860 5346 6916 5572
rect 6860 5294 6862 5346
rect 6914 5294 6916 5346
rect 6860 5180 6916 5294
rect 7084 5180 7140 5190
rect 6860 5114 6916 5124
rect 7028 5178 7140 5180
rect 7028 5126 7086 5178
rect 7138 5126 7140 5178
rect 7028 5114 7140 5126
rect 7252 5180 7308 5190
rect 6692 5058 6694 5110
rect 6746 5058 6748 5110
rect 6244 4620 6300 4630
rect 6076 4508 6132 4518
rect 5908 4506 6132 4508
rect 5908 4454 6078 4506
rect 6130 4454 6132 4506
rect 5908 4452 6132 4454
rect 5796 4442 5852 4452
rect 6076 4442 6132 4452
rect 5236 4342 5238 4394
rect 5290 4342 5292 4394
rect 5236 4330 5292 4342
rect 5684 4396 5740 4406
rect 5684 4338 5740 4340
rect 5684 4286 5686 4338
rect 5738 4286 5740 4338
rect 5236 4260 5292 4272
rect 5236 4208 5238 4260
rect 5290 4208 5292 4260
rect 5068 4172 5124 4182
rect 5236 4172 5292 4208
rect 4676 4116 4956 4172
rect 4564 3592 4620 3668
rect 4900 3722 4956 4116
rect 5068 4170 5180 4172
rect 5068 4118 5070 4170
rect 5122 4118 5180 4170
rect 5068 4106 5180 4118
rect 5236 4106 5292 4116
rect 4900 3670 4902 3722
rect 4954 3670 4956 3722
rect 4900 3658 4956 3670
rect 5124 3388 5180 4106
rect 5124 3322 5180 3332
rect 5460 3542 5516 3554
rect 5460 3490 5462 3542
rect 5514 3490 5516 3542
rect 4816 3164 5080 3174
rect 4872 3108 4920 3164
rect 4976 3108 5024 3164
rect 4816 3098 5080 3108
rect 4844 2658 4900 2670
rect 4844 2606 4846 2658
rect 4898 2606 4900 2658
rect 4844 2604 4900 2606
rect 3892 1990 3894 2042
rect 3946 1990 3948 2042
rect 3892 1932 3948 1990
rect 4788 2548 4900 2604
rect 4788 1942 4844 2548
rect 5348 2492 5404 2502
rect 4956 2156 5012 2166
rect 5348 2156 5404 2436
rect 4956 2154 5404 2156
rect 4956 2102 4958 2154
rect 5010 2102 5404 2154
rect 4956 2100 5404 2102
rect 4956 2090 5012 2100
rect 5348 1942 5404 2100
rect 5460 2156 5516 3490
rect 5684 3052 5740 4286
rect 6020 4340 6076 4350
rect 6244 4340 6300 4564
rect 6692 4620 6748 5058
rect 6692 4554 6748 4564
rect 6916 4956 6972 4966
rect 6916 4732 6972 4900
rect 6020 4338 6300 4340
rect 6020 4286 6022 4338
rect 6074 4286 6300 4338
rect 6020 4284 6300 4286
rect 6020 4274 6076 4284
rect 6916 4282 6972 4676
rect 6916 4230 6918 4282
rect 6970 4230 6972 4282
rect 6916 4218 6972 4230
rect 6188 4114 6244 4126
rect 6188 4062 6190 4114
rect 6242 4062 6244 4114
rect 6188 3836 6244 4062
rect 6188 3770 6244 3780
rect 6412 4114 6468 4126
rect 7028 4116 7084 5114
rect 7140 4998 7196 5010
rect 7140 4946 7142 4998
rect 7194 4956 7196 4998
rect 7252 4956 7308 5124
rect 7364 5122 7420 5686
rect 7364 5070 7366 5122
rect 7418 5070 7420 5122
rect 7364 5058 7420 5070
rect 7476 5684 7532 5740
rect 7476 5674 7588 5684
rect 7194 4946 7308 4956
rect 7140 4900 7308 4946
rect 7476 4844 7532 5674
rect 7700 5516 7756 6010
rect 8036 5740 8092 6132
rect 8036 5674 8092 5684
rect 8148 5964 8204 8372
rect 8260 8204 8316 8484
rect 8428 8316 8484 8326
rect 8428 8222 8484 8260
rect 8708 8258 8764 8270
rect 8260 7418 8316 8148
rect 8708 8206 8710 8258
rect 8762 8206 8764 8258
rect 8708 8092 8764 8206
rect 8708 8026 8764 8036
rect 8820 7980 8876 8810
rect 8932 8874 9156 8876
rect 8932 8822 9102 8874
rect 9154 8822 9156 8874
rect 8932 8820 9156 8822
rect 8932 8092 8988 8820
rect 9100 8810 9156 8820
rect 9324 8876 9380 8886
rect 9324 8782 9380 8820
rect 9772 8874 9828 8886
rect 9772 8822 9774 8874
rect 9826 8822 9828 8874
rect 9092 8652 9356 8662
rect 9148 8596 9196 8652
rect 9252 8596 9300 8652
rect 9092 8586 9356 8596
rect 9772 8540 9828 8822
rect 9772 8474 9828 8484
rect 9044 8428 9100 8438
rect 10388 8428 10444 9156
rect 10556 9146 10612 9156
rect 10724 9056 10780 9754
rect 10836 9548 10892 9940
rect 11172 9930 11228 9940
rect 11284 9996 11340 10006
rect 11284 9782 11340 9940
rect 11228 9772 11340 9782
rect 11172 9770 11340 9772
rect 11172 9718 11230 9770
rect 11282 9718 11340 9770
rect 11172 9716 11340 9718
rect 11452 9826 11508 10052
rect 12964 9996 13020 11396
rect 13132 11394 13188 11396
rect 13132 11342 13134 11394
rect 13186 11342 13188 11394
rect 13132 11330 13188 11342
rect 13972 11116 14028 11508
rect 13368 11004 13632 11014
rect 13424 10948 13472 11004
rect 13528 10948 13576 11004
rect 13368 10938 13632 10948
rect 13804 10780 13860 10790
rect 13804 10686 13860 10724
rect 13972 10332 14028 11060
rect 14196 11340 14252 11350
rect 14196 11116 14252 11284
rect 14196 11050 14252 11060
rect 14420 10778 14476 11844
rect 14644 10892 14700 11946
rect 14644 10826 14700 10836
rect 14756 11564 14812 11574
rect 14420 10726 14422 10778
rect 14474 10726 14476 10778
rect 14420 10714 14476 10726
rect 14084 10556 14140 10566
rect 14084 10462 14140 10500
rect 14756 10554 14812 11508
rect 15988 11562 16044 12068
rect 17668 12012 17724 12022
rect 17556 12010 17724 12012
rect 17556 11958 17670 12010
rect 17722 11958 17724 12010
rect 17556 11956 17724 11958
rect 17556 11900 17612 11956
rect 17668 11946 17724 11956
rect 17332 11844 17612 11900
rect 18004 11900 18060 13200
rect 21920 12572 22184 12582
rect 21976 12516 22024 12572
rect 22080 12516 22128 12572
rect 21920 12506 22184 12516
rect 18340 12348 18396 12358
rect 18340 12254 18396 12292
rect 21420 12348 21476 12358
rect 21420 12254 21476 12292
rect 22148 12236 22204 12246
rect 19740 12178 19796 12190
rect 18956 12124 19012 12134
rect 18956 12066 19012 12068
rect 18956 12014 18958 12066
rect 19010 12014 19012 12066
rect 19740 12126 19742 12178
rect 19794 12126 19796 12178
rect 23156 12236 23212 13200
rect 28308 12684 28364 13200
rect 28308 12628 28812 12684
rect 28308 12460 28364 12628
rect 28308 12394 28364 12404
rect 23380 12236 23436 12246
rect 23156 12234 23436 12236
rect 23156 12182 23382 12234
rect 23434 12182 23436 12234
rect 23156 12180 23436 12182
rect 18956 12002 19012 12014
rect 19404 12010 19460 12022
rect 17052 11676 17108 11686
rect 15988 11510 15990 11562
rect 16042 11510 16044 11562
rect 15988 11498 16044 11510
rect 16492 11564 16548 11574
rect 16492 11470 16548 11508
rect 17052 11562 17108 11620
rect 17052 11510 17054 11562
rect 17106 11510 17108 11562
rect 17052 11498 17108 11510
rect 17332 11676 17388 11844
rect 18004 11834 18060 11844
rect 19404 11958 19406 12010
rect 19458 11958 19460 12010
rect 17644 11788 17908 11798
rect 17700 11732 17748 11788
rect 17804 11732 17852 11788
rect 17644 11722 17908 11732
rect 16884 11450 16940 11462
rect 16268 11394 16324 11406
rect 16268 11342 16270 11394
rect 16322 11342 16324 11394
rect 14756 10502 14758 10554
rect 14810 10502 14812 10554
rect 14756 10490 14812 10502
rect 14868 10892 14924 10902
rect 16268 10892 16324 11342
rect 16884 11398 16886 11450
rect 16938 11398 16940 11450
rect 16436 11228 16492 11238
rect 16436 11134 16492 11172
rect 13692 10276 14028 10332
rect 14532 10332 14588 10342
rect 12852 9940 13020 9996
rect 13524 9996 13580 10006
rect 12180 9884 12236 9894
rect 11452 9774 11454 9826
rect 11506 9774 11508 9826
rect 11452 9772 11508 9774
rect 11732 9823 11788 9835
rect 11452 9716 11620 9772
rect 11172 9706 11284 9716
rect 10836 9492 10948 9548
rect 10500 9036 10556 9048
rect 10500 8988 10502 9036
rect 10554 8988 10556 9036
rect 10724 9000 10836 9056
rect 10500 8922 10556 8932
rect 10668 8818 10724 8830
rect 10668 8766 10670 8818
rect 10722 8766 10724 8818
rect 10668 8764 10724 8766
rect 10612 8708 10724 8764
rect 9044 8264 9100 8372
rect 10276 8372 10444 8428
rect 10500 8652 10556 8662
rect 9044 8212 9046 8264
rect 9098 8212 9100 8264
rect 9044 8200 9100 8212
rect 9212 8314 9268 8326
rect 9212 8262 9214 8314
rect 9266 8262 9268 8314
rect 9996 8316 10052 8354
rect 10276 8316 10332 8372
rect 9100 8092 9156 8102
rect 8932 8090 9156 8092
rect 8932 8038 9102 8090
rect 9154 8038 9156 8090
rect 8932 8036 9156 8038
rect 9100 8026 9156 8036
rect 8820 7914 8876 7924
rect 9212 7980 9268 8262
rect 9212 7914 9268 7924
rect 9436 8258 9492 8270
rect 9436 8206 9438 8258
rect 9490 8206 9492 8258
rect 9436 7756 9492 8206
rect 9772 8258 9828 8270
rect 9772 8206 9774 8258
rect 9826 8206 9828 8258
rect 9996 8250 10052 8260
rect 10220 8260 10332 8316
rect 10220 8258 10276 8260
rect 9772 8204 9828 8206
rect 10220 8206 10222 8258
rect 10274 8206 10276 8258
rect 10220 8194 10276 8206
rect 10388 8258 10444 8270
rect 10388 8206 10390 8258
rect 10442 8206 10444 8258
rect 9772 8138 9828 8148
rect 10052 8136 10108 8148
rect 9044 7700 9492 7756
rect 9940 8092 9996 8102
rect 9044 7642 9100 7700
rect 9044 7590 9046 7642
rect 9098 7590 9100 7642
rect 9044 7578 9100 7590
rect 9436 7532 9492 7542
rect 9436 7438 9492 7476
rect 9940 7430 9996 8036
rect 10052 8084 10054 8136
rect 10106 8084 10108 8136
rect 10052 7644 10108 8084
rect 10388 7868 10444 8206
rect 10388 7802 10444 7812
rect 10500 8204 10556 8596
rect 10052 7578 10108 7588
rect 10332 7644 10388 7654
rect 10500 7644 10556 8148
rect 10612 8316 10668 8708
rect 10780 8652 10836 9000
rect 10724 8596 10836 8652
rect 10892 8818 10948 9492
rect 11172 9100 11228 9706
rect 11564 9212 11620 9716
rect 11172 9042 11228 9044
rect 11172 8990 11174 9042
rect 11226 8990 11228 9042
rect 11172 8968 11228 8990
rect 11284 9148 11340 9160
rect 11284 9096 11286 9148
rect 11338 9096 11340 9148
rect 11284 8988 11340 9096
rect 11564 9080 11620 9156
rect 11732 9771 11734 9823
rect 11786 9771 11788 9823
rect 12180 9792 12182 9828
rect 12234 9792 12236 9828
rect 12180 9780 12236 9792
rect 11284 8922 11340 8932
rect 11732 8988 11788 9771
rect 12516 9772 12572 9782
rect 12516 9658 12572 9716
rect 12516 9606 12518 9658
rect 12570 9606 12572 9658
rect 11956 9324 12012 9334
rect 11956 9160 12012 9268
rect 12236 9324 12292 9334
rect 12236 9212 12292 9268
rect 11956 9108 11958 9160
rect 12010 9108 12012 9160
rect 11956 9096 12012 9108
rect 12180 9210 12292 9212
rect 12180 9158 12238 9210
rect 12290 9158 12292 9210
rect 12180 9146 12292 9158
rect 11732 8922 11788 8932
rect 12012 8988 12124 8998
rect 12012 8986 12068 8988
rect 12012 8934 12014 8986
rect 12066 8934 12068 8986
rect 12012 8932 12068 8934
rect 12012 8922 12124 8932
rect 10892 8766 10894 8818
rect 10946 8766 10948 8818
rect 10892 8652 10948 8766
rect 12180 8764 12236 9146
rect 10724 8438 10780 8596
rect 10892 8586 10948 8596
rect 12068 8708 12236 8764
rect 12404 8876 12460 8886
rect 12516 8876 12572 9606
rect 12684 9660 12740 9670
rect 12684 9100 12740 9604
rect 12852 9436 12908 9940
rect 13524 9902 13580 9940
rect 12684 9006 12740 9044
rect 12796 9380 12908 9436
rect 12964 9828 13300 9884
rect 12796 9056 12852 9380
rect 12964 9222 13020 9828
rect 13244 9826 13300 9828
rect 13244 9774 13246 9826
rect 13298 9774 13300 9826
rect 13692 9882 13748 10276
rect 14532 10076 14588 10276
rect 14868 10332 14924 10836
rect 16212 10836 16324 10892
rect 14980 10780 15036 10790
rect 14980 10610 15036 10724
rect 14980 10558 14982 10610
rect 15034 10558 15036 10610
rect 14980 10546 15036 10558
rect 16100 10610 16156 10622
rect 16100 10558 16102 10610
rect 16154 10558 16156 10610
rect 15764 10444 15820 10454
rect 16100 10444 16156 10558
rect 15764 10442 16156 10444
rect 15764 10390 15766 10442
rect 15818 10390 16156 10442
rect 15764 10388 16156 10390
rect 15764 10378 15820 10388
rect 14868 10266 14924 10276
rect 15484 10332 15540 10342
rect 14532 10024 14534 10076
rect 14586 10024 14588 10076
rect 14532 10012 14588 10024
rect 13692 9830 13694 9882
rect 13746 9830 13748 9882
rect 13692 9818 13748 9830
rect 14308 9996 14364 10006
rect 14308 9838 14364 9940
rect 14308 9786 14310 9838
rect 14362 9786 14364 9838
rect 14308 9774 14364 9786
rect 14532 9884 14588 9894
rect 13244 9762 13300 9774
rect 13132 9660 13188 9670
rect 13132 9566 13188 9604
rect 13916 9658 13972 9670
rect 13916 9606 13918 9658
rect 13970 9606 13972 9658
rect 12908 9212 13020 9222
rect 12964 9156 13020 9212
rect 13132 9436 13188 9446
rect 13132 9210 13188 9380
rect 13368 9436 13632 9446
rect 13424 9380 13472 9436
rect 13528 9380 13576 9436
rect 13368 9370 13632 9380
rect 13916 9324 13972 9606
rect 13916 9258 13972 9268
rect 14308 9660 14364 9670
rect 13132 9158 13134 9210
rect 13186 9158 13188 9210
rect 12908 9118 12964 9156
rect 13132 9146 13188 9158
rect 12796 9000 13020 9056
rect 14308 9054 14364 9604
rect 12516 8820 12684 8876
rect 11340 8540 11396 8550
rect 10724 8426 10836 8438
rect 10724 8374 10782 8426
rect 10834 8374 10836 8426
rect 10724 8372 10836 8374
rect 10780 8362 10836 8372
rect 10612 7980 10668 8260
rect 10612 7914 10668 7924
rect 10948 8316 11004 8326
rect 11340 8314 11396 8484
rect 12068 8540 12124 8708
rect 12068 8474 12124 8484
rect 12236 8540 12292 8550
rect 11732 8316 11788 8326
rect 10948 7868 11004 8260
rect 11116 8258 11172 8270
rect 11116 8206 11118 8258
rect 11170 8206 11172 8258
rect 11340 8262 11342 8314
rect 11394 8262 11396 8314
rect 11340 8250 11396 8262
rect 11620 8314 11788 8316
rect 11620 8262 11734 8314
rect 11786 8262 11788 8314
rect 11620 8260 11788 8262
rect 11116 7980 11172 8206
rect 11340 7980 11396 7990
rect 11116 7924 11228 7980
rect 10948 7812 11116 7868
rect 10332 7642 10556 7644
rect 10332 7590 10334 7642
rect 10386 7590 10556 7642
rect 10332 7588 10556 7590
rect 10948 7644 11004 7654
rect 10332 7578 10388 7588
rect 10948 7486 11004 7588
rect 10388 7474 10444 7486
rect 8260 7366 8262 7418
rect 8314 7366 8316 7418
rect 8260 7354 8316 7366
rect 8596 7420 8652 7430
rect 8596 7320 8598 7364
rect 8650 7320 8652 7364
rect 9660 7420 9716 7430
rect 9940 7418 10052 7430
rect 9940 7366 9998 7418
rect 10050 7366 10052 7418
rect 9940 7364 10052 7366
rect 9660 7326 9716 7364
rect 9996 7354 10052 7364
rect 10388 7422 10390 7474
rect 10442 7422 10444 7474
rect 10948 7434 10950 7486
rect 11002 7434 11004 7486
rect 10948 7422 11004 7434
rect 10388 7420 10444 7422
rect 10388 7354 10444 7364
rect 8596 7196 8652 7320
rect 10612 7308 10668 7318
rect 10500 7306 10668 7308
rect 10500 7254 10614 7306
rect 10666 7254 10668 7306
rect 10500 7252 10668 7254
rect 8316 7140 8652 7196
rect 9940 7196 9996 7206
rect 8316 6634 8372 7140
rect 9092 7084 9356 7094
rect 9148 7028 9196 7084
rect 9252 7028 9300 7084
rect 9092 7018 9356 7028
rect 9716 6748 9772 6758
rect 8316 6582 8318 6634
rect 8370 6582 8372 6634
rect 8316 6570 8372 6582
rect 8484 6678 8540 6690
rect 8484 6626 8486 6678
rect 8538 6626 8540 6678
rect 9044 6678 9100 6690
rect 8148 5908 8316 5964
rect 7252 4788 7532 4844
rect 7588 5460 7756 5516
rect 7252 4396 7308 4788
rect 7588 4732 7644 5460
rect 8148 5404 8204 5908
rect 8260 5906 8316 5908
rect 8260 5854 8262 5906
rect 8314 5854 8316 5906
rect 8260 5842 8316 5854
rect 7868 5348 8204 5404
rect 7868 5346 7924 5348
rect 7700 5292 7756 5302
rect 7868 5294 7870 5346
rect 7922 5294 7924 5346
rect 7868 5282 7924 5294
rect 8148 5292 8204 5348
rect 8316 5292 8372 5302
rect 8148 5236 8260 5292
rect 7700 5122 7756 5236
rect 7700 5070 7702 5122
rect 7754 5070 7756 5122
rect 7700 5058 7756 5070
rect 8092 5122 8148 5134
rect 8092 5070 8094 5122
rect 8146 5070 8148 5122
rect 7812 4956 7868 4966
rect 7812 4862 7868 4900
rect 7588 4676 7868 4732
rect 7364 4508 7420 4546
rect 7588 4508 7644 4518
rect 7364 4442 7420 4452
rect 7476 4452 7588 4508
rect 7308 4340 7364 4350
rect 7476 4340 7532 4452
rect 7588 4442 7644 4452
rect 7812 4340 7868 4676
rect 8092 4620 8148 5070
rect 8204 5068 8260 5236
rect 8316 5234 8372 5236
rect 8316 5182 8318 5234
rect 8370 5182 8372 5234
rect 8316 5170 8372 5182
rect 8484 5068 8540 6626
rect 8596 6636 8652 6646
rect 8596 5912 8652 6580
rect 9044 6626 9046 6678
rect 9098 6626 9100 6678
rect 9044 6076 9100 6626
rect 8596 5860 8598 5912
rect 8650 5860 8652 5912
rect 8708 6013 8764 6025
rect 8708 5964 8710 6013
rect 8762 5964 8764 6013
rect 9044 6010 9100 6020
rect 9716 6412 9772 6692
rect 8708 5898 8764 5908
rect 8596 5848 8652 5860
rect 9156 5852 9268 5862
rect 9212 5850 9268 5852
rect 9212 5798 9214 5850
rect 9266 5798 9268 5850
rect 9212 5796 9268 5798
rect 9156 5786 9268 5796
rect 9380 5850 9436 5862
rect 9380 5798 9382 5850
rect 9434 5798 9436 5850
rect 8764 5740 8820 5750
rect 9380 5740 9436 5798
rect 8764 5646 8820 5684
rect 8988 5682 9044 5694
rect 8988 5630 8990 5682
rect 9042 5630 9044 5682
rect 9380 5674 9436 5684
rect 9548 5738 9604 5750
rect 9548 5686 9550 5738
rect 9602 5686 9604 5738
rect 8988 5628 9044 5630
rect 8932 5572 9044 5628
rect 8932 5404 8988 5572
rect 9092 5516 9356 5526
rect 9148 5460 9196 5516
rect 9252 5460 9300 5516
rect 9092 5450 9356 5460
rect 8932 5348 9044 5404
rect 8652 5180 8708 5190
rect 8652 5086 8708 5124
rect 8876 5122 8932 5134
rect 8204 5012 8428 5068
rect 8372 4956 8428 5012
rect 8484 5002 8540 5012
rect 8764 5066 8820 5078
rect 8764 5014 8766 5066
rect 8818 5014 8820 5066
rect 8764 4956 8820 5014
rect 8036 4564 8148 4620
rect 8260 4732 8316 4742
rect 8036 4508 8092 4564
rect 8036 4442 8092 4452
rect 8260 4508 8316 4676
rect 8260 4442 8316 4452
rect 7252 4338 7364 4340
rect 7252 4286 7310 4338
rect 7362 4286 7364 4338
rect 7252 4274 7364 4286
rect 7420 4284 7532 4340
rect 7588 4284 7868 4340
rect 8260 4332 8316 4344
rect 7924 4284 8036 4294
rect 7252 4264 7308 4274
rect 7420 4172 7476 4284
rect 7588 4182 7644 4284
rect 7980 4282 8036 4284
rect 7980 4230 7982 4282
rect 8034 4230 8036 4282
rect 7980 4228 8036 4230
rect 7924 4218 8036 4228
rect 8260 4280 8262 4332
rect 8314 4280 8316 4332
rect 6412 4062 6414 4114
rect 6466 4062 6468 4114
rect 6412 3734 6468 4062
rect 6860 4060 7084 4116
rect 7364 4116 7476 4172
rect 7532 4170 7644 4182
rect 7532 4118 7534 4170
rect 7586 4118 7644 4170
rect 7532 4116 7644 4118
rect 7868 4116 7924 4126
rect 6412 3722 6524 3734
rect 6412 3670 6470 3722
rect 6522 3670 6524 3722
rect 6412 3668 6524 3670
rect 6468 3658 6524 3668
rect 6860 3500 6916 4060
rect 7364 3948 7420 4116
rect 7532 4106 7588 4116
rect 7700 4114 7924 4116
rect 7700 4062 7870 4114
rect 7922 4062 7924 4114
rect 7700 4060 7924 4062
rect 7588 3948 7644 3958
rect 7364 3892 7532 3948
rect 7252 3778 7308 3790
rect 7252 3726 7254 3778
rect 7306 3726 7308 3778
rect 5852 3442 5908 3454
rect 5852 3390 5854 3442
rect 5906 3390 5908 3442
rect 6860 3406 6916 3444
rect 7028 3542 7084 3554
rect 7028 3490 7030 3542
rect 7082 3490 7084 3542
rect 5852 3388 5908 3390
rect 5852 3322 5908 3332
rect 6076 3330 6132 3342
rect 6076 3278 6078 3330
rect 6130 3278 6132 3330
rect 6076 3164 6132 3278
rect 7028 3164 7084 3490
rect 6076 3108 6412 3164
rect 5684 2996 6132 3052
rect 6076 2938 6132 2996
rect 6076 2886 6078 2938
rect 6130 2886 6132 2938
rect 6076 2874 6132 2886
rect 6244 2876 6300 2888
rect 6244 2828 6246 2876
rect 6298 2828 6300 2876
rect 6244 2762 6300 2772
rect 6356 2772 6412 3108
rect 7028 3098 7084 3108
rect 7084 2940 7140 2950
rect 7084 2846 7140 2884
rect 6468 2772 6524 2782
rect 6356 2770 6524 2772
rect 5852 2716 5908 2726
rect 6356 2718 6470 2770
rect 6522 2718 6524 2770
rect 6356 2716 6524 2718
rect 5852 2622 5908 2660
rect 6468 2650 6524 2660
rect 6692 2716 6748 2726
rect 5460 2090 5516 2100
rect 6244 1986 6300 1998
rect 3892 1866 3948 1876
rect 4732 1932 4844 1942
rect 4788 1876 4844 1932
rect 5180 1932 5236 1942
rect 4732 1838 4788 1876
rect 4564 1820 4620 1830
rect 4564 1726 4620 1764
rect 5180 1708 5236 1876
rect 5180 1642 5236 1652
rect 5348 1930 5460 1942
rect 5348 1878 5406 1930
rect 5458 1878 5460 1930
rect 5348 1866 5460 1878
rect 5628 1930 5684 1942
rect 5628 1878 5630 1930
rect 5682 1878 5684 1930
rect 4816 1596 5080 1606
rect 4872 1540 4920 1596
rect 4976 1540 5024 1596
rect 4816 1530 5080 1540
rect 5348 1484 5404 1866
rect 5628 1708 5684 1878
rect 6244 1934 6246 1986
rect 6298 1934 6300 1986
rect 6244 1820 6300 1934
rect 6692 1930 6748 2660
rect 7252 2268 7308 3726
rect 7364 3542 7420 3554
rect 7364 3490 7366 3542
rect 7418 3490 7420 3542
rect 7364 3276 7420 3490
rect 7364 3210 7420 3220
rect 7476 3164 7532 3892
rect 7588 3566 7644 3892
rect 7588 3514 7590 3566
rect 7642 3514 7644 3566
rect 7588 3502 7644 3514
rect 7700 3387 7756 4060
rect 7868 4050 7924 4060
rect 8092 4114 8148 4126
rect 8092 4062 8094 4114
rect 8146 4062 8148 4114
rect 8092 3948 8148 4062
rect 7476 2940 7532 3108
rect 7476 2874 7532 2884
rect 7588 3331 7756 3387
rect 7812 3892 8148 3948
rect 7420 2772 7476 2782
rect 7420 2770 7532 2772
rect 7420 2718 7422 2770
rect 7474 2718 7532 2770
rect 7420 2706 7532 2718
rect 7476 2380 7532 2706
rect 7588 2604 7644 3331
rect 7588 2538 7644 2548
rect 7700 3164 7756 3174
rect 7476 2324 7588 2380
rect 7252 2212 7476 2268
rect 7420 2210 7476 2212
rect 6916 2179 6972 2194
rect 6916 2156 6918 2179
rect 6970 2156 6972 2179
rect 7420 2158 7422 2210
rect 7474 2158 7476 2210
rect 7420 2146 7476 2158
rect 7532 2154 7588 2324
rect 7700 2268 7756 3108
rect 7812 2940 7868 3892
rect 8260 3836 8316 4280
rect 8092 3780 8316 3836
rect 8092 3722 8148 3780
rect 8092 3670 8094 3722
rect 8146 3670 8148 3722
rect 8092 3658 8148 3670
rect 8204 3612 8260 3622
rect 8204 3610 8316 3612
rect 7980 3554 8036 3566
rect 7980 3502 7982 3554
rect 8034 3502 8036 3554
rect 8204 3558 8206 3610
rect 8258 3558 8316 3610
rect 8204 3546 8316 3558
rect 7980 3500 8036 3502
rect 7980 3434 8036 3444
rect 8260 3387 8316 3546
rect 8372 3560 8428 4900
rect 8708 4900 8820 4956
rect 8876 5070 8878 5122
rect 8930 5070 8932 5122
rect 8876 4956 8932 5070
rect 8988 5068 9044 5348
rect 9548 5292 9604 5686
rect 9716 5404 9772 6356
rect 9940 5918 9996 7140
rect 10500 5918 10556 7252
rect 10612 7242 10668 7252
rect 11060 7308 11116 7812
rect 11172 7532 11228 7924
rect 11340 7642 11396 7924
rect 11620 7980 11676 8260
rect 11732 8250 11788 8260
rect 11900 8316 11956 8326
rect 11900 8222 11956 8260
rect 12236 8258 12292 8484
rect 12404 8428 12460 8820
rect 12628 8428 12684 8820
rect 12404 8372 12572 8428
rect 12404 8336 12460 8372
rect 12404 8284 12406 8336
rect 12458 8284 12460 8336
rect 12404 8272 12460 8284
rect 12236 8206 12238 8258
rect 12290 8206 12292 8258
rect 12236 8204 12292 8206
rect 12236 8138 12292 8148
rect 12404 8204 12460 8214
rect 12404 8110 12460 8148
rect 11788 8092 11844 8102
rect 11620 7914 11676 7924
rect 11732 8090 11844 8092
rect 11732 8038 11790 8090
rect 11842 8038 11844 8090
rect 11732 8026 11844 8038
rect 11732 7868 11788 8026
rect 12068 7980 12124 7990
rect 11732 7802 11788 7812
rect 11956 7868 12012 7878
rect 11340 7590 11342 7642
rect 11394 7590 11396 7642
rect 11340 7578 11396 7590
rect 11452 7644 11508 7654
rect 11844 7644 11900 7654
rect 11956 7644 12012 7812
rect 11452 7642 12012 7644
rect 11452 7590 11454 7642
rect 11506 7590 11846 7642
rect 11898 7590 12012 7642
rect 11452 7588 12012 7590
rect 11452 7488 11508 7588
rect 11844 7578 11900 7588
rect 11228 7476 11508 7488
rect 11172 7432 11508 7476
rect 11172 7400 11228 7432
rect 11060 7242 11116 7252
rect 12068 7196 12124 7924
rect 12516 7868 12572 8372
rect 12628 8362 12684 8372
rect 12516 7802 12572 7812
rect 12964 8326 13020 9000
rect 13748 9030 13804 9042
rect 13748 8978 13750 9030
rect 13802 8978 13804 9030
rect 13524 8874 13580 8886
rect 13524 8822 13526 8874
rect 13578 8822 13580 8874
rect 12964 8314 13076 8326
rect 12964 8262 13022 8314
rect 13074 8262 13076 8314
rect 12964 8250 13076 8262
rect 13188 8316 13244 8326
rect 12628 7532 12684 7542
rect 12292 7530 12796 7532
rect 12292 7478 12630 7530
rect 12682 7478 12796 7530
rect 12292 7476 12796 7478
rect 12292 7430 12348 7476
rect 12628 7466 12684 7476
rect 12236 7418 12348 7430
rect 12236 7366 12238 7418
rect 12290 7366 12348 7418
rect 12236 7364 12348 7366
rect 12236 7354 12292 7364
rect 12068 7140 12292 7196
rect 12236 6858 12292 7140
rect 12236 6806 12238 6858
rect 12290 6806 12292 6858
rect 12236 6794 12292 6806
rect 11396 6748 11452 6758
rect 11396 6654 11452 6692
rect 12572 6636 12628 6646
rect 12572 6542 12628 6580
rect 9940 5866 9942 5918
rect 9994 5866 9996 5918
rect 9940 5854 9996 5866
rect 10444 5906 10556 5918
rect 10444 5854 10446 5906
rect 10498 5854 10556 5906
rect 10444 5840 10556 5854
rect 12068 6522 12124 6534
rect 12068 6470 12070 6522
rect 12122 6470 12124 6522
rect 11676 5628 11732 5638
rect 9380 5236 9604 5292
rect 9660 5348 9772 5404
rect 10108 5516 10164 5526
rect 9268 5180 9324 5190
rect 9268 5086 9324 5124
rect 8988 5012 9212 5068
rect 8876 4900 8988 4956
rect 8708 4844 8764 4900
rect 8708 4778 8764 4788
rect 8596 4732 8652 4742
rect 8596 4338 8652 4676
rect 8932 4732 8988 4900
rect 8932 4620 8988 4676
rect 8596 4286 8598 4338
rect 8650 4286 8652 4338
rect 8596 4274 8652 4286
rect 8820 4564 8988 4620
rect 8372 3508 8374 3560
rect 8426 3508 8428 3560
rect 8372 3496 8428 3508
rect 8484 4060 8540 4070
rect 8484 3387 8540 4004
rect 8708 3554 8764 3566
rect 8708 3502 8710 3554
rect 8762 3502 8764 3554
rect 8708 3500 8764 3502
rect 8708 3434 8764 3444
rect 8148 3331 8316 3387
rect 8372 3331 8540 3387
rect 8148 3276 8204 3331
rect 8036 3220 8204 3276
rect 8036 2940 8092 3220
rect 8372 3164 8428 3331
rect 8820 3276 8876 4564
rect 9044 4508 9100 4518
rect 9044 4294 9100 4452
rect 8988 4284 9100 4294
rect 8820 3210 8876 3220
rect 8932 4282 9100 4284
rect 8932 4230 8990 4282
rect 9042 4230 9100 4282
rect 8932 4228 9100 4230
rect 8932 4218 9044 4228
rect 7812 2884 8092 2940
rect 8148 3108 8428 3164
rect 7812 2714 7868 2726
rect 7812 2662 7814 2714
rect 7866 2662 7868 2714
rect 7812 2604 7868 2662
rect 7812 2538 7868 2548
rect 7700 2202 7756 2212
rect 6916 2090 6972 2100
rect 7532 2102 7534 2154
rect 7586 2102 7588 2154
rect 7532 2090 7588 2102
rect 7812 2156 7868 2166
rect 7644 2044 7700 2054
rect 7644 1950 7700 1988
rect 7812 2015 7868 2100
rect 7812 1963 7814 2015
rect 7866 1963 7868 2015
rect 7812 1951 7868 1963
rect 6692 1878 6694 1930
rect 6746 1878 6748 1930
rect 6692 1866 6748 1878
rect 6244 1754 6300 1764
rect 5628 1642 5684 1652
rect 5124 1428 5404 1484
rect 5124 1372 5180 1428
rect 4844 1316 5180 1372
rect 7924 1382 7980 2884
rect 8036 2716 8092 2726
rect 8036 2616 8038 2660
rect 8090 2616 8092 2660
rect 8036 2604 8092 2616
rect 8148 2054 8204 3108
rect 8596 3052 8652 3062
rect 8932 3052 8988 4218
rect 9156 4114 9212 5012
rect 9380 4732 9436 5236
rect 9660 5180 9716 5348
rect 10108 5346 10164 5460
rect 9884 5292 9940 5302
rect 10108 5294 10110 5346
rect 10162 5294 10164 5346
rect 10108 5282 10164 5294
rect 10836 5404 10892 5414
rect 10836 5302 10892 5348
rect 10836 5290 10948 5302
rect 10836 5238 10894 5290
rect 10946 5238 10948 5290
rect 10836 5236 10948 5238
rect 9884 5198 9940 5236
rect 10892 5226 10948 5236
rect 9548 5124 9716 5180
rect 9996 5180 10052 5190
rect 10388 5180 10444 5190
rect 9548 5066 9604 5124
rect 9996 5086 10052 5124
rect 10276 5116 10332 5128
rect 9548 5014 9550 5066
rect 9602 5014 9604 5066
rect 9548 5002 9604 5014
rect 10164 5068 10220 5078
rect 10276 5068 10278 5116
rect 10220 5064 10278 5068
rect 10330 5064 10332 5116
rect 10220 5012 10332 5064
rect 11060 5178 11116 5190
rect 10164 5002 10220 5012
rect 10388 4956 10444 5124
rect 10276 4900 10444 4956
rect 10500 5122 10556 5134
rect 10500 5070 10502 5122
rect 10554 5070 10556 5122
rect 10052 4844 10108 4854
rect 9380 4666 9436 4676
rect 9940 4732 9996 4742
rect 9940 4456 9996 4676
rect 9492 4396 9548 4406
rect 9940 4404 9942 4456
rect 9994 4404 9996 4456
rect 9940 4340 9996 4404
rect 9268 4326 9324 4338
rect 9268 4284 9270 4326
rect 9322 4284 9324 4326
rect 9492 4298 9494 4340
rect 9546 4298 9548 4340
rect 9492 4286 9548 4298
rect 9268 4218 9324 4228
rect 9828 4284 9996 4340
rect 10052 4396 10108 4788
rect 10276 4518 10332 4900
rect 10220 4506 10332 4518
rect 10220 4454 10222 4506
rect 10274 4454 10332 4506
rect 10220 4452 10332 4454
rect 10388 4732 10444 4742
rect 10220 4442 10276 4452
rect 10052 4330 10108 4340
rect 9156 4062 9158 4114
rect 9210 4062 9212 4114
rect 9156 4050 9212 4062
rect 9092 3948 9356 3958
rect 9148 3892 9196 3948
rect 9252 3892 9300 3948
rect 9092 3882 9356 3892
rect 9828 3948 9884 4284
rect 9996 4172 10052 4182
rect 9940 4170 10052 4172
rect 9940 4118 9998 4170
rect 10050 4118 10052 4170
rect 9940 4106 10052 4118
rect 9940 4060 9996 4106
rect 9940 3994 9996 4004
rect 9828 3882 9884 3892
rect 9548 3836 9604 3846
rect 10388 3836 10444 4676
rect 10500 4620 10556 5070
rect 11060 5126 11062 5178
rect 11114 5126 11116 5178
rect 11060 5068 11116 5126
rect 11060 5002 11116 5012
rect 11228 5122 11284 5134
rect 11228 5070 11230 5122
rect 11282 5070 11284 5122
rect 11228 4732 11284 5070
rect 11676 5010 11732 5572
rect 11676 4958 11678 5010
rect 11730 4958 11732 5010
rect 12068 5078 12124 6470
rect 12740 6300 12796 7476
rect 12852 7474 12908 7486
rect 12852 7422 12854 7474
rect 12906 7422 12908 7474
rect 12852 7420 12908 7422
rect 12852 7354 12908 7364
rect 12740 6234 12796 6244
rect 12852 6412 12908 6422
rect 12516 5964 12572 5974
rect 12180 5292 12236 5302
rect 12180 5198 12236 5236
rect 12292 5180 12348 5190
rect 12292 5099 12294 5124
rect 12346 5099 12348 5124
rect 12292 5086 12348 5099
rect 12068 5066 12180 5078
rect 12068 5014 12126 5066
rect 12178 5014 12180 5066
rect 12068 5002 12180 5014
rect 12404 5068 12460 5078
rect 11676 4946 11732 4958
rect 11900 4956 11956 4966
rect 11900 4862 11956 4900
rect 11228 4666 11284 4676
rect 11732 4732 11788 4742
rect 10500 4172 10556 4564
rect 11508 4620 11564 4630
rect 11172 4508 11228 4518
rect 11172 4414 11228 4452
rect 11508 4282 11564 4564
rect 11508 4230 11510 4282
rect 11562 4230 11564 4282
rect 11508 4218 11564 4230
rect 10500 4078 10556 4116
rect 10892 4172 10948 4182
rect 10892 4170 11004 4172
rect 10892 4118 10894 4170
rect 10946 4118 11004 4170
rect 10892 4106 11004 4118
rect 10948 3948 11004 4106
rect 11732 3948 11788 4676
rect 12068 4620 12124 5002
rect 12404 4732 12460 5012
rect 12068 4554 12124 4564
rect 12180 4676 12460 4732
rect 12180 4450 12236 4676
rect 12180 4398 12182 4450
rect 12234 4398 12236 4450
rect 12180 4386 12236 4398
rect 12516 4350 12572 5908
rect 12740 5852 12796 5862
rect 12852 5852 12908 6356
rect 12740 5850 12908 5852
rect 12740 5798 12742 5850
rect 12794 5798 12908 5850
rect 12740 5796 12908 5798
rect 12964 5852 13020 8250
rect 13188 6870 13244 8260
rect 13356 8316 13412 8326
rect 13356 8222 13412 8260
rect 13524 8092 13580 8822
rect 13748 8540 13804 8978
rect 14084 9030 14140 9042
rect 14084 8978 14086 9030
rect 14138 8978 14140 9030
rect 14084 8876 14140 8978
rect 14308 9002 14310 9054
rect 14362 9002 14364 9054
rect 14308 8988 14364 9002
rect 14308 8922 14364 8932
rect 14084 8810 14140 8820
rect 13972 8792 14028 8804
rect 13972 8740 13974 8792
rect 14026 8740 14028 8792
rect 13972 8540 14028 8740
rect 13972 8484 14084 8540
rect 13748 8474 13804 8484
rect 14028 8482 14084 8484
rect 14028 8430 14030 8482
rect 14082 8430 14084 8482
rect 14028 8418 14084 8430
rect 14532 8326 14588 9828
rect 14868 9884 14924 9894
rect 14644 9814 14700 9826
rect 14644 9772 14646 9814
rect 14698 9772 14700 9814
rect 14868 9786 14870 9828
rect 14922 9786 14924 9828
rect 15484 9882 15540 10276
rect 15484 9830 15486 9882
rect 15538 9830 15540 9882
rect 15484 9818 15540 9830
rect 15876 10220 15932 10230
rect 16212 10220 16268 10836
rect 16324 10720 16380 10732
rect 16324 10668 16326 10720
rect 16378 10668 16380 10720
rect 16324 10602 16380 10612
rect 16772 10598 16828 10610
rect 16772 10546 16774 10598
rect 16826 10546 16828 10598
rect 16380 10386 16436 10398
rect 16604 10388 16660 10398
rect 16380 10334 16382 10386
rect 16434 10334 16436 10386
rect 16380 10332 16436 10334
rect 16380 10266 16436 10276
rect 16548 10386 16660 10388
rect 16548 10334 16606 10386
rect 16658 10334 16660 10386
rect 16548 10322 16660 10334
rect 14868 9774 14924 9786
rect 14644 9706 14700 9716
rect 15092 9660 15148 9670
rect 15092 9210 15148 9604
rect 15260 9658 15316 9670
rect 15708 9660 15764 9670
rect 15260 9606 15262 9658
rect 15314 9606 15316 9658
rect 15260 9436 15316 9606
rect 15260 9370 15316 9380
rect 15652 9658 15764 9660
rect 15652 9606 15710 9658
rect 15762 9606 15764 9658
rect 15652 9594 15764 9606
rect 15092 9158 15094 9210
rect 15146 9158 15148 9210
rect 15092 9146 15148 9158
rect 15428 9212 15484 9222
rect 15428 9054 15484 9156
rect 15428 9002 15430 9054
rect 15482 9002 15484 9054
rect 15428 8990 15484 9002
rect 14700 8876 14756 8886
rect 13804 8316 13860 8326
rect 13636 8238 13692 8250
rect 13636 8186 13638 8238
rect 13690 8186 13692 8238
rect 13804 8222 13860 8260
rect 14196 8316 14252 8326
rect 13636 8092 13692 8186
rect 13916 8202 13972 8214
rect 13916 8150 13918 8202
rect 13970 8150 13972 8202
rect 13636 8036 13804 8092
rect 13524 8026 13580 8036
rect 13368 7868 13632 7878
rect 13424 7812 13472 7868
rect 13528 7812 13576 7868
rect 13368 7802 13632 7812
rect 13748 7644 13804 8036
rect 13916 7756 13972 8150
rect 13916 7690 13972 7700
rect 14084 8092 14140 8102
rect 13636 7588 13804 7644
rect 14084 7644 14140 8036
rect 14196 7756 14252 8260
rect 14476 8314 14588 8326
rect 14476 8262 14478 8314
rect 14530 8262 14588 8314
rect 14476 8260 14588 8262
rect 14644 8874 14756 8876
rect 14644 8822 14702 8874
rect 14754 8822 14756 8874
rect 14644 8810 14756 8822
rect 14476 8250 14532 8260
rect 14644 8102 14700 8810
rect 15652 8428 15708 9594
rect 15764 8876 15820 8886
rect 15764 8782 15820 8820
rect 15652 8362 15708 8372
rect 15148 8316 15204 8326
rect 15148 8314 15260 8316
rect 14924 8258 14980 8270
rect 14924 8206 14926 8258
rect 14978 8206 14980 8258
rect 15148 8262 15150 8314
rect 15202 8262 15260 8314
rect 15148 8250 15260 8262
rect 14924 8204 14980 8206
rect 14980 8148 15036 8204
rect 14924 8138 15036 8148
rect 14196 7690 14252 7700
rect 14308 8092 14364 8102
rect 13636 7542 13692 7588
rect 14084 7578 14140 7588
rect 14196 7586 14252 7598
rect 13580 7530 13692 7542
rect 13580 7478 13582 7530
rect 13634 7478 13692 7530
rect 13580 7476 13692 7478
rect 13916 7532 13972 7542
rect 13580 7466 13636 7476
rect 13916 7418 13972 7476
rect 14196 7534 14198 7586
rect 14250 7534 14252 7586
rect 14196 7532 14252 7534
rect 14196 7466 14252 7476
rect 14308 7488 14364 8036
rect 14588 8090 14700 8102
rect 14588 8038 14590 8090
rect 14642 8038 14700 8090
rect 14588 8036 14700 8038
rect 14588 7868 14644 8036
rect 14588 7802 14644 7812
rect 14308 7474 14420 7488
rect 14308 7432 14366 7474
rect 13916 7366 13918 7418
rect 13970 7366 13972 7418
rect 14364 7422 14366 7432
rect 14418 7422 14420 7474
rect 14364 7410 14420 7422
rect 14644 7462 14700 7474
rect 14644 7410 14646 7462
rect 14698 7410 14700 7462
rect 13916 7354 13972 7366
rect 14140 7250 14196 7262
rect 14140 7198 14142 7250
rect 14194 7198 14196 7250
rect 14140 6972 14196 7198
rect 14644 7196 14700 7410
rect 14980 7196 15036 8138
rect 15092 8092 15148 8102
rect 15092 7998 15148 8036
rect 15204 7980 15260 8250
rect 15540 8314 15596 8326
rect 15540 8262 15542 8314
rect 15594 8262 15596 8314
rect 15204 7924 15484 7980
rect 15204 7644 15260 7924
rect 15204 7578 15260 7588
rect 15316 7532 15372 7542
rect 15316 7434 15318 7476
rect 15370 7434 15372 7476
rect 15316 7422 15372 7434
rect 14980 7140 15316 7196
rect 14644 7130 14700 7140
rect 14140 6916 14924 6972
rect 13188 6858 13300 6870
rect 13188 6806 13246 6858
rect 13298 6806 13300 6858
rect 13188 6804 13300 6806
rect 13244 6794 13300 6804
rect 13580 6860 13636 6870
rect 13580 6766 13636 6804
rect 14868 6858 14924 6916
rect 14868 6806 14870 6858
rect 14922 6806 14924 6858
rect 14868 6794 14924 6806
rect 13076 6748 13132 6758
rect 13076 6654 13132 6692
rect 13804 6748 13860 6758
rect 14084 6748 14140 6758
rect 13804 6746 13916 6748
rect 13804 6694 13806 6746
rect 13858 6694 13916 6746
rect 13804 6682 13916 6694
rect 13076 6524 13188 6534
rect 13132 6522 13188 6524
rect 13132 6470 13134 6522
rect 13186 6470 13188 6522
rect 13132 6468 13188 6470
rect 13076 6458 13188 6468
rect 13748 6522 13804 6534
rect 13748 6470 13750 6522
rect 13802 6470 13804 6522
rect 13188 6300 13244 6310
rect 12740 5786 12796 5796
rect 12964 5786 13020 5796
rect 13076 6076 13132 6086
rect 13188 6076 13244 6244
rect 13368 6300 13632 6310
rect 13424 6244 13472 6300
rect 13528 6244 13576 6300
rect 13368 6234 13632 6244
rect 13412 6076 13468 6086
rect 13188 6074 13468 6076
rect 13188 6022 13414 6074
rect 13466 6022 13468 6074
rect 13188 6020 13468 6022
rect 13076 5140 13132 6020
rect 13412 6010 13468 6020
rect 13748 5964 13804 6470
rect 13748 5898 13804 5908
rect 13860 5896 13916 6682
rect 14084 6654 14140 6692
rect 14364 6636 14420 6646
rect 14588 6636 14644 6646
rect 14364 6634 14644 6636
rect 14364 6582 14366 6634
rect 14418 6582 14590 6634
rect 14642 6582 14644 6634
rect 14364 6580 14644 6582
rect 14364 6570 14420 6580
rect 14084 6524 14140 6534
rect 13972 6076 14028 6086
rect 13972 5982 14028 6020
rect 14084 5918 14140 6468
rect 14588 6412 14644 6580
rect 15260 6634 15316 7140
rect 15428 6758 15484 7924
rect 15540 7644 15596 8262
rect 15876 8214 15932 10164
rect 15988 10164 16268 10220
rect 15988 9660 16044 10164
rect 16548 10108 16604 10322
rect 16772 10108 16828 10546
rect 16100 10052 16604 10108
rect 16660 10052 16828 10108
rect 16884 10108 16940 11398
rect 16100 9994 16156 10052
rect 16100 9942 16102 9994
rect 16154 9942 16156 9994
rect 16100 9930 16156 9942
rect 16380 9884 16436 9894
rect 16660 9884 16716 10052
rect 16884 10042 16940 10052
rect 17052 10892 17108 10902
rect 17052 10666 17108 10836
rect 17052 10614 17054 10666
rect 17106 10614 17108 10666
rect 16436 9828 16716 9884
rect 17052 9884 17108 10614
rect 17332 10444 17388 11620
rect 17444 11562 17500 11574
rect 17444 11510 17446 11562
rect 17498 11510 17500 11562
rect 17444 11452 17500 11510
rect 17444 10892 17500 11396
rect 17892 11564 17948 11574
rect 17892 11450 17948 11508
rect 19404 11564 19460 11958
rect 19740 11788 19796 12126
rect 19740 11722 19796 11732
rect 20132 12122 20188 12134
rect 21084 12124 21140 12134
rect 20132 12070 20134 12122
rect 20186 12070 20188 12122
rect 19404 11498 19460 11508
rect 17892 11398 17894 11450
rect 17946 11398 17948 11450
rect 17892 11386 17948 11398
rect 18788 11452 18844 11462
rect 18788 11358 18844 11396
rect 19292 11452 19348 11462
rect 19292 11358 19348 11396
rect 20020 11452 20076 11462
rect 20020 11358 20076 11396
rect 20132 11452 20188 12070
rect 20468 12122 21140 12124
rect 20468 12070 21086 12122
rect 21138 12070 21140 12122
rect 20468 12068 21140 12070
rect 20468 12066 20580 12068
rect 20468 12014 20526 12066
rect 20578 12014 20580 12066
rect 21084 12058 21140 12068
rect 21812 12122 21868 12134
rect 21812 12070 21814 12122
rect 21866 12070 21868 12122
rect 20468 12002 20580 12014
rect 20468 11564 20524 12002
rect 21812 11900 21868 12070
rect 22148 12062 22204 12180
rect 23380 12170 23436 12180
rect 24164 12236 24220 12246
rect 24164 12138 24166 12180
rect 24218 12138 24220 12180
rect 28756 12178 28812 12628
rect 30472 12572 30736 12582
rect 30528 12516 30576 12572
rect 30632 12516 30680 12572
rect 30472 12506 30736 12516
rect 32676 12236 32732 12246
rect 24164 12126 24220 12138
rect 24724 12166 24780 12178
rect 22148 12012 22150 12062
rect 22202 12012 22204 12062
rect 24724 12114 24726 12166
rect 24778 12114 24780 12166
rect 22148 11946 22204 11956
rect 22652 12010 22708 12022
rect 22652 11958 22654 12010
rect 22706 11958 22708 12010
rect 21812 11834 21868 11844
rect 20412 11508 20524 11564
rect 20412 11506 20468 11508
rect 20412 11454 20414 11506
rect 20466 11454 20468 11506
rect 20412 11442 20468 11454
rect 20916 11452 20972 11462
rect 20132 11386 20188 11396
rect 20916 11338 20972 11396
rect 20916 11286 20918 11338
rect 20970 11286 20972 11338
rect 20916 11274 20972 11286
rect 21588 11450 21644 11462
rect 21588 11398 21590 11450
rect 21642 11398 21644 11450
rect 17444 10826 17500 10836
rect 18452 11226 18508 11238
rect 18452 11174 18454 11226
rect 18506 11174 18508 11226
rect 19796 11228 19852 11238
rect 17780 10668 17836 10678
rect 17332 10378 17388 10388
rect 17444 10592 17500 10604
rect 17444 10540 17446 10592
rect 17498 10540 17500 10592
rect 17780 10574 17836 10612
rect 18340 10592 18396 10604
rect 17444 10332 17500 10540
rect 18340 10540 18342 10592
rect 18394 10540 18396 10592
rect 17444 10266 17500 10276
rect 18004 10442 18060 10454
rect 18004 10390 18006 10442
rect 18058 10390 18060 10442
rect 17644 10220 17908 10230
rect 17700 10164 17748 10220
rect 17804 10164 17852 10220
rect 17644 10154 17908 10164
rect 18004 10108 18060 10390
rect 17948 10052 18060 10108
rect 17668 9996 17724 10006
rect 16380 9752 16436 9828
rect 17052 9818 17108 9828
rect 17556 9882 17612 9894
rect 17556 9830 17558 9882
rect 17610 9830 17612 9882
rect 16940 9772 16996 9782
rect 16940 9678 16996 9716
rect 17164 9772 17220 9782
rect 17556 9772 17612 9830
rect 17164 9770 17612 9772
rect 17164 9718 17166 9770
rect 17218 9718 17612 9770
rect 17164 9716 17612 9718
rect 17164 9706 17220 9716
rect 15988 9604 16156 9660
rect 16100 9054 16156 9604
rect 16716 9658 16772 9670
rect 16716 9606 16718 9658
rect 16770 9606 16772 9658
rect 16716 9548 16772 9606
rect 16716 9492 17388 9548
rect 17108 9212 17164 9222
rect 17332 9212 17388 9492
rect 17556 9436 17612 9716
rect 17668 9548 17724 9940
rect 17836 9884 17892 9894
rect 17836 9790 17892 9828
rect 17668 9482 17724 9492
rect 17780 9658 17836 9670
rect 17780 9606 17782 9658
rect 17834 9606 17836 9658
rect 17556 9370 17612 9380
rect 17780 9212 17836 9606
rect 17948 9660 18004 10052
rect 18340 9996 18396 10540
rect 18452 10556 18508 11174
rect 19628 11170 19684 11182
rect 19628 11118 19630 11170
rect 19682 11118 19684 11170
rect 19628 10780 19684 11118
rect 19628 10714 19684 10724
rect 18452 10490 18508 10500
rect 19012 10666 19068 10678
rect 19012 10614 19014 10666
rect 19066 10614 19068 10666
rect 18340 9930 18396 9940
rect 18060 9884 18116 9894
rect 18060 9790 18116 9828
rect 18452 9884 18508 9894
rect 18452 9790 18508 9828
rect 18788 9826 18844 9838
rect 18788 9774 18790 9826
rect 18842 9774 18844 9826
rect 18284 9660 18340 9670
rect 17948 9604 18060 9660
rect 17332 9156 17836 9212
rect 17892 9436 17948 9446
rect 17108 9118 17164 9156
rect 16100 9002 16102 9054
rect 16154 9002 16156 9054
rect 16100 8988 16156 9002
rect 16324 9100 16380 9110
rect 16324 9002 16326 9044
rect 16378 9002 16380 9044
rect 17220 9100 17276 9110
rect 16324 8990 16380 9002
rect 16660 9030 16716 9042
rect 15820 8202 15932 8214
rect 15820 8150 15822 8202
rect 15874 8150 15932 8202
rect 15820 8138 15932 8150
rect 15596 7588 15708 7644
rect 15540 7578 15596 7588
rect 15652 6758 15708 7588
rect 15428 6746 15540 6758
rect 15428 6694 15486 6746
rect 15538 6694 15540 6746
rect 15428 6692 15540 6694
rect 15652 6746 15764 6758
rect 15652 6694 15710 6746
rect 15762 6694 15764 6746
rect 15652 6692 15764 6694
rect 15484 6682 15540 6692
rect 15708 6682 15764 6692
rect 15260 6582 15262 6634
rect 15314 6582 15316 6634
rect 15260 6570 15316 6582
rect 14588 6346 14644 6356
rect 15876 6412 15932 8138
rect 15988 8932 16156 8988
rect 16436 8988 16492 8998
rect 15988 8204 16044 8932
rect 16436 8818 16492 8932
rect 16660 8978 16662 9030
rect 16714 8978 16716 9030
rect 17220 8998 17276 9044
rect 17780 9042 17836 9054
rect 16436 8766 16438 8818
rect 16490 8766 16492 8818
rect 16436 8754 16492 8766
rect 16548 8876 16604 8886
rect 15988 7532 16044 8148
rect 15988 7466 16044 7476
rect 16100 8316 16156 8328
rect 16548 8316 16604 8820
rect 16660 8764 16716 8978
rect 16660 8698 16716 8708
rect 16940 8986 16996 8998
rect 16940 8934 16942 8986
rect 16994 8934 16996 8986
rect 16940 8764 16996 8934
rect 17164 8986 17276 8998
rect 17164 8934 17166 8986
rect 17218 8934 17276 8986
rect 17164 8932 17276 8934
rect 17444 8988 17500 8998
rect 17164 8922 17220 8932
rect 17444 8894 17500 8932
rect 17780 8990 17782 9042
rect 17834 8990 17836 9042
rect 17780 8876 17836 8990
rect 17556 8820 17836 8876
rect 17892 8876 17948 9380
rect 18004 9324 18060 9604
rect 18004 9258 18060 9268
rect 18284 9266 18340 9604
rect 18284 9214 18286 9266
rect 18338 9214 18340 9266
rect 18284 9202 18340 9214
rect 18060 9154 18116 9166
rect 18060 9102 18062 9154
rect 18114 9102 18116 9154
rect 18060 9100 18116 9102
rect 17556 8764 17612 8820
rect 17892 8810 17948 8820
rect 18004 9044 18116 9100
rect 16940 8698 16996 8708
rect 17332 8708 17612 8764
rect 18004 8774 18060 9044
rect 18788 8886 18844 9774
rect 18340 8876 18396 8886
rect 18788 8876 18900 8886
rect 18788 8820 18844 8876
rect 18340 8782 18396 8820
rect 18844 8782 18900 8820
rect 18004 8764 18116 8774
rect 18004 8708 18060 8764
rect 17332 8316 17388 8708
rect 18060 8698 18116 8708
rect 17644 8652 17908 8662
rect 17700 8596 17748 8652
rect 17804 8596 17852 8652
rect 17644 8586 17908 8596
rect 16548 8260 16660 8316
rect 16100 8250 16156 8260
rect 16100 8198 16102 8250
rect 16154 8198 16156 8250
rect 16100 7196 16156 8198
rect 16604 8258 16660 8260
rect 16604 8206 16606 8258
rect 16658 8206 16660 8258
rect 17332 8250 17388 8260
rect 17444 8540 17500 8550
rect 16604 8194 16660 8206
rect 17220 7868 17276 7878
rect 16100 7130 16156 7140
rect 16660 7532 16716 7542
rect 16212 6914 16268 6926
rect 16212 6862 16214 6914
rect 16266 6862 16268 6914
rect 15876 6346 15932 6356
rect 15988 6678 16044 6690
rect 15988 6626 15990 6678
rect 16042 6626 16044 6678
rect 14028 5906 14140 5918
rect 13076 5088 13078 5140
rect 13130 5088 13132 5140
rect 13076 5076 13132 5088
rect 13188 5852 13244 5862
rect 13020 4508 13076 4518
rect 13188 4508 13244 5796
rect 13636 5852 13692 5862
rect 13860 5840 13972 5896
rect 14028 5854 14030 5906
rect 14082 5854 14140 5906
rect 14644 5964 14700 5974
rect 14644 5862 14646 5908
rect 14698 5862 14700 5908
rect 14028 5840 14140 5854
rect 14420 5852 14476 5862
rect 14644 5850 14700 5862
rect 15204 5894 15260 5906
rect 13636 5134 13692 5796
rect 13804 5740 13860 5760
rect 13916 5740 13972 5840
rect 14420 5758 14476 5796
rect 15204 5842 15206 5894
rect 15258 5842 15260 5894
rect 13916 5684 14028 5740
rect 13804 5682 13860 5684
rect 13804 5630 13806 5682
rect 13858 5630 13860 5682
rect 13804 5292 13860 5630
rect 13804 5226 13860 5236
rect 13636 5082 13638 5134
rect 13690 5082 13692 5134
rect 13636 5070 13692 5082
rect 13412 4956 13468 4966
rect 13412 4862 13468 4900
rect 13368 4732 13632 4742
rect 13424 4676 13472 4732
rect 13528 4676 13576 4732
rect 13368 4666 13632 4676
rect 13748 4620 13804 4630
rect 13972 4620 14028 5684
rect 14308 5110 14364 5122
rect 14308 5068 14310 5110
rect 14362 5068 14364 5110
rect 14308 5002 14364 5012
rect 15204 4956 15260 5842
rect 15988 5740 16044 6626
rect 16212 5852 16268 6862
rect 16324 6678 16380 6690
rect 16324 6626 16326 6678
rect 16378 6626 16380 6678
rect 16324 6524 16380 6626
rect 16324 6458 16380 6468
rect 16548 6678 16604 6690
rect 16548 6626 16550 6678
rect 16602 6626 16604 6678
rect 16212 5786 16268 5796
rect 15988 5674 16044 5684
rect 16548 5404 16604 6626
rect 16660 6636 16716 7476
rect 17220 6860 17276 7812
rect 17220 6708 17276 6804
rect 17220 6656 17222 6708
rect 17274 6656 17276 6708
rect 16884 6636 16940 6646
rect 17220 6644 17276 6656
rect 17332 7420 17388 7430
rect 16660 6634 16940 6636
rect 16660 6582 16886 6634
rect 16938 6582 16940 6634
rect 16660 6580 16940 6582
rect 16884 6570 16940 6580
rect 15204 4890 15260 4900
rect 16100 5348 16604 5404
rect 16660 6412 16716 6422
rect 17332 6412 17388 7364
rect 17444 6646 17500 8484
rect 17892 8428 17948 8438
rect 17556 7420 17612 7430
rect 17556 7338 17558 7364
rect 17610 7338 17612 7364
rect 17556 7326 17612 7338
rect 17892 7308 17948 8372
rect 18900 8246 18956 8258
rect 18900 8194 18902 8246
rect 18954 8194 18956 8246
rect 18508 7644 18564 7654
rect 18900 7644 18956 8194
rect 18508 7550 18564 7588
rect 18676 7588 18956 7644
rect 18676 7420 18732 7588
rect 17892 7252 18060 7308
rect 17644 7084 17908 7094
rect 17700 7028 17748 7084
rect 17804 7028 17852 7084
rect 17644 7018 17908 7028
rect 18004 6748 18060 7252
rect 17724 6692 18060 6748
rect 17444 6636 17556 6646
rect 17500 6634 17556 6636
rect 17500 6582 17502 6634
rect 17554 6582 17556 6634
rect 17500 6580 17556 6582
rect 17444 6570 17556 6580
rect 17724 6634 17780 6692
rect 18676 6646 18732 7364
rect 18844 7474 18900 7486
rect 18844 7422 18846 7474
rect 18898 7422 18900 7474
rect 18844 7196 18900 7422
rect 18844 6860 18900 7140
rect 17724 6582 17726 6634
rect 17778 6582 17780 6634
rect 17724 6570 17780 6582
rect 18396 6634 18452 6646
rect 18396 6582 18398 6634
rect 18450 6582 18452 6634
rect 17444 6504 17500 6570
rect 18004 6524 18116 6534
rect 18060 6522 18116 6524
rect 18060 6470 18062 6522
rect 18114 6470 18116 6522
rect 18060 6468 18116 6470
rect 18004 6458 18116 6468
rect 18172 6524 18228 6534
rect 18396 6524 18452 6582
rect 18172 6522 18284 6524
rect 18172 6470 18174 6522
rect 18226 6470 18284 6522
rect 18172 6458 18284 6470
rect 18396 6458 18452 6468
rect 18620 6634 18732 6646
rect 18620 6582 18622 6634
rect 18674 6582 18732 6634
rect 18620 6580 18732 6582
rect 18788 6858 18900 6860
rect 18788 6806 18846 6858
rect 18898 6806 18900 6858
rect 18788 6794 18900 6806
rect 19012 6860 19068 10614
rect 19684 10444 19740 10454
rect 19796 10444 19852 11172
rect 21588 11228 21644 11398
rect 22652 11452 22708 11958
rect 23940 11900 23996 11910
rect 22652 11396 22988 11452
rect 21588 11162 21644 11172
rect 22708 11116 22764 11126
rect 21920 11004 22184 11014
rect 21976 10948 22024 11004
rect 22080 10948 22128 11004
rect 21920 10938 22184 10948
rect 21812 10780 21868 10790
rect 21812 10556 21868 10724
rect 22036 10668 22092 10678
rect 22036 10570 22038 10612
rect 22090 10570 22092 10612
rect 22708 10668 22764 11060
rect 22036 10558 22092 10570
rect 22596 10598 22652 10610
rect 19740 10388 19852 10444
rect 21700 10500 21868 10556
rect 22596 10556 22598 10598
rect 22650 10556 22652 10598
rect 19684 10350 19740 10388
rect 21588 10332 21644 10342
rect 19684 10108 19740 10118
rect 19684 10006 19740 10052
rect 20692 10076 20748 10088
rect 20692 10024 20694 10076
rect 20746 10024 20748 10076
rect 19460 9996 19516 10006
rect 19684 9994 19796 10006
rect 19684 9942 19742 9994
rect 19794 9942 19796 9994
rect 19684 9940 19796 9942
rect 19460 9902 19516 9940
rect 19740 9930 19796 9940
rect 20076 9996 20132 10006
rect 20692 9996 20748 10024
rect 20692 9940 20860 9996
rect 20076 9902 20132 9940
rect 19908 9882 19964 9894
rect 19908 9830 19910 9882
rect 19962 9830 19964 9882
rect 19908 9772 19964 9830
rect 19908 9706 19964 9716
rect 20356 9814 20412 9826
rect 20356 9762 20358 9814
rect 20410 9762 20412 9814
rect 19908 9154 19964 9166
rect 19908 9102 19910 9154
rect 19962 9102 19964 9154
rect 19908 9100 19964 9102
rect 19572 9042 19628 9054
rect 19572 8990 19574 9042
rect 19626 8990 19628 9042
rect 19348 8316 19404 8326
rect 19124 7980 19180 7990
rect 19124 7756 19180 7924
rect 19124 7690 19180 7700
rect 19348 7308 19404 8260
rect 19572 7644 19628 8990
rect 19908 8426 19964 9044
rect 20244 8876 20300 8886
rect 20244 8782 20300 8820
rect 20356 8427 20412 9762
rect 20692 9814 20748 9826
rect 20692 9762 20694 9814
rect 20746 9762 20748 9814
rect 20692 9156 20748 9762
rect 20804 9660 20860 9940
rect 20972 9884 21028 9894
rect 20972 9882 21196 9884
rect 20972 9830 20974 9882
rect 21026 9830 21196 9882
rect 20972 9828 21196 9830
rect 20972 9818 21028 9828
rect 20804 9604 21028 9660
rect 20972 9266 21028 9604
rect 20972 9214 20974 9266
rect 21026 9214 21028 9266
rect 20972 9202 21028 9214
rect 19908 8374 19910 8426
rect 19962 8374 19964 8426
rect 19908 8362 19964 8374
rect 20244 8371 20412 8427
rect 20580 9100 20748 9156
rect 20580 8428 20636 9100
rect 20748 8988 20804 8998
rect 20748 8894 20804 8932
rect 20076 8204 20132 8214
rect 20020 8202 20132 8204
rect 20020 8150 20078 8202
rect 20130 8150 20132 8202
rect 20020 8138 20132 8150
rect 20020 8092 20076 8138
rect 19572 7578 19628 7588
rect 19684 7980 19740 7990
rect 19516 7474 19572 7486
rect 19516 7422 19518 7474
rect 19570 7422 19572 7474
rect 19516 7420 19572 7422
rect 19516 7364 19628 7420
rect 19348 6870 19404 7252
rect 19012 6794 19068 6804
rect 19292 6858 19404 6870
rect 19292 6806 19294 6858
rect 19346 6806 19404 6858
rect 19292 6804 19404 6806
rect 19292 6794 19348 6804
rect 17444 6412 17500 6422
rect 17332 6356 17444 6412
rect 13804 4564 14028 4620
rect 15260 4732 15316 4742
rect 13020 4414 13076 4452
rect 13132 4452 13244 4508
rect 13300 4508 13356 4518
rect 12460 4338 12572 4350
rect 13132 4340 13188 4452
rect 12348 4284 12404 4294
rect 12460 4286 12462 4338
rect 12514 4286 12572 4338
rect 12460 4284 12572 4286
rect 12964 4284 13188 4340
rect 13300 4294 13356 4452
rect 13468 4508 13524 4518
rect 13468 4414 13524 4452
rect 13748 4506 13804 4564
rect 13748 4454 13750 4506
rect 13802 4454 13804 4506
rect 13748 4442 13804 4454
rect 14756 4508 14812 4518
rect 12460 4274 12516 4284
rect 11900 4172 11956 4182
rect 11900 4078 11956 4116
rect 12124 4172 12180 4182
rect 12124 4078 12180 4116
rect 12068 3948 12124 3958
rect 11732 3892 12068 3948
rect 10948 3882 11004 3892
rect 9548 3778 9604 3780
rect 9044 3724 9100 3734
rect 9548 3726 9550 3778
rect 9602 3726 9604 3778
rect 10108 3780 10444 3836
rect 9548 3724 9604 3726
rect 9772 3724 9828 3734
rect 9548 3722 9828 3724
rect 9548 3670 9774 3722
rect 9826 3670 9828 3722
rect 9548 3668 9828 3670
rect 9044 3568 9100 3668
rect 9772 3658 9828 3668
rect 10108 3722 10164 3780
rect 10108 3670 10110 3722
rect 10162 3670 10164 3722
rect 10108 3658 10164 3670
rect 10388 3622 10444 3780
rect 11620 3836 11676 3846
rect 11284 3724 11340 3734
rect 10612 3722 11340 3724
rect 10612 3670 11286 3722
rect 11338 3670 11340 3722
rect 10612 3668 11340 3670
rect 11620 3724 11676 3780
rect 11620 3668 11732 3724
rect 9324 3612 9380 3622
rect 9044 3516 9046 3568
rect 9098 3516 9100 3568
rect 9044 3504 9100 3516
rect 9156 3610 9380 3612
rect 9156 3558 9326 3610
rect 9378 3558 9380 3610
rect 9156 3556 9380 3558
rect 8372 2940 8428 2950
rect 8092 2042 8204 2054
rect 8092 1990 8094 2042
rect 8146 1990 8204 2042
rect 8092 1988 8204 1990
rect 8260 2268 8316 2278
rect 8092 1978 8148 1988
rect 7924 1370 8036 1382
rect 7924 1318 7982 1370
rect 8034 1318 8036 1370
rect 7924 1316 8036 1318
rect 4844 1258 4900 1316
rect 7980 1306 8036 1316
rect 8260 1260 8316 2212
rect 8372 2166 8428 2884
rect 8596 2726 8652 2996
rect 8540 2714 8652 2726
rect 8540 2662 8542 2714
rect 8594 2662 8652 2714
rect 8540 2660 8652 2662
rect 8708 2996 8988 3052
rect 9044 3164 9100 3174
rect 8708 2714 8764 2996
rect 8708 2662 8710 2714
rect 8762 2662 8764 2714
rect 8876 2772 8932 2782
rect 9044 2772 9100 3108
rect 9156 3052 9212 3556
rect 9324 3546 9380 3556
rect 9940 3612 9996 3622
rect 9940 3518 9996 3556
rect 10276 3612 10332 3622
rect 10388 3610 10500 3622
rect 10388 3558 10446 3610
rect 10498 3558 10500 3610
rect 10388 3556 10500 3558
rect 9492 3500 9548 3510
rect 9716 3500 9772 3510
rect 9492 3442 9548 3444
rect 9492 3390 9494 3442
rect 9546 3390 9548 3442
rect 9492 3378 9548 3390
rect 9604 3444 9716 3500
rect 9156 2986 9212 2996
rect 9604 3276 9660 3444
rect 9716 3434 9772 3444
rect 10276 3387 10332 3556
rect 10444 3546 10500 3556
rect 8876 2770 9100 2772
rect 8876 2718 8878 2770
rect 8930 2718 9100 2770
rect 9268 2828 9324 2838
rect 9268 2730 9270 2772
rect 9322 2730 9324 2772
rect 9268 2718 9324 2730
rect 8876 2716 9100 2718
rect 8876 2706 8932 2716
rect 8540 2650 8596 2660
rect 8708 2650 8764 2662
rect 9092 2380 9356 2390
rect 9148 2324 9196 2380
rect 9252 2324 9300 2380
rect 9092 2314 9356 2324
rect 8596 2268 8652 2278
rect 9604 2268 9660 3220
rect 10164 3331 10332 3387
rect 9772 2772 9828 2782
rect 9772 2770 10108 2772
rect 9772 2718 9774 2770
rect 9826 2718 10108 2770
rect 9772 2716 10108 2718
rect 9772 2706 9828 2716
rect 8372 2154 8484 2166
rect 8372 2102 8430 2154
rect 8482 2102 8484 2154
rect 8372 2100 8484 2102
rect 8428 2090 8484 2100
rect 8596 2064 8652 2212
rect 9492 2212 9828 2268
rect 9100 2156 9156 2166
rect 9492 2156 9548 2212
rect 9100 2154 9548 2156
rect 9100 2102 9102 2154
rect 9154 2102 9548 2154
rect 9100 2100 9548 2102
rect 9772 2154 9828 2212
rect 9772 2102 9774 2154
rect 9826 2102 9828 2154
rect 9100 2090 9156 2100
rect 9772 2090 9828 2102
rect 10052 2154 10108 2716
rect 10164 2268 10220 3331
rect 10164 2202 10220 2212
rect 10052 2102 10054 2154
rect 10106 2102 10108 2154
rect 10052 2090 10108 2102
rect 10444 2156 10500 2166
rect 10612 2156 10668 3668
rect 11284 3658 11340 3668
rect 11396 3612 11452 3622
rect 10836 3554 10892 3566
rect 10724 3500 10780 3510
rect 10724 3396 10726 3444
rect 10778 3396 10780 3444
rect 10724 3384 10780 3396
rect 10836 3502 10838 3554
rect 10890 3502 10892 3554
rect 11396 3510 11452 3556
rect 10836 3387 10892 3502
rect 11116 3498 11172 3510
rect 11116 3446 11118 3498
rect 11170 3446 11172 3498
rect 11116 3388 11172 3446
rect 11340 3498 11452 3510
rect 11340 3446 11342 3498
rect 11394 3446 11452 3498
rect 11340 3444 11452 3446
rect 11508 3500 11620 3510
rect 11564 3498 11620 3500
rect 11564 3446 11566 3498
rect 11618 3446 11620 3498
rect 11564 3444 11620 3446
rect 11340 3434 11396 3444
rect 11508 3434 11620 3444
rect 10836 3331 11004 3387
rect 10948 2940 11004 3331
rect 11116 3322 11172 3332
rect 11676 3276 11732 3668
rect 11788 3612 11844 3622
rect 11788 3610 11900 3612
rect 11788 3558 11790 3610
rect 11842 3558 11900 3610
rect 11788 3546 11900 3558
rect 11844 3500 11900 3546
rect 12068 3566 12124 3892
rect 12348 3722 12404 4228
rect 12628 4172 12684 4182
rect 12628 4078 12684 4116
rect 12964 3734 13020 4284
rect 13244 4282 13356 4294
rect 13244 4230 13246 4282
rect 13298 4230 13356 4282
rect 13860 4396 13916 4406
rect 13860 4338 13916 4340
rect 13860 4286 13862 4338
rect 13914 4286 13916 4338
rect 13860 4274 13916 4286
rect 14644 4396 14700 4406
rect 14644 4282 14700 4340
rect 13244 4228 13356 4230
rect 13244 4218 13300 4228
rect 14420 4226 14476 4238
rect 12348 3670 12350 3722
rect 12402 3670 12404 3722
rect 12348 3658 12404 3670
rect 12908 3722 13020 3734
rect 12908 3670 12910 3722
rect 12962 3670 13020 3722
rect 12908 3658 13020 3670
rect 13132 4172 13188 4182
rect 13132 3722 13188 4116
rect 13132 3670 13134 3722
rect 13186 3670 13188 3722
rect 13132 3658 13188 3670
rect 13524 4172 13580 4182
rect 13524 3836 13580 4116
rect 12068 3514 12070 3566
rect 12122 3514 12124 3566
rect 12068 3502 12124 3514
rect 11844 3434 11900 3444
rect 11956 3388 12012 3398
rect 12460 3388 12516 3426
rect 12012 3332 12236 3387
rect 11956 3331 12236 3332
rect 11956 3322 12012 3331
rect 10948 2874 11004 2884
rect 11620 3220 11732 3276
rect 11396 2604 11452 2614
rect 10444 2154 10668 2156
rect 10444 2102 10446 2154
rect 10498 2102 10668 2154
rect 10444 2100 10668 2102
rect 10724 2268 10780 2278
rect 10444 2090 10500 2100
rect 8596 2012 8598 2064
rect 8650 2012 8652 2064
rect 8596 2000 8652 2012
rect 8988 2044 9044 2054
rect 8988 1950 9044 1988
rect 10724 1942 10780 2212
rect 11396 2166 11452 2548
rect 11396 2154 11508 2166
rect 11396 2102 11454 2154
rect 11506 2102 11508 2154
rect 11396 2100 11508 2102
rect 11452 2090 11508 2100
rect 11620 2042 11676 3220
rect 12068 2602 12124 2614
rect 12068 2550 12070 2602
rect 12122 2550 12124 2602
rect 12068 2380 12124 2550
rect 12068 2314 12124 2324
rect 11788 2156 11844 2166
rect 12180 2156 12236 3331
rect 12460 3322 12516 3332
rect 12964 3052 13020 3658
rect 13524 3610 13580 3780
rect 14420 4174 14422 4226
rect 14474 4174 14476 4226
rect 14644 4230 14646 4282
rect 14698 4230 14700 4282
rect 14644 4218 14700 4230
rect 14420 3836 14476 4174
rect 14420 3770 14476 3780
rect 13524 3558 13526 3610
rect 13578 3558 13580 3610
rect 13524 3546 13580 3558
rect 13804 3612 13860 3622
rect 14196 3612 14252 3622
rect 13804 3518 13860 3556
rect 14028 3554 14084 3566
rect 14028 3502 14030 3554
rect 14082 3502 14084 3554
rect 13860 3388 13916 3426
rect 14028 3387 14084 3502
rect 13860 3322 13916 3332
rect 13972 3331 14084 3387
rect 11788 2154 12236 2156
rect 11788 2102 11790 2154
rect 11842 2102 12236 2154
rect 11788 2100 12236 2102
rect 12292 2940 12348 2950
rect 11788 2090 11844 2100
rect 12292 2044 12348 2884
rect 12740 2940 12796 2950
rect 12740 2846 12796 2884
rect 12964 2828 13020 2996
rect 12516 2716 12572 2726
rect 11620 1990 11622 2042
rect 11674 1990 11676 2042
rect 11620 1978 11676 1990
rect 12124 1988 12348 2044
rect 12404 2492 12460 2502
rect 8596 1932 8652 1942
rect 8596 1838 8652 1876
rect 9324 1932 9380 1942
rect 9548 1932 9604 1942
rect 9324 1930 9604 1932
rect 9324 1878 9326 1930
rect 9378 1878 9550 1930
rect 9602 1878 9604 1930
rect 9324 1876 9604 1878
rect 9324 1708 9380 1876
rect 9548 1866 9604 1876
rect 10668 1930 10780 1942
rect 10668 1878 10670 1930
rect 10722 1878 10780 1930
rect 10668 1876 10780 1878
rect 11228 1930 11284 1942
rect 11228 1878 11230 1930
rect 11282 1878 11284 1930
rect 10668 1866 10724 1876
rect 9324 1642 9380 1652
rect 11228 1708 11284 1878
rect 12124 1930 12180 1988
rect 12124 1878 12126 1930
rect 12178 1878 12180 1930
rect 12124 1866 12180 1878
rect 12404 1880 12460 2436
rect 12516 1986 12572 2660
rect 12516 1934 12518 1986
rect 12570 1934 12572 1986
rect 12516 1922 12572 1934
rect 12404 1828 12406 1880
rect 12458 1828 12460 1880
rect 12404 1816 12460 1828
rect 12964 1820 13020 2772
rect 13188 3164 13244 3174
rect 13188 2790 13244 3108
rect 13368 3164 13632 3174
rect 13424 3108 13472 3164
rect 13528 3108 13576 3164
rect 13368 3098 13632 3108
rect 13356 2940 13412 2950
rect 13356 2846 13412 2884
rect 13188 2738 13190 2790
rect 13242 2738 13244 2790
rect 13076 2716 13132 2726
rect 13076 2054 13132 2660
rect 13188 2604 13244 2738
rect 13580 2770 13636 2782
rect 13972 2772 14028 3331
rect 13580 2718 13582 2770
rect 13634 2718 13636 2770
rect 13580 2716 13636 2718
rect 13580 2650 13636 2660
rect 13748 2716 14028 2772
rect 14084 2716 14140 2726
rect 13188 2538 13244 2548
rect 13300 2602 13356 2614
rect 13300 2550 13302 2602
rect 13354 2550 13356 2602
rect 13300 2156 13356 2550
rect 13748 2166 13804 2716
rect 13972 2604 14028 2614
rect 13972 2510 14028 2548
rect 13300 2090 13356 2100
rect 13692 2154 13804 2166
rect 13692 2102 13694 2154
rect 13746 2102 13804 2154
rect 13692 2100 13804 2102
rect 13692 2090 13748 2100
rect 13076 2042 13188 2054
rect 13076 1990 13134 2042
rect 13186 1990 13188 2042
rect 13076 1988 13188 1990
rect 13132 1978 13188 1988
rect 14084 1994 14140 2660
rect 14196 2166 14252 3556
rect 14420 3554 14476 3566
rect 14420 3502 14422 3554
rect 14474 3502 14476 3554
rect 14308 3276 14364 3286
rect 14308 2782 14364 3220
rect 14308 2730 14310 2782
rect 14362 2730 14364 2782
rect 14308 2718 14364 2730
rect 14420 2604 14476 3502
rect 14756 3548 14812 4452
rect 15092 4396 15148 4406
rect 14924 4060 14980 4070
rect 15092 4060 15148 4340
rect 15260 4338 15316 4676
rect 16100 4620 16156 5348
rect 16660 5292 16716 6356
rect 17444 5918 17500 6356
rect 17444 5866 17446 5918
rect 17498 5866 17500 5918
rect 17444 5854 17500 5866
rect 17644 5516 17908 5526
rect 17700 5460 17748 5516
rect 17804 5460 17852 5516
rect 17644 5450 17908 5460
rect 18004 5292 18060 6458
rect 18228 6076 18284 6458
rect 18620 6412 18676 6580
rect 18620 6346 18676 6356
rect 18452 6076 18508 6086
rect 18788 6076 18844 6794
rect 19572 6748 19628 7364
rect 19572 6682 19628 6692
rect 19684 6646 19740 7924
rect 20020 7196 20076 8036
rect 20244 7980 20300 8371
rect 20580 8362 20636 8372
rect 20916 8764 20972 8774
rect 20916 8270 20972 8708
rect 21140 8540 21196 9828
rect 21364 9882 21420 9894
rect 21364 9830 21366 9882
rect 21418 9830 21420 9882
rect 21364 9164 21420 9830
rect 21364 9112 21366 9164
rect 21418 9112 21420 9164
rect 21364 9100 21420 9112
rect 21476 9772 21532 9782
rect 21252 9022 21308 9034
rect 21252 8970 21254 9022
rect 21306 8970 21308 9022
rect 21476 8998 21532 9716
rect 21588 9324 21644 10276
rect 21700 9994 21756 10500
rect 22596 10490 22652 10500
rect 22428 9996 22484 10006
rect 21700 9942 21702 9994
rect 21754 9942 21756 9994
rect 21700 9548 21756 9942
rect 22036 9940 22428 9996
rect 22036 9660 22092 9940
rect 22428 9864 22484 9940
rect 22596 9884 22652 9894
rect 22204 9826 22260 9838
rect 22204 9774 22206 9826
rect 22258 9774 22260 9826
rect 22204 9660 22260 9774
rect 22372 9660 22428 9670
rect 22204 9604 22316 9660
rect 22036 9594 22092 9604
rect 21700 9482 21756 9492
rect 21920 9436 22184 9446
rect 21976 9380 22024 9436
rect 22080 9380 22128 9436
rect 21920 9370 22184 9380
rect 21588 9268 21868 9324
rect 21812 9212 21868 9268
rect 22092 9212 22148 9222
rect 21812 9210 22148 9212
rect 21812 9158 22094 9210
rect 22146 9158 22148 9210
rect 21812 9156 22148 9158
rect 22092 9146 22148 9156
rect 21252 8652 21308 8970
rect 21420 8986 21532 8998
rect 21420 8934 21422 8986
rect 21474 8934 21532 8986
rect 21420 8932 21532 8934
rect 22148 9034 22204 9046
rect 22148 8988 22150 9034
rect 22202 8988 22204 9034
rect 21420 8922 21476 8932
rect 22148 8922 22204 8932
rect 21644 8876 21700 8886
rect 21644 8782 21700 8820
rect 21252 8596 21532 8652
rect 21476 8540 21532 8596
rect 21028 8482 21084 8494
rect 21140 8484 21420 8540
rect 21028 8430 21030 8482
rect 21082 8430 21084 8482
rect 21028 8428 21084 8430
rect 21028 8362 21084 8372
rect 20244 7914 20300 7924
rect 20580 8246 20636 8258
rect 20580 8194 20582 8246
rect 20634 8194 20636 8246
rect 20916 8218 20918 8270
rect 20970 8218 20972 8270
rect 21196 8316 21252 8326
rect 21196 8222 21252 8260
rect 20580 7980 20636 8194
rect 20748 8204 20860 8214
rect 20916 8206 20972 8218
rect 20748 8202 20804 8204
rect 20748 8150 20750 8202
rect 20802 8150 20804 8202
rect 20748 8148 20804 8150
rect 20748 8138 20860 8148
rect 20580 7914 20636 7924
rect 20020 7130 20076 7140
rect 21364 7532 21420 8484
rect 20916 6883 20972 6895
rect 20524 6860 20580 6870
rect 20916 6860 20918 6883
rect 20524 6858 20918 6860
rect 20524 6806 20526 6858
rect 20578 6831 20918 6858
rect 20970 6831 20972 6883
rect 20578 6806 20972 6831
rect 20524 6804 20972 6806
rect 20524 6794 20580 6804
rect 20132 6748 20188 6758
rect 20132 6654 20188 6692
rect 21364 6690 21420 7476
rect 19404 6636 19460 6646
rect 19684 6634 19796 6646
rect 19684 6582 19742 6634
rect 19794 6582 19796 6634
rect 21364 6638 21366 6690
rect 21418 6638 21420 6690
rect 21476 6748 21532 8484
rect 22260 8427 22316 9604
rect 22372 9566 22428 9604
rect 22596 9436 22652 9828
rect 22428 9380 22652 9436
rect 22428 9210 22484 9380
rect 22428 9158 22430 9210
rect 22482 9158 22484 9210
rect 22428 9146 22484 9158
rect 22708 9100 22764 10612
rect 22820 10444 22876 10454
rect 22820 10350 22876 10388
rect 22708 9034 22764 9044
rect 22820 9882 22876 9894
rect 22820 9830 22822 9882
rect 22874 9830 22876 9882
rect 22820 9772 22876 9830
rect 22932 9782 22988 11396
rect 23940 11382 23996 11844
rect 23940 11340 23942 11382
rect 23994 11340 23996 11382
rect 24500 11564 24556 11574
rect 24500 11406 24556 11508
rect 24500 11354 24502 11406
rect 24554 11354 24556 11406
rect 24500 11342 24556 11354
rect 24724 11452 24780 12114
rect 25396 12166 25452 12178
rect 25396 12124 25398 12166
rect 25450 12124 25452 12166
rect 28756 12126 28758 12178
rect 28810 12126 28812 12178
rect 28756 12114 28812 12126
rect 30660 12166 30716 12178
rect 30660 12114 30662 12166
rect 30714 12114 30716 12166
rect 25396 12058 25452 12068
rect 27636 12056 27692 12068
rect 27636 12004 27638 12056
rect 27690 12004 27692 12056
rect 26068 11900 26124 11910
rect 23940 11274 23996 11284
rect 24724 10892 24780 11396
rect 25116 11452 25172 11462
rect 26068 11452 26124 11844
rect 26196 11788 26460 11798
rect 26252 11732 26300 11788
rect 26356 11732 26404 11788
rect 26196 11722 26460 11732
rect 25116 11450 25228 11452
rect 25116 11398 25118 11450
rect 25170 11398 25228 11450
rect 25116 11386 25228 11398
rect 25004 11228 25060 11238
rect 24724 10826 24780 10836
rect 24836 11226 25060 11228
rect 24836 11174 25006 11226
rect 25058 11174 25060 11226
rect 24836 11172 25060 11174
rect 23492 10444 23548 10454
rect 22932 9772 23044 9782
rect 22820 9716 22988 9772
rect 22652 8874 22708 8886
rect 22652 8822 22654 8874
rect 22706 8822 22708 8874
rect 22652 8427 22708 8822
rect 22820 8876 22876 9716
rect 22988 9678 23044 9716
rect 23492 9770 23548 10388
rect 24836 10220 24892 11172
rect 25004 11162 25060 11172
rect 25172 11228 25228 11386
rect 26068 11354 26070 11396
rect 26122 11354 26124 11396
rect 26068 11342 26124 11354
rect 26740 11452 26796 11462
rect 26740 11354 26742 11396
rect 26794 11354 26796 11396
rect 26740 11342 26796 11354
rect 27188 11340 27244 11350
rect 24276 10164 24892 10220
rect 25004 10498 25060 10510
rect 25004 10446 25006 10498
rect 25058 10446 25060 10498
rect 25004 10444 25060 10446
rect 23492 9718 23494 9770
rect 23546 9718 23548 9770
rect 23492 9706 23548 9718
rect 23716 9826 23772 9838
rect 23716 9774 23718 9826
rect 23770 9774 23772 9826
rect 23044 9548 23100 9558
rect 23044 9054 23100 9492
rect 23716 9212 23772 9774
rect 23716 9146 23772 9156
rect 23044 9002 23046 9054
rect 23098 9002 23100 9054
rect 23044 8990 23100 9002
rect 23604 9030 23660 9042
rect 22820 8810 22876 8820
rect 23604 8978 23606 9030
rect 23658 8978 23660 9030
rect 23604 8540 23660 8978
rect 23604 8474 23660 8484
rect 22260 8371 22372 8427
rect 22652 8371 23100 8427
rect 21588 8246 21644 8258
rect 21588 8194 21590 8246
rect 21642 8194 21644 8246
rect 21588 8092 21644 8194
rect 21588 8026 21644 8036
rect 22316 8146 22372 8371
rect 22316 8094 22318 8146
rect 22370 8094 22372 8146
rect 21920 7868 22184 7878
rect 21976 7812 22024 7868
rect 22080 7812 22128 7868
rect 21920 7802 22184 7812
rect 22316 7644 22372 8094
rect 22708 8092 22764 8371
rect 22708 8026 22764 8036
rect 22260 7588 22372 7644
rect 21700 7462 21756 7474
rect 21700 7420 21702 7462
rect 21754 7420 21756 7462
rect 21700 7354 21756 7364
rect 21476 6682 21532 6692
rect 21364 6626 21420 6638
rect 21812 6634 21868 6646
rect 19684 6580 19796 6582
rect 19404 6542 19460 6580
rect 19740 6570 19796 6580
rect 21812 6582 21814 6634
rect 21866 6582 21868 6634
rect 19852 6524 19908 6534
rect 19852 6430 19908 6468
rect 18228 6074 18508 6076
rect 18228 6022 18454 6074
rect 18506 6022 18508 6074
rect 18228 6020 18508 6022
rect 18452 6010 18508 6020
rect 18564 6020 18844 6076
rect 19684 6412 19740 6422
rect 15428 4508 15484 4518
rect 15428 4414 15484 4452
rect 16100 4506 16156 4564
rect 16100 4454 16102 4506
rect 16154 4454 16156 4506
rect 16100 4442 16156 4454
rect 16436 5236 16716 5292
rect 17892 5236 18060 5292
rect 18340 5292 18396 5302
rect 15260 4286 15262 4338
rect 15314 4286 15316 4338
rect 16436 4334 16492 5236
rect 16604 5234 16660 5236
rect 16604 5182 16606 5234
rect 16658 5182 16660 5234
rect 16604 5170 16660 5182
rect 17780 5068 17836 5078
rect 17892 5068 17948 5236
rect 17780 5066 17948 5068
rect 17780 5014 17782 5066
rect 17834 5014 17948 5066
rect 17780 5012 17948 5014
rect 18004 5122 18060 5134
rect 18004 5070 18006 5122
rect 18058 5070 18060 5122
rect 17780 5002 17836 5012
rect 17500 4954 17556 4966
rect 17500 4902 17502 4954
rect 17554 4902 17556 4954
rect 17500 4844 17556 4902
rect 17500 4778 17556 4788
rect 18004 4844 18060 5070
rect 18004 4778 18060 4788
rect 17892 4732 17948 4742
rect 15260 4274 15316 4286
rect 15876 4284 15932 4294
rect 15484 4114 15540 4126
rect 15484 4062 15486 4114
rect 15538 4062 15540 4114
rect 15484 4060 15540 4062
rect 15092 4004 15204 4060
rect 14924 3836 14980 4004
rect 15148 3948 15204 4004
rect 15484 3994 15540 4004
rect 15876 3948 15932 4228
rect 15148 3892 15260 3948
rect 14924 3778 14980 3780
rect 14924 3726 14926 3778
rect 14978 3726 14980 3778
rect 14924 3714 14980 3726
rect 15204 3622 15260 3892
rect 15876 3882 15932 3892
rect 16380 4278 16492 4334
rect 17332 4396 17388 4406
rect 17332 4298 17334 4340
rect 17386 4298 17388 4340
rect 16716 4284 16772 4294
rect 17332 4286 17388 4298
rect 17892 4338 17948 4676
rect 18340 4518 18396 5236
rect 18284 4506 18396 4518
rect 17892 4286 17894 4338
rect 17946 4286 17948 4338
rect 18004 4444 18060 4456
rect 18004 4396 18006 4444
rect 18058 4396 18060 4444
rect 18284 4454 18286 4506
rect 18338 4454 18396 4506
rect 18284 4452 18396 4454
rect 18284 4442 18340 4452
rect 18004 4330 18060 4340
rect 14756 3500 14758 3548
rect 14810 3500 14812 3548
rect 15148 3610 15260 3622
rect 15148 3558 15150 3610
rect 15202 3558 15260 3610
rect 15148 3556 15260 3558
rect 16380 3722 16436 4278
rect 17892 4274 17948 4286
rect 16716 4190 16772 4228
rect 16492 4172 16548 4182
rect 16940 4172 16996 4182
rect 16492 4170 16604 4172
rect 16492 4118 16494 4170
rect 16546 4118 16604 4170
rect 16492 4106 16604 4118
rect 16380 3670 16382 3722
rect 16434 3670 16436 3722
rect 15148 3546 15204 3556
rect 14756 3434 14812 3444
rect 15036 3500 15092 3510
rect 15036 3406 15092 3444
rect 15708 3500 15764 3510
rect 15708 3406 15764 3444
rect 15484 3388 15540 3398
rect 16044 3388 16100 3398
rect 15484 3294 15540 3332
rect 15876 3386 16100 3388
rect 16380 3387 16436 3670
rect 15876 3334 16046 3386
rect 16098 3334 16100 3386
rect 15876 3332 16100 3334
rect 14756 3052 14812 3062
rect 14420 2538 14476 2548
rect 14532 2940 14588 2950
rect 14532 2390 14588 2884
rect 14756 2778 14812 2996
rect 14756 2726 14758 2778
rect 14810 2726 14812 2778
rect 14756 2714 14812 2726
rect 15372 2770 15428 2782
rect 15372 2718 15374 2770
rect 15426 2718 15428 2770
rect 15372 2716 15428 2718
rect 15372 2660 15484 2716
rect 14532 2380 14644 2390
rect 14532 2324 14588 2380
rect 14196 2154 14308 2166
rect 14196 2102 14254 2154
rect 14306 2102 14308 2154
rect 14196 2100 14308 2102
rect 14252 2090 14308 2100
rect 14588 2154 14644 2324
rect 14588 2102 14590 2154
rect 14642 2102 14644 2154
rect 14588 2090 14644 2102
rect 15316 2156 15372 2166
rect 15428 2156 15484 2660
rect 15764 2156 15820 2166
rect 15428 2154 15820 2156
rect 15428 2102 15766 2154
rect 15818 2102 15820 2154
rect 15428 2100 15820 2102
rect 14084 1942 14086 1994
rect 14138 1942 14140 1994
rect 15316 1996 15372 2100
rect 15764 2090 15820 2100
rect 13356 1932 13412 1942
rect 14084 1930 14140 1942
rect 14364 1932 14420 1942
rect 15316 1940 15652 1996
rect 13356 1838 13412 1876
rect 14364 1838 14420 1876
rect 15540 1930 15652 1940
rect 15540 1878 15598 1930
rect 15650 1878 15652 1930
rect 15540 1866 15652 1878
rect 12964 1764 13188 1820
rect 11228 1642 11284 1652
rect 4844 1206 4846 1258
rect 4898 1206 4900 1258
rect 4844 1194 4900 1206
rect 8148 1204 8316 1260
rect 12908 1596 12964 1606
rect 12908 1258 12964 1540
rect 12908 1206 12910 1258
rect 12962 1206 12964 1258
rect 7868 1148 7924 1158
rect 8148 1148 8204 1204
rect 12908 1194 12964 1206
rect 13132 1258 13188 1764
rect 15372 1818 15428 1830
rect 15372 1766 15374 1818
rect 15426 1766 15428 1818
rect 15372 1708 15428 1766
rect 15540 1820 15596 1866
rect 15540 1754 15596 1764
rect 15372 1642 15428 1652
rect 15876 1708 15932 3332
rect 16044 3322 16100 3332
rect 16324 3331 16436 3387
rect 16548 3388 16604 4106
rect 16884 4170 16996 4172
rect 16884 4118 16942 4170
rect 16994 4118 16996 4170
rect 16884 4106 16996 4118
rect 17668 4172 17724 4182
rect 17668 4170 18060 4172
rect 17668 4118 17670 4170
rect 17722 4118 18060 4170
rect 17668 4116 18060 4118
rect 17668 4106 17724 4116
rect 16660 3724 16716 3734
rect 16660 3630 16716 3668
rect 16884 3724 16940 4106
rect 17644 3948 17908 3958
rect 17700 3892 17748 3948
rect 17804 3892 17852 3948
rect 17644 3882 17908 3892
rect 16884 3668 17388 3724
rect 16324 2940 16380 3331
rect 16548 3322 16604 3332
rect 16324 2874 16380 2884
rect 16884 3052 16940 3668
rect 17332 3566 17388 3668
rect 18004 3566 18060 4116
rect 15988 2828 16044 2838
rect 15988 2002 16044 2772
rect 15988 1950 15990 2002
rect 16042 1950 16044 2002
rect 16156 2604 16212 2614
rect 16156 2042 16212 2548
rect 16884 2156 16940 2996
rect 16996 3542 17052 3554
rect 16996 3490 16998 3542
rect 17050 3490 17052 3542
rect 17332 3514 17334 3566
rect 17386 3514 17388 3566
rect 17332 3502 17388 3514
rect 17948 3554 18060 3566
rect 17948 3502 17950 3554
rect 18002 3502 18060 3554
rect 17948 3500 18060 3502
rect 17948 3490 18004 3500
rect 16996 2828 17052 3490
rect 18564 3387 18620 6020
rect 19460 5898 19516 5910
rect 18844 5852 18900 5862
rect 18844 5758 18900 5796
rect 19180 5850 19236 5862
rect 19180 5798 19182 5850
rect 19234 5798 19236 5850
rect 18676 5315 18732 5327
rect 18676 5263 18678 5315
rect 18730 5263 18732 5315
rect 18676 4956 18732 5263
rect 19180 5292 19236 5798
rect 19460 5852 19462 5898
rect 19514 5852 19516 5898
rect 19460 5786 19516 5796
rect 19292 5740 19348 5750
rect 19292 5738 19404 5740
rect 19292 5686 19294 5738
rect 19346 5686 19404 5738
rect 19292 5674 19404 5686
rect 19348 5628 19404 5674
rect 19684 5628 19740 6356
rect 21812 6412 21868 6582
rect 22092 6634 22148 6646
rect 22092 6582 22094 6634
rect 22146 6582 22148 6634
rect 22092 6524 22148 6582
rect 22260 6524 22316 7588
rect 22708 7532 22764 7542
rect 22708 7438 22764 7476
rect 23044 7461 23100 8371
rect 24276 8316 24332 10164
rect 25004 10108 25060 10388
rect 25004 10042 25060 10052
rect 24388 10019 24444 10034
rect 24388 9996 24390 10019
rect 24442 9996 24444 10019
rect 24388 9930 24444 9940
rect 25060 9772 25116 9782
rect 24500 9770 25116 9772
rect 24500 9718 25062 9770
rect 25114 9718 25116 9770
rect 24500 9716 25116 9718
rect 24500 8426 24556 9716
rect 25060 9706 25116 9716
rect 25172 9548 25228 11172
rect 25340 11228 25396 11238
rect 25340 11226 25564 11228
rect 25340 11174 25342 11226
rect 25394 11174 25564 11226
rect 25340 11172 25564 11174
rect 25340 11162 25396 11172
rect 25508 10108 25564 11172
rect 25676 11226 25732 11238
rect 25676 11174 25678 11226
rect 25730 11174 25732 11226
rect 25676 10780 25732 11174
rect 25788 11228 25844 11238
rect 25788 11134 25844 11172
rect 26964 11228 27020 11238
rect 25676 10724 25900 10780
rect 24948 9492 25228 9548
rect 25284 9826 25340 9838
rect 25284 9774 25286 9826
rect 25338 9774 25340 9826
rect 24948 8427 25004 9492
rect 25284 8764 25340 9774
rect 25284 8698 25340 8708
rect 25396 8482 25452 8494
rect 24500 8374 24502 8426
rect 24554 8374 24556 8426
rect 24500 8362 24556 8374
rect 24836 8371 25004 8427
rect 25060 8428 25116 8438
rect 24276 8250 24332 8260
rect 24836 7644 24892 8371
rect 25060 8270 25116 8372
rect 25060 8218 25062 8270
rect 25114 8218 25116 8270
rect 25396 8430 25398 8482
rect 25450 8430 25452 8482
rect 25060 8206 25116 8218
rect 25284 8246 25340 8258
rect 25172 8204 25228 8214
rect 23044 7409 23046 7461
rect 23098 7409 23100 7461
rect 23044 7196 23100 7409
rect 23044 7130 23100 7140
rect 23492 7462 23548 7474
rect 23492 7410 23494 7462
rect 23546 7410 23548 7462
rect 23380 6690 23436 6702
rect 22148 6468 22316 6524
rect 22092 6458 22148 6468
rect 21812 6346 21868 6356
rect 21920 6300 22184 6310
rect 21976 6244 22024 6300
rect 22080 6244 22128 6300
rect 21920 6234 22184 6244
rect 19908 5894 19964 5906
rect 19908 5852 19910 5894
rect 19962 5852 19964 5894
rect 19964 5796 20076 5852
rect 19908 5786 19964 5796
rect 19348 5572 19572 5628
rect 19684 5572 19964 5628
rect 19516 5346 19572 5572
rect 19516 5294 19518 5346
rect 19570 5294 19572 5346
rect 19180 5236 19292 5292
rect 19516 5282 19572 5294
rect 19740 5404 19796 5414
rect 19740 5346 19796 5348
rect 19740 5294 19742 5346
rect 19794 5294 19796 5346
rect 19740 5282 19796 5294
rect 19068 4956 19124 4966
rect 18676 4954 19124 4956
rect 18676 4902 19070 4954
rect 19122 4902 19124 4954
rect 18676 4900 19124 4902
rect 19068 4890 19124 4900
rect 19012 4732 19068 4742
rect 18844 4620 18900 4630
rect 18844 4396 18900 4564
rect 18844 4302 18900 4340
rect 19012 3724 19068 4676
rect 19124 4620 19180 4630
rect 19124 4294 19180 4564
rect 19236 4508 19292 5236
rect 19348 5102 19404 5114
rect 19348 5068 19350 5102
rect 19402 5068 19404 5102
rect 19348 5002 19404 5012
rect 19628 5066 19684 5078
rect 19628 5014 19630 5066
rect 19682 5014 19684 5066
rect 19628 4732 19684 5014
rect 19908 4956 19964 5572
rect 20020 5078 20076 5796
rect 20636 5794 20692 5806
rect 20636 5742 20638 5794
rect 20690 5742 20692 5794
rect 20636 5292 20692 5742
rect 22260 5628 22316 6468
rect 22484 6678 22540 6690
rect 22484 6626 22486 6678
rect 22538 6626 22540 6678
rect 22484 6524 22540 6626
rect 22820 6636 22876 6646
rect 22820 6542 22876 6580
rect 23156 6634 23212 6646
rect 23156 6582 23158 6634
rect 23210 6582 23212 6634
rect 22484 6458 22540 6468
rect 22820 5852 22876 5862
rect 22820 5758 22876 5796
rect 22260 5562 22316 5572
rect 20580 5236 20692 5292
rect 20132 5124 20468 5180
rect 20132 5078 20188 5124
rect 20020 5066 20188 5078
rect 20020 5014 20078 5066
rect 20130 5014 20188 5066
rect 20412 5122 20468 5124
rect 20412 5070 20414 5122
rect 20466 5070 20468 5122
rect 20412 5058 20468 5070
rect 20020 5012 20188 5014
rect 20076 4936 20188 5012
rect 19908 4890 19964 4900
rect 19236 4442 19292 4452
rect 19460 4676 19684 4732
rect 19124 4282 19236 4294
rect 19124 4230 19182 4282
rect 19234 4230 19236 4282
rect 19124 4228 19236 4230
rect 19180 4218 19236 4228
rect 19460 4282 19516 4676
rect 19796 4620 19852 4630
rect 20020 4620 20076 4630
rect 19796 4506 19852 4564
rect 19796 4454 19798 4506
rect 19850 4454 19852 4506
rect 19796 4442 19852 4454
rect 19908 4564 20020 4620
rect 19908 4396 19964 4564
rect 20020 4554 20076 4564
rect 19908 4330 19964 4340
rect 19460 4230 19462 4282
rect 19514 4230 19516 4282
rect 19460 4218 19516 4230
rect 19012 3387 19068 3668
rect 20132 4192 20188 4936
rect 20356 4956 20412 4966
rect 20132 4170 20244 4192
rect 20132 4118 20190 4170
rect 20242 4118 20244 4170
rect 20132 4106 20244 4118
rect 20356 4182 20412 4900
rect 20580 4396 20636 5236
rect 21196 5010 21252 5022
rect 21196 4958 21198 5010
rect 21250 4958 21252 5010
rect 21196 4620 21252 4958
rect 22932 4956 22988 4966
rect 21920 4732 22184 4742
rect 21976 4676 22024 4732
rect 22080 4676 22128 4732
rect 21920 4666 22184 4676
rect 21196 4564 21364 4620
rect 20692 4508 20748 4518
rect 20692 4414 20748 4452
rect 20580 4330 20636 4340
rect 21084 4396 21140 4406
rect 21084 4302 21140 4340
rect 21308 4226 21364 4564
rect 22708 4508 22764 4518
rect 22708 4506 22876 4508
rect 22708 4454 22710 4506
rect 22762 4454 22876 4506
rect 22708 4452 22876 4454
rect 22708 4442 22764 4452
rect 20356 4172 20468 4182
rect 20356 4116 20412 4172
rect 18564 3331 18732 3387
rect 19012 3331 19180 3387
rect 16996 2762 17052 2772
rect 17556 2940 17612 2950
rect 17556 2686 17612 2884
rect 17556 2634 17558 2686
rect 17610 2634 17612 2686
rect 17556 2622 17612 2634
rect 18116 2940 18172 2950
rect 18116 2492 18172 2884
rect 18508 2828 18564 2838
rect 18452 2826 18564 2828
rect 18452 2774 18510 2826
rect 18562 2774 18564 2826
rect 18452 2762 18564 2774
rect 18452 2716 18508 2762
rect 18452 2650 18508 2660
rect 17644 2380 17908 2390
rect 17700 2324 17748 2380
rect 17804 2324 17852 2380
rect 18116 2380 18172 2436
rect 18116 2324 18228 2380
rect 17644 2314 17908 2324
rect 16884 2090 16940 2100
rect 17724 2156 17780 2166
rect 16156 1990 16158 2042
rect 16210 1990 16212 2042
rect 16156 1978 16212 1990
rect 17612 2044 17668 2054
rect 17612 1950 17668 1988
rect 15988 1938 16044 1950
rect 15876 1642 15932 1652
rect 17724 1708 17780 2100
rect 18060 2156 18116 2166
rect 18060 2062 18116 2100
rect 18172 2154 18228 2324
rect 18676 2166 18732 3331
rect 19124 2940 19180 3331
rect 19404 3164 19460 3174
rect 19124 2884 19236 2940
rect 19180 2770 19236 2884
rect 19012 2716 19068 2726
rect 19180 2718 19182 2770
rect 19234 2718 19236 2770
rect 19180 2706 19236 2718
rect 19012 2622 19068 2660
rect 18788 2604 18900 2614
rect 18844 2602 18900 2604
rect 18844 2550 18846 2602
rect 18898 2550 18900 2602
rect 18844 2548 18900 2550
rect 18788 2538 18900 2548
rect 19404 2602 19460 3108
rect 20132 3164 20188 4106
rect 20356 4078 20468 4116
rect 21308 4174 21310 4226
rect 21362 4174 21364 4226
rect 20244 3724 20300 3734
rect 20356 3724 20412 4078
rect 21308 3836 21364 4174
rect 21308 3770 21364 3780
rect 21700 4320 21756 4332
rect 21700 4268 21702 4320
rect 21754 4268 21756 4320
rect 20244 3722 20412 3724
rect 20244 3670 20246 3722
rect 20298 3670 20412 3722
rect 20244 3668 20412 3670
rect 20244 3658 20300 3668
rect 21700 3612 21756 4268
rect 22036 4284 22092 4294
rect 22428 4284 22484 4294
rect 22092 4228 22316 4284
rect 22036 4190 22092 4228
rect 22260 3724 22316 4228
rect 22428 4190 22484 4228
rect 22652 4114 22708 4126
rect 22652 4062 22654 4114
rect 22706 4062 22708 4114
rect 22652 4060 22708 4062
rect 22484 4004 22708 4060
rect 22484 3836 22540 4004
rect 22820 3836 22876 4452
rect 22484 3770 22540 3780
rect 22596 3780 22876 3836
rect 22260 3668 22428 3724
rect 21700 3546 21756 3556
rect 21980 3612 22036 3622
rect 21980 3518 22036 3556
rect 21308 3500 21364 3510
rect 21308 3406 21364 3444
rect 22204 3500 22260 3510
rect 22204 3406 22260 3444
rect 20916 3388 20972 3398
rect 20916 3294 20972 3332
rect 21196 3388 21252 3398
rect 21644 3387 21700 3398
rect 21196 3294 21252 3332
rect 21588 3386 21700 3387
rect 21588 3334 21646 3386
rect 21698 3334 21700 3386
rect 21588 3322 21700 3334
rect 21476 3276 21532 3286
rect 20132 3098 20188 3108
rect 20580 3164 20636 3174
rect 20132 2940 20188 2950
rect 20132 2938 20524 2940
rect 20132 2886 20134 2938
rect 20186 2886 20524 2938
rect 20132 2884 20524 2886
rect 20132 2874 20188 2884
rect 20020 2828 20076 2838
rect 20020 2726 20076 2772
rect 19404 2550 19406 2602
rect 19458 2550 19460 2602
rect 19068 2492 19124 2502
rect 18172 2102 18174 2154
rect 18226 2102 18228 2154
rect 18172 2090 18228 2102
rect 18508 2156 18564 2166
rect 18508 2062 18564 2100
rect 18620 2154 18732 2166
rect 18620 2102 18622 2154
rect 18674 2102 18732 2154
rect 18620 2100 18732 2102
rect 18844 2380 18900 2390
rect 18620 2090 18676 2100
rect 17724 1642 17780 1652
rect 18844 1930 18900 2324
rect 19068 2156 19124 2436
rect 19404 2380 19460 2550
rect 19404 2314 19460 2324
rect 19684 2714 19740 2726
rect 19684 2662 19686 2714
rect 19738 2662 19740 2714
rect 19292 2156 19348 2166
rect 19516 2156 19572 2166
rect 18844 1878 18846 1930
rect 18898 1878 18900 1930
rect 18844 1708 18900 1878
rect 18844 1642 18900 1652
rect 19012 2154 19572 2156
rect 19012 2102 19070 2154
rect 19122 2102 19294 2154
rect 19346 2102 19518 2154
rect 19570 2102 19572 2154
rect 19012 2100 19572 2102
rect 19012 2090 19124 2100
rect 19292 2090 19348 2100
rect 19516 2090 19572 2100
rect 19684 2156 19740 2662
rect 20020 2714 20132 2726
rect 20020 2662 20078 2714
rect 20130 2662 20132 2714
rect 20020 2660 20132 2662
rect 20076 2650 20132 2660
rect 20300 2548 20356 2558
rect 20300 2546 20412 2548
rect 19684 2090 19740 2100
rect 19964 2492 20020 2502
rect 20300 2494 20302 2546
rect 20354 2494 20412 2546
rect 20300 2482 20412 2494
rect 19964 2156 20020 2436
rect 20188 2156 20244 2166
rect 19964 2154 20244 2156
rect 19964 2102 19966 2154
rect 20018 2102 20190 2154
rect 20242 2102 20244 2154
rect 19964 2100 20244 2102
rect 19964 2090 20020 2100
rect 13368 1596 13632 1606
rect 13424 1540 13472 1596
rect 13528 1540 13576 1596
rect 13368 1530 13632 1540
rect 13132 1206 13134 1258
rect 13186 1206 13188 1258
rect 13132 1194 13188 1206
rect 17724 1260 17780 1270
rect 17724 1166 17780 1204
rect 18844 1260 18900 1270
rect 19012 1260 19068 2090
rect 19740 1930 19796 1942
rect 19740 1878 19742 1930
rect 19794 1878 19796 1930
rect 18844 1258 19068 1260
rect 18844 1206 18846 1258
rect 18898 1206 19068 1258
rect 18844 1204 19068 1206
rect 19180 1708 19236 1718
rect 19180 1258 19236 1652
rect 19572 1708 19628 1718
rect 19572 1484 19628 1652
rect 19740 1708 19796 1878
rect 19740 1642 19796 1652
rect 20188 1932 20244 2100
rect 20188 1484 20244 1876
rect 20356 1820 20412 2482
rect 20468 2054 20524 2884
rect 20580 2782 20636 3108
rect 20580 2730 20582 2782
rect 20634 2730 20636 2782
rect 20580 2380 20636 2730
rect 20580 2314 20636 2324
rect 20692 2828 20748 2838
rect 20468 2042 20580 2054
rect 20468 1990 20526 2042
rect 20578 1990 20580 2042
rect 20468 1988 20580 1990
rect 20524 1978 20580 1988
rect 20692 2002 20748 2772
rect 21084 2770 21140 2782
rect 21084 2718 21086 2770
rect 21138 2718 21140 2770
rect 21084 2716 21140 2718
rect 21028 2660 21140 2716
rect 20692 1950 20694 2002
rect 20746 1950 20748 2002
rect 20692 1938 20748 1950
rect 20804 2268 20860 2278
rect 20804 1820 20860 2212
rect 20916 2156 20972 2166
rect 21028 2156 21084 2660
rect 20916 2154 21084 2156
rect 20916 2102 20918 2154
rect 20970 2102 21084 2154
rect 20916 2100 21084 2102
rect 20916 2090 20972 2100
rect 21308 2044 21364 2054
rect 21308 1950 21364 1988
rect 21084 1820 21140 1830
rect 20804 1764 21028 1820
rect 20356 1754 20412 1764
rect 19572 1428 19908 1484
rect 19180 1206 19182 1258
rect 19234 1206 19236 1258
rect 18844 1194 18900 1204
rect 19180 1194 19236 1206
rect 19628 1260 19684 1270
rect 19628 1166 19684 1204
rect 19852 1258 19908 1428
rect 20188 1418 20244 1428
rect 20300 1596 20356 1606
rect 19852 1206 19854 1258
rect 19906 1206 19908 1258
rect 19852 1194 19908 1206
rect 20076 1372 20132 1382
rect 20076 1258 20132 1316
rect 20076 1206 20078 1258
rect 20130 1206 20132 1258
rect 20076 1194 20132 1206
rect 20300 1258 20356 1540
rect 20300 1206 20302 1258
rect 20354 1206 20356 1258
rect 7868 1146 8204 1148
rect 7868 1094 7870 1146
rect 7922 1094 8204 1146
rect 7868 1092 8204 1094
rect 19404 1148 19460 1158
rect 7868 1082 7924 1092
rect 19404 1054 19460 1092
rect 17500 1034 17556 1046
rect 17500 982 17502 1034
rect 17554 982 17556 1034
rect 9092 812 9356 822
rect 9148 756 9196 812
rect 9252 756 9300 812
rect 9092 746 9356 756
rect 17500 700 17556 982
rect 17948 1036 18004 1046
rect 17948 942 18004 980
rect 18172 1034 18228 1046
rect 18172 982 18174 1034
rect 18226 982 18228 1034
rect 18172 924 18228 982
rect 18172 858 18228 868
rect 18396 1034 18452 1046
rect 18396 982 18398 1034
rect 18450 982 18452 1034
rect 17644 812 17908 822
rect 17700 756 17748 812
rect 17804 756 17852 812
rect 17644 746 17908 756
rect 17500 634 17556 644
rect 18396 588 18452 982
rect 18396 522 18452 532
rect 20300 586 20356 1206
rect 20412 1484 20468 1494
rect 20412 1258 20468 1428
rect 20412 1206 20414 1258
rect 20466 1206 20468 1258
rect 20412 1194 20468 1206
rect 20748 1372 20804 1382
rect 20748 1258 20804 1316
rect 20748 1206 20750 1258
rect 20802 1206 20804 1258
rect 20748 1194 20804 1206
rect 20972 1258 21028 1764
rect 21084 1726 21140 1764
rect 21476 1596 21532 3220
rect 21588 2828 21644 3322
rect 21920 3164 22184 3174
rect 21976 3108 22024 3164
rect 22080 3108 22128 3164
rect 21920 3098 22184 3108
rect 21588 2762 21644 2772
rect 22260 2828 22316 2838
rect 22260 2716 22316 2772
rect 22204 2660 22316 2716
rect 21868 2604 21924 2614
rect 20972 1206 20974 1258
rect 21026 1206 21028 1258
rect 20300 534 20302 586
rect 20354 534 20356 586
rect 20300 522 20356 534
rect 20972 474 21028 1206
rect 21196 1540 21532 1596
rect 21644 2380 21700 2390
rect 21644 2154 21700 2324
rect 21644 2102 21646 2154
rect 21698 2102 21700 2154
rect 21196 1258 21252 1540
rect 21644 1484 21700 2102
rect 21868 1932 21924 2548
rect 22204 2210 22260 2660
rect 22372 2492 22428 3668
rect 22596 3612 22652 3780
rect 22932 3722 22988 4900
rect 23156 4620 23212 6582
rect 23380 6638 23382 6690
rect 23434 6638 23436 6690
rect 23380 6076 23436 6638
rect 23492 6636 23548 7410
rect 23492 6570 23548 6580
rect 23940 6883 23996 6895
rect 23940 6831 23942 6883
rect 23994 6831 23996 6883
rect 23268 6020 23436 6076
rect 23268 4954 23324 6020
rect 23828 5964 23884 5974
rect 23604 5962 23884 5964
rect 23380 5906 23436 5918
rect 23380 5854 23382 5906
rect 23434 5854 23436 5906
rect 23380 5852 23436 5854
rect 23380 5786 23436 5796
rect 23604 5910 23830 5962
rect 23882 5910 23884 5962
rect 23604 5908 23884 5910
rect 23268 4902 23270 4954
rect 23322 4902 23324 4954
rect 23268 4890 23324 4902
rect 23156 4554 23212 4564
rect 23604 4508 23660 5908
rect 23828 5898 23884 5908
rect 23716 5678 23772 5690
rect 23716 5626 23718 5678
rect 23770 5626 23772 5678
rect 23716 5151 23772 5626
rect 23828 5292 23884 5302
rect 23828 5198 23884 5236
rect 23716 5099 23718 5151
rect 23770 5099 23772 5151
rect 23716 5087 23772 5099
rect 23940 5068 23996 6831
rect 24332 6636 24388 6712
rect 24836 6680 24892 7588
rect 24276 6580 24332 6636
rect 24276 6570 24388 6580
rect 24556 6636 24612 6646
rect 24276 5180 24332 6570
rect 24388 6412 24444 6422
rect 24388 5740 24444 6356
rect 24556 6130 24612 6580
rect 24556 6078 24558 6130
rect 24610 6078 24612 6130
rect 24556 6066 24612 6078
rect 24780 6624 24892 6680
rect 25060 8092 25116 8102
rect 24780 6130 24836 6624
rect 24948 6522 25004 6534
rect 24948 6470 24950 6522
rect 25002 6470 25004 6522
rect 24948 6412 25004 6470
rect 24780 6078 24782 6130
rect 24834 6078 24836 6130
rect 24780 6066 24836 6078
rect 24892 6356 25004 6412
rect 24892 5964 24948 6356
rect 25060 6300 25116 8036
rect 25004 6244 25116 6300
rect 25172 7420 25228 8148
rect 25284 8194 25286 8246
rect 25338 8194 25340 8246
rect 25284 7980 25340 8194
rect 25284 7914 25340 7924
rect 25004 6130 25060 6244
rect 25004 6078 25006 6130
rect 25058 6078 25060 6130
rect 25004 6066 25060 6078
rect 24836 5908 24948 5964
rect 25172 5927 25228 7364
rect 25396 6524 25452 8430
rect 25508 8092 25564 10052
rect 25732 10598 25788 10610
rect 25732 10556 25734 10598
rect 25786 10556 25788 10598
rect 25620 8246 25676 8258
rect 25620 8204 25622 8246
rect 25674 8204 25676 8246
rect 25620 8138 25676 8148
rect 25508 8026 25564 8036
rect 25732 7756 25788 10500
rect 25620 7700 25788 7756
rect 25396 6458 25452 6468
rect 25508 7196 25564 7206
rect 25620 7196 25676 7700
rect 25564 7140 25676 7196
rect 25732 7532 25788 7542
rect 25732 7434 25734 7476
rect 25786 7434 25788 7476
rect 24612 5740 24668 5750
rect 24388 5738 24668 5740
rect 24388 5686 24614 5738
rect 24666 5686 24668 5738
rect 24388 5684 24668 5686
rect 24612 5674 24668 5684
rect 24276 5114 24332 5124
rect 23884 5012 23996 5068
rect 23884 5010 23940 5012
rect 23884 4958 23886 5010
rect 23938 4958 23940 5010
rect 23884 4946 23940 4958
rect 24108 4956 24164 4966
rect 24108 4862 24164 4900
rect 24332 4956 24388 4966
rect 24332 4862 24388 4900
rect 24500 4620 24556 4630
rect 23604 4452 23772 4508
rect 23044 4396 23100 4406
rect 23044 4282 23100 4340
rect 23044 4230 23046 4282
rect 23098 4230 23100 4282
rect 23044 4218 23100 4230
rect 23604 4326 23660 4338
rect 23604 4274 23606 4326
rect 23658 4274 23660 4326
rect 23212 4172 23268 4182
rect 23212 4078 23268 4116
rect 23492 3747 23548 3759
rect 22932 3670 22934 3722
rect 22986 3670 22988 3722
rect 22932 3658 22988 3670
rect 23380 3724 23436 3734
rect 22596 3520 22598 3556
rect 22650 3520 22652 3556
rect 22596 3480 22652 3520
rect 22372 2436 22484 2492
rect 22204 2158 22206 2210
rect 22258 2158 22260 2210
rect 22204 2146 22260 2158
rect 22428 2268 22484 2436
rect 23380 2268 23436 3668
rect 23492 3695 23494 3747
rect 23546 3695 23548 3747
rect 23492 2828 23548 3695
rect 23492 2762 23548 2772
rect 23604 2716 23660 4274
rect 23604 2650 23660 2660
rect 23716 3500 23772 4452
rect 24332 4396 24388 4406
rect 24332 4302 24388 4340
rect 24052 4172 24108 4182
rect 24052 3554 24108 4116
rect 24052 3502 24054 3554
rect 24106 3502 24108 3554
rect 24052 3490 24108 3502
rect 24276 3836 24332 3846
rect 24276 3498 24332 3780
rect 23716 3276 23772 3444
rect 24276 3446 24278 3498
rect 24330 3446 24332 3498
rect 24276 3434 24332 3446
rect 24500 3387 24556 4564
rect 24836 4284 24892 5908
rect 25172 5875 25174 5927
rect 25226 5875 25228 5927
rect 25172 5134 25228 5875
rect 25508 5750 25564 7140
rect 25620 6860 25676 6870
rect 25732 6860 25788 7434
rect 25620 6858 25788 6860
rect 25620 6806 25622 6858
rect 25674 6806 25788 6858
rect 25620 6804 25788 6806
rect 25620 6794 25676 6804
rect 25844 6748 25900 10724
rect 26012 10668 26068 10678
rect 26012 10574 26068 10612
rect 26292 10666 26348 10678
rect 26292 10614 26294 10666
rect 26346 10614 26348 10666
rect 26068 10444 26124 10454
rect 25956 10019 26012 10031
rect 25956 9967 25958 10019
rect 26010 9967 26012 10019
rect 25956 9772 26012 9967
rect 25956 9706 26012 9716
rect 25956 8988 26012 8998
rect 25956 8894 26012 8932
rect 26068 8876 26124 10388
rect 26292 10444 26348 10614
rect 26964 10554 27020 11172
rect 26964 10502 26966 10554
rect 27018 10502 27020 10554
rect 26964 10490 27020 10502
rect 26292 10378 26348 10388
rect 26196 10220 26460 10230
rect 26252 10164 26300 10220
rect 26356 10164 26404 10220
rect 26196 10154 26460 10164
rect 26404 9996 26460 10006
rect 26404 9855 26460 9940
rect 26516 9996 26572 10006
rect 26628 9996 26684 10006
rect 26516 9994 26628 9996
rect 26516 9942 26518 9994
rect 26570 9942 26628 9994
rect 26516 9940 26628 9942
rect 26516 9930 26572 9940
rect 26628 9930 26684 9940
rect 26404 9803 26406 9855
rect 26458 9803 26460 9855
rect 26404 9791 26460 9803
rect 27020 9884 27076 9894
rect 27020 9826 27076 9828
rect 26572 9772 26628 9782
rect 27020 9774 27022 9826
rect 27074 9774 27076 9826
rect 27020 9762 27076 9774
rect 26572 9678 26628 9716
rect 26796 9602 26852 9614
rect 26796 9550 26798 9602
rect 26850 9550 26852 9602
rect 26796 9436 26852 9550
rect 26740 9380 26852 9436
rect 26740 9324 26796 9380
rect 26740 9258 26796 9268
rect 26628 9212 26684 9222
rect 26628 9118 26684 9156
rect 26852 9212 26908 9222
rect 27188 9212 27244 11284
rect 27636 11340 27692 12004
rect 28588 12010 28644 12022
rect 28588 11958 28590 12010
rect 28642 11958 28644 12010
rect 28588 11452 28644 11958
rect 29428 12010 29484 12022
rect 29428 11958 29430 12010
rect 29482 11958 29484 12010
rect 29428 11564 29484 11958
rect 30268 12012 30324 12022
rect 29932 11788 29988 11798
rect 29484 11508 29596 11564
rect 29428 11498 29484 11508
rect 28588 11386 28644 11396
rect 28980 11478 29036 11490
rect 28980 11426 28982 11478
rect 29034 11426 29036 11478
rect 27636 11274 27692 11284
rect 28980 11340 29036 11426
rect 28980 11274 29036 11284
rect 29428 11340 29484 11350
rect 29316 10598 29372 10610
rect 29316 10546 29318 10598
rect 29370 10546 29372 10598
rect 28196 10108 28252 10118
rect 27916 9884 27972 9894
rect 27916 9882 28140 9884
rect 27692 9826 27748 9838
rect 27468 9772 27524 9782
rect 26852 9210 27244 9212
rect 26852 9158 26854 9210
rect 26906 9158 27244 9210
rect 26852 9156 27244 9158
rect 27412 9770 27524 9772
rect 27412 9718 27470 9770
rect 27522 9718 27524 9770
rect 27412 9706 27524 9718
rect 27692 9774 27694 9826
rect 27746 9774 27748 9826
rect 27916 9830 27918 9882
rect 27970 9830 28140 9882
rect 27916 9828 28140 9830
rect 27916 9818 27972 9828
rect 26852 9146 26908 9156
rect 26068 8810 26124 8820
rect 26516 8988 26572 8998
rect 26196 8652 26460 8662
rect 26252 8596 26300 8652
rect 26356 8596 26404 8652
rect 26196 8586 26460 8596
rect 26404 8428 26460 8466
rect 26404 8362 26460 8372
rect 26012 8092 26068 8102
rect 25452 5738 25564 5750
rect 25452 5686 25454 5738
rect 25506 5686 25564 5738
rect 25452 5674 25564 5686
rect 25508 5628 25564 5674
rect 25732 6692 25900 6748
rect 25956 8090 26068 8092
rect 25956 8038 26014 8090
rect 26066 8038 26068 8090
rect 25956 8026 26068 8038
rect 26236 8092 26292 8102
rect 25508 5572 25676 5628
rect 25172 5082 25174 5134
rect 25226 5082 25228 5134
rect 25172 5070 25228 5082
rect 25396 5516 25452 5526
rect 25396 5134 25452 5460
rect 25508 5404 25564 5414
rect 25508 5320 25510 5348
rect 25562 5320 25564 5348
rect 25508 5308 25564 5320
rect 25620 5180 25676 5572
rect 25396 5082 25398 5134
rect 25450 5082 25452 5134
rect 25396 5068 25452 5082
rect 24836 3612 24892 4228
rect 25284 5012 25396 5068
rect 24948 4060 25004 4070
rect 24948 3734 25004 4004
rect 24948 3722 25060 3734
rect 24948 3670 25006 3722
rect 25058 3670 25060 3722
rect 24948 3668 25060 3670
rect 25004 3658 25060 3668
rect 24836 3546 24892 3556
rect 23492 2604 23548 2614
rect 23492 2380 23548 2548
rect 23716 2604 23772 3220
rect 24388 3331 24556 3387
rect 24164 2938 24220 2950
rect 24164 2886 24166 2938
rect 24218 2886 24220 2938
rect 23716 2538 23772 2548
rect 23940 2716 23996 2726
rect 23492 2314 23548 2324
rect 23604 2492 23660 2502
rect 22428 2212 23156 2268
rect 22428 2210 22484 2212
rect 22428 2158 22430 2210
rect 22482 2158 22484 2210
rect 22428 2146 22484 2158
rect 23100 2154 23156 2212
rect 23380 2202 23436 2212
rect 23604 2166 23660 2436
rect 23100 2102 23102 2154
rect 23154 2102 23156 2154
rect 23100 2090 23156 2102
rect 23268 2156 23324 2166
rect 23268 2064 23324 2100
rect 23548 2154 23660 2166
rect 23548 2102 23550 2154
rect 23602 2102 23660 2154
rect 23548 2100 23660 2102
rect 23772 2268 23828 2278
rect 23772 2154 23828 2212
rect 23772 2102 23774 2154
rect 23826 2102 23828 2154
rect 23548 2090 23604 2100
rect 23772 2090 23828 2102
rect 21812 1876 21868 1932
rect 21812 1838 21924 1876
rect 22372 2044 22428 2054
rect 21812 1820 21868 1838
rect 21644 1418 21700 1428
rect 21756 1764 21868 1820
rect 22372 1818 22428 1988
rect 22708 2044 22764 2054
rect 22372 1766 22374 1818
rect 22426 1766 22428 1818
rect 21196 1206 21198 1258
rect 21250 1206 21252 1258
rect 21196 1194 21252 1206
rect 21420 1372 21476 1382
rect 21420 1258 21476 1316
rect 21420 1206 21422 1258
rect 21474 1206 21476 1258
rect 21420 1194 21476 1206
rect 21756 1258 21812 1764
rect 22372 1754 22428 1766
rect 22540 1820 22596 1830
rect 22260 1708 22316 1718
rect 21920 1596 22184 1606
rect 21976 1540 22024 1596
rect 22080 1540 22128 1596
rect 21920 1530 22184 1540
rect 22260 1372 22316 1652
rect 21756 1206 21758 1258
rect 21810 1206 21812 1258
rect 21756 1194 21812 1206
rect 22148 1316 22316 1372
rect 22148 1158 22204 1316
rect 22092 1148 22204 1158
rect 22148 1092 22204 1148
rect 22092 1054 22148 1092
rect 21644 1034 21700 1046
rect 21644 982 21646 1034
rect 21698 982 21700 1034
rect 21644 586 21700 982
rect 21644 534 21646 586
rect 21698 534 21700 586
rect 21644 522 21700 534
rect 22316 1034 22372 1046
rect 22316 982 22318 1034
rect 22370 982 22372 1034
rect 20972 422 20974 474
rect 21026 422 21028 474
rect 20972 410 21028 422
rect 22316 474 22372 982
rect 22540 1034 22596 1764
rect 22708 1270 22764 1988
rect 22820 2042 22876 2054
rect 22820 1990 22822 2042
rect 22874 1990 22876 2042
rect 23268 2012 23270 2064
rect 23322 2012 23324 2064
rect 23268 2000 23324 2012
rect 23940 2064 23996 2660
rect 24164 2156 24220 2886
rect 24388 2838 24444 3331
rect 24332 2826 24444 2838
rect 24332 2774 24334 2826
rect 24386 2774 24444 2826
rect 24332 2772 24444 2774
rect 24332 2762 24388 2772
rect 24164 2090 24220 2100
rect 24332 2604 24388 2614
rect 24332 2154 24388 2548
rect 24556 2602 24612 2614
rect 24556 2550 24558 2602
rect 24610 2550 24612 2602
rect 24556 2380 24612 2550
rect 24556 2314 24612 2324
rect 24892 2602 24948 2614
rect 25116 2604 25172 2614
rect 24892 2550 24894 2602
rect 24946 2550 24948 2602
rect 24892 2268 24948 2550
rect 24892 2202 24948 2212
rect 25060 2548 25116 2604
rect 25060 2472 25172 2548
rect 24332 2102 24334 2154
rect 24386 2102 24388 2154
rect 24332 2090 24388 2102
rect 23940 2044 24052 2064
rect 22820 1932 22876 1990
rect 23940 1988 23996 2044
rect 22820 1866 22876 1876
rect 23268 1932 23324 1942
rect 23268 1838 23324 1876
rect 23940 1912 24052 1988
rect 24948 2044 25004 2054
rect 24948 1946 24950 1988
rect 25002 1946 25004 1988
rect 22652 1258 22764 1270
rect 22652 1206 22654 1258
rect 22706 1206 22764 1258
rect 22652 1194 22764 1206
rect 22988 1484 23044 1494
rect 22988 1258 23044 1428
rect 22988 1206 22990 1258
rect 23042 1206 23044 1258
rect 22988 1194 23044 1206
rect 23436 1484 23492 1494
rect 23436 1258 23492 1428
rect 23940 1484 23996 1912
rect 23940 1418 23996 1428
rect 24948 1708 25004 1946
rect 25060 1820 25116 2472
rect 25060 1754 25116 1764
rect 23436 1206 23438 1258
rect 23490 1206 23492 1258
rect 23436 1194 23492 1206
rect 23660 1260 23716 1270
rect 22540 982 22542 1034
rect 22594 982 22596 1034
rect 22540 586 22596 982
rect 22708 1036 22764 1194
rect 23660 1166 23716 1204
rect 24108 1260 24164 1270
rect 24108 1166 24164 1204
rect 24780 1260 24836 1270
rect 24780 1166 24836 1204
rect 24948 1046 25004 1652
rect 25284 1270 25340 5012
rect 25396 5002 25452 5012
rect 25508 5124 25676 5180
rect 25732 5134 25788 6692
rect 25396 3724 25452 3734
rect 25396 3630 25452 3668
rect 25508 3500 25564 5124
rect 25732 5082 25734 5134
rect 25786 5082 25788 5134
rect 25732 5070 25788 5082
rect 25844 5964 25900 5974
rect 25844 5862 25846 5908
rect 25898 5862 25900 5908
rect 25396 3444 25564 3500
rect 25620 4060 25676 4070
rect 25620 3722 25676 4004
rect 25620 3670 25622 3722
rect 25674 3670 25676 3722
rect 25396 2268 25452 3444
rect 25620 3388 25676 3670
rect 25620 3322 25676 3332
rect 25564 2828 25620 2838
rect 25564 2734 25620 2772
rect 25676 2716 25732 2726
rect 25676 2622 25732 2660
rect 25844 2604 25900 5862
rect 25956 5404 26012 8026
rect 26236 7998 26292 8036
rect 26516 7532 26572 8932
rect 27188 8876 27244 8886
rect 26796 8316 26852 8326
rect 26628 8246 26684 8258
rect 26628 8204 26630 8246
rect 26682 8204 26684 8246
rect 26796 8222 26852 8260
rect 26628 7980 26684 8148
rect 27020 8204 27076 8214
rect 27020 8092 27076 8148
rect 26628 7914 26684 7924
rect 26852 8036 27076 8092
rect 26516 7466 26572 7476
rect 26740 7308 26796 7318
rect 26740 7214 26796 7252
rect 26196 7084 26460 7094
rect 26252 7028 26300 7084
rect 26356 7028 26404 7084
rect 26196 7018 26460 7028
rect 26852 6860 26908 8036
rect 27188 7980 27244 8820
rect 26852 6794 26908 6804
rect 26964 7924 27244 7980
rect 27300 8246 27356 8258
rect 27300 8194 27302 8246
rect 27354 8194 27356 8246
rect 26404 5894 26460 5906
rect 26404 5852 26406 5894
rect 26458 5852 26460 5894
rect 26404 5786 26460 5796
rect 25956 5338 26012 5348
rect 26068 5628 26124 5638
rect 26068 5178 26124 5572
rect 26196 5516 26460 5526
rect 26252 5460 26300 5516
rect 26356 5460 26404 5516
rect 26196 5450 26460 5460
rect 26964 5290 27020 7924
rect 27300 7644 27356 8194
rect 27076 7588 27356 7644
rect 27412 8204 27468 9706
rect 27692 9324 27748 9774
rect 27636 9268 27748 9324
rect 27860 9660 27916 9670
rect 27524 8876 27580 8886
rect 27524 8782 27580 8820
rect 27076 7462 27132 7588
rect 27076 7410 27078 7462
rect 27130 7410 27132 7462
rect 27076 7196 27132 7410
rect 27076 7130 27132 7140
rect 27412 6748 27468 8148
rect 27636 7308 27692 9268
rect 27860 9212 27916 9604
rect 27748 9156 27916 9212
rect 27972 9658 28028 9670
rect 27972 9606 27974 9658
rect 28026 9606 28028 9658
rect 27748 8540 27804 9156
rect 27748 8092 27804 8484
rect 27860 8428 27916 8438
rect 27860 8270 27916 8372
rect 27860 8218 27862 8270
rect 27914 8218 27916 8270
rect 27972 8316 28028 9606
rect 27972 8250 28028 8260
rect 27860 8206 27916 8218
rect 27748 8036 27860 8092
rect 27804 7586 27860 8036
rect 27804 7534 27806 7586
rect 27858 7534 27860 7586
rect 27804 7522 27860 7534
rect 27636 7242 27692 7252
rect 28084 6860 28140 9828
rect 28196 9882 28252 10052
rect 28532 10108 28588 10118
rect 28532 9994 28588 10052
rect 28532 9942 28534 9994
rect 28586 9942 28588 9994
rect 28532 9930 28588 9942
rect 28196 9830 28198 9882
rect 28250 9830 28252 9882
rect 28196 9818 28252 9830
rect 29316 9212 29372 10546
rect 29428 9826 29484 11284
rect 29428 9774 29430 9826
rect 29482 9774 29484 9826
rect 29428 9772 29484 9774
rect 29428 9706 29484 9716
rect 29316 9146 29372 9156
rect 29540 9100 29596 11508
rect 29932 11562 29988 11732
rect 29932 11510 29934 11562
rect 29986 11510 29988 11562
rect 29932 11498 29988 11510
rect 30268 11562 30324 11956
rect 30660 11900 30716 12114
rect 30660 11834 30716 11844
rect 31332 12166 31388 12178
rect 31332 12114 31334 12166
rect 31386 12114 31388 12166
rect 31332 11788 31388 12114
rect 31332 11722 31388 11732
rect 30268 11510 30270 11562
rect 30322 11510 30324 11562
rect 30268 11498 30324 11510
rect 30828 11394 31052 11408
rect 30044 11340 30100 11350
rect 30828 11342 30830 11394
rect 30882 11352 31052 11394
rect 30882 11342 30884 11352
rect 30828 11330 30884 11342
rect 30044 11246 30100 11284
rect 30472 11004 30736 11014
rect 30528 10948 30576 11004
rect 30632 10948 30680 11004
rect 30472 10938 30736 10948
rect 29764 10780 29820 10790
rect 29764 10598 29820 10724
rect 29764 10556 29766 10598
rect 29818 10556 29820 10598
rect 29764 10490 29820 10500
rect 30996 10598 31052 11352
rect 30996 10556 30998 10598
rect 31050 10556 31052 10598
rect 30996 10490 31052 10500
rect 31220 11382 31276 11394
rect 31220 11330 31222 11382
rect 31274 11330 31276 11382
rect 30156 10444 30212 10454
rect 29876 10442 30212 10444
rect 29876 10390 30158 10442
rect 30210 10390 30212 10442
rect 29876 10388 30212 10390
rect 29876 9884 29932 10388
rect 30156 10378 30212 10388
rect 30268 10442 30324 10454
rect 30268 10390 30270 10442
rect 30322 10390 30324 10442
rect 30268 10108 30324 10390
rect 29876 9818 29932 9828
rect 29988 10052 30324 10108
rect 31220 10108 31276 11330
rect 31388 10610 31444 10622
rect 31388 10558 31390 10610
rect 31442 10558 31444 10610
rect 31388 10556 31444 10558
rect 29540 9034 29596 9044
rect 29876 9030 29932 9042
rect 29876 8978 29878 9030
rect 29930 8978 29932 9030
rect 29876 8428 29932 8978
rect 29876 8362 29932 8372
rect 29316 8204 29372 8214
rect 28084 6794 28140 6804
rect 28756 7308 28812 7318
rect 27412 6682 27468 6692
rect 27972 6678 28028 6690
rect 27972 6626 27974 6678
rect 28026 6626 28028 6678
rect 27972 6076 28028 6626
rect 27972 6010 28028 6020
rect 28420 6678 28476 6690
rect 28420 6626 28422 6678
rect 28474 6626 28476 6678
rect 28420 5964 28476 6626
rect 28420 5898 28476 5908
rect 28644 6300 28700 6310
rect 28644 5918 28700 6244
rect 28644 5866 28646 5918
rect 28698 5866 28700 5918
rect 28644 5854 28700 5866
rect 26964 5238 26966 5290
rect 27018 5238 27020 5290
rect 26964 5226 27020 5238
rect 27972 5292 28028 5302
rect 26068 5126 26070 5178
rect 26122 5126 26124 5178
rect 25956 4396 26012 4406
rect 25956 3722 26012 4340
rect 26068 4172 26124 5126
rect 26404 5180 26460 5190
rect 26404 4954 26460 5124
rect 27860 5178 27916 5190
rect 27860 5126 27862 5178
rect 27914 5126 27916 5178
rect 26628 5068 26684 5078
rect 26628 4974 26684 5012
rect 26404 4902 26406 4954
rect 26458 4902 26460 4954
rect 26404 4844 26460 4902
rect 27356 4956 27412 4966
rect 27356 4862 27412 4900
rect 27468 4954 27524 4966
rect 27468 4902 27470 4954
rect 27522 4902 27524 4954
rect 26404 4778 26460 4788
rect 26516 4508 26572 4518
rect 26516 4414 26572 4452
rect 27468 4508 27524 4902
rect 27860 4732 27916 5126
rect 27972 4956 28028 5236
rect 28140 5180 28196 5190
rect 28140 5086 28196 5124
rect 28364 5122 28420 5134
rect 28364 5070 28366 5122
rect 28418 5070 28420 5122
rect 28084 4956 28140 4966
rect 27972 4954 28140 4956
rect 27972 4902 28086 4954
rect 28138 4902 28140 4954
rect 27972 4900 28140 4902
rect 28084 4890 28140 4900
rect 27860 4676 28084 4732
rect 27468 4442 27524 4452
rect 27916 4508 27972 4518
rect 27916 4414 27972 4452
rect 27524 4282 27580 4294
rect 27524 4230 27526 4282
rect 27578 4230 27580 4282
rect 26684 4172 26740 4182
rect 26068 4170 26740 4172
rect 26068 4118 26686 4170
rect 26738 4118 26740 4170
rect 27132 4170 27188 4182
rect 26068 4116 26740 4118
rect 26628 4106 26740 4116
rect 27020 4114 27076 4126
rect 26196 3948 26460 3958
rect 26252 3892 26300 3948
rect 26356 3892 26404 3948
rect 26196 3882 26460 3892
rect 25956 3670 25958 3722
rect 26010 3670 26012 3722
rect 25956 3658 26012 3670
rect 26404 3612 26460 3622
rect 26124 3388 26180 3398
rect 26124 2994 26180 3332
rect 26404 3388 26460 3556
rect 26404 3322 26460 3332
rect 26516 3500 26572 3510
rect 26516 3164 26572 3444
rect 26628 3276 26684 4106
rect 26852 4060 26908 4070
rect 27020 4062 27022 4114
rect 27074 4062 27076 4114
rect 27020 4060 27076 4062
rect 26908 4004 27076 4060
rect 27132 4118 27134 4170
rect 27186 4118 27188 4170
rect 26740 3500 26796 3510
rect 26740 3406 26796 3444
rect 26628 3220 26796 3276
rect 26516 3098 26572 3108
rect 26124 2942 26126 2994
rect 26178 2942 26180 2994
rect 26628 3052 26684 3062
rect 26124 2930 26180 2942
rect 26348 2940 26404 2950
rect 26348 2846 26404 2884
rect 26628 2773 26684 2996
rect 26628 2721 26630 2773
rect 26682 2721 26684 2773
rect 26628 2709 26684 2721
rect 25844 2538 25900 2548
rect 26404 2604 26460 2642
rect 26404 2538 26460 2548
rect 26740 2492 26796 3220
rect 26852 3052 26908 4004
rect 27132 3948 27188 4118
rect 27020 3892 27188 3948
rect 27244 4114 27300 4126
rect 27244 4062 27246 4114
rect 27298 4062 27300 4114
rect 27020 3610 27076 3892
rect 27020 3558 27022 3610
rect 27074 3558 27076 3610
rect 27020 3546 27076 3558
rect 27244 3612 27300 4062
rect 27244 3518 27300 3556
rect 27412 3722 27468 3734
rect 27412 3670 27414 3722
rect 27466 3670 27468 3722
rect 26852 2986 26908 2996
rect 27412 3052 27468 3670
rect 27412 2986 27468 2996
rect 27524 3510 27580 4230
rect 28028 4172 28084 4676
rect 28364 4620 28420 5070
rect 28756 5122 28812 7252
rect 28756 5070 28758 5122
rect 28810 5070 28812 5122
rect 28756 5058 28812 5070
rect 28868 6522 28924 6534
rect 28868 6470 28870 6522
rect 28922 6470 28924 6522
rect 28868 5740 28924 6470
rect 28028 4078 28084 4116
rect 28308 4564 28420 4620
rect 28532 4620 28588 4630
rect 28308 3836 28364 4564
rect 28420 4396 28476 4406
rect 28420 4282 28476 4340
rect 28420 4230 28422 4282
rect 28474 4230 28476 4282
rect 28420 4218 28476 4230
rect 28308 3780 28476 3836
rect 27748 3724 27804 3734
rect 27748 3612 27804 3668
rect 28196 3724 28252 3734
rect 28252 3668 28308 3724
rect 28196 3666 28308 3668
rect 28196 3658 28254 3666
rect 27692 3556 27804 3612
rect 28252 3614 28254 3658
rect 28306 3614 28308 3666
rect 28252 3602 28308 3614
rect 27524 3498 27636 3510
rect 27524 3446 27582 3498
rect 27634 3446 27636 3498
rect 27524 3434 27636 3446
rect 27524 2940 27580 3434
rect 27692 3164 27748 3556
rect 27804 3387 27860 3398
rect 28420 3387 28476 3780
rect 28532 3566 28588 4564
rect 28868 3836 28924 5684
rect 29316 5290 29372 8148
rect 29988 7642 30044 10052
rect 31220 10042 31276 10052
rect 31332 10500 31444 10556
rect 32340 10556 32396 10566
rect 29988 7590 29990 7642
rect 30042 7590 30044 7642
rect 29988 7578 30044 7590
rect 30100 9772 30156 9782
rect 30100 8876 30156 9716
rect 30472 9436 30736 9446
rect 30528 9380 30576 9436
rect 30632 9380 30680 9436
rect 30472 9370 30736 9380
rect 30884 9212 30940 9222
rect 31332 9212 31388 10500
rect 30884 9210 31388 9212
rect 30884 9158 30886 9210
rect 30938 9158 31388 9210
rect 30884 9156 31388 9158
rect 31556 10108 31612 10118
rect 30884 9146 30940 9156
rect 30324 9100 30380 9110
rect 30324 9002 30326 9044
rect 30378 9002 30380 9044
rect 30324 8990 30380 9002
rect 30100 8428 30156 8820
rect 31108 8988 31164 8998
rect 30212 8428 30268 8438
rect 30100 8372 30212 8428
rect 30100 7420 30156 8372
rect 30212 8334 30268 8372
rect 30884 8092 30940 8102
rect 30884 7998 30940 8036
rect 30472 7868 30736 7878
rect 30528 7812 30576 7868
rect 30632 7812 30680 7868
rect 30472 7802 30736 7812
rect 30884 7644 30940 7654
rect 30884 7550 30940 7588
rect 29876 7364 30156 7420
rect 30268 7420 30324 7430
rect 29876 6702 29932 7364
rect 30268 7326 30324 7364
rect 30380 7308 30436 7318
rect 30380 7214 30436 7252
rect 29876 6650 29878 6702
rect 29930 6650 29932 6702
rect 29876 6300 29932 6650
rect 30996 6636 31052 6646
rect 29876 6234 29932 6244
rect 30472 6300 30736 6310
rect 30528 6244 30576 6300
rect 30632 6244 30680 6300
rect 30472 6234 30736 6244
rect 29652 6188 29708 6198
rect 29652 6074 29708 6132
rect 29652 6022 29654 6074
rect 29706 6022 29708 6074
rect 29652 6010 29708 6022
rect 30884 6076 30940 6086
rect 30884 5982 30940 6020
rect 29316 5238 29318 5290
rect 29370 5238 29372 5290
rect 29316 5226 29372 5238
rect 29764 5964 29820 5974
rect 29764 5134 29820 5908
rect 29764 5082 29766 5134
rect 29818 5082 29820 5134
rect 29764 5068 29820 5082
rect 29652 5012 29820 5068
rect 29876 5738 29932 5750
rect 29876 5686 29878 5738
rect 29930 5686 29932 5738
rect 29036 4956 29092 4966
rect 29036 4862 29092 4900
rect 29260 4956 29316 4966
rect 29260 4862 29316 4900
rect 29092 4338 29148 4350
rect 29092 4286 29094 4338
rect 29146 4286 29148 4338
rect 29092 4284 29148 4286
rect 29092 4218 29148 4228
rect 29428 4172 29484 4182
rect 29428 4170 29596 4172
rect 29428 4118 29430 4170
rect 29482 4118 29596 4170
rect 29428 4116 29596 4118
rect 29428 4106 29484 4116
rect 28532 3514 28534 3566
rect 28586 3514 28588 3566
rect 28532 3502 28588 3514
rect 28700 3612 28756 3622
rect 28700 3498 28756 3556
rect 28700 3446 28702 3498
rect 28754 3446 28756 3498
rect 28700 3387 28756 3446
rect 27804 3386 28364 3387
rect 27804 3334 27806 3386
rect 27858 3334 28364 3386
rect 27804 3331 28364 3334
rect 28420 3331 28588 3387
rect 27804 3322 27860 3331
rect 27188 2826 27244 2838
rect 27188 2774 27190 2826
rect 27242 2774 27244 2826
rect 26908 2604 26964 2614
rect 26740 2426 26796 2436
rect 26852 2602 26964 2604
rect 26852 2550 26910 2602
rect 26962 2550 26964 2602
rect 26852 2538 26964 2550
rect 27188 2604 27244 2774
rect 27188 2538 27244 2548
rect 27412 2828 27468 2838
rect 27412 2770 27468 2772
rect 27412 2718 27414 2770
rect 27466 2718 27468 2770
rect 25396 2202 25452 2212
rect 25956 2380 26012 2390
rect 25452 1986 25508 1998
rect 25452 1934 25454 1986
rect 25506 1934 25508 1986
rect 25452 1932 25508 1934
rect 25396 1876 25508 1932
rect 25956 1932 26012 2324
rect 26196 2380 26460 2390
rect 26252 2324 26300 2380
rect 26356 2324 26404 2380
rect 26196 2314 26460 2324
rect 25396 1370 25452 1876
rect 25396 1318 25398 1370
rect 25450 1318 25452 1370
rect 25396 1306 25452 1318
rect 25732 1596 25788 1606
rect 25228 1260 25340 1270
rect 25284 1204 25340 1260
rect 25732 1214 25788 1540
rect 25228 1128 25284 1204
rect 25732 1162 25734 1214
rect 25786 1162 25788 1214
rect 25956 1270 26012 1876
rect 26740 1932 26796 1942
rect 26572 1820 26628 1830
rect 25956 1258 26068 1270
rect 25956 1206 26014 1258
rect 26066 1206 26068 1258
rect 25956 1204 26068 1206
rect 26012 1194 26068 1204
rect 26572 1258 26628 1764
rect 26740 1270 26796 1876
rect 26852 1596 26908 2538
rect 27412 1932 27468 2718
rect 27412 1866 27468 1876
rect 26852 1530 26908 1540
rect 27524 1382 27580 2884
rect 27468 1370 27580 1382
rect 27468 1318 27470 1370
rect 27522 1318 27580 1370
rect 27468 1316 27580 1318
rect 27636 3108 27748 3164
rect 28196 3164 28252 3174
rect 27636 1320 27692 3108
rect 28196 2782 28252 3108
rect 28308 2940 28364 3331
rect 28532 3276 28588 3331
rect 28532 3210 28588 3220
rect 28644 3331 28756 3387
rect 28308 2884 28476 2940
rect 28196 2730 28198 2782
rect 28250 2730 28252 2782
rect 28196 2718 28252 2730
rect 28420 2546 28476 2884
rect 28532 2758 28588 2770
rect 28532 2716 28534 2758
rect 28586 2716 28588 2758
rect 28532 2650 28588 2660
rect 28308 2492 28364 2502
rect 28420 2494 28422 2546
rect 28474 2494 28476 2546
rect 28420 2482 28476 2494
rect 28084 2268 28140 2278
rect 27860 2044 27916 2054
rect 27860 1950 27916 1988
rect 27468 1306 27524 1316
rect 26572 1206 26574 1258
rect 26626 1206 26628 1258
rect 26572 1194 26628 1206
rect 26684 1258 26796 1270
rect 26684 1206 26686 1258
rect 26738 1206 26796 1258
rect 26684 1204 26796 1206
rect 26908 1260 26964 1270
rect 26684 1194 26740 1204
rect 26908 1166 26964 1204
rect 27132 1260 27188 1270
rect 27636 1268 27638 1320
rect 27690 1268 27692 1320
rect 27636 1256 27692 1268
rect 27748 1932 27804 1942
rect 27132 1166 27188 1204
rect 27748 1210 27804 1876
rect 25732 1150 25788 1162
rect 27748 1158 27750 1210
rect 27802 1158 27804 1210
rect 28084 1270 28140 2212
rect 28308 1270 28364 2436
rect 28532 1932 28588 1942
rect 28532 1838 28588 1876
rect 28644 1270 28700 3331
rect 28868 3164 28924 3780
rect 28980 3724 29036 3734
rect 28980 3722 29372 3724
rect 28980 3670 28982 3722
rect 29034 3670 29372 3722
rect 28980 3668 29372 3670
rect 28980 3658 29036 3668
rect 29316 3622 29372 3668
rect 29316 3610 29428 3622
rect 28868 3098 28924 3108
rect 28980 3542 29036 3576
rect 29316 3558 29374 3610
rect 29426 3558 29428 3610
rect 29316 3556 29428 3558
rect 29372 3546 29428 3556
rect 28980 3500 28982 3542
rect 29034 3500 29036 3542
rect 28812 2716 28868 2726
rect 28980 2716 29036 3444
rect 29092 3388 29148 3398
rect 29148 3332 29204 3387
rect 29092 3322 29204 3332
rect 29148 2938 29204 3322
rect 29148 2886 29150 2938
rect 29202 2886 29204 2938
rect 29148 2874 29204 2886
rect 29316 3276 29372 3286
rect 29316 2888 29372 3220
rect 29316 2836 29318 2888
rect 29370 2836 29372 2888
rect 29316 2824 29372 2836
rect 29428 3164 29484 3174
rect 28812 2714 29036 2716
rect 29428 2778 29484 3108
rect 29428 2726 29430 2778
rect 29482 2726 29484 2778
rect 29428 2714 29484 2726
rect 29540 2716 29596 4116
rect 29652 3836 29708 5012
rect 29876 4620 29932 5686
rect 30212 5740 30268 5750
rect 30212 5646 30268 5684
rect 29876 4554 29932 4564
rect 30212 5110 30268 5122
rect 30212 5058 30214 5110
rect 30266 5058 30268 5110
rect 29764 4450 29820 4462
rect 29764 4398 29766 4450
rect 29818 4398 29820 4450
rect 29764 4396 29820 4398
rect 29764 4330 29820 4340
rect 29820 4172 29876 4182
rect 29820 4078 29876 4116
rect 30044 4114 30100 4126
rect 30044 4062 30046 4114
rect 30098 4062 30100 4114
rect 30044 4060 30100 4062
rect 30044 3836 30100 4004
rect 29652 3770 29708 3780
rect 29764 3778 29820 3790
rect 29764 3726 29766 3778
rect 29818 3726 29820 3778
rect 29652 3612 29708 3622
rect 29652 3514 29654 3556
rect 29706 3514 29708 3556
rect 29652 3502 29708 3514
rect 29764 3388 29820 3726
rect 29764 3322 29820 3332
rect 29876 3780 30100 3836
rect 28812 2662 28814 2714
rect 28866 2662 29036 2714
rect 28812 2660 29036 2662
rect 28812 2154 28868 2660
rect 29540 2650 29596 2660
rect 29652 3276 29708 3286
rect 29652 2166 29708 3220
rect 29876 3164 29932 3780
rect 30212 3724 30268 5058
rect 30472 4732 30736 4742
rect 30528 4676 30576 4732
rect 30632 4676 30680 4732
rect 30472 4666 30736 4676
rect 30884 4508 30940 4518
rect 30884 4414 30940 4452
rect 30100 3668 30268 3724
rect 30324 4324 30380 4336
rect 30324 4272 30326 4324
rect 30378 4272 30380 4324
rect 30324 3724 30380 4272
rect 29988 3542 30044 3554
rect 29988 3500 29990 3542
rect 30042 3500 30044 3542
rect 29988 3434 30044 3444
rect 30100 3276 30156 3668
rect 30324 3658 30380 3668
rect 30436 3836 30492 3846
rect 30996 3836 31052 6580
rect 30436 3567 30492 3780
rect 30436 3515 30438 3567
rect 30490 3515 30492 3567
rect 30268 3498 30324 3510
rect 30436 3503 30492 3515
rect 30548 3780 31052 3836
rect 31108 3836 31164 8932
rect 31556 8874 31612 10052
rect 31780 9814 31836 9826
rect 31780 9762 31782 9814
rect 31834 9762 31836 9814
rect 31780 8988 31836 9762
rect 32340 9818 32396 10500
rect 32340 9772 32342 9818
rect 32394 9772 32396 9818
rect 32340 9706 32396 9716
rect 31780 8922 31836 8932
rect 32564 9658 32620 9670
rect 32564 9606 32566 9658
rect 32618 9606 32620 9658
rect 31556 8822 31558 8874
rect 31610 8822 31612 8874
rect 31556 8428 31612 8822
rect 32452 8652 32508 8662
rect 31444 8258 31500 8270
rect 31220 8204 31276 8214
rect 31220 8110 31276 8148
rect 31444 8206 31446 8258
rect 31498 8206 31500 8258
rect 31444 7644 31500 8206
rect 31444 7578 31500 7588
rect 31556 7306 31612 8372
rect 31780 8482 31836 8494
rect 31780 8430 31782 8482
rect 31834 8430 31836 8482
rect 31780 8428 31836 8430
rect 31780 8362 31836 8372
rect 31556 7254 31558 7306
rect 31610 7254 31612 7306
rect 31556 5738 31612 7254
rect 32116 6678 32172 6690
rect 32116 6626 32118 6678
rect 32170 6626 32172 6678
rect 32116 6188 32172 6626
rect 32116 6122 32172 6132
rect 31556 5686 31558 5738
rect 31610 5686 31612 5738
rect 31556 4172 31612 5686
rect 31556 4078 31612 4116
rect 30268 3446 30270 3498
rect 30322 3446 30324 3498
rect 30268 3388 30324 3446
rect 30548 3388 30604 3780
rect 30940 3554 30996 3566
rect 30940 3502 30942 3554
rect 30994 3502 30996 3554
rect 30940 3500 30996 3502
rect 30268 3332 30604 3388
rect 30884 3444 30996 3500
rect 30100 3220 30268 3276
rect 28812 2102 28814 2154
rect 28866 2102 28868 2154
rect 28812 2090 28868 2102
rect 28924 2156 28980 2166
rect 28924 2062 28980 2100
rect 29596 2154 29708 2166
rect 29596 2102 29598 2154
rect 29650 2102 29708 2154
rect 29596 2100 29708 2102
rect 29764 3108 29932 3164
rect 29764 2156 29820 3108
rect 29876 2716 29988 2726
rect 29932 2714 29988 2716
rect 29932 2662 29934 2714
rect 29986 2662 29988 2714
rect 29932 2660 29988 2662
rect 29876 2650 29988 2660
rect 30212 2604 30268 3220
rect 30472 3164 30736 3174
rect 30528 3108 30576 3164
rect 30632 3108 30680 3164
rect 30472 3098 30736 3108
rect 30884 3052 30940 3444
rect 30772 2996 30940 3052
rect 30996 3276 31052 3286
rect 30324 2940 30380 2950
rect 30772 2940 30828 2996
rect 30324 2938 30828 2940
rect 30324 2886 30326 2938
rect 30378 2886 30828 2938
rect 30324 2884 30828 2886
rect 30324 2874 30380 2884
rect 30884 2828 30940 2838
rect 30884 2730 30886 2772
rect 30938 2730 30940 2772
rect 30212 2548 30492 2604
rect 29596 2090 29652 2100
rect 29764 2090 29820 2100
rect 29988 2492 30044 2502
rect 29148 2044 29204 2054
rect 29148 1932 29204 1988
rect 29372 1932 29428 1942
rect 29148 1930 29428 1932
rect 29148 1878 29150 1930
rect 29202 1878 29374 1930
rect 29426 1878 29428 1930
rect 29148 1876 29428 1878
rect 29148 1866 29204 1876
rect 28084 1260 28196 1270
rect 28084 1204 28140 1260
rect 28308 1258 28420 1270
rect 28308 1206 28366 1258
rect 28418 1206 28420 1258
rect 28308 1204 28420 1206
rect 28140 1166 28196 1204
rect 28364 1194 28420 1204
rect 28588 1258 28700 1270
rect 28588 1206 28590 1258
rect 28642 1206 28700 1258
rect 28588 1204 28700 1206
rect 28812 1708 28868 1718
rect 28812 1258 28868 1652
rect 28812 1206 28814 1258
rect 28866 1206 28868 1258
rect 28588 1194 28644 1204
rect 28812 1194 28868 1206
rect 28924 1484 28980 1494
rect 28924 1258 28980 1428
rect 29372 1484 29428 1876
rect 29372 1418 29428 1428
rect 29988 1708 30044 2436
rect 30436 2154 30492 2548
rect 30436 2102 30438 2154
rect 30490 2102 30492 2154
rect 30436 2090 30492 2102
rect 30884 2044 30940 2730
rect 30828 1986 30940 2044
rect 30100 1974 30156 1986
rect 30100 1922 30102 1974
rect 30154 1922 30156 1974
rect 30828 1934 30830 1986
rect 30882 1934 30940 1986
rect 30828 1922 30940 1934
rect 30100 1708 30156 1922
rect 29988 1652 30156 1708
rect 30884 1708 30940 1922
rect 28924 1206 28926 1258
rect 28978 1206 28980 1258
rect 28924 1194 28980 1206
rect 29372 1260 29428 1270
rect 29764 1260 29820 1270
rect 29372 1258 29820 1260
rect 29372 1206 29374 1258
rect 29426 1206 29766 1258
rect 29818 1206 29820 1258
rect 29372 1204 29820 1206
rect 29372 1194 29428 1204
rect 29764 1194 29820 1204
rect 26348 1148 26404 1158
rect 27748 1146 27804 1158
rect 26348 1054 26404 1092
rect 23100 1036 23156 1046
rect 23772 1036 23828 1046
rect 24220 1036 24276 1046
rect 22708 1034 24276 1036
rect 22708 982 23102 1034
rect 23154 982 23774 1034
rect 23826 982 24222 1034
rect 24274 982 24276 1034
rect 22708 980 24276 982
rect 24948 1034 25060 1046
rect 24948 982 25006 1034
rect 25058 982 25060 1034
rect 24948 980 25060 982
rect 23100 970 23156 980
rect 23772 970 23828 980
rect 24220 970 24276 980
rect 25004 970 25060 980
rect 29484 1036 29540 1046
rect 29484 942 29540 980
rect 26196 812 26460 822
rect 26252 756 26300 812
rect 26356 756 26404 812
rect 26196 746 26460 756
rect 22540 534 22542 586
rect 22594 534 22596 586
rect 22540 522 22596 534
rect 29988 588 30044 1652
rect 30884 1642 30940 1652
rect 30472 1596 30736 1606
rect 30528 1540 30576 1596
rect 30632 1540 30680 1596
rect 30472 1530 30736 1540
rect 30716 1260 30772 1270
rect 30100 1184 30156 1196
rect 30100 1132 30102 1184
rect 30154 1132 30156 1184
rect 30100 924 30156 1132
rect 30716 1036 30772 1204
rect 30996 1214 31052 3220
rect 31108 2828 31164 3780
rect 31108 2762 31164 2772
rect 31444 3052 31500 3062
rect 31444 2782 31500 2996
rect 31444 2730 31446 2782
rect 31498 2730 31500 2782
rect 31444 2718 31500 2730
rect 31276 1986 31332 1998
rect 31276 1934 31278 1986
rect 31330 1934 31332 1986
rect 31276 1932 31332 1934
rect 31276 1876 31388 1932
rect 31332 1370 31388 1876
rect 31332 1318 31334 1370
rect 31386 1318 31388 1370
rect 31332 1306 31388 1318
rect 31500 1596 31556 1606
rect 30996 1162 30998 1214
rect 31050 1162 31052 1214
rect 31500 1258 31556 1540
rect 32452 1370 32508 8596
rect 32564 8316 32620 9606
rect 32564 8224 32566 8260
rect 32618 8224 32620 8260
rect 32564 8184 32620 8224
rect 32564 6682 32620 6694
rect 32564 6630 32566 6682
rect 32618 6630 32620 6682
rect 32564 5964 32620 6630
rect 32564 5898 32620 5908
rect 32564 5740 32620 5750
rect 32564 5178 32620 5684
rect 32676 5292 32732 12180
rect 33460 11564 33516 13200
rect 33348 11508 33516 11564
rect 33572 12056 33628 12068
rect 33572 12004 33574 12056
rect 33626 12004 33628 12056
rect 32956 9996 33012 10006
rect 33180 9996 33236 10006
rect 32956 9994 33180 9996
rect 32956 9942 32958 9994
rect 33010 9942 33180 9994
rect 32956 9940 33180 9942
rect 32956 9930 33068 9940
rect 33012 8540 33068 9930
rect 33180 9902 33236 9940
rect 33348 9884 33404 11508
rect 33572 11394 33628 12004
rect 34524 12012 34580 12022
rect 34524 12010 34748 12012
rect 34524 11958 34526 12010
rect 34578 11958 34748 12010
rect 34524 11956 34748 11958
rect 34524 11946 34580 11956
rect 33572 11342 33574 11394
rect 33626 11342 33628 11394
rect 33572 10444 33628 11342
rect 34468 11228 34524 11238
rect 34244 11226 34524 11228
rect 34244 11174 34470 11226
rect 34522 11174 34524 11226
rect 34244 11172 34524 11174
rect 33796 10444 33852 10454
rect 33572 10442 33852 10444
rect 33572 10390 33798 10442
rect 33850 10390 33852 10442
rect 33572 10388 33852 10390
rect 33796 10108 33852 10388
rect 33796 10042 33852 10052
rect 33348 9818 33404 9828
rect 33684 9884 33740 9894
rect 33684 9790 33740 9828
rect 33964 9042 34020 9054
rect 33012 8474 33068 8484
rect 33348 8988 33404 8998
rect 33964 8990 33966 9042
rect 34018 8990 34020 9042
rect 33964 8988 34020 8990
rect 33964 8932 34076 8988
rect 32788 8428 32844 8438
rect 32788 6860 32844 8372
rect 33348 8314 33404 8932
rect 34020 8426 34076 8932
rect 34020 8374 34022 8426
rect 34074 8374 34076 8426
rect 34020 8362 34076 8374
rect 33348 8262 33350 8314
rect 33402 8262 33404 8314
rect 33348 8250 33404 8262
rect 33684 8246 33740 8258
rect 32900 8204 32956 8214
rect 33068 8204 33124 8214
rect 33684 8204 33686 8246
rect 33738 8204 33740 8246
rect 32900 8202 33180 8204
rect 32900 8150 32902 8202
rect 32954 8150 33070 8202
rect 33122 8150 33180 8202
rect 32900 8148 33180 8150
rect 32900 8138 32956 8148
rect 33068 8138 33180 8148
rect 33684 8138 33740 8148
rect 32956 6860 33012 6870
rect 32788 6858 33012 6860
rect 32788 6806 32958 6858
rect 33010 6806 33012 6858
rect 32788 6804 33012 6806
rect 32956 6794 33012 6804
rect 33124 6748 33180 8138
rect 33908 7462 33964 7474
rect 33908 7410 33910 7462
rect 33962 7410 33964 7462
rect 33124 6682 33180 6692
rect 33348 6748 33404 6758
rect 33348 6634 33404 6692
rect 33908 6748 33964 7410
rect 33908 6682 33964 6692
rect 33348 6582 33350 6634
rect 33402 6582 33404 6634
rect 33348 6570 33404 6582
rect 33516 6636 33572 6646
rect 33740 6636 33796 6646
rect 34132 6636 34188 6646
rect 33516 6634 33628 6636
rect 33516 6582 33518 6634
rect 33570 6582 33628 6634
rect 33516 6570 33628 6582
rect 33740 6634 33852 6636
rect 33740 6582 33742 6634
rect 33794 6582 33852 6634
rect 33740 6570 33852 6582
rect 33572 6524 33628 6570
rect 33460 5292 33516 5302
rect 32676 5290 33516 5292
rect 32676 5238 33462 5290
rect 33514 5238 33516 5290
rect 32676 5236 33516 5238
rect 33460 5226 33516 5236
rect 32564 5126 32566 5178
rect 32618 5126 32620 5178
rect 32564 4172 32620 5126
rect 33348 5068 33404 5078
rect 33236 4956 33292 4966
rect 33236 4862 33292 4900
rect 32564 4106 32620 4116
rect 33236 4172 33292 4182
rect 33236 3542 33292 4116
rect 33236 3490 33238 3542
rect 33290 3490 33292 3542
rect 33236 2716 33292 3490
rect 33236 2650 33292 2660
rect 32452 1318 32454 1370
rect 32506 1318 32508 1370
rect 32452 1306 32508 1318
rect 33348 1320 33404 5012
rect 33572 3387 33628 6468
rect 33684 5852 33740 5862
rect 33684 4844 33740 5796
rect 33796 5740 33852 6570
rect 34020 6522 34076 6534
rect 34020 6470 34022 6522
rect 34074 6470 34076 6522
rect 34020 5964 34076 6470
rect 33964 5908 34076 5964
rect 33964 5906 34020 5908
rect 33964 5854 33966 5906
rect 34018 5854 34020 5906
rect 33964 5842 34020 5854
rect 33796 5674 33852 5684
rect 34132 5302 34188 6580
rect 34244 5628 34300 11172
rect 34468 11162 34524 11172
rect 34468 10668 34524 10678
rect 34468 10666 34636 10668
rect 34468 10614 34470 10666
rect 34522 10614 34636 10666
rect 34468 10612 34636 10614
rect 34468 10602 34524 10612
rect 34580 9996 34636 10612
rect 34356 9772 34412 9782
rect 34356 9054 34412 9716
rect 34356 9002 34358 9054
rect 34410 9002 34412 9054
rect 34356 8990 34412 9002
rect 34468 9658 34524 9670
rect 34468 9606 34470 9658
rect 34522 9606 34524 9658
rect 34356 8246 34412 8258
rect 34356 8194 34358 8246
rect 34410 8194 34412 8246
rect 34356 7868 34412 8194
rect 34356 7802 34412 7812
rect 34468 7462 34524 9606
rect 34468 7410 34470 7462
rect 34522 7410 34524 7462
rect 34356 6678 34412 6690
rect 34356 6636 34358 6678
rect 34410 6636 34412 6678
rect 34356 6570 34412 6580
rect 34468 6524 34524 7410
rect 34468 6458 34524 6468
rect 34244 5562 34300 5572
rect 34356 5964 34412 5974
rect 34356 5894 34412 5908
rect 34356 5842 34358 5894
rect 34410 5842 34412 5894
rect 34356 5516 34412 5842
rect 34356 5460 34524 5516
rect 34076 5290 34188 5302
rect 34076 5238 34078 5290
rect 34130 5238 34188 5290
rect 34076 5236 34188 5238
rect 34300 5292 34356 5302
rect 34076 5226 34132 5236
rect 34300 5198 34356 5236
rect 33796 5110 33852 5122
rect 33796 5068 33798 5110
rect 33850 5068 33852 5110
rect 33796 5002 33852 5012
rect 33908 4956 33964 4966
rect 33684 4788 33852 4844
rect 33796 3387 33852 4788
rect 33908 4350 33964 4900
rect 33908 4298 33910 4350
rect 33962 4298 33964 4350
rect 33908 4286 33964 4298
rect 34468 4350 34524 5460
rect 34580 5292 34636 9940
rect 34580 5226 34636 5236
rect 34468 4298 34470 4350
rect 34522 4298 34524 4350
rect 34244 4284 34300 4294
rect 34468 4286 34524 4298
rect 34580 4396 34636 4406
rect 34244 3722 34300 4228
rect 34244 3670 34246 3722
rect 34298 3670 34300 3722
rect 34244 3658 34300 3670
rect 34412 3612 34468 3622
rect 34412 3518 34468 3556
rect 33572 3331 33740 3387
rect 33796 3331 34076 3387
rect 33460 2716 33516 2726
rect 33460 1998 33516 2660
rect 33460 1946 33462 1998
rect 33514 1946 33516 1998
rect 33460 1708 33516 1946
rect 33460 1642 33516 1652
rect 31500 1206 31502 1258
rect 31554 1206 31556 1258
rect 31500 1194 31556 1206
rect 32788 1260 32844 1270
rect 33348 1268 33350 1320
rect 33402 1268 33404 1320
rect 33516 1372 33572 1382
rect 33516 1278 33572 1316
rect 33348 1256 33404 1268
rect 30996 1150 31052 1162
rect 31892 1184 31948 1196
rect 31892 1148 31894 1184
rect 31946 1148 31948 1184
rect 32788 1162 32790 1204
rect 32842 1162 32844 1204
rect 31892 1082 31948 1092
rect 32228 1148 32284 1158
rect 32788 1150 32844 1162
rect 33124 1202 33180 1214
rect 33124 1150 33126 1202
rect 33178 1150 33180 1202
rect 32228 1054 32284 1092
rect 33124 1148 33180 1150
rect 33124 1082 33180 1092
rect 30716 942 30772 980
rect 33684 1036 33740 3331
rect 33796 2716 33852 2726
rect 33796 2622 33852 2660
rect 34020 1370 34076 3331
rect 34468 2940 34524 2950
rect 34468 2846 34524 2884
rect 34468 2156 34524 2166
rect 34468 2062 34524 2100
rect 34020 1318 34022 1370
rect 34074 1318 34076 1370
rect 34020 1306 34076 1318
rect 34580 1260 34636 4340
rect 34692 1372 34748 11956
rect 34692 1306 34748 1316
rect 34468 1204 34636 1260
rect 34468 1158 34524 1204
rect 34412 1146 34524 1158
rect 34412 1094 34414 1146
rect 34466 1094 34524 1146
rect 34412 1082 34524 1094
rect 33684 970 33740 980
rect 33852 1036 33908 1046
rect 33852 942 33908 980
rect 30100 858 30156 868
rect 34468 700 34524 1082
rect 34468 634 34524 644
rect 29988 522 30044 532
rect 22316 422 22318 474
rect 22370 422 22372 474
rect 22316 410 22372 422
<< via2 >>
rect 1820 12234 1876 12236
rect 1820 12182 1822 12234
rect 1822 12182 1874 12234
rect 1874 12182 1876 12234
rect 1820 12180 1876 12182
rect 4816 12570 4872 12572
rect 4816 12518 4818 12570
rect 4818 12518 4870 12570
rect 4870 12518 4872 12570
rect 4816 12516 4872 12518
rect 4920 12570 4976 12572
rect 4920 12518 4922 12570
rect 4922 12518 4974 12570
rect 4974 12518 4976 12570
rect 4920 12516 4976 12518
rect 5024 12570 5080 12572
rect 5024 12518 5026 12570
rect 5026 12518 5078 12570
rect 5078 12518 5080 12570
rect 5024 12516 5080 12518
rect 2548 12180 2604 12236
rect 1092 11396 1148 11452
rect 1372 11450 1428 11452
rect 1372 11398 1374 11450
rect 1374 11398 1426 11450
rect 1426 11398 1428 11450
rect 1372 11396 1428 11398
rect 1708 10836 1764 10892
rect 1540 10388 1596 10444
rect 2156 11620 2212 11676
rect 2828 11620 2884 11676
rect 3892 11620 3948 11676
rect 2604 11450 2660 11452
rect 2604 11398 2606 11450
rect 2606 11398 2658 11450
rect 2658 11398 2660 11450
rect 2604 11396 2660 11398
rect 3276 11450 3332 11452
rect 3276 11398 3278 11450
rect 3278 11398 3330 11450
rect 3330 11398 3332 11450
rect 3276 11396 3332 11398
rect 2212 9604 2268 9660
rect 1316 9044 1372 9100
rect 2492 9492 2548 9548
rect 980 8932 1036 8988
rect 1484 8596 1540 8652
rect 1932 9098 1988 9100
rect 1932 9046 1934 9098
rect 1934 9046 1986 9098
rect 1986 9046 1988 9098
rect 1932 9044 1988 9046
rect 3668 10276 3724 10332
rect 4340 11396 4396 11452
rect 4004 11338 4060 11340
rect 4004 11286 4006 11338
rect 4006 11286 4058 11338
rect 4058 11286 4060 11338
rect 4004 11284 4060 11286
rect 3892 11172 3948 11228
rect 4788 11330 4790 11340
rect 4790 11330 4842 11340
rect 4842 11330 4844 11340
rect 4788 11284 4844 11330
rect 6916 11508 6972 11564
rect 4900 11172 4956 11228
rect 7140 11172 7196 11228
rect 12404 12346 12460 12348
rect 12404 12294 12406 12346
rect 12406 12294 12458 12346
rect 12458 12294 12460 12346
rect 12404 12292 12460 12294
rect 13368 12570 13424 12572
rect 13368 12518 13370 12570
rect 13370 12518 13422 12570
rect 13422 12518 13424 12570
rect 13368 12516 13424 12518
rect 13472 12570 13528 12572
rect 13472 12518 13474 12570
rect 13474 12518 13526 12570
rect 13526 12518 13528 12570
rect 13472 12516 13528 12518
rect 13576 12570 13632 12572
rect 13576 12518 13578 12570
rect 13578 12518 13630 12570
rect 13630 12518 13632 12570
rect 13576 12516 13632 12518
rect 12852 12292 12908 12348
rect 13356 12180 13412 12236
rect 7700 11732 7756 11788
rect 9092 11786 9148 11788
rect 9092 11734 9094 11786
rect 9094 11734 9146 11786
rect 9146 11734 9148 11786
rect 9092 11732 9148 11734
rect 9196 11786 9252 11788
rect 9196 11734 9198 11786
rect 9198 11734 9250 11786
rect 9250 11734 9252 11786
rect 9196 11732 9252 11734
rect 9300 11786 9356 11788
rect 9300 11734 9302 11786
rect 9302 11734 9354 11786
rect 9354 11734 9356 11786
rect 9300 11732 9356 11734
rect 10388 12114 10390 12124
rect 10390 12114 10442 12124
rect 10442 12114 10444 12124
rect 10388 12068 10444 12114
rect 9940 11732 9996 11788
rect 10276 11620 10332 11676
rect 8372 11510 8428 11564
rect 8372 11508 8374 11510
rect 8374 11508 8426 11510
rect 8426 11508 8428 11510
rect 9940 11508 9996 11564
rect 7588 11172 7644 11228
rect 4816 11002 4872 11004
rect 4816 10950 4818 11002
rect 4818 10950 4870 11002
rect 4870 10950 4872 11002
rect 4816 10948 4872 10950
rect 4920 11002 4976 11004
rect 4920 10950 4922 11002
rect 4922 10950 4974 11002
rect 4974 10950 4976 11002
rect 4920 10948 4976 10950
rect 5024 11002 5080 11004
rect 5024 10950 5026 11002
rect 5026 10950 5078 11002
rect 5078 10950 5080 11002
rect 5024 10948 5080 10950
rect 7252 10948 7308 11004
rect 5964 10836 6020 10892
rect 4340 10612 4396 10668
rect 2996 9492 3052 9548
rect 5068 10442 5124 10444
rect 5068 10390 5070 10442
rect 5070 10390 5122 10442
rect 5122 10390 5124 10442
rect 5068 10388 5124 10390
rect 4788 10164 4844 10220
rect 6412 10666 6468 10668
rect 6412 10614 6414 10666
rect 6414 10614 6466 10666
rect 6466 10614 6468 10666
rect 6412 10612 6468 10614
rect 5012 9940 5068 9996
rect 4564 9770 4620 9772
rect 4564 9718 4566 9770
rect 4566 9718 4618 9770
rect 4618 9718 4620 9770
rect 4564 9716 4620 9718
rect 3108 9268 3164 9324
rect 2492 9044 2548 9100
rect 2660 9098 2716 9100
rect 2660 9046 2662 9098
rect 2662 9046 2714 9098
rect 2714 9046 2716 9098
rect 2660 9044 2716 9046
rect 2660 8820 2716 8876
rect 2996 8874 3052 8876
rect 2996 8822 2998 8874
rect 2998 8822 3050 8874
rect 3050 8822 3052 8874
rect 2996 8820 3052 8822
rect 2268 8708 2324 8764
rect 2660 8596 2716 8652
rect 3332 8972 3334 8988
rect 3334 8972 3386 8988
rect 3386 8972 3388 8988
rect 3332 8932 3388 8972
rect 2660 6804 2716 6860
rect 3500 7140 3556 7196
rect 3500 6858 3556 6860
rect 3500 6806 3502 6858
rect 3502 6806 3554 6858
rect 3554 6806 3556 6858
rect 3500 6804 3556 6806
rect 1092 6580 1148 6636
rect 3892 9044 3948 9100
rect 5124 9658 5180 9660
rect 5124 9606 5126 9658
rect 5126 9606 5178 9658
rect 5178 9606 5180 9658
rect 5124 9604 5180 9606
rect 5236 9492 5292 9548
rect 4816 9434 4872 9436
rect 4816 9382 4818 9434
rect 4818 9382 4870 9434
rect 4870 9382 4872 9434
rect 4816 9380 4872 9382
rect 4920 9434 4976 9436
rect 4920 9382 4922 9434
rect 4922 9382 4974 9434
rect 4974 9382 4976 9434
rect 4920 9380 4976 9382
rect 5024 9434 5080 9436
rect 5024 9382 5026 9434
rect 5026 9382 5078 9434
rect 5078 9382 5080 9434
rect 5024 9380 5080 9382
rect 5124 9156 5180 9212
rect 4956 8986 5012 8988
rect 4956 8934 4958 8986
rect 4958 8934 5010 8986
rect 5010 8934 5012 8986
rect 4956 8932 5012 8934
rect 6132 10388 6188 10444
rect 5740 9828 5796 9884
rect 6076 10164 6132 10220
rect 5852 9770 5908 9772
rect 5852 9718 5854 9770
rect 5854 9718 5906 9770
rect 5906 9718 5908 9770
rect 5852 9716 5908 9718
rect 7476 10388 7532 10444
rect 7252 10164 7308 10220
rect 7532 10164 7588 10220
rect 6916 10052 6972 10108
rect 7140 10052 7196 10108
rect 6468 9940 6524 9996
rect 6636 9940 6692 9996
rect 8708 11450 8764 11452
rect 8708 11398 8710 11450
rect 8710 11398 8762 11450
rect 8762 11398 8764 11450
rect 8708 11396 8764 11398
rect 9436 11338 9492 11340
rect 9436 11286 9438 11338
rect 9438 11286 9490 11338
rect 9490 11286 9492 11338
rect 9436 11284 9492 11286
rect 9100 11226 9156 11228
rect 9100 11174 9102 11226
rect 9102 11174 9154 11226
rect 9154 11174 9156 11226
rect 9100 11172 9156 11174
rect 8372 11060 8428 11116
rect 9548 10778 9604 10780
rect 9548 10726 9550 10778
rect 9550 10726 9602 10778
rect 9602 10726 9604 10778
rect 9548 10724 9604 10726
rect 10500 11508 10556 11564
rect 10612 11396 10668 11452
rect 8764 10666 8820 10668
rect 8764 10614 8766 10666
rect 8766 10614 8818 10666
rect 8818 10614 8820 10666
rect 8764 10612 8820 10614
rect 8036 10500 8092 10556
rect 8988 10554 9044 10556
rect 8988 10502 8990 10554
rect 8990 10502 9042 10554
rect 9042 10502 9044 10554
rect 8988 10500 9044 10502
rect 9156 10442 9212 10444
rect 7924 10052 7980 10108
rect 9156 10390 9158 10442
rect 9158 10390 9210 10442
rect 9210 10390 9212 10442
rect 9156 10388 9212 10390
rect 8092 9940 8148 9996
rect 6972 9882 7028 9884
rect 6972 9830 6974 9882
rect 6974 9830 7026 9882
rect 7026 9830 7028 9882
rect 6972 9828 7028 9830
rect 5460 8932 5516 8988
rect 4396 8708 4452 8764
rect 5236 8820 5292 8876
rect 4172 8260 4228 8316
rect 4732 8596 4788 8652
rect 7476 9716 7532 9772
rect 6468 9380 6524 9436
rect 6972 9380 7028 9436
rect 6188 9210 6244 9212
rect 6188 9158 6190 9210
rect 6190 9158 6242 9210
rect 6242 9158 6244 9210
rect 6188 9156 6244 9158
rect 6524 9098 6580 9100
rect 6524 9046 6526 9098
rect 6526 9046 6578 9098
rect 6578 9046 6580 9098
rect 6524 9044 6580 9046
rect 5908 8982 5910 8988
rect 5910 8982 5962 8988
rect 5962 8982 5964 8988
rect 5908 8932 5964 8982
rect 6860 8932 6916 8988
rect 5572 8372 5628 8428
rect 7252 9210 7308 9212
rect 7252 9158 7254 9210
rect 7254 9158 7306 9210
rect 7306 9158 7308 9210
rect 7252 9156 7308 9158
rect 7756 9716 7812 9772
rect 7700 9380 7756 9436
rect 7140 8820 7196 8876
rect 8260 9716 8316 9772
rect 9092 10218 9148 10220
rect 9092 10166 9094 10218
rect 9094 10166 9146 10218
rect 9146 10166 9148 10218
rect 9092 10164 9148 10166
rect 9196 10218 9252 10220
rect 9196 10166 9198 10218
rect 9198 10166 9250 10218
rect 9250 10166 9252 10218
rect 9196 10164 9252 10166
rect 9300 10218 9356 10220
rect 9300 10166 9302 10218
rect 9302 10166 9354 10218
rect 9354 10166 9356 10218
rect 9300 10164 9356 10166
rect 9940 10164 9996 10220
rect 8484 9940 8540 9996
rect 8876 9994 8932 9996
rect 8876 9942 8878 9994
rect 8878 9942 8930 9994
rect 8930 9942 8932 9994
rect 8876 9940 8932 9942
rect 11844 12068 11900 12124
rect 10836 11508 10892 11564
rect 11396 12010 11452 12012
rect 11396 11958 11398 12010
rect 11398 11958 11450 12010
rect 11450 11958 11452 12010
rect 11396 11956 11452 11958
rect 11004 11620 11060 11676
rect 11172 11732 11228 11788
rect 11732 11732 11788 11788
rect 13020 12010 13076 12012
rect 13020 11958 13022 12010
rect 13022 11958 13074 12010
rect 13074 11958 13076 12010
rect 13020 11956 13076 11958
rect 13188 11956 13244 12012
rect 12068 11620 12124 11676
rect 11396 11508 11452 11564
rect 11004 11396 11060 11452
rect 10724 10724 10780 10780
rect 10612 10388 10668 10444
rect 10948 10500 11004 10556
rect 10276 9940 10332 9996
rect 11956 11508 12012 11564
rect 12852 11508 12908 11564
rect 11508 11330 11510 11340
rect 11510 11330 11562 11340
rect 11562 11330 11564 11340
rect 11508 11284 11564 11330
rect 12404 10724 12460 10780
rect 13356 11844 13412 11900
rect 14084 12076 14140 12124
rect 14084 12068 14086 12076
rect 14086 12068 14138 12076
rect 14138 12068 14140 12076
rect 15316 12114 15318 12124
rect 15318 12114 15370 12124
rect 15370 12114 15372 12124
rect 15316 12068 15372 12114
rect 15988 12068 16044 12124
rect 14756 11956 14812 12012
rect 14420 11844 14476 11900
rect 13636 11508 13692 11564
rect 13804 11732 13860 11788
rect 13972 11508 14028 11564
rect 8708 9604 8764 9660
rect 9212 9882 9268 9884
rect 9212 9830 9214 9882
rect 9214 9830 9266 9882
rect 9266 9830 9268 9882
rect 9212 9828 9268 9830
rect 8820 9156 8876 9212
rect 9044 9268 9100 9324
rect 8372 9044 8428 9100
rect 8596 9044 8652 9100
rect 10164 9716 10220 9772
rect 9436 9492 9492 9548
rect 9212 9044 9268 9100
rect 10164 9268 10220 9324
rect 10276 9156 10332 9212
rect 7924 8820 7980 8876
rect 8036 8708 8092 8764
rect 3780 8036 3836 8092
rect 4004 7476 4060 7532
rect 4172 7140 4228 7196
rect 4788 8090 4844 8092
rect 4788 8038 4790 8090
rect 4790 8038 4842 8090
rect 4842 8038 4844 8090
rect 4788 8036 4844 8038
rect 7028 8260 7084 8316
rect 4816 7866 4872 7868
rect 4816 7814 4818 7866
rect 4818 7814 4870 7866
rect 4870 7814 4872 7866
rect 4816 7812 4872 7814
rect 4920 7866 4976 7868
rect 4920 7814 4922 7866
rect 4922 7814 4974 7866
rect 4974 7814 4976 7866
rect 4920 7812 4976 7814
rect 5024 7866 5080 7868
rect 5024 7814 5026 7866
rect 5026 7814 5078 7866
rect 5078 7814 5080 7866
rect 5024 7812 5080 7814
rect 5180 7476 5236 7532
rect 4564 7140 4620 7196
rect 3276 6634 3332 6636
rect 3276 6582 3278 6634
rect 3278 6582 3330 6634
rect 3330 6582 3332 6634
rect 3276 6580 3332 6582
rect 4676 7252 4732 7308
rect 5460 7306 5516 7308
rect 5460 7254 5462 7306
rect 5462 7254 5514 7306
rect 5514 7254 5516 7306
rect 5460 7252 5516 7254
rect 6020 7588 6076 7644
rect 6132 8036 6188 8092
rect 7700 8260 7756 8316
rect 7868 8148 7924 8204
rect 8036 8202 8092 8204
rect 8036 8150 8038 8202
rect 8038 8150 8090 8202
rect 8090 8150 8092 8202
rect 8036 8148 8092 8150
rect 6412 7306 6468 7308
rect 6412 7254 6414 7306
rect 6414 7254 6466 7306
rect 6466 7254 6468 7306
rect 6412 7252 6468 7254
rect 7084 7306 7140 7308
rect 7084 7254 7086 7306
rect 7086 7254 7138 7306
rect 7138 7254 7140 7306
rect 7084 7252 7140 7254
rect 6860 7140 6916 7196
rect 7084 6692 7140 6748
rect 4816 6298 4872 6300
rect 4816 6246 4818 6298
rect 4818 6246 4870 6298
rect 4870 6246 4872 6298
rect 4816 6244 4872 6246
rect 4920 6298 4976 6300
rect 4920 6246 4922 6298
rect 4922 6246 4974 6298
rect 4974 6246 4976 6298
rect 4920 6244 4976 6246
rect 5024 6298 5080 6300
rect 5024 6246 5026 6298
rect 5026 6246 5078 6298
rect 5078 6246 5080 6298
rect 5024 6244 5080 6246
rect 7140 6132 7196 6188
rect 6244 6020 6300 6076
rect 6468 5918 6524 5964
rect 6468 5908 6470 5918
rect 6470 5908 6522 5918
rect 6522 5908 6524 5918
rect 6188 5850 6244 5852
rect 6188 5798 6190 5850
rect 6190 5798 6242 5850
rect 6242 5798 6244 5850
rect 6188 5796 6244 5798
rect 2100 4788 2156 4844
rect 1764 4452 1820 4508
rect 1540 3780 1596 3836
rect 5572 5738 5628 5740
rect 5572 5686 5574 5738
rect 5574 5686 5626 5738
rect 5626 5686 5628 5738
rect 5572 5684 5628 5686
rect 6076 5348 6132 5404
rect 5572 5236 5628 5292
rect 5348 5124 5404 5180
rect 2212 4228 2268 4284
rect 4172 3892 4228 3948
rect 1092 2996 1148 3052
rect 2100 2996 2156 3052
rect 2884 2884 2940 2940
rect 3556 2996 3612 3052
rect 3556 2436 3612 2492
rect 4060 3722 4116 3724
rect 4060 3670 4062 3722
rect 4062 3670 4114 3722
rect 4114 3670 4116 3722
rect 4060 3668 4116 3670
rect 4676 4900 4732 4956
rect 5460 4900 5516 4956
rect 4816 4730 4872 4732
rect 4816 4678 4818 4730
rect 4818 4678 4870 4730
rect 4870 4678 4872 4730
rect 4816 4676 4872 4678
rect 4920 4730 4976 4732
rect 4920 4678 4922 4730
rect 4922 4678 4974 4730
rect 4974 4678 4976 4730
rect 4920 4676 4976 4678
rect 5024 4730 5080 4732
rect 5024 4678 5026 4730
rect 5026 4678 5078 4730
rect 5078 4678 5080 4730
rect 5024 4676 5080 4678
rect 4788 4340 4844 4396
rect 5796 4452 5852 4508
rect 6356 5058 6358 5068
rect 6358 5058 6410 5068
rect 6410 5058 6412 5068
rect 6356 5012 6412 5058
rect 7532 7642 7588 7644
rect 7532 7590 7534 7642
rect 7534 7590 7586 7642
rect 7586 7590 7588 7642
rect 7532 7588 7588 7590
rect 7364 6722 7366 6748
rect 7366 6722 7418 6748
rect 7418 6722 7420 6748
rect 7364 6692 7420 6722
rect 7868 7700 7924 7756
rect 7700 6580 7756 6636
rect 6860 5124 6916 5180
rect 7252 5124 7308 5180
rect 6244 4564 6300 4620
rect 5684 4340 5740 4396
rect 4564 3722 4620 3724
rect 4564 3670 4566 3722
rect 4566 3670 4618 3722
rect 4618 3670 4620 3722
rect 4564 3668 4620 3670
rect 5236 4116 5292 4172
rect 5124 3386 5180 3388
rect 5124 3334 5126 3386
rect 5126 3334 5178 3386
rect 5178 3334 5180 3386
rect 5124 3332 5180 3334
rect 4816 3162 4872 3164
rect 4816 3110 4818 3162
rect 4818 3110 4870 3162
rect 4870 3110 4872 3162
rect 4816 3108 4872 3110
rect 4920 3162 4976 3164
rect 4920 3110 4922 3162
rect 4922 3110 4974 3162
rect 4974 3110 4976 3162
rect 4920 3108 4976 3110
rect 5024 3162 5080 3164
rect 5024 3110 5026 3162
rect 5026 3110 5078 3162
rect 5078 3110 5080 3162
rect 5024 3108 5080 3110
rect 5348 2436 5404 2492
rect 6692 4564 6748 4620
rect 6916 4900 6972 4956
rect 6916 4676 6972 4732
rect 6188 3780 6244 3836
rect 7532 5684 7588 5740
rect 8036 5684 8092 5740
rect 8428 8314 8484 8316
rect 8428 8262 8430 8314
rect 8430 8262 8482 8314
rect 8482 8262 8484 8314
rect 8428 8260 8484 8262
rect 8260 8148 8316 8204
rect 8708 8036 8764 8092
rect 9324 8874 9380 8876
rect 9324 8822 9326 8874
rect 9326 8822 9378 8874
rect 9378 8822 9380 8874
rect 9324 8820 9380 8822
rect 9092 8650 9148 8652
rect 9092 8598 9094 8650
rect 9094 8598 9146 8650
rect 9146 8598 9148 8650
rect 9092 8596 9148 8598
rect 9196 8650 9252 8652
rect 9196 8598 9198 8650
rect 9198 8598 9250 8650
rect 9250 8598 9252 8650
rect 9196 8596 9252 8598
rect 9300 8650 9356 8652
rect 9300 8598 9302 8650
rect 9302 8598 9354 8650
rect 9354 8598 9356 8650
rect 9300 8596 9356 8598
rect 9772 8484 9828 8540
rect 11284 9940 11340 9996
rect 13972 11060 14028 11116
rect 13368 11002 13424 11004
rect 13368 10950 13370 11002
rect 13370 10950 13422 11002
rect 13422 10950 13424 11002
rect 13368 10948 13424 10950
rect 13472 11002 13528 11004
rect 13472 10950 13474 11002
rect 13474 10950 13526 11002
rect 13526 10950 13528 11002
rect 13472 10948 13528 10950
rect 13576 11002 13632 11004
rect 13576 10950 13578 11002
rect 13578 10950 13630 11002
rect 13630 10950 13632 11002
rect 13576 10948 13632 10950
rect 13804 10778 13860 10780
rect 13804 10726 13806 10778
rect 13806 10726 13858 10778
rect 13858 10726 13860 10778
rect 13804 10724 13860 10726
rect 14196 11284 14252 11340
rect 14196 11060 14252 11116
rect 14644 10836 14700 10892
rect 14756 11508 14812 11564
rect 14084 10554 14140 10556
rect 14084 10502 14086 10554
rect 14086 10502 14138 10554
rect 14138 10502 14140 10554
rect 14084 10500 14140 10502
rect 21920 12570 21976 12572
rect 21920 12518 21922 12570
rect 21922 12518 21974 12570
rect 21974 12518 21976 12570
rect 21920 12516 21976 12518
rect 22024 12570 22080 12572
rect 22024 12518 22026 12570
rect 22026 12518 22078 12570
rect 22078 12518 22080 12570
rect 22024 12516 22080 12518
rect 22128 12570 22184 12572
rect 22128 12518 22130 12570
rect 22130 12518 22182 12570
rect 22182 12518 22184 12570
rect 22128 12516 22184 12518
rect 18340 12346 18396 12348
rect 18340 12294 18342 12346
rect 18342 12294 18394 12346
rect 18394 12294 18396 12346
rect 18340 12292 18396 12294
rect 21420 12346 21476 12348
rect 21420 12294 21422 12346
rect 21422 12294 21474 12346
rect 21474 12294 21476 12346
rect 21420 12292 21476 12294
rect 18956 12068 19012 12124
rect 22148 12180 22204 12236
rect 28308 12404 28364 12460
rect 18004 11844 18060 11900
rect 17052 11620 17108 11676
rect 16492 11562 16548 11564
rect 16492 11510 16494 11562
rect 16494 11510 16546 11562
rect 16546 11510 16548 11562
rect 16492 11508 16548 11510
rect 17644 11786 17700 11788
rect 17644 11734 17646 11786
rect 17646 11734 17698 11786
rect 17698 11734 17700 11786
rect 17644 11732 17700 11734
rect 17748 11786 17804 11788
rect 17748 11734 17750 11786
rect 17750 11734 17802 11786
rect 17802 11734 17804 11786
rect 17748 11732 17804 11734
rect 17852 11786 17908 11788
rect 17852 11734 17854 11786
rect 17854 11734 17906 11786
rect 17906 11734 17908 11786
rect 17852 11732 17908 11734
rect 17332 11620 17388 11676
rect 16436 11226 16492 11228
rect 16436 11174 16438 11226
rect 16438 11174 16490 11226
rect 16490 11174 16492 11226
rect 16436 11172 16492 11174
rect 14868 10836 14924 10892
rect 14532 10276 14588 10332
rect 13524 9994 13580 9996
rect 13524 9942 13526 9994
rect 13526 9942 13578 9994
rect 13578 9942 13580 9994
rect 13524 9940 13580 9942
rect 12180 9844 12236 9884
rect 10500 8984 10502 8988
rect 10502 8984 10554 8988
rect 10554 8984 10556 8988
rect 10500 8932 10556 8984
rect 9044 8372 9100 8428
rect 10500 8596 10556 8652
rect 9996 8314 10052 8316
rect 8820 7924 8876 7980
rect 9212 7924 9268 7980
rect 9996 8262 9998 8314
rect 9998 8262 10050 8314
rect 10050 8262 10052 8314
rect 9996 8260 10052 8262
rect 9772 8148 9828 8204
rect 9940 8036 9996 8092
rect 9436 7530 9492 7532
rect 9436 7478 9438 7530
rect 9438 7478 9490 7530
rect 9490 7478 9492 7530
rect 9436 7476 9492 7478
rect 10388 7812 10444 7868
rect 10500 8148 10556 8204
rect 10052 7588 10108 7644
rect 11564 9210 11620 9212
rect 11172 9044 11228 9100
rect 11564 9158 11566 9210
rect 11566 9158 11618 9210
rect 11618 9158 11620 9210
rect 11564 9156 11620 9158
rect 12180 9828 12182 9844
rect 12182 9828 12234 9844
rect 12234 9828 12236 9844
rect 11284 8932 11340 8988
rect 12516 9716 12572 9772
rect 11956 9268 12012 9324
rect 12236 9268 12292 9324
rect 11732 8932 11788 8988
rect 12068 8932 12124 8988
rect 10892 8596 10948 8652
rect 12404 8820 12460 8876
rect 12684 9604 12740 9660
rect 12684 9098 12740 9100
rect 12684 9046 12686 9098
rect 12686 9046 12738 9098
rect 12738 9046 12740 9098
rect 12684 9044 12740 9046
rect 14980 10724 15036 10780
rect 14868 10276 14924 10332
rect 15484 10276 15540 10332
rect 14308 9940 14364 9996
rect 14532 9828 14588 9884
rect 13132 9658 13188 9660
rect 13132 9606 13134 9658
rect 13134 9606 13186 9658
rect 13186 9606 13188 9658
rect 13132 9604 13188 9606
rect 12908 9210 12964 9212
rect 12908 9158 12910 9210
rect 12910 9158 12962 9210
rect 12962 9158 12964 9210
rect 12908 9156 12964 9158
rect 13132 9380 13188 9436
rect 13368 9434 13424 9436
rect 13368 9382 13370 9434
rect 13370 9382 13422 9434
rect 13422 9382 13424 9434
rect 13368 9380 13424 9382
rect 13472 9434 13528 9436
rect 13472 9382 13474 9434
rect 13474 9382 13526 9434
rect 13526 9382 13528 9434
rect 13472 9380 13528 9382
rect 13576 9434 13632 9436
rect 13576 9382 13578 9434
rect 13578 9382 13630 9434
rect 13630 9382 13632 9434
rect 13576 9380 13632 9382
rect 13916 9268 13972 9324
rect 14308 9604 14364 9660
rect 11340 8484 11396 8540
rect 10612 8260 10668 8316
rect 10612 7924 10668 7980
rect 10948 8314 11004 8316
rect 10948 8262 10950 8314
rect 10950 8262 11002 8314
rect 11002 8262 11004 8314
rect 12068 8484 12124 8540
rect 12236 8484 12292 8540
rect 10948 8260 11004 8262
rect 10948 7588 11004 7644
rect 8596 7372 8652 7420
rect 8596 7364 8598 7372
rect 8598 7364 8650 7372
rect 8650 7364 8652 7372
rect 9660 7418 9716 7420
rect 9660 7366 9662 7418
rect 9662 7366 9714 7418
rect 9714 7366 9716 7418
rect 9660 7364 9716 7366
rect 10388 7364 10444 7420
rect 9940 7140 9996 7196
rect 9092 7082 9148 7084
rect 9092 7030 9094 7082
rect 9094 7030 9146 7082
rect 9146 7030 9148 7082
rect 9092 7028 9148 7030
rect 9196 7082 9252 7084
rect 9196 7030 9198 7082
rect 9198 7030 9250 7082
rect 9250 7030 9252 7082
rect 9196 7028 9252 7030
rect 9300 7082 9356 7084
rect 9300 7030 9302 7082
rect 9302 7030 9354 7082
rect 9354 7030 9356 7082
rect 9300 7028 9356 7030
rect 9716 6692 9772 6748
rect 7700 5236 7756 5292
rect 7812 4954 7868 4956
rect 7812 4902 7814 4954
rect 7814 4902 7866 4954
rect 7866 4902 7868 4954
rect 7812 4900 7868 4902
rect 7364 4506 7420 4508
rect 7364 4454 7366 4506
rect 7366 4454 7418 4506
rect 7418 4454 7420 4506
rect 7364 4452 7420 4454
rect 7588 4452 7644 4508
rect 7252 4340 7308 4396
rect 8316 5236 8372 5292
rect 8596 6580 8652 6636
rect 9044 6020 9100 6076
rect 9716 6356 9772 6412
rect 8708 5961 8710 5964
rect 8710 5961 8762 5964
rect 8762 5961 8764 5964
rect 8708 5908 8764 5961
rect 9156 5796 9212 5852
rect 8764 5738 8820 5740
rect 8764 5686 8766 5738
rect 8766 5686 8818 5738
rect 8818 5686 8820 5738
rect 8764 5684 8820 5686
rect 9380 5684 9436 5740
rect 9092 5514 9148 5516
rect 9092 5462 9094 5514
rect 9094 5462 9146 5514
rect 9146 5462 9148 5514
rect 9092 5460 9148 5462
rect 9196 5514 9252 5516
rect 9196 5462 9198 5514
rect 9198 5462 9250 5514
rect 9250 5462 9252 5514
rect 9196 5460 9252 5462
rect 9300 5514 9356 5516
rect 9300 5462 9302 5514
rect 9302 5462 9354 5514
rect 9354 5462 9356 5514
rect 9300 5460 9356 5462
rect 8652 5178 8708 5180
rect 8652 5126 8654 5178
rect 8654 5126 8706 5178
rect 8706 5126 8708 5178
rect 8652 5124 8708 5126
rect 8484 5012 8540 5068
rect 8372 4900 8428 4956
rect 8260 4676 8316 4732
rect 8036 4452 8092 4508
rect 8260 4452 8316 4508
rect 7924 4228 7980 4284
rect 6860 3498 6916 3500
rect 6860 3446 6862 3498
rect 6862 3446 6914 3498
rect 6914 3446 6916 3498
rect 6860 3444 6916 3446
rect 5852 3332 5908 3388
rect 6244 2824 6246 2828
rect 6246 2824 6298 2828
rect 6298 2824 6300 2828
rect 6244 2772 6300 2824
rect 7028 3108 7084 3164
rect 7084 2938 7140 2940
rect 7084 2886 7086 2938
rect 7086 2886 7138 2938
rect 7138 2886 7140 2938
rect 7084 2884 7140 2886
rect 5852 2714 5908 2716
rect 5852 2662 5854 2714
rect 5854 2662 5906 2714
rect 5906 2662 5908 2714
rect 5852 2660 5908 2662
rect 6468 2660 6524 2716
rect 6692 2660 6748 2716
rect 5460 2100 5516 2156
rect 3892 1876 3948 1932
rect 4732 1930 4788 1932
rect 4732 1878 4734 1930
rect 4734 1878 4786 1930
rect 4786 1878 4788 1930
rect 4732 1876 4788 1878
rect 5180 1930 5236 1932
rect 5180 1878 5182 1930
rect 5182 1878 5234 1930
rect 5234 1878 5236 1930
rect 5180 1876 5236 1878
rect 4564 1818 4620 1820
rect 4564 1766 4566 1818
rect 4566 1766 4618 1818
rect 4618 1766 4620 1818
rect 4564 1764 4620 1766
rect 5180 1652 5236 1708
rect 4816 1594 4872 1596
rect 4816 1542 4818 1594
rect 4818 1542 4870 1594
rect 4870 1542 4872 1594
rect 4816 1540 4872 1542
rect 4920 1594 4976 1596
rect 4920 1542 4922 1594
rect 4922 1542 4974 1594
rect 4974 1542 4976 1594
rect 4920 1540 4976 1542
rect 5024 1594 5080 1596
rect 5024 1542 5026 1594
rect 5026 1542 5078 1594
rect 5078 1542 5080 1594
rect 5024 1540 5080 1542
rect 7364 3220 7420 3276
rect 7588 3892 7644 3948
rect 7476 3108 7532 3164
rect 7476 2884 7532 2940
rect 7588 2548 7644 2604
rect 7700 3108 7756 3164
rect 6916 2127 6918 2156
rect 6918 2127 6970 2156
rect 6970 2127 6972 2156
rect 7980 3444 8036 3500
rect 11340 7924 11396 7980
rect 11900 8314 11956 8316
rect 11900 8262 11902 8314
rect 11902 8262 11954 8314
rect 11954 8262 11956 8314
rect 11900 8260 11956 8262
rect 12236 8148 12292 8204
rect 12404 8202 12460 8204
rect 12404 8150 12406 8202
rect 12406 8150 12458 8202
rect 12458 8150 12460 8202
rect 12404 8148 12460 8150
rect 11620 7924 11676 7980
rect 12068 7924 12124 7980
rect 11732 7812 11788 7868
rect 11956 7812 12012 7868
rect 11172 7476 11228 7532
rect 11060 7252 11116 7308
rect 12628 8372 12684 8428
rect 12516 7812 12572 7868
rect 13188 8260 13244 8316
rect 11396 6746 11452 6748
rect 11396 6694 11398 6746
rect 11398 6694 11450 6746
rect 11450 6694 11452 6746
rect 11396 6692 11452 6694
rect 12572 6634 12628 6636
rect 12572 6582 12574 6634
rect 12574 6582 12626 6634
rect 12626 6582 12628 6634
rect 12572 6580 12628 6582
rect 11676 5572 11732 5628
rect 10108 5460 10164 5516
rect 9268 5178 9324 5180
rect 9268 5126 9270 5178
rect 9270 5126 9322 5178
rect 9322 5126 9324 5178
rect 9268 5124 9324 5126
rect 8708 4788 8764 4844
rect 8596 4676 8652 4732
rect 8932 4676 8988 4732
rect 8484 4004 8540 4060
rect 8708 3444 8764 3500
rect 9044 4452 9100 4508
rect 8820 3220 8876 3276
rect 7812 2548 7868 2604
rect 7700 2212 7756 2268
rect 6916 2100 6972 2127
rect 7812 2100 7868 2156
rect 7644 2042 7700 2044
rect 7644 1990 7646 2042
rect 7646 1990 7698 2042
rect 7698 1990 7700 2042
rect 7644 1988 7700 1990
rect 6244 1764 6300 1820
rect 5628 1652 5684 1708
rect 8036 2668 8092 2716
rect 8036 2660 8038 2668
rect 8038 2660 8090 2668
rect 8090 2660 8092 2668
rect 9884 5290 9940 5292
rect 9884 5238 9886 5290
rect 9886 5238 9938 5290
rect 9938 5238 9940 5290
rect 10836 5348 10892 5404
rect 9884 5236 9940 5238
rect 9996 5178 10052 5180
rect 9996 5126 9998 5178
rect 9998 5126 10050 5178
rect 10050 5126 10052 5178
rect 9996 5124 10052 5126
rect 10164 5012 10220 5068
rect 10388 5124 10444 5180
rect 10052 4788 10108 4844
rect 9380 4676 9436 4732
rect 9940 4676 9996 4732
rect 9492 4350 9548 4396
rect 9492 4340 9494 4350
rect 9494 4340 9546 4350
rect 9546 4340 9548 4350
rect 9268 4274 9270 4284
rect 9270 4274 9322 4284
rect 9322 4274 9324 4284
rect 9268 4228 9324 4274
rect 10388 4676 10444 4732
rect 10052 4340 10108 4396
rect 9092 3946 9148 3948
rect 9092 3894 9094 3946
rect 9094 3894 9146 3946
rect 9146 3894 9148 3946
rect 9092 3892 9148 3894
rect 9196 3946 9252 3948
rect 9196 3894 9198 3946
rect 9198 3894 9250 3946
rect 9250 3894 9252 3946
rect 9196 3892 9252 3894
rect 9300 3946 9356 3948
rect 9300 3894 9302 3946
rect 9302 3894 9354 3946
rect 9354 3894 9356 3946
rect 9300 3892 9356 3894
rect 9940 4004 9996 4060
rect 9828 3892 9884 3948
rect 11060 5012 11116 5068
rect 12852 7364 12908 7420
rect 12740 6244 12796 6300
rect 12852 6356 12908 6412
rect 12516 5908 12572 5964
rect 12180 5290 12236 5292
rect 12180 5238 12182 5290
rect 12182 5238 12234 5290
rect 12234 5238 12236 5290
rect 12180 5236 12236 5238
rect 12292 5151 12348 5180
rect 12292 5124 12294 5151
rect 12294 5124 12346 5151
rect 12346 5124 12348 5151
rect 12404 5012 12460 5068
rect 11900 4954 11956 4956
rect 11900 4902 11902 4954
rect 11902 4902 11954 4954
rect 11954 4902 11956 4954
rect 11900 4900 11956 4902
rect 11228 4676 11284 4732
rect 11732 4676 11788 4732
rect 10500 4564 10556 4620
rect 11508 4564 11564 4620
rect 11172 4506 11228 4508
rect 11172 4454 11174 4506
rect 11174 4454 11226 4506
rect 11226 4454 11228 4506
rect 11172 4452 11228 4454
rect 10500 4170 10556 4172
rect 10500 4118 10502 4170
rect 10502 4118 10554 4170
rect 10554 4118 10556 4170
rect 10500 4116 10556 4118
rect 10948 3892 11004 3948
rect 12068 4564 12124 4620
rect 13356 8314 13412 8316
rect 13356 8262 13358 8314
rect 13358 8262 13410 8314
rect 13410 8262 13412 8314
rect 13356 8260 13412 8262
rect 14308 8932 14364 8988
rect 14084 8820 14140 8876
rect 13748 8484 13804 8540
rect 14868 9838 14924 9884
rect 14868 9828 14870 9838
rect 14870 9828 14922 9838
rect 14922 9828 14924 9838
rect 16324 10612 16380 10668
rect 16380 10276 16436 10332
rect 15876 10164 15932 10220
rect 14644 9762 14646 9772
rect 14646 9762 14698 9772
rect 14698 9762 14700 9772
rect 14644 9716 14700 9762
rect 15092 9604 15148 9660
rect 15260 9380 15316 9436
rect 15428 9156 15484 9212
rect 13804 8314 13860 8316
rect 13804 8262 13806 8314
rect 13806 8262 13858 8314
rect 13858 8262 13860 8314
rect 13804 8260 13860 8262
rect 13524 8036 13580 8092
rect 14196 8260 14252 8316
rect 13368 7866 13424 7868
rect 13368 7814 13370 7866
rect 13370 7814 13422 7866
rect 13422 7814 13424 7866
rect 13368 7812 13424 7814
rect 13472 7866 13528 7868
rect 13472 7814 13474 7866
rect 13474 7814 13526 7866
rect 13526 7814 13528 7866
rect 13472 7812 13528 7814
rect 13576 7866 13632 7868
rect 13576 7814 13578 7866
rect 13578 7814 13630 7866
rect 13630 7814 13632 7866
rect 13576 7812 13632 7814
rect 13916 7700 13972 7756
rect 14084 8036 14140 8092
rect 15764 8874 15820 8876
rect 15764 8822 15766 8874
rect 15766 8822 15818 8874
rect 15818 8822 15820 8874
rect 15764 8820 15820 8822
rect 15652 8372 15708 8428
rect 14924 8148 14980 8204
rect 14196 7700 14252 7756
rect 14308 8036 14364 8092
rect 14084 7588 14140 7644
rect 13916 7476 13972 7532
rect 14196 7476 14252 7532
rect 14588 7812 14644 7868
rect 14644 7140 14700 7196
rect 15092 8090 15148 8092
rect 15092 8038 15094 8090
rect 15094 8038 15146 8090
rect 15146 8038 15148 8090
rect 15092 8036 15148 8038
rect 15204 7588 15260 7644
rect 15316 7486 15372 7532
rect 15316 7476 15318 7486
rect 15318 7476 15370 7486
rect 15370 7476 15372 7486
rect 13580 6858 13636 6860
rect 13580 6806 13582 6858
rect 13582 6806 13634 6858
rect 13634 6806 13636 6858
rect 13580 6804 13636 6806
rect 13076 6746 13132 6748
rect 13076 6694 13078 6746
rect 13078 6694 13130 6746
rect 13130 6694 13132 6746
rect 13076 6692 13132 6694
rect 13076 6468 13132 6524
rect 13188 6244 13244 6300
rect 12964 5796 13020 5852
rect 13076 6020 13132 6076
rect 13368 6298 13424 6300
rect 13368 6246 13370 6298
rect 13370 6246 13422 6298
rect 13422 6246 13424 6298
rect 13368 6244 13424 6246
rect 13472 6298 13528 6300
rect 13472 6246 13474 6298
rect 13474 6246 13526 6298
rect 13526 6246 13528 6298
rect 13472 6244 13528 6246
rect 13576 6298 13632 6300
rect 13576 6246 13578 6298
rect 13578 6246 13630 6298
rect 13630 6246 13632 6298
rect 13576 6244 13632 6246
rect 13748 5908 13804 5964
rect 14084 6746 14140 6748
rect 14084 6694 14086 6746
rect 14086 6694 14138 6746
rect 14138 6694 14140 6746
rect 14084 6692 14140 6694
rect 14084 6468 14140 6524
rect 13972 6074 14028 6076
rect 13972 6022 13974 6074
rect 13974 6022 14026 6074
rect 14026 6022 14028 6074
rect 13972 6020 14028 6022
rect 16884 10052 16940 10108
rect 17052 10836 17108 10892
rect 16380 9882 16436 9884
rect 16380 9830 16382 9882
rect 16382 9830 16434 9882
rect 16434 9830 16436 9882
rect 16380 9828 16436 9830
rect 17444 11396 17500 11452
rect 17892 11508 17948 11564
rect 19740 11732 19796 11788
rect 19404 11508 19460 11564
rect 18788 11450 18844 11452
rect 18788 11398 18790 11450
rect 18790 11398 18842 11450
rect 18842 11398 18844 11450
rect 18788 11396 18844 11398
rect 19292 11450 19348 11452
rect 19292 11398 19294 11450
rect 19294 11398 19346 11450
rect 19346 11398 19348 11450
rect 19292 11396 19348 11398
rect 20020 11450 20076 11452
rect 20020 11398 20022 11450
rect 20022 11398 20074 11450
rect 20074 11398 20076 11450
rect 20020 11396 20076 11398
rect 24164 12190 24220 12236
rect 24164 12180 24166 12190
rect 24166 12180 24218 12190
rect 24218 12180 24220 12190
rect 30472 12570 30528 12572
rect 30472 12518 30474 12570
rect 30474 12518 30526 12570
rect 30526 12518 30528 12570
rect 30472 12516 30528 12518
rect 30576 12570 30632 12572
rect 30576 12518 30578 12570
rect 30578 12518 30630 12570
rect 30630 12518 30632 12570
rect 30576 12516 30632 12518
rect 30680 12570 30736 12572
rect 30680 12518 30682 12570
rect 30682 12518 30734 12570
rect 30734 12518 30736 12570
rect 30680 12516 30736 12518
rect 32676 12180 32732 12236
rect 22148 12010 22150 12012
rect 22150 12010 22202 12012
rect 22202 12010 22204 12012
rect 22148 11956 22204 12010
rect 21812 11844 21868 11900
rect 20132 11396 20188 11452
rect 20916 11396 20972 11452
rect 17444 10836 17500 10892
rect 17780 10666 17836 10668
rect 17780 10614 17782 10666
rect 17782 10614 17834 10666
rect 17834 10614 17836 10666
rect 17780 10612 17836 10614
rect 17332 10388 17388 10444
rect 17444 10276 17500 10332
rect 17644 10218 17700 10220
rect 17644 10166 17646 10218
rect 17646 10166 17698 10218
rect 17698 10166 17700 10218
rect 17644 10164 17700 10166
rect 17748 10218 17804 10220
rect 17748 10166 17750 10218
rect 17750 10166 17802 10218
rect 17802 10166 17804 10218
rect 17748 10164 17804 10166
rect 17852 10218 17908 10220
rect 17852 10166 17854 10218
rect 17854 10166 17906 10218
rect 17906 10166 17908 10218
rect 17852 10164 17908 10166
rect 17668 9940 17724 9996
rect 17052 9828 17108 9884
rect 16940 9770 16996 9772
rect 16940 9718 16942 9770
rect 16942 9718 16994 9770
rect 16994 9718 16996 9770
rect 16940 9716 16996 9718
rect 17108 9210 17164 9212
rect 17108 9158 17110 9210
rect 17110 9158 17162 9210
rect 17162 9158 17164 9210
rect 17108 9156 17164 9158
rect 17836 9882 17892 9884
rect 17836 9830 17838 9882
rect 17838 9830 17890 9882
rect 17890 9830 17892 9882
rect 17836 9828 17892 9830
rect 17668 9492 17724 9548
rect 17556 9380 17612 9436
rect 19628 10724 19684 10780
rect 19796 11172 19852 11228
rect 18452 10500 18508 10556
rect 18340 9940 18396 9996
rect 18060 9882 18116 9884
rect 18060 9830 18062 9882
rect 18062 9830 18114 9882
rect 18114 9830 18116 9882
rect 18060 9828 18116 9830
rect 18452 9882 18508 9884
rect 18452 9830 18454 9882
rect 18454 9830 18506 9882
rect 18506 9830 18508 9882
rect 18452 9828 18508 9830
rect 17892 9380 17948 9436
rect 16324 9054 16380 9100
rect 16324 9044 16326 9054
rect 16326 9044 16378 9054
rect 16378 9044 16380 9054
rect 17220 9044 17276 9100
rect 15540 7588 15596 7644
rect 14588 6356 14644 6412
rect 16436 8932 16492 8988
rect 16548 8820 16604 8876
rect 15988 8148 16044 8204
rect 15988 7476 16044 7532
rect 16100 8260 16156 8316
rect 16660 8708 16716 8764
rect 17444 8986 17500 8988
rect 17444 8934 17446 8986
rect 17446 8934 17498 8986
rect 17498 8934 17500 8986
rect 17444 8932 17500 8934
rect 18004 9268 18060 9324
rect 18284 9604 18340 9660
rect 17892 8820 17948 8876
rect 16940 8708 16996 8764
rect 18340 8874 18396 8876
rect 18340 8822 18342 8874
rect 18342 8822 18394 8874
rect 18394 8822 18396 8874
rect 18340 8820 18396 8822
rect 18844 8874 18900 8876
rect 18844 8822 18846 8874
rect 18846 8822 18898 8874
rect 18898 8822 18900 8874
rect 18844 8820 18900 8822
rect 18060 8708 18116 8764
rect 17644 8650 17700 8652
rect 17644 8598 17646 8650
rect 17646 8598 17698 8650
rect 17698 8598 17700 8650
rect 17644 8596 17700 8598
rect 17748 8650 17804 8652
rect 17748 8598 17750 8650
rect 17750 8598 17802 8650
rect 17802 8598 17804 8650
rect 17748 8596 17804 8598
rect 17852 8650 17908 8652
rect 17852 8598 17854 8650
rect 17854 8598 17906 8650
rect 17906 8598 17908 8650
rect 17852 8596 17908 8598
rect 17332 8260 17388 8316
rect 17444 8484 17500 8540
rect 17220 7812 17276 7868
rect 16100 7140 16156 7196
rect 16660 7476 16716 7532
rect 15876 6356 15932 6412
rect 13188 5796 13244 5852
rect 13636 5796 13692 5852
rect 14644 5914 14700 5964
rect 14644 5908 14646 5914
rect 14646 5908 14698 5914
rect 14698 5908 14700 5914
rect 14420 5850 14476 5852
rect 13804 5684 13860 5740
rect 14420 5798 14422 5850
rect 14422 5798 14474 5850
rect 14474 5798 14476 5850
rect 14420 5796 14476 5798
rect 13804 5236 13860 5292
rect 13412 4954 13468 4956
rect 13412 4902 13414 4954
rect 13414 4902 13466 4954
rect 13466 4902 13468 4954
rect 13412 4900 13468 4902
rect 13368 4730 13424 4732
rect 13368 4678 13370 4730
rect 13370 4678 13422 4730
rect 13422 4678 13424 4730
rect 13368 4676 13424 4678
rect 13472 4730 13528 4732
rect 13472 4678 13474 4730
rect 13474 4678 13526 4730
rect 13526 4678 13528 4730
rect 13472 4676 13528 4678
rect 13576 4730 13632 4732
rect 13576 4678 13578 4730
rect 13578 4678 13630 4730
rect 13630 4678 13632 4730
rect 13576 4676 13632 4678
rect 14308 5058 14310 5068
rect 14310 5058 14362 5068
rect 14362 5058 14364 5068
rect 14308 5012 14364 5058
rect 16324 6468 16380 6524
rect 16212 5796 16268 5852
rect 15988 5684 16044 5740
rect 17220 6804 17276 6860
rect 17332 7364 17388 7420
rect 15204 4900 15260 4956
rect 16660 6356 16716 6412
rect 17892 8372 17948 8428
rect 17556 7390 17612 7420
rect 17556 7364 17558 7390
rect 17558 7364 17610 7390
rect 17610 7364 17612 7390
rect 18508 7642 18564 7644
rect 18508 7590 18510 7642
rect 18510 7590 18562 7642
rect 18562 7590 18564 7642
rect 18508 7588 18564 7590
rect 18676 7364 18732 7420
rect 17644 7082 17700 7084
rect 17644 7030 17646 7082
rect 17646 7030 17698 7082
rect 17698 7030 17700 7082
rect 17644 7028 17700 7030
rect 17748 7082 17804 7084
rect 17748 7030 17750 7082
rect 17750 7030 17802 7082
rect 17802 7030 17804 7082
rect 17748 7028 17804 7030
rect 17852 7082 17908 7084
rect 17852 7030 17854 7082
rect 17854 7030 17906 7082
rect 17906 7030 17908 7082
rect 17852 7028 17908 7030
rect 17444 6580 17500 6636
rect 18844 7140 18900 7196
rect 18004 6468 18060 6524
rect 18396 6468 18452 6524
rect 23940 11844 23996 11900
rect 21588 11172 21644 11228
rect 22708 11060 22764 11116
rect 21920 11002 21976 11004
rect 21920 10950 21922 11002
rect 21922 10950 21974 11002
rect 21974 10950 21976 11002
rect 21920 10948 21976 10950
rect 22024 11002 22080 11004
rect 22024 10950 22026 11002
rect 22026 10950 22078 11002
rect 22078 10950 22080 11002
rect 22024 10948 22080 10950
rect 22128 11002 22184 11004
rect 22128 10950 22130 11002
rect 22130 10950 22182 11002
rect 22182 10950 22184 11002
rect 22128 10948 22184 10950
rect 21812 10724 21868 10780
rect 22036 10622 22092 10668
rect 22036 10612 22038 10622
rect 22038 10612 22090 10622
rect 22090 10612 22092 10622
rect 22708 10612 22764 10668
rect 19684 10442 19740 10444
rect 19684 10390 19686 10442
rect 19686 10390 19738 10442
rect 19738 10390 19740 10442
rect 19684 10388 19740 10390
rect 22596 10546 22598 10556
rect 22598 10546 22650 10556
rect 22650 10546 22652 10556
rect 22596 10500 22652 10546
rect 21588 10276 21644 10332
rect 19684 10052 19740 10108
rect 19460 9994 19516 9996
rect 19460 9942 19462 9994
rect 19462 9942 19514 9994
rect 19514 9942 19516 9994
rect 19460 9940 19516 9942
rect 20076 9994 20132 9996
rect 20076 9942 20078 9994
rect 20078 9942 20130 9994
rect 20130 9942 20132 9994
rect 20076 9940 20132 9942
rect 19908 9716 19964 9772
rect 19348 8260 19404 8316
rect 19124 7924 19180 7980
rect 19124 7700 19180 7756
rect 19908 9044 19964 9100
rect 20244 8874 20300 8876
rect 20244 8822 20246 8874
rect 20246 8822 20298 8874
rect 20298 8822 20300 8874
rect 20244 8820 20300 8822
rect 20748 8986 20804 8988
rect 20748 8934 20750 8986
rect 20750 8934 20802 8986
rect 20802 8934 20804 8986
rect 20748 8932 20804 8934
rect 20580 8372 20636 8428
rect 20020 8036 20076 8092
rect 19572 7588 19628 7644
rect 19684 7924 19740 7980
rect 19348 7252 19404 7308
rect 19012 6804 19068 6860
rect 17444 6356 17500 6412
rect 13748 4564 13804 4620
rect 15260 4676 15316 4732
rect 13020 4506 13076 4508
rect 13020 4454 13022 4506
rect 13022 4454 13074 4506
rect 13074 4454 13076 4506
rect 13020 4452 13076 4454
rect 13300 4452 13356 4508
rect 12348 4228 12404 4284
rect 13468 4506 13524 4508
rect 13468 4454 13470 4506
rect 13470 4454 13522 4506
rect 13522 4454 13524 4506
rect 13468 4452 13524 4454
rect 14756 4452 14812 4508
rect 11900 4170 11956 4172
rect 11900 4118 11902 4170
rect 11902 4118 11954 4170
rect 11954 4118 11956 4170
rect 11900 4116 11956 4118
rect 12124 4170 12180 4172
rect 12124 4118 12126 4170
rect 12126 4118 12178 4170
rect 12178 4118 12180 4170
rect 12124 4116 12180 4118
rect 12068 3892 12124 3948
rect 9548 3780 9604 3836
rect 9044 3668 9100 3724
rect 11620 3780 11676 3836
rect 8596 2996 8652 3052
rect 8372 2884 8428 2940
rect 8260 2212 8316 2268
rect 9044 3108 9100 3164
rect 9940 3610 9996 3612
rect 9940 3558 9942 3610
rect 9942 3558 9994 3610
rect 9994 3558 9996 3610
rect 9940 3556 9996 3558
rect 10276 3556 10332 3612
rect 9492 3444 9548 3500
rect 9716 3444 9772 3500
rect 9156 2996 9212 3052
rect 9604 3220 9660 3276
rect 9268 2782 9324 2828
rect 9268 2772 9270 2782
rect 9270 2772 9322 2782
rect 9322 2772 9324 2782
rect 9092 2378 9148 2380
rect 9092 2326 9094 2378
rect 9094 2326 9146 2378
rect 9146 2326 9148 2378
rect 9092 2324 9148 2326
rect 9196 2378 9252 2380
rect 9196 2326 9198 2378
rect 9198 2326 9250 2378
rect 9250 2326 9252 2378
rect 9196 2324 9252 2326
rect 9300 2378 9356 2380
rect 9300 2326 9302 2378
rect 9302 2326 9354 2378
rect 9354 2326 9356 2378
rect 9300 2324 9356 2326
rect 8596 2212 8652 2268
rect 10164 2212 10220 2268
rect 10724 3448 10780 3500
rect 10724 3444 10726 3448
rect 10726 3444 10778 3448
rect 10778 3444 10780 3448
rect 11396 3556 11452 3612
rect 11508 3444 11564 3500
rect 11116 3332 11172 3388
rect 12628 4170 12684 4172
rect 12628 4118 12630 4170
rect 12630 4118 12682 4170
rect 12682 4118 12684 4170
rect 12628 4116 12684 4118
rect 13860 4340 13916 4396
rect 14644 4340 14700 4396
rect 13132 4116 13188 4172
rect 13524 4116 13580 4172
rect 13524 3780 13580 3836
rect 11844 3444 11900 3500
rect 11956 3332 12012 3388
rect 10948 2884 11004 2940
rect 11396 2548 11452 2604
rect 10724 2212 10780 2268
rect 8988 2042 9044 2044
rect 8988 1990 8990 2042
rect 8990 1990 9042 2042
rect 9042 1990 9044 2042
rect 8988 1988 9044 1990
rect 12068 2324 12124 2380
rect 12460 3386 12516 3388
rect 12460 3334 12462 3386
rect 12462 3334 12514 3386
rect 12514 3334 12516 3386
rect 12460 3332 12516 3334
rect 14420 3780 14476 3836
rect 13804 3610 13860 3612
rect 13804 3558 13806 3610
rect 13806 3558 13858 3610
rect 13858 3558 13860 3610
rect 13804 3556 13860 3558
rect 13860 3386 13916 3388
rect 13860 3334 13862 3386
rect 13862 3334 13914 3386
rect 13914 3334 13916 3386
rect 13860 3332 13916 3334
rect 14196 3556 14252 3612
rect 12964 2996 13020 3052
rect 12292 2884 12348 2940
rect 12740 2938 12796 2940
rect 12740 2886 12742 2938
rect 12742 2886 12794 2938
rect 12794 2886 12796 2938
rect 12740 2884 12796 2886
rect 12964 2772 13020 2828
rect 12516 2660 12572 2716
rect 12404 2436 12460 2492
rect 8596 1930 8652 1932
rect 8596 1878 8598 1930
rect 8598 1878 8650 1930
rect 8650 1878 8652 1930
rect 8596 1876 8652 1878
rect 9324 1652 9380 1708
rect 13188 3108 13244 3164
rect 13368 3162 13424 3164
rect 13368 3110 13370 3162
rect 13370 3110 13422 3162
rect 13422 3110 13424 3162
rect 13368 3108 13424 3110
rect 13472 3162 13528 3164
rect 13472 3110 13474 3162
rect 13474 3110 13526 3162
rect 13526 3110 13528 3162
rect 13472 3108 13528 3110
rect 13576 3162 13632 3164
rect 13576 3110 13578 3162
rect 13578 3110 13630 3162
rect 13630 3110 13632 3162
rect 13576 3108 13632 3110
rect 13356 2938 13412 2940
rect 13356 2886 13358 2938
rect 13358 2886 13410 2938
rect 13410 2886 13412 2938
rect 13356 2884 13412 2886
rect 13076 2660 13132 2716
rect 13580 2660 13636 2716
rect 13188 2548 13244 2604
rect 14084 2660 14140 2716
rect 13972 2602 14028 2604
rect 13972 2550 13974 2602
rect 13974 2550 14026 2602
rect 14026 2550 14028 2602
rect 13972 2548 14028 2550
rect 13300 2100 13356 2156
rect 14308 3220 14364 3276
rect 15092 4340 15148 4396
rect 14924 4004 14980 4060
rect 17644 5514 17700 5516
rect 17644 5462 17646 5514
rect 17646 5462 17698 5514
rect 17698 5462 17700 5514
rect 17644 5460 17700 5462
rect 17748 5514 17804 5516
rect 17748 5462 17750 5514
rect 17750 5462 17802 5514
rect 17802 5462 17804 5514
rect 17748 5460 17804 5462
rect 17852 5514 17908 5516
rect 17852 5462 17854 5514
rect 17854 5462 17906 5514
rect 17906 5462 17908 5514
rect 17852 5460 17908 5462
rect 18620 6356 18676 6412
rect 19572 6692 19628 6748
rect 20916 8708 20972 8764
rect 21476 9716 21532 9772
rect 22428 9994 22484 9996
rect 22428 9942 22430 9994
rect 22430 9942 22482 9994
rect 22482 9942 22484 9994
rect 22428 9940 22484 9942
rect 22036 9604 22092 9660
rect 22596 9828 22652 9884
rect 21700 9492 21756 9548
rect 21920 9434 21976 9436
rect 21920 9382 21922 9434
rect 21922 9382 21974 9434
rect 21974 9382 21976 9434
rect 21920 9380 21976 9382
rect 22024 9434 22080 9436
rect 22024 9382 22026 9434
rect 22026 9382 22078 9434
rect 22078 9382 22080 9434
rect 22024 9380 22080 9382
rect 22128 9434 22184 9436
rect 22128 9382 22130 9434
rect 22130 9382 22182 9434
rect 22182 9382 22184 9434
rect 22128 9380 22184 9382
rect 22148 8982 22150 8988
rect 22150 8982 22202 8988
rect 22202 8982 22204 8988
rect 22148 8932 22204 8982
rect 21644 8874 21700 8876
rect 21644 8822 21646 8874
rect 21646 8822 21698 8874
rect 21698 8822 21700 8874
rect 21644 8820 21700 8822
rect 21028 8372 21084 8428
rect 20244 7924 20300 7980
rect 21196 8314 21252 8316
rect 21196 8262 21198 8314
rect 21198 8262 21250 8314
rect 21250 8262 21252 8314
rect 21196 8260 21252 8262
rect 20804 8148 20860 8204
rect 20580 7924 20636 7980
rect 20020 7140 20076 7196
rect 21364 7476 21420 7532
rect 20132 6746 20188 6748
rect 20132 6694 20134 6746
rect 20134 6694 20186 6746
rect 20186 6694 20188 6746
rect 20132 6692 20188 6694
rect 19404 6634 19460 6636
rect 19404 6582 19406 6634
rect 19406 6582 19458 6634
rect 19458 6582 19460 6634
rect 19404 6580 19460 6582
rect 21476 8484 21532 8540
rect 22372 9658 22428 9660
rect 22372 9606 22374 9658
rect 22374 9606 22426 9658
rect 22426 9606 22428 9658
rect 22372 9604 22428 9606
rect 22820 10442 22876 10444
rect 22820 10390 22822 10442
rect 22822 10390 22874 10442
rect 22874 10390 22876 10442
rect 22820 10388 22876 10390
rect 22708 9044 22764 9100
rect 24500 11508 24556 11564
rect 25396 12114 25398 12124
rect 25398 12114 25450 12124
rect 25450 12114 25452 12124
rect 25396 12068 25452 12114
rect 26068 11844 26124 11900
rect 24724 11396 24780 11452
rect 23940 11330 23942 11340
rect 23942 11330 23994 11340
rect 23994 11330 23996 11340
rect 23940 11284 23996 11330
rect 26196 11786 26252 11788
rect 26196 11734 26198 11786
rect 26198 11734 26250 11786
rect 26250 11734 26252 11786
rect 26196 11732 26252 11734
rect 26300 11786 26356 11788
rect 26300 11734 26302 11786
rect 26302 11734 26354 11786
rect 26354 11734 26356 11786
rect 26300 11732 26356 11734
rect 26404 11786 26460 11788
rect 26404 11734 26406 11786
rect 26406 11734 26458 11786
rect 26458 11734 26460 11786
rect 26404 11732 26460 11734
rect 24724 10836 24780 10892
rect 23492 10388 23548 10444
rect 22988 9770 23044 9772
rect 22988 9718 22990 9770
rect 22990 9718 23042 9770
rect 23042 9718 23044 9770
rect 22988 9716 23044 9718
rect 26068 11406 26124 11452
rect 26068 11396 26070 11406
rect 26070 11396 26122 11406
rect 26122 11396 26124 11406
rect 26740 11406 26796 11452
rect 26740 11396 26742 11406
rect 26742 11396 26794 11406
rect 26794 11396 26796 11406
rect 27188 11284 27244 11340
rect 25172 11172 25228 11228
rect 25004 10388 25060 10444
rect 23044 9492 23100 9548
rect 23716 9156 23772 9212
rect 22820 8820 22876 8876
rect 23604 8484 23660 8540
rect 21588 8036 21644 8092
rect 21920 7866 21976 7868
rect 21920 7814 21922 7866
rect 21922 7814 21974 7866
rect 21974 7814 21976 7866
rect 21920 7812 21976 7814
rect 22024 7866 22080 7868
rect 22024 7814 22026 7866
rect 22026 7814 22078 7866
rect 22078 7814 22080 7866
rect 22024 7812 22080 7814
rect 22128 7866 22184 7868
rect 22128 7814 22130 7866
rect 22130 7814 22182 7866
rect 22182 7814 22184 7866
rect 22128 7812 22184 7814
rect 22708 8036 22764 8092
rect 21700 7410 21702 7420
rect 21702 7410 21754 7420
rect 21754 7410 21756 7420
rect 21700 7364 21756 7410
rect 21476 6692 21532 6748
rect 19852 6522 19908 6524
rect 19852 6470 19854 6522
rect 19854 6470 19906 6522
rect 19906 6470 19908 6522
rect 19852 6468 19908 6470
rect 19684 6356 19740 6412
rect 16100 4564 16156 4620
rect 15428 4506 15484 4508
rect 15428 4454 15430 4506
rect 15430 4454 15482 4506
rect 15482 4454 15484 4506
rect 15428 4452 15484 4454
rect 18340 5236 18396 5292
rect 17500 4788 17556 4844
rect 18004 4788 18060 4844
rect 17892 4676 17948 4732
rect 15876 4282 15932 4284
rect 15876 4230 15878 4282
rect 15878 4230 15930 4282
rect 15930 4230 15932 4282
rect 15876 4228 15932 4230
rect 15484 4004 15540 4060
rect 14924 3780 14980 3836
rect 15876 3892 15932 3948
rect 17332 4350 17388 4396
rect 17332 4340 17334 4350
rect 17334 4340 17386 4350
rect 17386 4340 17388 4350
rect 18004 4392 18006 4396
rect 18006 4392 18058 4396
rect 18058 4392 18060 4396
rect 18004 4340 18060 4392
rect 16716 4282 16772 4284
rect 16716 4230 16718 4282
rect 16718 4230 16770 4282
rect 16770 4230 16772 4282
rect 16716 4228 16772 4230
rect 14756 3496 14758 3500
rect 14758 3496 14810 3500
rect 14810 3496 14812 3500
rect 14756 3444 14812 3496
rect 15036 3498 15092 3500
rect 15036 3446 15038 3498
rect 15038 3446 15090 3498
rect 15090 3446 15092 3498
rect 15036 3444 15092 3446
rect 15708 3498 15764 3500
rect 15708 3446 15710 3498
rect 15710 3446 15762 3498
rect 15762 3446 15764 3498
rect 15708 3444 15764 3446
rect 15484 3386 15540 3388
rect 15484 3334 15486 3386
rect 15486 3334 15538 3386
rect 15538 3334 15540 3386
rect 15484 3332 15540 3334
rect 14756 2996 14812 3052
rect 14420 2548 14476 2604
rect 14532 2884 14588 2940
rect 14588 2324 14644 2380
rect 15316 2100 15372 2156
rect 13356 1930 13412 1932
rect 14364 1930 14420 1932
rect 13356 1878 13358 1930
rect 13358 1878 13410 1930
rect 13410 1878 13412 1930
rect 13356 1876 13412 1878
rect 14364 1878 14366 1930
rect 14366 1878 14418 1930
rect 14418 1878 14420 1930
rect 14364 1876 14420 1878
rect 11228 1652 11284 1708
rect 12908 1540 12964 1596
rect 15540 1764 15596 1820
rect 15372 1652 15428 1708
rect 16660 3722 16716 3724
rect 16660 3670 16662 3722
rect 16662 3670 16714 3722
rect 16714 3670 16716 3722
rect 16660 3668 16716 3670
rect 17644 3946 17700 3948
rect 17644 3894 17646 3946
rect 17646 3894 17698 3946
rect 17698 3894 17700 3946
rect 17644 3892 17700 3894
rect 17748 3946 17804 3948
rect 17748 3894 17750 3946
rect 17750 3894 17802 3946
rect 17802 3894 17804 3946
rect 17748 3892 17804 3894
rect 17852 3946 17908 3948
rect 17852 3894 17854 3946
rect 17854 3894 17906 3946
rect 17906 3894 17908 3946
rect 17852 3892 17908 3894
rect 16548 3332 16604 3388
rect 16324 2884 16380 2940
rect 16884 2996 16940 3052
rect 15988 2772 16044 2828
rect 16156 2548 16212 2604
rect 18844 5850 18900 5852
rect 18844 5798 18846 5850
rect 18846 5798 18898 5850
rect 18898 5798 18900 5850
rect 18844 5796 18900 5798
rect 19460 5846 19462 5852
rect 19462 5846 19514 5852
rect 19514 5846 19516 5852
rect 19460 5796 19516 5846
rect 22708 7530 22764 7532
rect 22708 7478 22710 7530
rect 22710 7478 22762 7530
rect 22762 7478 22764 7530
rect 22708 7476 22764 7478
rect 25004 10052 25060 10108
rect 24388 9967 24390 9996
rect 24390 9967 24442 9996
rect 24442 9967 24444 9996
rect 24388 9940 24444 9967
rect 25788 11226 25844 11228
rect 25788 11174 25790 11226
rect 25790 11174 25842 11226
rect 25842 11174 25844 11226
rect 25788 11172 25844 11174
rect 26964 11172 27020 11228
rect 25508 10052 25564 10108
rect 25284 8708 25340 8764
rect 25060 8372 25116 8428
rect 24276 8260 24332 8316
rect 25172 8148 25228 8204
rect 24836 7588 24892 7644
rect 23044 7140 23100 7196
rect 22092 6468 22148 6524
rect 21812 6356 21868 6412
rect 21920 6298 21976 6300
rect 21920 6246 21922 6298
rect 21922 6246 21974 6298
rect 21974 6246 21976 6298
rect 21920 6244 21976 6246
rect 22024 6298 22080 6300
rect 22024 6246 22026 6298
rect 22026 6246 22078 6298
rect 22078 6246 22080 6298
rect 22024 6244 22080 6246
rect 22128 6298 22184 6300
rect 22128 6246 22130 6298
rect 22130 6246 22182 6298
rect 22182 6246 22184 6298
rect 22128 6244 22184 6246
rect 19908 5842 19910 5852
rect 19910 5842 19962 5852
rect 19962 5842 19964 5852
rect 19908 5796 19964 5842
rect 19740 5348 19796 5404
rect 19012 4676 19068 4732
rect 18844 4564 18900 4620
rect 18844 4394 18900 4396
rect 18844 4342 18846 4394
rect 18846 4342 18898 4394
rect 18898 4342 18900 4394
rect 18844 4340 18900 4342
rect 19124 4564 19180 4620
rect 19348 5050 19350 5068
rect 19350 5050 19402 5068
rect 19402 5050 19404 5068
rect 19348 5012 19404 5050
rect 22820 6634 22876 6636
rect 22820 6582 22822 6634
rect 22822 6582 22874 6634
rect 22874 6582 22876 6634
rect 22820 6580 22876 6582
rect 22484 6468 22540 6524
rect 22820 5850 22876 5852
rect 22820 5798 22822 5850
rect 22822 5798 22874 5850
rect 22874 5798 22876 5850
rect 22820 5796 22876 5798
rect 22260 5572 22316 5628
rect 19908 4900 19964 4956
rect 19236 4452 19292 4508
rect 19796 4564 19852 4620
rect 20020 4564 20076 4620
rect 19908 4340 19964 4396
rect 19012 3668 19068 3724
rect 20356 4900 20412 4956
rect 22932 4900 22988 4956
rect 21920 4730 21976 4732
rect 21920 4678 21922 4730
rect 21922 4678 21974 4730
rect 21974 4678 21976 4730
rect 21920 4676 21976 4678
rect 22024 4730 22080 4732
rect 22024 4678 22026 4730
rect 22026 4678 22078 4730
rect 22078 4678 22080 4730
rect 22024 4676 22080 4678
rect 22128 4730 22184 4732
rect 22128 4678 22130 4730
rect 22130 4678 22182 4730
rect 22182 4678 22184 4730
rect 22128 4676 22184 4678
rect 20692 4506 20748 4508
rect 20692 4454 20694 4506
rect 20694 4454 20746 4506
rect 20746 4454 20748 4506
rect 20692 4452 20748 4454
rect 20580 4340 20636 4396
rect 21084 4394 21140 4396
rect 21084 4342 21086 4394
rect 21086 4342 21138 4394
rect 21138 4342 21140 4394
rect 21084 4340 21140 4342
rect 20412 4170 20468 4172
rect 20412 4118 20414 4170
rect 20414 4118 20466 4170
rect 20466 4118 20468 4170
rect 20412 4116 20468 4118
rect 16996 2772 17052 2828
rect 17556 2884 17612 2940
rect 18116 2884 18172 2940
rect 18452 2660 18508 2716
rect 18116 2436 18172 2492
rect 17644 2378 17700 2380
rect 17644 2326 17646 2378
rect 17646 2326 17698 2378
rect 17698 2326 17700 2378
rect 17644 2324 17700 2326
rect 17748 2378 17804 2380
rect 17748 2326 17750 2378
rect 17750 2326 17802 2378
rect 17802 2326 17804 2378
rect 17748 2324 17804 2326
rect 17852 2378 17908 2380
rect 17852 2326 17854 2378
rect 17854 2326 17906 2378
rect 17906 2326 17908 2378
rect 17852 2324 17908 2326
rect 16884 2100 16940 2156
rect 17724 2154 17780 2156
rect 17724 2102 17726 2154
rect 17726 2102 17778 2154
rect 17778 2102 17780 2154
rect 17724 2100 17780 2102
rect 17612 2042 17668 2044
rect 17612 1990 17614 2042
rect 17614 1990 17666 2042
rect 17666 1990 17668 2042
rect 17612 1988 17668 1990
rect 15876 1652 15932 1708
rect 18060 2154 18116 2156
rect 18060 2102 18062 2154
rect 18062 2102 18114 2154
rect 18114 2102 18116 2154
rect 18060 2100 18116 2102
rect 19404 3108 19460 3164
rect 19012 2714 19068 2716
rect 19012 2662 19014 2714
rect 19014 2662 19066 2714
rect 19066 2662 19068 2714
rect 19012 2660 19068 2662
rect 18788 2548 18844 2604
rect 21308 3780 21364 3836
rect 22036 4282 22092 4284
rect 22036 4230 22038 4282
rect 22038 4230 22090 4282
rect 22090 4230 22092 4282
rect 22036 4228 22092 4230
rect 22428 4282 22484 4284
rect 22428 4230 22430 4282
rect 22430 4230 22482 4282
rect 22482 4230 22484 4282
rect 22428 4228 22484 4230
rect 22484 3780 22540 3836
rect 21700 3556 21756 3612
rect 21980 3610 22036 3612
rect 21980 3558 21982 3610
rect 21982 3558 22034 3610
rect 22034 3558 22036 3610
rect 21980 3556 22036 3558
rect 21308 3498 21364 3500
rect 21308 3446 21310 3498
rect 21310 3446 21362 3498
rect 21362 3446 21364 3498
rect 21308 3444 21364 3446
rect 22204 3498 22260 3500
rect 22204 3446 22206 3498
rect 22206 3446 22258 3498
rect 22258 3446 22260 3498
rect 22204 3444 22260 3446
rect 20916 3386 20972 3388
rect 20916 3334 20918 3386
rect 20918 3334 20970 3386
rect 20970 3334 20972 3386
rect 20916 3332 20972 3334
rect 21196 3386 21252 3388
rect 21196 3334 21198 3386
rect 21198 3334 21250 3386
rect 21250 3334 21252 3386
rect 21196 3332 21252 3334
rect 21476 3220 21532 3276
rect 20132 3108 20188 3164
rect 20580 3108 20636 3164
rect 20020 2772 20076 2828
rect 19068 2436 19124 2492
rect 18508 2154 18564 2156
rect 18508 2102 18510 2154
rect 18510 2102 18562 2154
rect 18562 2102 18564 2154
rect 18508 2100 18564 2102
rect 18844 2324 18900 2380
rect 17724 1652 17780 1708
rect 19404 2324 19460 2380
rect 18844 1652 18900 1708
rect 19684 2100 19740 2156
rect 19964 2436 20020 2492
rect 13368 1594 13424 1596
rect 13368 1542 13370 1594
rect 13370 1542 13422 1594
rect 13422 1542 13424 1594
rect 13368 1540 13424 1542
rect 13472 1594 13528 1596
rect 13472 1542 13474 1594
rect 13474 1542 13526 1594
rect 13526 1542 13528 1594
rect 13472 1540 13528 1542
rect 13576 1594 13632 1596
rect 13576 1542 13578 1594
rect 13578 1542 13630 1594
rect 13630 1542 13632 1594
rect 13576 1540 13632 1542
rect 17724 1258 17780 1260
rect 17724 1206 17726 1258
rect 17726 1206 17778 1258
rect 17778 1206 17780 1258
rect 17724 1204 17780 1206
rect 19180 1652 19236 1708
rect 19572 1652 19628 1708
rect 19740 1652 19796 1708
rect 20188 1876 20244 1932
rect 20580 2324 20636 2380
rect 20692 2772 20748 2828
rect 20804 2212 20860 2268
rect 20356 1764 20412 1820
rect 21308 2042 21364 2044
rect 21308 1990 21310 2042
rect 21310 1990 21362 2042
rect 21362 1990 21364 2042
rect 21308 1988 21364 1990
rect 19628 1258 19684 1260
rect 19628 1206 19630 1258
rect 19630 1206 19682 1258
rect 19682 1206 19684 1258
rect 19628 1204 19684 1206
rect 20188 1428 20244 1484
rect 20300 1540 20356 1596
rect 20076 1316 20132 1372
rect 19404 1146 19460 1148
rect 19404 1094 19406 1146
rect 19406 1094 19458 1146
rect 19458 1094 19460 1146
rect 19404 1092 19460 1094
rect 9092 810 9148 812
rect 9092 758 9094 810
rect 9094 758 9146 810
rect 9146 758 9148 810
rect 9092 756 9148 758
rect 9196 810 9252 812
rect 9196 758 9198 810
rect 9198 758 9250 810
rect 9250 758 9252 810
rect 9196 756 9252 758
rect 9300 810 9356 812
rect 9300 758 9302 810
rect 9302 758 9354 810
rect 9354 758 9356 810
rect 9300 756 9356 758
rect 17948 1034 18004 1036
rect 17948 982 17950 1034
rect 17950 982 18002 1034
rect 18002 982 18004 1034
rect 17948 980 18004 982
rect 18172 868 18228 924
rect 17644 810 17700 812
rect 17644 758 17646 810
rect 17646 758 17698 810
rect 17698 758 17700 810
rect 17644 756 17700 758
rect 17748 810 17804 812
rect 17748 758 17750 810
rect 17750 758 17802 810
rect 17802 758 17804 810
rect 17748 756 17804 758
rect 17852 810 17908 812
rect 17852 758 17854 810
rect 17854 758 17906 810
rect 17906 758 17908 810
rect 17852 756 17908 758
rect 17500 644 17556 700
rect 18396 532 18452 588
rect 20412 1428 20468 1484
rect 20748 1316 20804 1372
rect 21084 1818 21140 1820
rect 21084 1766 21086 1818
rect 21086 1766 21138 1818
rect 21138 1766 21140 1818
rect 21084 1764 21140 1766
rect 21920 3162 21976 3164
rect 21920 3110 21922 3162
rect 21922 3110 21974 3162
rect 21974 3110 21976 3162
rect 21920 3108 21976 3110
rect 22024 3162 22080 3164
rect 22024 3110 22026 3162
rect 22026 3110 22078 3162
rect 22078 3110 22080 3162
rect 22024 3108 22080 3110
rect 22128 3162 22184 3164
rect 22128 3110 22130 3162
rect 22130 3110 22182 3162
rect 22182 3110 22184 3162
rect 22128 3108 22184 3110
rect 21588 2772 21644 2828
rect 22260 2772 22316 2828
rect 21868 2548 21924 2604
rect 21644 2324 21700 2380
rect 23492 6580 23548 6636
rect 23380 5796 23436 5852
rect 23156 4564 23212 4620
rect 23828 5290 23884 5292
rect 23828 5238 23830 5290
rect 23830 5238 23882 5290
rect 23882 5238 23884 5290
rect 23828 5236 23884 5238
rect 24332 6634 24388 6636
rect 24332 6582 24334 6634
rect 24334 6582 24386 6634
rect 24386 6582 24388 6634
rect 24332 6580 24388 6582
rect 24556 6580 24612 6636
rect 24388 6356 24444 6412
rect 25060 8036 25116 8092
rect 25284 7924 25340 7980
rect 25172 7364 25228 7420
rect 25732 10546 25734 10556
rect 25734 10546 25786 10556
rect 25786 10546 25788 10556
rect 25732 10500 25788 10546
rect 25620 8194 25622 8204
rect 25622 8194 25674 8204
rect 25674 8194 25676 8204
rect 25620 8148 25676 8194
rect 25508 8036 25564 8092
rect 25396 6468 25452 6524
rect 25508 7140 25564 7196
rect 25732 7486 25788 7532
rect 25732 7476 25734 7486
rect 25734 7476 25786 7486
rect 25786 7476 25788 7486
rect 24276 5124 24332 5180
rect 24108 4954 24164 4956
rect 24108 4902 24110 4954
rect 24110 4902 24162 4954
rect 24162 4902 24164 4954
rect 24108 4900 24164 4902
rect 24332 4954 24388 4956
rect 24332 4902 24334 4954
rect 24334 4902 24386 4954
rect 24386 4902 24388 4954
rect 24332 4900 24388 4902
rect 24500 4564 24556 4620
rect 23044 4340 23100 4396
rect 23212 4170 23268 4172
rect 23212 4118 23214 4170
rect 23214 4118 23266 4170
rect 23266 4118 23268 4170
rect 23212 4116 23268 4118
rect 23380 3668 23436 3724
rect 22596 3572 22652 3612
rect 22596 3556 22598 3572
rect 22598 3556 22650 3572
rect 22650 3556 22652 3572
rect 23492 2772 23548 2828
rect 23604 2660 23660 2716
rect 24332 4394 24388 4396
rect 24332 4342 24334 4394
rect 24334 4342 24386 4394
rect 24386 4342 24388 4394
rect 24332 4340 24388 4342
rect 23716 3444 23772 3500
rect 24052 4116 24108 4172
rect 24276 3780 24332 3836
rect 26012 10666 26068 10668
rect 26012 10614 26014 10666
rect 26014 10614 26066 10666
rect 26066 10614 26068 10666
rect 26012 10612 26068 10614
rect 26068 10388 26124 10444
rect 25956 9716 26012 9772
rect 25956 8986 26012 8988
rect 25956 8934 25958 8986
rect 25958 8934 26010 8986
rect 26010 8934 26012 8986
rect 25956 8932 26012 8934
rect 26292 10388 26348 10444
rect 26196 10218 26252 10220
rect 26196 10166 26198 10218
rect 26198 10166 26250 10218
rect 26250 10166 26252 10218
rect 26196 10164 26252 10166
rect 26300 10218 26356 10220
rect 26300 10166 26302 10218
rect 26302 10166 26354 10218
rect 26354 10166 26356 10218
rect 26300 10164 26356 10166
rect 26404 10218 26460 10220
rect 26404 10166 26406 10218
rect 26406 10166 26458 10218
rect 26458 10166 26460 10218
rect 26404 10164 26460 10166
rect 26404 9940 26460 9996
rect 26628 9940 26684 9996
rect 27020 9828 27076 9884
rect 26572 9770 26628 9772
rect 26572 9718 26574 9770
rect 26574 9718 26626 9770
rect 26626 9718 26628 9770
rect 26572 9716 26628 9718
rect 26740 9268 26796 9324
rect 26628 9210 26684 9212
rect 26628 9158 26630 9210
rect 26630 9158 26682 9210
rect 26682 9158 26684 9210
rect 26628 9156 26684 9158
rect 30268 11956 30324 12012
rect 29932 11732 29988 11788
rect 29428 11508 29484 11564
rect 28588 11396 28644 11452
rect 27636 11284 27692 11340
rect 28980 11284 29036 11340
rect 29428 11284 29484 11340
rect 28196 10052 28252 10108
rect 26068 8820 26124 8876
rect 26516 8932 26572 8988
rect 26196 8650 26252 8652
rect 26196 8598 26198 8650
rect 26198 8598 26250 8650
rect 26250 8598 26252 8650
rect 26196 8596 26252 8598
rect 26300 8650 26356 8652
rect 26300 8598 26302 8650
rect 26302 8598 26354 8650
rect 26354 8598 26356 8650
rect 26300 8596 26356 8598
rect 26404 8650 26460 8652
rect 26404 8598 26406 8650
rect 26406 8598 26458 8650
rect 26458 8598 26460 8650
rect 26404 8596 26460 8598
rect 26404 8426 26460 8428
rect 26404 8374 26406 8426
rect 26406 8374 26458 8426
rect 26458 8374 26460 8426
rect 26404 8372 26460 8374
rect 26236 8090 26292 8092
rect 26236 8038 26238 8090
rect 26238 8038 26290 8090
rect 26290 8038 26292 8090
rect 26236 8036 26292 8038
rect 25396 5460 25452 5516
rect 25508 5372 25564 5404
rect 25508 5348 25510 5372
rect 25510 5348 25562 5372
rect 25562 5348 25564 5372
rect 24836 4228 24892 4284
rect 25396 5012 25452 5068
rect 24948 4004 25004 4060
rect 24836 3556 24892 3612
rect 23716 3220 23772 3276
rect 23492 2602 23548 2604
rect 23492 2550 23494 2602
rect 23494 2550 23546 2602
rect 23546 2550 23548 2602
rect 23492 2548 23548 2550
rect 23716 2548 23772 2604
rect 23940 2660 23996 2716
rect 23492 2324 23548 2380
rect 23604 2436 23660 2492
rect 23380 2212 23436 2268
rect 23268 2100 23324 2156
rect 23772 2212 23828 2268
rect 21868 1930 21924 1932
rect 21868 1878 21870 1930
rect 21870 1878 21922 1930
rect 21922 1878 21924 1930
rect 21868 1876 21924 1878
rect 22372 1988 22428 2044
rect 21644 1428 21700 1484
rect 22708 1988 22764 2044
rect 21420 1316 21476 1372
rect 22540 1764 22596 1820
rect 22260 1652 22316 1708
rect 21920 1594 21976 1596
rect 21920 1542 21922 1594
rect 21922 1542 21974 1594
rect 21974 1542 21976 1594
rect 21920 1540 21976 1542
rect 22024 1594 22080 1596
rect 22024 1542 22026 1594
rect 22026 1542 22078 1594
rect 22078 1542 22080 1594
rect 22024 1540 22080 1542
rect 22128 1594 22184 1596
rect 22128 1542 22130 1594
rect 22130 1542 22182 1594
rect 22182 1542 22184 1594
rect 22128 1540 22184 1542
rect 22092 1146 22148 1148
rect 22092 1094 22094 1146
rect 22094 1094 22146 1146
rect 22146 1094 22148 1146
rect 22092 1092 22148 1094
rect 24164 2100 24220 2156
rect 24332 2548 24388 2604
rect 24556 2324 24612 2380
rect 24892 2212 24948 2268
rect 25116 2602 25172 2604
rect 25116 2550 25118 2602
rect 25118 2550 25170 2602
rect 25170 2550 25172 2602
rect 25116 2548 25172 2550
rect 23996 2042 24052 2044
rect 23996 1990 23998 2042
rect 23998 1990 24050 2042
rect 24050 1990 24052 2042
rect 23996 1988 24052 1990
rect 22820 1876 22876 1932
rect 23268 1930 23324 1932
rect 23268 1878 23270 1930
rect 23270 1878 23322 1930
rect 23322 1878 23324 1930
rect 23268 1876 23324 1878
rect 24948 1998 25004 2044
rect 24948 1988 24950 1998
rect 24950 1988 25002 1998
rect 25002 1988 25004 1998
rect 22988 1428 23044 1484
rect 23436 1428 23492 1484
rect 23940 1428 23996 1484
rect 25060 1764 25116 1820
rect 24948 1652 25004 1708
rect 23660 1258 23716 1260
rect 23660 1206 23662 1258
rect 23662 1206 23714 1258
rect 23714 1206 23716 1258
rect 23660 1204 23716 1206
rect 24108 1258 24164 1260
rect 24108 1206 24110 1258
rect 24110 1206 24162 1258
rect 24162 1206 24164 1258
rect 24108 1204 24164 1206
rect 24780 1258 24836 1260
rect 24780 1206 24782 1258
rect 24782 1206 24834 1258
rect 24834 1206 24836 1258
rect 24780 1204 24836 1206
rect 25396 3722 25452 3724
rect 25396 3670 25398 3722
rect 25398 3670 25450 3722
rect 25450 3670 25452 3722
rect 25396 3668 25452 3670
rect 25844 5914 25900 5964
rect 25844 5908 25846 5914
rect 25846 5908 25898 5914
rect 25898 5908 25900 5914
rect 25620 4004 25676 4060
rect 25620 3332 25676 3388
rect 25564 2826 25620 2828
rect 25564 2774 25566 2826
rect 25566 2774 25618 2826
rect 25618 2774 25620 2826
rect 25564 2772 25620 2774
rect 25676 2714 25732 2716
rect 25676 2662 25678 2714
rect 25678 2662 25730 2714
rect 25730 2662 25732 2714
rect 25676 2660 25732 2662
rect 27188 8820 27244 8876
rect 26796 8314 26852 8316
rect 26796 8262 26798 8314
rect 26798 8262 26850 8314
rect 26850 8262 26852 8314
rect 26796 8260 26852 8262
rect 26628 8194 26630 8204
rect 26630 8194 26682 8204
rect 26682 8194 26684 8204
rect 26628 8148 26684 8194
rect 27020 8202 27076 8204
rect 27020 8150 27022 8202
rect 27022 8150 27074 8202
rect 27074 8150 27076 8202
rect 27020 8148 27076 8150
rect 26628 7924 26684 7980
rect 26516 7476 26572 7532
rect 26740 7306 26796 7308
rect 26740 7254 26742 7306
rect 26742 7254 26794 7306
rect 26794 7254 26796 7306
rect 26740 7252 26796 7254
rect 26196 7082 26252 7084
rect 26196 7030 26198 7082
rect 26198 7030 26250 7082
rect 26250 7030 26252 7082
rect 26196 7028 26252 7030
rect 26300 7082 26356 7084
rect 26300 7030 26302 7082
rect 26302 7030 26354 7082
rect 26354 7030 26356 7082
rect 26300 7028 26356 7030
rect 26404 7082 26460 7084
rect 26404 7030 26406 7082
rect 26406 7030 26458 7082
rect 26458 7030 26460 7082
rect 26404 7028 26460 7030
rect 26852 6804 26908 6860
rect 26404 5842 26406 5852
rect 26406 5842 26458 5852
rect 26458 5842 26460 5852
rect 26404 5796 26460 5842
rect 25956 5348 26012 5404
rect 26068 5572 26124 5628
rect 26196 5514 26252 5516
rect 26196 5462 26198 5514
rect 26198 5462 26250 5514
rect 26250 5462 26252 5514
rect 26196 5460 26252 5462
rect 26300 5514 26356 5516
rect 26300 5462 26302 5514
rect 26302 5462 26354 5514
rect 26354 5462 26356 5514
rect 26300 5460 26356 5462
rect 26404 5514 26460 5516
rect 26404 5462 26406 5514
rect 26406 5462 26458 5514
rect 26458 5462 26460 5514
rect 26404 5460 26460 5462
rect 27860 9604 27916 9660
rect 27524 8874 27580 8876
rect 27524 8822 27526 8874
rect 27526 8822 27578 8874
rect 27578 8822 27580 8874
rect 27524 8820 27580 8822
rect 27412 8148 27468 8204
rect 27076 7140 27132 7196
rect 27748 8484 27804 8540
rect 27860 8372 27916 8428
rect 27972 8260 28028 8316
rect 27636 7252 27692 7308
rect 28532 10052 28588 10108
rect 29428 9716 29484 9772
rect 29316 9156 29372 9212
rect 30660 11844 30716 11900
rect 31332 11732 31388 11788
rect 30044 11338 30100 11340
rect 30044 11286 30046 11338
rect 30046 11286 30098 11338
rect 30098 11286 30100 11338
rect 30044 11284 30100 11286
rect 30472 11002 30528 11004
rect 30472 10950 30474 11002
rect 30474 10950 30526 11002
rect 30526 10950 30528 11002
rect 30472 10948 30528 10950
rect 30576 11002 30632 11004
rect 30576 10950 30578 11002
rect 30578 10950 30630 11002
rect 30630 10950 30632 11002
rect 30576 10948 30632 10950
rect 30680 11002 30736 11004
rect 30680 10950 30682 11002
rect 30682 10950 30734 11002
rect 30734 10950 30736 11002
rect 30680 10948 30736 10950
rect 29764 10724 29820 10780
rect 29764 10546 29766 10556
rect 29766 10546 29818 10556
rect 29818 10546 29820 10556
rect 29764 10500 29820 10546
rect 30996 10546 30998 10556
rect 30998 10546 31050 10556
rect 31050 10546 31052 10556
rect 30996 10500 31052 10546
rect 29876 9828 29932 9884
rect 31220 10052 31276 10108
rect 29540 9044 29596 9100
rect 29876 8372 29932 8428
rect 29316 8148 29372 8204
rect 28084 6804 28140 6860
rect 28756 7252 28812 7308
rect 27412 6692 27468 6748
rect 27972 6020 28028 6076
rect 28420 5908 28476 5964
rect 28644 6244 28700 6300
rect 27972 5236 28028 5292
rect 25956 4340 26012 4396
rect 26404 5124 26460 5180
rect 26628 5066 26684 5068
rect 26628 5014 26630 5066
rect 26630 5014 26682 5066
rect 26682 5014 26684 5066
rect 26628 5012 26684 5014
rect 27356 4954 27412 4956
rect 27356 4902 27358 4954
rect 27358 4902 27410 4954
rect 27410 4902 27412 4954
rect 27356 4900 27412 4902
rect 26404 4788 26460 4844
rect 26516 4506 26572 4508
rect 26516 4454 26518 4506
rect 26518 4454 26570 4506
rect 26570 4454 26572 4506
rect 26516 4452 26572 4454
rect 28140 5178 28196 5180
rect 28140 5126 28142 5178
rect 28142 5126 28194 5178
rect 28194 5126 28196 5178
rect 28140 5124 28196 5126
rect 27468 4452 27524 4508
rect 27916 4506 27972 4508
rect 27916 4454 27918 4506
rect 27918 4454 27970 4506
rect 27970 4454 27972 4506
rect 27916 4452 27972 4454
rect 26196 3946 26252 3948
rect 26196 3894 26198 3946
rect 26198 3894 26250 3946
rect 26250 3894 26252 3946
rect 26196 3892 26252 3894
rect 26300 3946 26356 3948
rect 26300 3894 26302 3946
rect 26302 3894 26354 3946
rect 26354 3894 26356 3946
rect 26300 3892 26356 3894
rect 26404 3946 26460 3948
rect 26404 3894 26406 3946
rect 26406 3894 26458 3946
rect 26458 3894 26460 3946
rect 26404 3892 26460 3894
rect 26404 3610 26460 3612
rect 26404 3558 26406 3610
rect 26406 3558 26458 3610
rect 26458 3558 26460 3610
rect 26404 3556 26460 3558
rect 26124 3332 26180 3388
rect 26404 3332 26460 3388
rect 26516 3444 26572 3500
rect 26852 4004 26908 4060
rect 26740 3498 26796 3500
rect 26740 3446 26742 3498
rect 26742 3446 26794 3498
rect 26794 3446 26796 3498
rect 26740 3444 26796 3446
rect 26516 3108 26572 3164
rect 26628 2996 26684 3052
rect 26348 2938 26404 2940
rect 26348 2886 26350 2938
rect 26350 2886 26402 2938
rect 26402 2886 26404 2938
rect 26348 2884 26404 2886
rect 25844 2548 25900 2604
rect 26404 2602 26460 2604
rect 26404 2550 26406 2602
rect 26406 2550 26458 2602
rect 26458 2550 26460 2602
rect 26404 2548 26460 2550
rect 27244 3610 27300 3612
rect 27244 3558 27246 3610
rect 27246 3558 27298 3610
rect 27298 3558 27300 3610
rect 27244 3556 27300 3558
rect 26852 2996 26908 3052
rect 27412 2996 27468 3052
rect 28868 5684 28924 5740
rect 28028 4170 28084 4172
rect 28028 4118 28030 4170
rect 28030 4118 28082 4170
rect 28082 4118 28084 4170
rect 28028 4116 28084 4118
rect 28532 4564 28588 4620
rect 28420 4340 28476 4396
rect 27748 3668 27804 3724
rect 28196 3668 28252 3724
rect 32340 10500 32396 10556
rect 30100 9716 30156 9772
rect 30472 9434 30528 9436
rect 30472 9382 30474 9434
rect 30474 9382 30526 9434
rect 30526 9382 30528 9434
rect 30472 9380 30528 9382
rect 30576 9434 30632 9436
rect 30576 9382 30578 9434
rect 30578 9382 30630 9434
rect 30630 9382 30632 9434
rect 30576 9380 30632 9382
rect 30680 9434 30736 9436
rect 30680 9382 30682 9434
rect 30682 9382 30734 9434
rect 30734 9382 30736 9434
rect 30680 9380 30736 9382
rect 31556 10052 31612 10108
rect 30324 9054 30380 9100
rect 30324 9044 30326 9054
rect 30326 9044 30378 9054
rect 30378 9044 30380 9054
rect 30100 8820 30156 8876
rect 31108 8932 31164 8988
rect 30212 8426 30268 8428
rect 30212 8374 30214 8426
rect 30214 8374 30266 8426
rect 30266 8374 30268 8426
rect 30212 8372 30268 8374
rect 30884 8090 30940 8092
rect 30884 8038 30886 8090
rect 30886 8038 30938 8090
rect 30938 8038 30940 8090
rect 30884 8036 30940 8038
rect 30472 7866 30528 7868
rect 30472 7814 30474 7866
rect 30474 7814 30526 7866
rect 30526 7814 30528 7866
rect 30472 7812 30528 7814
rect 30576 7866 30632 7868
rect 30576 7814 30578 7866
rect 30578 7814 30630 7866
rect 30630 7814 30632 7866
rect 30576 7812 30632 7814
rect 30680 7866 30736 7868
rect 30680 7814 30682 7866
rect 30682 7814 30734 7866
rect 30734 7814 30736 7866
rect 30680 7812 30736 7814
rect 30884 7642 30940 7644
rect 30884 7590 30886 7642
rect 30886 7590 30938 7642
rect 30938 7590 30940 7642
rect 30884 7588 30940 7590
rect 30268 7418 30324 7420
rect 30268 7366 30270 7418
rect 30270 7366 30322 7418
rect 30322 7366 30324 7418
rect 30268 7364 30324 7366
rect 30380 7306 30436 7308
rect 30380 7254 30382 7306
rect 30382 7254 30434 7306
rect 30434 7254 30436 7306
rect 30380 7252 30436 7254
rect 30996 6580 31052 6636
rect 29876 6244 29932 6300
rect 30472 6298 30528 6300
rect 30472 6246 30474 6298
rect 30474 6246 30526 6298
rect 30526 6246 30528 6298
rect 30472 6244 30528 6246
rect 30576 6298 30632 6300
rect 30576 6246 30578 6298
rect 30578 6246 30630 6298
rect 30630 6246 30632 6298
rect 30576 6244 30632 6246
rect 30680 6298 30736 6300
rect 30680 6246 30682 6298
rect 30682 6246 30734 6298
rect 30734 6246 30736 6298
rect 30680 6244 30736 6246
rect 29652 6132 29708 6188
rect 30884 6074 30940 6076
rect 30884 6022 30886 6074
rect 30886 6022 30938 6074
rect 30938 6022 30940 6074
rect 30884 6020 30940 6022
rect 29764 5908 29820 5964
rect 29036 4954 29092 4956
rect 29036 4902 29038 4954
rect 29038 4902 29090 4954
rect 29090 4902 29092 4954
rect 29036 4900 29092 4902
rect 29260 4954 29316 4956
rect 29260 4902 29262 4954
rect 29262 4902 29314 4954
rect 29314 4902 29316 4954
rect 29260 4900 29316 4902
rect 29092 4228 29148 4284
rect 28868 3780 28924 3836
rect 28700 3556 28756 3612
rect 27524 2884 27580 2940
rect 26740 2436 26796 2492
rect 27188 2548 27244 2604
rect 27412 2772 27468 2828
rect 25396 2212 25452 2268
rect 25956 2324 26012 2380
rect 26196 2378 26252 2380
rect 26196 2326 26198 2378
rect 26198 2326 26250 2378
rect 26250 2326 26252 2378
rect 26196 2324 26252 2326
rect 26300 2378 26356 2380
rect 26300 2326 26302 2378
rect 26302 2326 26354 2378
rect 26354 2326 26356 2378
rect 26300 2324 26356 2326
rect 26404 2378 26460 2380
rect 26404 2326 26406 2378
rect 26406 2326 26458 2378
rect 26458 2326 26460 2378
rect 26404 2324 26460 2326
rect 25956 1876 26012 1932
rect 25732 1540 25788 1596
rect 25228 1258 25284 1260
rect 25228 1206 25230 1258
rect 25230 1206 25282 1258
rect 25282 1206 25284 1258
rect 25228 1204 25284 1206
rect 26740 1876 26796 1932
rect 26572 1764 26628 1820
rect 27412 1876 27468 1932
rect 26852 1540 26908 1596
rect 28196 3108 28252 3164
rect 28532 3220 28588 3276
rect 28532 2706 28534 2716
rect 28534 2706 28586 2716
rect 28586 2706 28588 2716
rect 28532 2660 28588 2706
rect 28308 2436 28364 2492
rect 28084 2212 28140 2268
rect 27860 2042 27916 2044
rect 27860 1990 27862 2042
rect 27862 1990 27914 2042
rect 27914 1990 27916 2042
rect 27860 1988 27916 1990
rect 26908 1258 26964 1260
rect 26908 1206 26910 1258
rect 26910 1206 26962 1258
rect 26962 1206 26964 1258
rect 26908 1204 26964 1206
rect 27132 1258 27188 1260
rect 27132 1206 27134 1258
rect 27134 1206 27186 1258
rect 27186 1206 27188 1258
rect 27748 1876 27804 1932
rect 27132 1204 27188 1206
rect 28532 1930 28588 1932
rect 28532 1878 28534 1930
rect 28534 1878 28586 1930
rect 28586 1878 28588 1930
rect 28532 1876 28588 1878
rect 28868 3108 28924 3164
rect 28980 3490 28982 3500
rect 28982 3490 29034 3500
rect 29034 3490 29036 3500
rect 28980 3444 29036 3490
rect 29092 3332 29148 3388
rect 29316 3220 29372 3276
rect 29428 3108 29484 3164
rect 30212 5738 30268 5740
rect 30212 5686 30214 5738
rect 30214 5686 30266 5738
rect 30266 5686 30268 5738
rect 30212 5684 30268 5686
rect 29876 4564 29932 4620
rect 29764 4340 29820 4396
rect 29820 4170 29876 4172
rect 29820 4118 29822 4170
rect 29822 4118 29874 4170
rect 29874 4118 29876 4170
rect 29820 4116 29876 4118
rect 30044 4004 30100 4060
rect 29652 3780 29708 3836
rect 29652 3566 29708 3612
rect 29652 3556 29654 3566
rect 29654 3556 29706 3566
rect 29706 3556 29708 3566
rect 29764 3332 29820 3388
rect 29540 2660 29596 2716
rect 29652 3220 29708 3276
rect 30472 4730 30528 4732
rect 30472 4678 30474 4730
rect 30474 4678 30526 4730
rect 30526 4678 30528 4730
rect 30472 4676 30528 4678
rect 30576 4730 30632 4732
rect 30576 4678 30578 4730
rect 30578 4678 30630 4730
rect 30630 4678 30632 4730
rect 30576 4676 30632 4678
rect 30680 4730 30736 4732
rect 30680 4678 30682 4730
rect 30682 4678 30734 4730
rect 30734 4678 30736 4730
rect 30680 4676 30736 4678
rect 30884 4506 30940 4508
rect 30884 4454 30886 4506
rect 30886 4454 30938 4506
rect 30938 4454 30940 4506
rect 30884 4452 30940 4454
rect 30324 3668 30380 3724
rect 29988 3490 29990 3500
rect 29990 3490 30042 3500
rect 30042 3490 30044 3500
rect 29988 3444 30044 3490
rect 30436 3780 30492 3836
rect 32340 9766 32342 9772
rect 32342 9766 32394 9772
rect 32394 9766 32396 9772
rect 32340 9716 32396 9766
rect 31780 8932 31836 8988
rect 32452 8596 32508 8652
rect 31556 8372 31612 8428
rect 31220 8202 31276 8204
rect 31220 8150 31222 8202
rect 31222 8150 31274 8202
rect 31274 8150 31276 8202
rect 31220 8148 31276 8150
rect 31444 7588 31500 7644
rect 31780 8372 31836 8428
rect 32116 6132 32172 6188
rect 31556 4170 31612 4172
rect 31556 4118 31558 4170
rect 31558 4118 31610 4170
rect 31610 4118 31612 4170
rect 31556 4116 31612 4118
rect 31108 3780 31164 3836
rect 28924 2154 28980 2156
rect 28924 2102 28926 2154
rect 28926 2102 28978 2154
rect 28978 2102 28980 2154
rect 28924 2100 28980 2102
rect 29876 2660 29932 2716
rect 30472 3162 30528 3164
rect 30472 3110 30474 3162
rect 30474 3110 30526 3162
rect 30526 3110 30528 3162
rect 30472 3108 30528 3110
rect 30576 3162 30632 3164
rect 30576 3110 30578 3162
rect 30578 3110 30630 3162
rect 30630 3110 30632 3162
rect 30576 3108 30632 3110
rect 30680 3162 30736 3164
rect 30680 3110 30682 3162
rect 30682 3110 30734 3162
rect 30734 3110 30736 3162
rect 30680 3108 30736 3110
rect 30996 3220 31052 3276
rect 30884 2782 30940 2828
rect 30884 2772 30886 2782
rect 30886 2772 30938 2782
rect 30938 2772 30940 2782
rect 29764 2100 29820 2156
rect 29988 2436 30044 2492
rect 29148 1988 29204 2044
rect 28140 1258 28196 1260
rect 28140 1206 28142 1258
rect 28142 1206 28194 1258
rect 28194 1206 28196 1258
rect 28140 1204 28196 1206
rect 28812 1652 28868 1708
rect 28924 1428 28980 1484
rect 29372 1428 29428 1484
rect 30884 1652 30940 1708
rect 26348 1146 26404 1148
rect 26348 1094 26350 1146
rect 26350 1094 26402 1146
rect 26402 1094 26404 1146
rect 26348 1092 26404 1094
rect 29484 1034 29540 1036
rect 29484 982 29486 1034
rect 29486 982 29538 1034
rect 29538 982 29540 1034
rect 29484 980 29540 982
rect 26196 810 26252 812
rect 26196 758 26198 810
rect 26198 758 26250 810
rect 26250 758 26252 810
rect 26196 756 26252 758
rect 26300 810 26356 812
rect 26300 758 26302 810
rect 26302 758 26354 810
rect 26354 758 26356 810
rect 26300 756 26356 758
rect 26404 810 26460 812
rect 26404 758 26406 810
rect 26406 758 26458 810
rect 26458 758 26460 810
rect 26404 756 26460 758
rect 30472 1594 30528 1596
rect 30472 1542 30474 1594
rect 30474 1542 30526 1594
rect 30526 1542 30528 1594
rect 30472 1540 30528 1542
rect 30576 1594 30632 1596
rect 30576 1542 30578 1594
rect 30578 1542 30630 1594
rect 30630 1542 30632 1594
rect 30576 1540 30632 1542
rect 30680 1594 30736 1596
rect 30680 1542 30682 1594
rect 30682 1542 30734 1594
rect 30734 1542 30736 1594
rect 30680 1540 30736 1542
rect 30716 1204 30772 1260
rect 31108 2772 31164 2828
rect 31444 2996 31500 3052
rect 31500 1540 31556 1596
rect 32564 8276 32620 8316
rect 32564 8260 32566 8276
rect 32566 8260 32618 8276
rect 32618 8260 32620 8276
rect 32564 5908 32620 5964
rect 32564 5684 32620 5740
rect 33180 9994 33236 9996
rect 33180 9942 33182 9994
rect 33182 9942 33234 9994
rect 33234 9942 33236 9994
rect 33180 9940 33236 9942
rect 33796 10052 33852 10108
rect 33348 9828 33404 9884
rect 33684 9882 33740 9884
rect 33684 9830 33686 9882
rect 33686 9830 33738 9882
rect 33738 9830 33740 9882
rect 33684 9828 33740 9830
rect 33012 8484 33068 8540
rect 33348 8932 33404 8988
rect 32788 8372 32844 8428
rect 33684 8194 33686 8204
rect 33686 8194 33738 8204
rect 33738 8194 33740 8204
rect 33684 8148 33740 8194
rect 33124 6692 33180 6748
rect 33348 6692 33404 6748
rect 33908 6692 33964 6748
rect 33572 6468 33628 6524
rect 33348 5012 33404 5068
rect 33236 4954 33292 4956
rect 33236 4902 33238 4954
rect 33238 4902 33290 4954
rect 33290 4902 33292 4954
rect 33236 4900 33292 4902
rect 32564 4116 32620 4172
rect 33236 4116 33292 4172
rect 33236 2660 33292 2716
rect 33684 5796 33740 5852
rect 34132 6580 34188 6636
rect 33796 5684 33852 5740
rect 34580 9940 34636 9996
rect 34356 9716 34412 9772
rect 34356 7812 34412 7868
rect 34356 6626 34358 6636
rect 34358 6626 34410 6636
rect 34410 6626 34412 6636
rect 34356 6580 34412 6626
rect 34468 6468 34524 6524
rect 34244 5572 34300 5628
rect 34356 5908 34412 5964
rect 34300 5290 34356 5292
rect 34300 5238 34302 5290
rect 34302 5238 34354 5290
rect 34354 5238 34356 5290
rect 34300 5236 34356 5238
rect 33796 5058 33798 5068
rect 33798 5058 33850 5068
rect 33850 5058 33852 5068
rect 33796 5012 33852 5058
rect 33908 4900 33964 4956
rect 34580 5236 34636 5292
rect 34580 4340 34636 4396
rect 34244 4228 34300 4284
rect 34412 3610 34468 3612
rect 34412 3558 34414 3610
rect 34414 3558 34466 3610
rect 34466 3558 34468 3610
rect 34412 3556 34468 3558
rect 33460 2660 33516 2716
rect 33460 1652 33516 1708
rect 32788 1214 32844 1260
rect 33516 1370 33572 1372
rect 33516 1318 33518 1370
rect 33518 1318 33570 1370
rect 33570 1318 33572 1370
rect 33516 1316 33572 1318
rect 32788 1204 32790 1214
rect 32790 1204 32842 1214
rect 32842 1204 32844 1214
rect 31892 1132 31894 1148
rect 31894 1132 31946 1148
rect 31946 1132 31948 1148
rect 31892 1092 31948 1132
rect 32228 1146 32284 1148
rect 32228 1094 32230 1146
rect 32230 1094 32282 1146
rect 32282 1094 32284 1146
rect 32228 1092 32284 1094
rect 33124 1092 33180 1148
rect 30716 1034 30772 1036
rect 30716 982 30718 1034
rect 30718 982 30770 1034
rect 30770 982 30772 1034
rect 30716 980 30772 982
rect 33796 2714 33852 2716
rect 33796 2662 33798 2714
rect 33798 2662 33850 2714
rect 33850 2662 33852 2714
rect 33796 2660 33852 2662
rect 34468 2938 34524 2940
rect 34468 2886 34470 2938
rect 34470 2886 34522 2938
rect 34522 2886 34524 2938
rect 34468 2884 34524 2886
rect 34468 2154 34524 2156
rect 34468 2102 34470 2154
rect 34470 2102 34522 2154
rect 34522 2102 34524 2154
rect 34468 2100 34524 2102
rect 34692 1316 34748 1372
rect 33684 980 33740 1036
rect 33852 1034 33908 1036
rect 33852 982 33854 1034
rect 33854 982 33906 1034
rect 33906 982 33908 1034
rect 33852 980 33908 982
rect 30100 868 30156 924
rect 34468 644 34524 700
rect 29988 532 30044 588
<< metal3 >>
rect 35200 13132 36000 13160
rect 31994 13076 32004 13132
rect 32060 13076 36000 13132
rect 35200 13048 36000 13076
rect 4806 12516 4816 12572
rect 4872 12516 4920 12572
rect 4976 12516 5024 12572
rect 5080 12516 5090 12572
rect 13358 12516 13368 12572
rect 13424 12516 13472 12572
rect 13528 12516 13576 12572
rect 13632 12516 13642 12572
rect 21910 12516 21920 12572
rect 21976 12516 22024 12572
rect 22080 12516 22128 12572
rect 22184 12516 22194 12572
rect 30462 12516 30472 12572
rect 30528 12516 30576 12572
rect 30632 12516 30680 12572
rect 30736 12516 30746 12572
rect 21466 12404 21476 12460
rect 21532 12404 28308 12460
rect 28364 12404 28374 12460
rect 12394 12292 12404 12348
rect 12460 12292 12852 12348
rect 12908 12292 12918 12348
rect 18330 12292 18340 12348
rect 18396 12292 21420 12348
rect 21476 12292 21486 12348
rect 1810 12180 1820 12236
rect 1876 12180 2548 12236
rect 2604 12180 2614 12236
rect 13346 12180 13356 12236
rect 13412 12180 22148 12236
rect 22204 12180 22214 12236
rect 24154 12180 24164 12236
rect 24220 12180 32676 12236
rect 32732 12180 32742 12236
rect 9930 12068 9940 12124
rect 9996 12068 10388 12124
rect 10444 12068 10454 12124
rect 11834 12068 11844 12124
rect 11900 12068 13244 12124
rect 14074 12068 14084 12124
rect 14140 12068 15316 12124
rect 15372 12068 15988 12124
rect 16044 12068 16054 12124
rect 18946 12068 18956 12124
rect 19012 12068 25396 12124
rect 25452 12068 25462 12124
rect 13188 12012 13244 12068
rect 11386 11956 11396 12012
rect 11452 11956 13020 12012
rect 13076 11956 13086 12012
rect 13178 11956 13188 12012
rect 13244 11956 14756 12012
rect 14812 11956 14822 12012
rect 22138 11956 22148 12012
rect 22204 11956 30268 12012
rect 30324 11956 30334 12012
rect 8372 11844 13356 11900
rect 13412 11844 13422 11900
rect 14410 11844 14420 11900
rect 14476 11844 18004 11900
rect 18060 11844 18070 11900
rect 21802 11844 21812 11900
rect 21868 11844 23940 11900
rect 23996 11844 24006 11900
rect 26058 11844 26068 11900
rect 26124 11844 30660 11900
rect 30716 11844 30726 11900
rect 8372 11788 8428 11844
rect 7690 11732 7700 11788
rect 7756 11732 8372 11788
rect 8428 11732 8438 11788
rect 9082 11732 9092 11788
rect 9148 11732 9196 11788
rect 9252 11732 9300 11788
rect 9356 11732 9366 11788
rect 9930 11732 9940 11788
rect 9996 11732 11172 11788
rect 11228 11732 11238 11788
rect 11722 11732 11732 11788
rect 11788 11732 13804 11788
rect 13860 11732 13870 11788
rect 17634 11732 17644 11788
rect 17700 11732 17748 11788
rect 17804 11732 17852 11788
rect 17908 11732 17918 11788
rect 19730 11732 19740 11788
rect 19852 11732 19862 11788
rect 26186 11732 26196 11788
rect 26252 11732 26300 11788
rect 26356 11732 26404 11788
rect 26460 11732 26470 11788
rect 29922 11732 29932 11788
rect 29988 11732 31332 11788
rect 31388 11732 31398 11788
rect 2146 11620 2156 11676
rect 2212 11620 2828 11676
rect 2884 11620 3892 11676
rect 3948 11620 3958 11676
rect 10266 11620 10276 11676
rect 10332 11620 11004 11676
rect 11060 11620 11070 11676
rect 12030 11620 12068 11676
rect 12124 11620 12134 11676
rect 13636 11620 17052 11676
rect 17108 11620 17332 11676
rect 17388 11620 17398 11676
rect 13636 11564 13692 11620
rect 6906 11508 6916 11564
rect 6972 11508 8372 11564
rect 8428 11508 8438 11564
rect 9930 11508 9940 11564
rect 9996 11508 10500 11564
rect 10556 11508 10566 11564
rect 10826 11508 10836 11564
rect 10892 11508 11396 11564
rect 11452 11508 11956 11564
rect 12012 11508 12022 11564
rect 12842 11508 12852 11564
rect 12908 11508 13636 11564
rect 13692 11508 13702 11564
rect 13962 11508 13972 11564
rect 14028 11508 14756 11564
rect 14812 11508 16492 11564
rect 16548 11508 16558 11564
rect 17882 11508 17892 11564
rect 17948 11508 19404 11564
rect 19460 11508 19470 11564
rect 24490 11508 24500 11564
rect 24556 11508 29428 11564
rect 29484 11508 29494 11564
rect 1082 11396 1092 11452
rect 1148 11396 1372 11452
rect 1428 11396 2604 11452
rect 2660 11396 3276 11452
rect 3332 11396 4340 11452
rect 4396 11396 4406 11452
rect 8698 11396 8708 11452
rect 8764 11396 10612 11452
rect 10668 11396 10678 11452
rect 10994 11396 11004 11452
rect 11060 11396 11788 11452
rect 12058 11396 12068 11452
rect 12124 11396 17444 11452
rect 17500 11396 17510 11452
rect 18778 11396 18788 11452
rect 18844 11396 19292 11452
rect 19348 11396 19358 11452
rect 20010 11396 20020 11452
rect 20076 11396 20132 11452
rect 20188 11396 20916 11452
rect 20972 11396 20982 11452
rect 24714 11396 24724 11452
rect 24780 11396 26068 11452
rect 26124 11396 26134 11452
rect 26730 11396 26740 11452
rect 26796 11396 28588 11452
rect 28644 11396 28654 11452
rect 11732 11340 11788 11396
rect 35200 11340 36000 11368
rect 3994 11284 4004 11340
rect 4060 11284 4788 11340
rect 4844 11284 4854 11340
rect 9426 11284 9436 11340
rect 9492 11284 11508 11340
rect 11564 11284 11574 11340
rect 11732 11284 14196 11340
rect 14252 11284 14262 11340
rect 23930 11284 23940 11340
rect 23996 11284 27188 11340
rect 27244 11284 27254 11340
rect 27626 11284 27636 11340
rect 27692 11284 28980 11340
rect 29036 11284 29428 11340
rect 29484 11284 30044 11340
rect 30100 11284 30110 11340
rect 32778 11284 32788 11340
rect 32844 11284 36000 11340
rect 27636 11228 27692 11284
rect 35200 11256 36000 11284
rect 3882 11172 3892 11228
rect 3948 11172 4900 11228
rect 4956 11172 7140 11228
rect 7196 11172 7588 11228
rect 7644 11172 7654 11228
rect 9090 11172 9100 11228
rect 9156 11172 16436 11228
rect 16492 11172 16502 11228
rect 19786 11172 19796 11228
rect 19852 11172 21588 11228
rect 21644 11172 21654 11228
rect 25162 11172 25172 11228
rect 25228 11172 25788 11228
rect 25844 11172 25854 11228
rect 26954 11172 26964 11228
rect 27020 11172 27692 11228
rect 8362 11060 8372 11116
rect 8428 11060 13972 11116
rect 14028 11060 14038 11116
rect 14186 11060 14196 11116
rect 14252 11060 22708 11116
rect 22764 11060 22774 11116
rect 4806 10948 4816 11004
rect 4872 10948 4920 11004
rect 4976 10948 5024 11004
rect 5080 10948 5090 11004
rect 7242 10948 7252 11004
rect 7308 10948 10948 11004
rect 11004 10948 11014 11004
rect 13358 10948 13368 11004
rect 13424 10948 13472 11004
rect 13528 10948 13576 11004
rect 13632 10948 13642 11004
rect 21910 10948 21920 11004
rect 21976 10948 22024 11004
rect 22080 10948 22128 11004
rect 22184 10948 22194 11004
rect 30462 10948 30472 11004
rect 30528 10948 30576 11004
rect 30632 10948 30680 11004
rect 30736 10948 30746 11004
rect 1698 10836 1708 10892
rect 1764 10836 5964 10892
rect 6020 10836 14644 10892
rect 14700 10836 14868 10892
rect 14924 10836 17052 10892
rect 17108 10836 17118 10892
rect 17434 10836 17444 10892
rect 17500 10836 20020 10892
rect 20076 10836 24724 10892
rect 24780 10836 24790 10892
rect 9538 10724 9548 10780
rect 9604 10724 10724 10780
rect 10780 10724 10790 10780
rect 12394 10724 12404 10780
rect 12460 10724 13804 10780
rect 13860 10724 14980 10780
rect 15036 10724 15046 10780
rect 19618 10724 19628 10780
rect 19684 10724 21812 10780
rect 21868 10724 29764 10780
rect 29820 10724 29830 10780
rect 4330 10612 4340 10668
rect 4396 10612 6412 10668
rect 6468 10612 6478 10668
rect 8754 10612 8764 10668
rect 8820 10612 16324 10668
rect 16380 10612 16390 10668
rect 17770 10612 17780 10668
rect 17836 10612 22036 10668
rect 22092 10612 22102 10668
rect 22698 10612 22708 10668
rect 22764 10612 26012 10668
rect 26068 10612 26078 10668
rect 1540 10500 8036 10556
rect 8092 10500 8102 10556
rect 8978 10500 8988 10556
rect 9044 10500 10948 10556
rect 11004 10500 11014 10556
rect 14074 10500 14084 10556
rect 14140 10500 18452 10556
rect 18508 10500 18518 10556
rect 22586 10500 22596 10556
rect 22652 10500 25732 10556
rect 25788 10500 25798 10556
rect 29754 10500 29764 10556
rect 29820 10500 30996 10556
rect 31052 10500 32340 10556
rect 32396 10500 32406 10556
rect 1540 10444 1596 10500
rect 1530 10388 1540 10444
rect 1596 10388 1606 10444
rect 3322 10388 3332 10444
rect 3388 10388 5068 10444
rect 5124 10388 5134 10444
rect 6122 10388 6132 10444
rect 6188 10388 7476 10444
rect 7532 10388 7542 10444
rect 9146 10388 9156 10444
rect 9212 10388 10612 10444
rect 10668 10388 10678 10444
rect 15988 10388 17332 10444
rect 17388 10388 19684 10444
rect 19740 10388 19750 10444
rect 22810 10388 22820 10444
rect 22876 10388 23492 10444
rect 23548 10388 23558 10444
rect 24994 10388 25004 10444
rect 25060 10388 26068 10444
rect 26124 10388 26292 10444
rect 26348 10388 26358 10444
rect 3658 10276 3668 10332
rect 3724 10276 14532 10332
rect 14588 10276 14598 10332
rect 14858 10276 14868 10332
rect 14924 10276 15484 10332
rect 15540 10276 15550 10332
rect 15988 10220 16044 10388
rect 4778 10164 4788 10220
rect 4844 10164 6076 10220
rect 6132 10164 6142 10220
rect 7242 10164 7252 10220
rect 7308 10164 7532 10220
rect 7588 10164 7598 10220
rect 9082 10164 9092 10220
rect 9148 10164 9196 10220
rect 9252 10164 9300 10220
rect 9356 10164 9366 10220
rect 9902 10164 9940 10220
rect 9996 10164 10006 10220
rect 15866 10164 15876 10220
rect 15932 10164 16044 10220
rect 5898 10052 5908 10108
rect 5964 10052 6916 10108
rect 6972 10052 6982 10108
rect 7130 10052 7140 10108
rect 7196 10052 7234 10108
rect 7914 10052 7924 10108
rect 7980 10052 11340 10108
rect 11284 9996 11340 10052
rect 16324 9996 16380 10332
rect 16436 10276 16446 10332
rect 17434 10276 17444 10332
rect 17500 10276 21588 10332
rect 21644 10276 21654 10332
rect 17634 10164 17644 10220
rect 17700 10164 17748 10220
rect 17804 10164 17852 10220
rect 17908 10164 17918 10220
rect 26186 10164 26196 10220
rect 26252 10164 26300 10220
rect 26356 10164 26404 10220
rect 26460 10164 26470 10220
rect 16874 10052 16884 10108
rect 16940 10052 19684 10108
rect 19740 10052 19750 10108
rect 24164 10052 25004 10108
rect 25060 10052 25070 10108
rect 25498 10052 25508 10108
rect 25564 10052 28196 10108
rect 28252 10052 28262 10108
rect 28522 10052 28532 10108
rect 28588 10052 31220 10108
rect 31276 10052 31286 10108
rect 31546 10052 31556 10108
rect 31612 10052 33796 10108
rect 33852 10052 33862 10108
rect 24164 9996 24220 10052
rect 5002 9940 5012 9996
rect 5068 9940 6468 9996
rect 6524 9940 6534 9996
rect 6626 9940 6636 9996
rect 6692 9940 7196 9996
rect 8082 9940 8092 9996
rect 8148 9940 8484 9996
rect 8540 9940 8550 9996
rect 8866 9940 8876 9996
rect 8932 9940 10276 9996
rect 10332 9940 10342 9996
rect 11274 9940 11284 9996
rect 11340 9940 11350 9996
rect 13514 9940 13524 9996
rect 13580 9940 14308 9996
rect 14364 9940 14374 9996
rect 14532 9940 16380 9996
rect 17658 9940 17668 9996
rect 17724 9940 18340 9996
rect 18396 9940 18732 9996
rect 19450 9940 19460 9996
rect 19516 9940 20076 9996
rect 20132 9940 20142 9996
rect 22418 9940 22428 9996
rect 22484 9940 24220 9996
rect 24378 9940 24388 9996
rect 24444 9940 26404 9996
rect 26460 9940 26470 9996
rect 26618 9940 26628 9996
rect 26684 9940 26694 9996
rect 33170 9940 33180 9996
rect 33236 9940 34580 9996
rect 34636 9940 34646 9996
rect 7140 9884 7196 9940
rect 14532 9884 14588 9940
rect 18676 9884 18732 9940
rect 26628 9884 26684 9940
rect 5730 9828 5740 9884
rect 5796 9828 6972 9884
rect 7028 9828 7038 9884
rect 7140 9828 9212 9884
rect 9268 9828 12180 9884
rect 12236 9828 14532 9884
rect 14588 9828 14598 9884
rect 14858 9828 14868 9884
rect 14924 9828 16380 9884
rect 16436 9828 16446 9884
rect 17042 9828 17052 9884
rect 17108 9828 17444 9884
rect 17500 9828 17836 9884
rect 17892 9828 17902 9884
rect 18050 9828 18060 9884
rect 18116 9828 18452 9884
rect 18508 9828 18518 9884
rect 18676 9828 20187 9884
rect 22586 9828 22596 9884
rect 22652 9828 26684 9884
rect 27010 9828 27020 9884
rect 27076 9828 29876 9884
rect 29932 9828 29942 9884
rect 31882 9828 31892 9884
rect 31948 9828 33348 9884
rect 33404 9828 33684 9884
rect 33740 9828 33750 9884
rect 20131 9772 20187 9828
rect 4554 9716 4564 9772
rect 4620 9716 5852 9772
rect 5908 9716 7140 9772
rect 7196 9716 7476 9772
rect 7532 9716 7756 9772
rect 7812 9716 7822 9772
rect 8250 9716 8260 9772
rect 8316 9716 10164 9772
rect 10220 9716 10230 9772
rect 12506 9716 12516 9772
rect 12572 9716 14644 9772
rect 14700 9716 14710 9772
rect 16930 9716 16940 9772
rect 7756 9660 7812 9716
rect 16996 9660 17052 9772
rect 18004 9716 19908 9772
rect 19964 9716 19974 9772
rect 20131 9716 21476 9772
rect 21532 9716 22428 9772
rect 22978 9716 22988 9772
rect 18004 9660 18060 9716
rect 22372 9660 22428 9716
rect 23044 9660 23100 9772
rect 25946 9716 25956 9772
rect 26012 9716 26572 9772
rect 26628 9716 26638 9772
rect 29418 9716 29428 9772
rect 29484 9716 30100 9772
rect 30156 9716 30166 9772
rect 32330 9716 32340 9772
rect 32396 9716 34356 9772
rect 34412 9716 34422 9772
rect 35200 9660 36000 9688
rect 2202 9604 2212 9660
rect 2268 9604 5124 9660
rect 5180 9604 5190 9660
rect 7756 9604 8708 9660
rect 8764 9604 8774 9660
rect 12674 9604 12684 9660
rect 12740 9604 13132 9660
rect 13188 9604 13198 9660
rect 14298 9604 14308 9660
rect 14364 9604 15092 9660
rect 15148 9604 18060 9660
rect 18274 9604 18284 9660
rect 18340 9604 19460 9660
rect 19516 9604 22036 9660
rect 22092 9604 22102 9660
rect 22362 9604 22372 9660
rect 22428 9604 22438 9660
rect 23044 9604 27860 9660
rect 27916 9604 27926 9660
rect 33674 9604 33684 9660
rect 33740 9604 36000 9660
rect 35200 9576 36000 9604
rect 2482 9492 2492 9548
rect 2548 9492 2996 9548
rect 3052 9492 5236 9548
rect 5292 9492 5302 9548
rect 7700 9492 9436 9548
rect 9492 9492 17668 9548
rect 17724 9492 17734 9548
rect 21690 9492 21700 9548
rect 21756 9492 23044 9548
rect 23100 9492 23110 9548
rect 7700 9436 7756 9492
rect 4806 9380 4816 9436
rect 4872 9380 4920 9436
rect 4976 9380 5024 9436
rect 5080 9380 5090 9436
rect 6458 9380 6468 9436
rect 6524 9380 6972 9436
rect 7028 9380 7038 9436
rect 7690 9380 7700 9436
rect 7756 9380 7766 9436
rect 13122 9380 13132 9436
rect 13188 9380 13244 9492
rect 13358 9380 13368 9436
rect 13424 9380 13472 9436
rect 13528 9380 13576 9436
rect 13632 9380 13642 9436
rect 15250 9380 15260 9436
rect 15316 9380 17556 9436
rect 17612 9380 17892 9436
rect 17948 9380 21700 9436
rect 21756 9380 21766 9436
rect 21910 9380 21920 9436
rect 21976 9380 22024 9436
rect 22080 9380 22128 9436
rect 22184 9380 22194 9436
rect 30462 9380 30472 9436
rect 30528 9380 30576 9436
rect 30632 9380 30680 9436
rect 30736 9380 30746 9436
rect 3098 9268 3108 9324
rect 3164 9268 9044 9324
rect 9100 9268 9110 9324
rect 10154 9268 10164 9324
rect 10220 9268 11956 9324
rect 12012 9268 12022 9324
rect 12226 9268 12236 9324
rect 12292 9268 13916 9324
rect 13972 9268 18004 9324
rect 18060 9268 26740 9324
rect 26796 9268 26852 9324
rect 26908 9268 26918 9324
rect 5114 9156 5124 9212
rect 5180 9156 6188 9212
rect 6244 9156 7252 9212
rect 7308 9156 7318 9212
rect 7476 9156 8820 9212
rect 8876 9156 8886 9212
rect 10266 9156 10276 9212
rect 10332 9156 10342 9212
rect 11554 9156 11564 9212
rect 11620 9156 12908 9212
rect 12964 9156 12974 9212
rect 15418 9156 15428 9212
rect 15484 9156 17108 9212
rect 17164 9156 17174 9212
rect 17434 9156 17444 9212
rect 17500 9156 18004 9212
rect 18060 9156 18070 9212
rect 18442 9156 18452 9212
rect 18508 9156 20187 9212
rect 21690 9156 21700 9212
rect 21756 9156 23716 9212
rect 23772 9156 23782 9212
rect 26618 9156 26628 9212
rect 26684 9156 29316 9212
rect 29372 9156 29382 9212
rect 1306 9044 1316 9100
rect 1372 9044 1932 9100
rect 1988 9044 2492 9100
rect 2548 9044 2558 9100
rect 2650 9044 2660 9100
rect 2716 9044 3892 9100
rect 3948 9044 3958 9100
rect 6514 9044 6524 9100
rect 6636 9044 6646 9100
rect 7476 8988 7532 9156
rect 8362 9044 8372 9100
rect 8428 9044 8438 9100
rect 8586 9044 8596 9100
rect 8652 9044 9212 9100
rect 9268 9044 9278 9100
rect 970 8932 980 8988
rect 1036 8932 3332 8988
rect 3388 8932 3464 8988
rect 4900 8876 4956 8988
rect 5012 8932 5460 8988
rect 5516 8932 5908 8988
rect 5964 8932 5974 8988
rect 6132 8932 6860 8988
rect 6916 8932 7532 8988
rect 6132 8876 6188 8932
rect 8372 8876 8428 9044
rect 10276 8988 10332 9156
rect 20131 9100 20187 9156
rect 11162 9044 11172 9100
rect 11228 9044 12684 9100
rect 12740 9044 12750 9100
rect 16314 9044 16324 9100
rect 16380 9044 17220 9100
rect 17276 9044 19908 9100
rect 19964 9044 19974 9100
rect 20131 9044 21868 9100
rect 22698 9044 22708 9100
rect 22764 9044 22774 9100
rect 29530 9044 29540 9100
rect 29596 9044 30324 9100
rect 30380 9044 31164 9100
rect 10276 8932 10500 8988
rect 10556 8932 11284 8988
rect 11340 8932 11350 8988
rect 11722 8932 11732 8988
rect 11788 8932 12068 8988
rect 12124 8932 14308 8988
rect 14364 8932 14374 8988
rect 16426 8932 16436 8988
rect 16492 8932 17444 8988
rect 17500 8932 17510 8988
rect 18340 8932 20748 8988
rect 20804 8932 20814 8988
rect 18340 8876 18396 8932
rect 21812 8876 21868 9044
rect 22708 8988 22764 9044
rect 31108 8988 31164 9044
rect 22138 8932 22148 8988
rect 22204 8932 22764 8988
rect 25946 8932 25956 8988
rect 26012 8932 26516 8988
rect 26572 8932 27580 8988
rect 31098 8932 31108 8988
rect 31164 8932 31174 8988
rect 31770 8932 31780 8988
rect 31836 8932 33348 8988
rect 33404 8932 33414 8988
rect 27524 8876 27580 8932
rect 2650 8820 2660 8876
rect 2716 8820 2996 8876
rect 3052 8820 4956 8876
rect 5226 8820 5236 8876
rect 5292 8820 6188 8876
rect 7130 8820 7140 8876
rect 7196 8820 7924 8876
rect 7980 8820 7990 8876
rect 8372 8820 9324 8876
rect 9380 8820 11732 8876
rect 11788 8820 11798 8876
rect 12394 8820 12404 8876
rect 12460 8820 14084 8876
rect 14140 8820 14150 8876
rect 15754 8820 15764 8876
rect 15820 8820 16548 8876
rect 16604 8820 16614 8876
rect 17882 8820 17892 8876
rect 17948 8820 17958 8876
rect 18330 8820 18340 8876
rect 18396 8820 18406 8876
rect 18564 8820 18844 8876
rect 18900 8820 19684 8876
rect 19740 8820 19750 8876
rect 20234 8820 20244 8876
rect 20300 8820 21644 8876
rect 21700 8820 21710 8876
rect 21812 8820 22820 8876
rect 22876 8820 22886 8876
rect 26058 8820 26068 8876
rect 26124 8820 27188 8876
rect 27244 8820 27254 8876
rect 27514 8820 27524 8876
rect 27580 8820 30100 8876
rect 30156 8820 30166 8876
rect 17892 8764 17948 8820
rect 18564 8764 18620 8820
rect 2258 8708 2268 8764
rect 2324 8708 3387 8764
rect 4386 8708 4396 8764
rect 4452 8708 8036 8764
rect 8092 8708 16660 8764
rect 16716 8708 16940 8764
rect 16996 8708 17006 8764
rect 17444 8708 17948 8764
rect 18050 8708 18060 8764
rect 18116 8708 18620 8764
rect 20131 8708 20916 8764
rect 20972 8708 24388 8764
rect 24444 8708 25284 8764
rect 25340 8708 25350 8764
rect 3331 8652 3387 8708
rect 1474 8596 1484 8652
rect 1540 8596 2660 8652
rect 2716 8596 2726 8652
rect 3331 8596 4732 8652
rect 4788 8596 4798 8652
rect 9082 8596 9092 8652
rect 9148 8596 9196 8652
rect 9252 8596 9300 8652
rect 9356 8596 9366 8652
rect 10490 8596 10500 8652
rect 10556 8596 10892 8652
rect 10948 8596 10958 8652
rect 17444 8540 17500 8708
rect 20131 8652 20187 8708
rect 17634 8596 17644 8652
rect 17700 8596 17748 8652
rect 17804 8596 17852 8652
rect 17908 8596 17918 8652
rect 17994 8596 18004 8652
rect 18060 8596 20187 8652
rect 26186 8596 26196 8652
rect 26252 8596 26300 8652
rect 26356 8596 26404 8652
rect 26460 8596 26470 8652
rect 26851 8596 32452 8652
rect 32508 8596 32518 8652
rect 26851 8540 26907 8596
rect 8474 8484 8484 8540
rect 8540 8484 9772 8540
rect 9828 8484 11340 8540
rect 11396 8484 12068 8540
rect 12124 8484 12134 8540
rect 12226 8484 12236 8540
rect 12292 8484 13748 8540
rect 13804 8484 13814 8540
rect 17434 8484 17444 8540
rect 17500 8484 17510 8540
rect 20356 8484 21476 8540
rect 21532 8484 21542 8540
rect 23594 8484 23604 8540
rect 23660 8484 26907 8540
rect 27738 8484 27748 8540
rect 27804 8484 33012 8540
rect 33068 8484 33078 8540
rect 20356 8428 20412 8484
rect 5562 8372 5572 8428
rect 5628 8372 9044 8428
rect 9100 8372 12628 8428
rect 12684 8372 13188 8428
rect 13244 8372 13254 8428
rect 13636 8372 14476 8428
rect 15642 8372 15652 8428
rect 15708 8372 17892 8428
rect 17948 8372 20412 8428
rect 20570 8372 20580 8428
rect 20636 8372 20646 8428
rect 21018 8372 21028 8428
rect 21084 8372 25060 8428
rect 25116 8372 25126 8428
rect 26394 8372 26404 8428
rect 26460 8372 27860 8428
rect 27916 8372 27926 8428
rect 29838 8372 29876 8428
rect 29932 8372 29942 8428
rect 30202 8372 30212 8428
rect 30268 8372 31556 8428
rect 31612 8372 31622 8428
rect 31770 8372 31780 8428
rect 31836 8372 32788 8428
rect 32844 8372 32854 8428
rect 13636 8316 13692 8372
rect 14420 8316 14476 8372
rect 20580 8316 20636 8372
rect 4162 8260 4172 8316
rect 4228 8260 5964 8316
rect 7018 8260 7028 8316
rect 7084 8260 7700 8316
rect 7756 8260 7766 8316
rect 8362 8260 8372 8316
rect 8484 8260 8494 8316
rect 9986 8260 9996 8316
rect 10052 8260 10612 8316
rect 10668 8260 10678 8316
rect 10910 8260 10948 8316
rect 11004 8260 11014 8316
rect 11890 8260 11900 8316
rect 11956 8260 13188 8316
rect 13244 8260 13356 8316
rect 13412 8260 13692 8316
rect 13794 8260 13804 8316
rect 13860 8260 14196 8316
rect 14252 8260 14262 8316
rect 14420 8260 15147 8316
rect 16090 8260 16100 8316
rect 16156 8260 17332 8316
rect 17388 8260 17398 8316
rect 19338 8260 19348 8316
rect 19404 8260 20636 8316
rect 21186 8260 21196 8316
rect 21252 8260 24276 8316
rect 24332 8260 24342 8316
rect 26786 8260 26796 8316
rect 26852 8260 27972 8316
rect 28028 8260 28038 8316
rect 28196 8260 29316 8316
rect 29372 8260 32564 8316
rect 32620 8260 32630 8316
rect 3770 8036 3780 8092
rect 3836 8036 4788 8092
rect 4844 8036 4854 8092
rect 5908 7868 5964 8260
rect 15091 8204 15147 8260
rect 28196 8204 28252 8260
rect 7354 8148 7364 8204
rect 7420 8148 7868 8204
rect 7924 8148 7934 8204
rect 8026 8148 8036 8204
rect 8092 8148 8130 8204
rect 8250 8148 8260 8204
rect 8316 8148 9772 8204
rect 9828 8148 9838 8204
rect 10490 8148 10500 8204
rect 10556 8148 12236 8204
rect 12292 8148 12302 8204
rect 12394 8148 12404 8204
rect 12460 8148 14924 8204
rect 14980 8148 14990 8204
rect 15091 8148 15988 8204
rect 16044 8148 16054 8204
rect 20794 8148 20804 8204
rect 20860 8148 25172 8204
rect 25228 8148 25620 8204
rect 25676 8148 25686 8204
rect 26618 8148 26628 8204
rect 26684 8148 27020 8204
rect 27076 8148 27086 8204
rect 27402 8148 27412 8204
rect 27468 8148 28252 8204
rect 29306 8148 29316 8204
rect 29372 8148 31220 8204
rect 31276 8148 31286 8204
rect 33646 8148 33684 8204
rect 33740 8148 33750 8204
rect 6122 8036 6132 8092
rect 6188 8036 8708 8092
rect 8764 8036 9940 8092
rect 9996 8036 10006 8092
rect 10164 8036 13524 8092
rect 13580 8036 14084 8092
rect 14140 8036 14150 8092
rect 14298 8036 14308 8092
rect 14364 8036 15092 8092
rect 15148 8036 15158 8092
rect 20010 8036 20020 8092
rect 20076 8036 21588 8092
rect 21644 8036 22708 8092
rect 22764 8036 22774 8092
rect 25050 8036 25060 8092
rect 25116 8036 25508 8092
rect 25564 8036 26236 8092
rect 26292 8036 28980 8092
rect 29036 8036 30884 8092
rect 30940 8036 30950 8092
rect 10164 7980 10220 8036
rect 8810 7924 8820 7980
rect 8876 7924 9212 7980
rect 9268 7924 10220 7980
rect 10602 7924 10612 7980
rect 10668 7924 11340 7980
rect 11396 7924 11406 7980
rect 11610 7924 11620 7980
rect 11676 7924 12068 7980
rect 12124 7924 17500 7980
rect 19114 7924 19124 7980
rect 19180 7924 19684 7980
rect 19740 7924 20244 7980
rect 20300 7924 20310 7980
rect 20570 7924 20580 7980
rect 20636 7924 25284 7980
rect 25340 7924 26628 7980
rect 26684 7924 26694 7980
rect 17444 7868 17500 7924
rect 20580 7868 20636 7924
rect 35200 7868 36000 7896
rect 4806 7812 4816 7868
rect 4872 7812 4920 7868
rect 4976 7812 5024 7868
rect 5080 7812 5090 7868
rect 5908 7812 10388 7868
rect 10444 7812 11732 7868
rect 11788 7812 11798 7868
rect 11946 7812 11956 7868
rect 12012 7812 12516 7868
rect 12572 7812 12582 7868
rect 13358 7812 13368 7868
rect 13424 7812 13472 7868
rect 13528 7812 13576 7868
rect 13632 7812 13642 7868
rect 14578 7812 14588 7868
rect 14644 7812 17220 7868
rect 17276 7812 17286 7868
rect 17444 7812 20636 7868
rect 21910 7812 21920 7868
rect 21976 7812 22024 7868
rect 22080 7812 22128 7868
rect 22184 7812 22194 7868
rect 30462 7812 30472 7868
rect 30528 7812 30576 7868
rect 30632 7812 30680 7868
rect 30736 7812 30746 7868
rect 33786 7812 33796 7868
rect 33852 7812 34356 7868
rect 34412 7812 36000 7868
rect 35200 7784 36000 7812
rect 7858 7700 7868 7756
rect 7924 7700 13916 7756
rect 13972 7700 13982 7756
rect 14186 7700 14196 7756
rect 14252 7700 19124 7756
rect 19180 7700 19190 7756
rect 6010 7588 6020 7644
rect 6076 7588 7532 7644
rect 7588 7588 7598 7644
rect 10042 7588 10052 7644
rect 10108 7588 10948 7644
rect 11004 7588 11014 7644
rect 14074 7588 14084 7644
rect 14140 7588 15204 7644
rect 15260 7588 15270 7644
rect 15530 7588 15540 7644
rect 15596 7588 18508 7644
rect 18564 7588 19572 7644
rect 19628 7588 19638 7644
rect 24826 7588 24836 7644
rect 24892 7588 30884 7644
rect 30940 7588 31444 7644
rect 31500 7588 31510 7644
rect 3994 7476 4004 7532
rect 4060 7476 5180 7532
rect 5236 7476 8484 7532
rect 8540 7476 8550 7532
rect 9426 7476 9436 7532
rect 9492 7476 11172 7532
rect 11228 7476 11238 7532
rect 13178 7476 13188 7532
rect 13244 7476 13916 7532
rect 13972 7476 13982 7532
rect 14186 7476 14196 7532
rect 14252 7476 15316 7532
rect 15372 7476 15382 7532
rect 15978 7476 15988 7532
rect 16044 7476 16660 7532
rect 16716 7476 16726 7532
rect 21354 7476 21364 7532
rect 21420 7476 22708 7532
rect 22764 7476 22774 7532
rect 25722 7476 25732 7532
rect 25788 7476 26516 7532
rect 26572 7476 26582 7532
rect 8586 7364 8596 7420
rect 8652 7364 9660 7420
rect 9716 7364 10388 7420
rect 10444 7364 12852 7420
rect 12908 7364 12918 7420
rect 17322 7364 17332 7420
rect 17388 7364 17556 7420
rect 17612 7364 17622 7420
rect 18666 7364 18676 7420
rect 18732 7364 21700 7420
rect 21756 7364 21766 7420
rect 25162 7364 25172 7420
rect 25228 7364 30268 7420
rect 30324 7364 30334 7420
rect 4666 7252 4676 7308
rect 4732 7252 5460 7308
rect 5516 7252 6412 7308
rect 6468 7252 7084 7308
rect 7140 7252 7150 7308
rect 11050 7252 11060 7308
rect 11116 7252 19348 7308
rect 19404 7252 19414 7308
rect 26730 7252 26740 7308
rect 26796 7252 27636 7308
rect 27692 7252 28756 7308
rect 28812 7252 30380 7308
rect 30436 7252 30446 7308
rect 3490 7140 3500 7196
rect 3556 7140 4172 7196
rect 4228 7140 4564 7196
rect 4620 7140 6860 7196
rect 6916 7140 9940 7196
rect 9996 7140 13188 7196
rect 13244 7140 14644 7196
rect 14700 7140 16100 7196
rect 16156 7140 18844 7196
rect 18900 7140 20020 7196
rect 20076 7140 20086 7196
rect 23034 7140 23044 7196
rect 23100 7140 25508 7196
rect 25564 7140 27076 7196
rect 27132 7140 27142 7196
rect 9082 7028 9092 7084
rect 9148 7028 9196 7084
rect 9252 7028 9300 7084
rect 9356 7028 9366 7084
rect 17634 7028 17644 7084
rect 17700 7028 17748 7084
rect 17804 7028 17852 7084
rect 17908 7028 17918 7084
rect 26186 7028 26196 7084
rect 26252 7028 26300 7084
rect 26356 7028 26404 7084
rect 26460 7028 26470 7084
rect 2650 6804 2660 6860
rect 2716 6804 3500 6860
rect 3556 6804 3566 6860
rect 13066 6804 13076 6860
rect 13132 6804 13580 6860
rect 13636 6804 13646 6860
rect 17210 6804 17220 6860
rect 17276 6804 19012 6860
rect 19068 6804 19078 6860
rect 26842 6804 26852 6860
rect 26908 6804 28084 6860
rect 28140 6804 31052 6860
rect 7074 6692 7084 6748
rect 7140 6692 7364 6748
rect 7420 6692 9716 6748
rect 9772 6692 9782 6748
rect 11386 6692 11396 6748
rect 11452 6692 11462 6748
rect 13066 6692 13076 6748
rect 13132 6692 13142 6748
rect 14046 6692 14084 6748
rect 14140 6692 14150 6748
rect 19562 6692 19572 6748
rect 19628 6692 20132 6748
rect 20188 6692 20198 6748
rect 21466 6692 21476 6748
rect 21532 6692 23492 6748
rect 23548 6692 27412 6748
rect 27468 6692 27478 6748
rect 1082 6580 1092 6636
rect 1148 6580 3276 6636
rect 3332 6580 3342 6636
rect 7690 6580 7700 6636
rect 7756 6580 8596 6636
rect 8652 6580 8662 6636
rect 11396 6412 11452 6692
rect 13076 6636 13132 6692
rect 12562 6580 12572 6636
rect 12628 6580 17444 6636
rect 17500 6580 17510 6636
rect 19394 6580 19404 6636
rect 19516 6580 19526 6636
rect 22810 6580 22820 6636
rect 22876 6580 23492 6636
rect 23548 6580 23558 6636
rect 24322 6580 24332 6636
rect 24444 6580 24454 6636
rect 24546 6580 24556 6636
rect 24612 6580 24668 6692
rect 30996 6636 31052 6804
rect 33114 6692 33124 6748
rect 33180 6692 33190 6748
rect 33338 6692 33348 6748
rect 33404 6692 33908 6748
rect 33964 6692 33974 6748
rect 33124 6636 33180 6692
rect 30986 6580 30996 6636
rect 31052 6580 34132 6636
rect 34188 6580 34198 6636
rect 34318 6580 34356 6636
rect 34412 6580 34422 6636
rect 11722 6468 11732 6524
rect 11788 6468 13076 6524
rect 13132 6468 13142 6524
rect 14074 6468 14084 6524
rect 14140 6468 16324 6524
rect 16380 6468 18004 6524
rect 18060 6468 18070 6524
rect 18386 6468 18396 6524
rect 18452 6468 19684 6524
rect 19740 6468 19852 6524
rect 19908 6468 22092 6524
rect 22148 6468 22158 6524
rect 22474 6468 22484 6524
rect 22540 6468 25396 6524
rect 25452 6468 25462 6524
rect 33562 6468 33572 6524
rect 33628 6468 34468 6524
rect 34524 6468 34534 6524
rect 9706 6356 9716 6412
rect 9772 6356 12852 6412
rect 12908 6356 14588 6412
rect 14644 6356 15876 6412
rect 15932 6356 16660 6412
rect 16716 6356 17444 6412
rect 17500 6356 18620 6412
rect 18676 6356 19684 6412
rect 19740 6356 19750 6412
rect 21802 6356 21812 6412
rect 21868 6356 24388 6412
rect 24444 6356 24454 6412
rect 4806 6244 4816 6300
rect 4872 6244 4920 6300
rect 4976 6244 5024 6300
rect 5080 6244 5090 6300
rect 12730 6244 12740 6300
rect 12796 6244 13188 6300
rect 13244 6244 13254 6300
rect 13358 6244 13368 6300
rect 13424 6244 13472 6300
rect 13528 6244 13576 6300
rect 13632 6244 13642 6300
rect 21910 6244 21920 6300
rect 21976 6244 22024 6300
rect 22080 6244 22128 6300
rect 22184 6244 22194 6300
rect 28634 6244 28644 6300
rect 28700 6244 29876 6300
rect 29932 6244 29942 6300
rect 30462 6244 30472 6300
rect 30528 6244 30576 6300
rect 30632 6244 30680 6300
rect 30736 6244 30746 6300
rect 7102 6132 7140 6188
rect 7196 6132 7206 6188
rect 29642 6132 29652 6188
rect 29708 6132 32116 6188
rect 32172 6132 32182 6188
rect 35200 6076 36000 6104
rect 6234 6020 6244 6076
rect 6300 6020 9044 6076
rect 9100 6020 9110 6076
rect 13066 6020 13076 6076
rect 13132 6020 13972 6076
rect 14028 6020 14038 6076
rect 27962 6020 27972 6076
rect 28028 6020 30884 6076
rect 30940 6020 30950 6076
rect 34346 6020 34356 6076
rect 34412 6020 36000 6076
rect 35200 5992 36000 6020
rect 6458 5908 6468 5964
rect 6524 5908 8708 5964
rect 8764 5908 8774 5964
rect 12506 5908 12516 5964
rect 12572 5908 13748 5964
rect 13804 5908 13814 5964
rect 14196 5908 14644 5964
rect 14700 5908 14710 5964
rect 25834 5908 25844 5964
rect 25900 5908 28420 5964
rect 28476 5908 29764 5964
rect 29820 5908 32564 5964
rect 32620 5908 34356 5964
rect 34412 5908 34422 5964
rect 14196 5852 14252 5908
rect 6178 5796 6188 5852
rect 6244 5796 9156 5852
rect 9212 5796 9222 5852
rect 12954 5796 12964 5852
rect 13020 5796 13188 5852
rect 13244 5796 13636 5852
rect 13692 5796 14252 5852
rect 14410 5796 14420 5852
rect 14476 5796 16212 5852
rect 16268 5796 16278 5852
rect 18834 5796 18844 5852
rect 18900 5796 19460 5852
rect 19516 5796 19908 5852
rect 19964 5796 19974 5852
rect 22810 5796 22820 5852
rect 22876 5796 23380 5852
rect 23436 5796 23446 5852
rect 26394 5796 26404 5852
rect 26460 5796 33684 5852
rect 33740 5796 33750 5852
rect 5562 5684 5572 5740
rect 5628 5684 7532 5740
rect 7588 5684 7598 5740
rect 8026 5684 8036 5740
rect 8092 5684 8764 5740
rect 8820 5684 9380 5740
rect 9436 5684 9940 5740
rect 9996 5684 10006 5740
rect 13794 5684 13804 5740
rect 13860 5684 15988 5740
rect 16044 5684 16054 5740
rect 28858 5684 28868 5740
rect 28924 5684 30212 5740
rect 30268 5684 30278 5740
rect 32554 5684 32564 5740
rect 32620 5684 33796 5740
rect 33852 5684 33862 5740
rect 7130 5572 7140 5628
rect 7196 5572 11676 5628
rect 11732 5572 11742 5628
rect 22250 5572 22260 5628
rect 22316 5572 26068 5628
rect 26124 5572 34244 5628
rect 34300 5572 34310 5628
rect 9082 5460 9092 5516
rect 9148 5460 9196 5516
rect 9252 5460 9300 5516
rect 9356 5460 9366 5516
rect 9594 5460 9604 5516
rect 9660 5460 10108 5516
rect 10164 5460 10174 5516
rect 17634 5460 17644 5516
rect 17700 5460 17748 5516
rect 17804 5460 17852 5516
rect 17908 5460 17918 5516
rect 23706 5460 23716 5516
rect 23772 5460 25396 5516
rect 25452 5460 25462 5516
rect 26186 5460 26196 5516
rect 26252 5460 26300 5516
rect 26356 5460 26404 5516
rect 26460 5460 26470 5516
rect 6066 5348 6076 5404
rect 6132 5348 10836 5404
rect 10892 5348 10902 5404
rect 19730 5348 19740 5404
rect 19796 5348 24108 5404
rect 25498 5348 25508 5404
rect 25564 5348 25956 5404
rect 26012 5348 26022 5404
rect 24052 5292 24108 5348
rect 5562 5236 5572 5292
rect 5628 5236 7700 5292
rect 7756 5236 7766 5292
rect 8306 5236 8316 5292
rect 8372 5236 8708 5292
rect 8764 5236 8774 5292
rect 9874 5236 9884 5292
rect 9940 5236 10332 5292
rect 12170 5236 12180 5292
rect 12236 5236 13804 5292
rect 13860 5236 13870 5292
rect 18330 5236 18340 5292
rect 18396 5236 23828 5292
rect 23884 5236 23894 5292
rect 24052 5236 27972 5292
rect 28028 5236 28038 5292
rect 34290 5236 34300 5292
rect 34356 5236 34580 5292
rect 34636 5236 34646 5292
rect 10276 5180 10332 5236
rect 5338 5124 5348 5180
rect 5404 5124 6860 5180
rect 6916 5124 6926 5180
rect 7242 5124 7252 5180
rect 7308 5124 8652 5180
rect 8708 5124 8718 5180
rect 9258 5124 9268 5180
rect 9324 5124 9996 5180
rect 10052 5124 10062 5180
rect 10276 5124 10388 5180
rect 10444 5124 12292 5180
rect 12348 5124 19404 5180
rect 24266 5124 24276 5180
rect 24332 5124 26404 5180
rect 26460 5124 26470 5180
rect 28130 5124 28140 5180
rect 28196 5124 29092 5180
rect 29148 5124 29158 5180
rect 19348 5068 19404 5124
rect 6346 5012 6356 5068
rect 6412 5012 7868 5068
rect 8446 5012 8484 5068
rect 8540 5012 8550 5068
rect 10154 5012 10164 5068
rect 10220 5012 10230 5068
rect 11050 5012 11060 5068
rect 11116 5012 12180 5068
rect 12236 5012 12246 5068
rect 12394 5012 12404 5068
rect 12460 5012 14308 5068
rect 14364 5012 14374 5068
rect 19338 5012 19348 5068
rect 19404 5012 23436 5068
rect 25386 5012 25396 5068
rect 25452 5012 26628 5068
rect 26684 5012 26694 5068
rect 33338 5012 33348 5068
rect 33404 5012 33796 5068
rect 33852 5012 33862 5068
rect 7812 4956 7868 5012
rect 10164 4956 10220 5012
rect 22932 4956 22988 5012
rect 23380 4956 23436 5012
rect 4666 4900 4676 4956
rect 4732 4900 5460 4956
rect 5516 4900 6916 4956
rect 6972 4900 6982 4956
rect 7802 4900 7812 4956
rect 7868 4900 7878 4956
rect 8362 4900 8372 4956
rect 8428 4900 9884 4956
rect 2090 4788 2100 4844
rect 2156 4788 8708 4844
rect 8764 4788 8774 4844
rect 9828 4732 9884 4900
rect 10052 4900 11900 4956
rect 11956 4900 11966 4956
rect 13402 4900 13412 4956
rect 13468 4900 15204 4956
rect 15260 4900 15270 4956
rect 19898 4900 19908 4956
rect 19964 4900 20356 4956
rect 20412 4900 20422 4956
rect 22922 4900 22932 4956
rect 22988 4900 22998 4956
rect 23380 4900 24108 4956
rect 24164 4900 24174 4956
rect 24322 4900 24332 4956
rect 24388 4900 27356 4956
rect 27412 4900 27422 4956
rect 28970 4900 28980 4956
rect 29092 4900 29102 4956
rect 29250 4900 29260 4956
rect 29372 4900 29382 4956
rect 33226 4900 33236 4956
rect 33292 4900 33908 4956
rect 33964 4900 33974 4956
rect 10052 4844 10108 4900
rect 10042 4788 10052 4844
rect 10108 4788 10118 4844
rect 10378 4788 10388 4844
rect 10444 4788 13804 4844
rect 14074 4788 14084 4844
rect 14140 4788 17500 4844
rect 17556 4788 18004 4844
rect 18060 4788 18070 4844
rect 26394 4788 26404 4844
rect 26460 4788 27076 4844
rect 27132 4788 27142 4844
rect 13748 4732 13804 4788
rect 4806 4676 4816 4732
rect 4872 4676 4920 4732
rect 4976 4676 5024 4732
rect 5080 4676 5090 4732
rect 6906 4676 6916 4732
rect 6972 4676 8260 4732
rect 8316 4676 8326 4732
rect 8558 4676 8596 4732
rect 8652 4676 8662 4732
rect 8922 4676 8932 4732
rect 8988 4676 9380 4732
rect 9436 4676 9446 4732
rect 9828 4676 9940 4732
rect 9996 4676 10006 4732
rect 10378 4676 10388 4732
rect 10444 4676 11228 4732
rect 11284 4676 11732 4732
rect 11788 4676 11798 4732
rect 11946 4676 11956 4732
rect 12012 4676 13244 4732
rect 13358 4676 13368 4732
rect 13424 4676 13472 4732
rect 13528 4676 13576 4732
rect 13632 4676 13642 4732
rect 13748 4676 15260 4732
rect 15316 4676 16380 4732
rect 17882 4676 17892 4732
rect 17948 4676 19012 4732
rect 19068 4676 19078 4732
rect 21910 4676 21920 4732
rect 21976 4676 22024 4732
rect 22080 4676 22128 4732
rect 22184 4676 22194 4732
rect 30462 4676 30472 4732
rect 30528 4676 30576 4732
rect 30632 4676 30680 4732
rect 30736 4676 30746 4732
rect 13188 4620 13244 4676
rect 16324 4620 16380 4676
rect 6234 4564 6244 4620
rect 6300 4564 6692 4620
rect 6748 4564 10500 4620
rect 10556 4564 10566 4620
rect 11498 4564 11508 4620
rect 11564 4564 12068 4620
rect 12124 4564 12134 4620
rect 13188 4564 13748 4620
rect 13804 4564 13814 4620
rect 14308 4564 16100 4620
rect 16156 4564 16166 4620
rect 16324 4564 18844 4620
rect 18900 4564 18910 4620
rect 19114 4564 19124 4620
rect 19180 4564 19796 4620
rect 19852 4564 19862 4620
rect 20010 4564 20020 4620
rect 20076 4564 20692 4620
rect 20748 4564 23156 4620
rect 23212 4564 24500 4620
rect 24556 4564 28532 4620
rect 28588 4564 29876 4620
rect 29932 4564 29942 4620
rect 13300 4508 13356 4564
rect 1754 4452 1764 4508
rect 1820 4452 5796 4508
rect 5852 4452 5862 4508
rect 7326 4452 7364 4508
rect 7420 4452 7430 4508
rect 7578 4452 7588 4508
rect 7644 4452 8036 4508
rect 8092 4452 8102 4508
rect 8250 4452 8260 4508
rect 8316 4452 9044 4508
rect 9100 4452 9604 4508
rect 9660 4452 9670 4508
rect 9930 4452 9940 4508
rect 9996 4452 11172 4508
rect 11228 4452 11238 4508
rect 13010 4452 13020 4508
rect 13132 4452 13142 4508
rect 13290 4452 13300 4508
rect 13356 4452 13366 4508
rect 13458 4452 13468 4508
rect 13524 4452 14084 4508
rect 14140 4452 14150 4508
rect 4778 4340 4788 4396
rect 4844 4340 5684 4396
rect 5740 4340 5750 4396
rect 7242 4340 7252 4396
rect 7308 4340 9492 4396
rect 9548 4340 10052 4396
rect 10108 4340 10118 4396
rect 10266 4340 10276 4396
rect 10332 4340 12404 4396
rect 12460 4340 13860 4396
rect 13916 4340 13926 4396
rect 14308 4284 14364 4564
rect 14746 4452 14756 4508
rect 14812 4452 15428 4508
rect 15484 4452 15494 4508
rect 15652 4452 19236 4508
rect 19292 4452 20692 4508
rect 20748 4452 20758 4508
rect 26506 4452 26516 4508
rect 26572 4452 27468 4508
rect 27524 4452 27534 4508
rect 15652 4396 15708 4452
rect 27860 4396 27916 4508
rect 27972 4452 30884 4508
rect 30940 4452 30950 4508
rect 35200 4396 36000 4424
rect 14634 4340 14644 4396
rect 14700 4340 15092 4396
rect 15148 4340 15708 4396
rect 17322 4340 17332 4396
rect 17388 4340 18004 4396
rect 18060 4340 18070 4396
rect 18834 4340 18844 4396
rect 18900 4340 19908 4396
rect 19964 4340 19974 4396
rect 20131 4340 20356 4396
rect 20412 4340 20422 4396
rect 20570 4340 20580 4396
rect 20636 4340 21084 4396
rect 21140 4340 22428 4396
rect 23034 4340 23044 4396
rect 23100 4340 24332 4396
rect 24388 4340 25956 4396
rect 26012 4340 27916 4396
rect 28410 4340 28420 4396
rect 28476 4340 29764 4396
rect 29820 4340 29830 4396
rect 34570 4340 34580 4396
rect 34636 4340 36000 4396
rect 20131 4284 20187 4340
rect 2202 4228 2212 4284
rect 2268 4228 7924 4284
rect 7980 4228 7990 4284
rect 9258 4228 9268 4284
rect 9324 4228 12348 4284
rect 12404 4228 12414 4284
rect 12964 4228 14364 4284
rect 15866 4228 15876 4284
rect 15932 4228 16716 4284
rect 16772 4228 20187 4284
rect 20244 4228 22036 4284
rect 22092 4228 22102 4284
rect 22372 4228 22428 4340
rect 35200 4312 36000 4340
rect 22484 4228 24836 4284
rect 24892 4228 24902 4284
rect 29016 4228 29092 4284
rect 29148 4228 34244 4284
rect 34300 4228 34310 4284
rect 9268 4172 9324 4228
rect 5226 4116 5236 4172
rect 5292 4116 9324 4172
rect 10490 4116 10500 4172
rect 10556 4116 11900 4172
rect 11956 4116 11966 4172
rect 12114 4116 12124 4172
rect 12180 4116 12628 4172
rect 12684 4116 12694 4172
rect 7588 4004 8484 4060
rect 8540 4004 9940 4060
rect 9996 4004 12740 4060
rect 12796 4004 12806 4060
rect 7588 3948 7644 4004
rect 12964 3948 13020 4228
rect 20244 4172 20300 4228
rect 13122 4116 13132 4172
rect 13244 4116 13254 4172
rect 13514 4116 13524 4172
rect 13580 4116 20300 4172
rect 20402 4116 20412 4172
rect 20468 4116 23212 4172
rect 23268 4116 23278 4172
rect 24042 4116 24052 4172
rect 24108 4116 28028 4172
rect 28084 4116 29820 4172
rect 29876 4116 29886 4172
rect 31546 4116 31556 4172
rect 31612 4116 32564 4172
rect 32620 4116 33236 4172
rect 33292 4116 33302 4172
rect 14914 4004 14924 4060
rect 14980 4004 15484 4060
rect 15540 4004 24948 4060
rect 25004 4004 25620 4060
rect 25676 4004 25686 4060
rect 26842 4004 26852 4060
rect 26908 4004 30044 4060
rect 30100 4004 30110 4060
rect 4162 3892 4172 3948
rect 4228 3892 7140 3948
rect 7196 3892 7206 3948
rect 7578 3892 7588 3948
rect 7644 3892 7654 3948
rect 9082 3892 9092 3948
rect 9148 3892 9196 3948
rect 9252 3892 9300 3948
rect 9356 3892 9366 3948
rect 9818 3892 9828 3948
rect 9884 3892 9894 3948
rect 10938 3892 10948 3948
rect 11004 3892 11676 3948
rect 12058 3892 12068 3948
rect 12124 3892 13020 3948
rect 13178 3892 13188 3948
rect 13244 3892 15876 3948
rect 15932 3892 15942 3948
rect 17634 3892 17644 3948
rect 17700 3892 17748 3948
rect 17804 3892 17852 3948
rect 17908 3892 17918 3948
rect 26186 3892 26196 3948
rect 26252 3892 26300 3948
rect 26356 3892 26404 3948
rect 26460 3892 26470 3948
rect 1530 3780 1540 3836
rect 1596 3780 3387 3836
rect 6178 3780 6188 3836
rect 6244 3780 8372 3836
rect 8428 3780 8438 3836
rect 8586 3780 8596 3836
rect 8652 3780 9548 3836
rect 9604 3780 9614 3836
rect 3331 3612 3387 3780
rect 9828 3724 9884 3892
rect 11620 3836 11676 3892
rect 11610 3780 11620 3836
rect 11676 3780 13524 3836
rect 13580 3780 13590 3836
rect 14410 3780 14420 3836
rect 14476 3780 14924 3836
rect 14980 3780 14990 3836
rect 21298 3780 21308 3836
rect 21364 3780 22484 3836
rect 22540 3780 24276 3836
rect 24332 3780 28868 3836
rect 28924 3780 28934 3836
rect 29614 3780 29652 3836
rect 29708 3780 29718 3836
rect 30426 3780 30436 3836
rect 30492 3780 31108 3836
rect 31164 3780 31174 3836
rect 4050 3668 4060 3724
rect 4116 3668 4564 3724
rect 4620 3668 4630 3724
rect 8026 3668 8036 3724
rect 8092 3668 9044 3724
rect 9100 3668 9110 3724
rect 9828 3668 10556 3724
rect 11722 3668 11732 3724
rect 11788 3668 16660 3724
rect 16716 3668 19012 3724
rect 19068 3668 19078 3724
rect 23370 3668 23380 3724
rect 23436 3668 25396 3724
rect 25452 3668 26907 3724
rect 27738 3668 27748 3724
rect 27804 3668 28196 3724
rect 28252 3668 30324 3724
rect 30380 3668 30390 3724
rect 3331 3556 9548 3612
rect 9930 3556 9940 3612
rect 9996 3556 10276 3612
rect 10332 3556 10342 3612
rect 9492 3500 9548 3556
rect 6850 3444 6860 3500
rect 6916 3444 7756 3500
rect 7970 3444 7980 3500
rect 8092 3444 8102 3500
rect 8632 3444 8708 3500
rect 8764 3444 9212 3500
rect 9482 3444 9492 3500
rect 9548 3444 9558 3500
rect 9706 3444 9716 3500
rect 9772 3444 10276 3500
rect 10332 3444 10342 3500
rect 7700 3388 7756 3444
rect 9156 3388 9212 3444
rect 10500 3388 10556 3668
rect 26851 3612 26907 3668
rect 11386 3556 11396 3612
rect 11452 3556 13804 3612
rect 13860 3556 14196 3612
rect 14252 3556 14262 3612
rect 21690 3556 21700 3612
rect 21756 3556 21766 3612
rect 21970 3556 21980 3612
rect 22036 3556 22596 3612
rect 22652 3556 22662 3612
rect 24826 3556 24836 3612
rect 24892 3556 26404 3612
rect 26460 3556 26470 3612
rect 26851 3556 27244 3612
rect 27300 3556 28700 3612
rect 28756 3556 29652 3612
rect 29708 3556 34412 3612
rect 34468 3556 34478 3612
rect 21700 3500 21756 3556
rect 10714 3444 10724 3500
rect 10780 3444 11508 3500
rect 11564 3444 11574 3500
rect 11834 3444 11844 3500
rect 11900 3444 14756 3500
rect 14812 3444 14822 3500
rect 15026 3444 15036 3500
rect 15092 3444 15708 3500
rect 15764 3444 15774 3500
rect 21298 3444 21308 3500
rect 21364 3444 22204 3500
rect 22260 3444 22270 3500
rect 23706 3444 23716 3500
rect 23772 3444 26516 3500
rect 26572 3444 26740 3500
rect 26796 3444 26806 3500
rect 28970 3444 28980 3500
rect 29036 3444 29988 3500
rect 30044 3444 30054 3500
rect 5114 3332 5124 3388
rect 5180 3332 5852 3388
rect 5908 3332 7420 3388
rect 7700 3332 9100 3388
rect 9156 3332 9940 3388
rect 9996 3332 10006 3388
rect 10500 3332 11116 3388
rect 11172 3332 11182 3388
rect 11722 3332 11732 3388
rect 11788 3332 11798 3388
rect 11946 3332 11956 3388
rect 12012 3332 12050 3388
rect 12170 3332 12180 3388
rect 12236 3332 12460 3388
rect 12516 3332 13076 3388
rect 13132 3332 13142 3388
rect 13850 3332 13860 3388
rect 13916 3332 15484 3388
rect 15540 3332 15550 3388
rect 16538 3332 16548 3388
rect 16604 3332 20916 3388
rect 20972 3332 21196 3388
rect 21252 3332 21262 3388
rect 25610 3332 25620 3388
rect 25676 3332 26124 3388
rect 26180 3332 26190 3388
rect 26394 3332 26404 3388
rect 26460 3332 29092 3388
rect 29148 3332 29158 3388
rect 29754 3332 29764 3388
rect 29820 3332 31052 3388
rect 7364 3276 7420 3332
rect 9044 3276 9100 3332
rect 7354 3220 7364 3276
rect 7420 3220 7756 3276
rect 8810 3220 8820 3276
rect 8876 3220 8886 3276
rect 9044 3220 9604 3276
rect 9660 3220 9670 3276
rect 7700 3164 7756 3220
rect 8820 3164 8876 3220
rect 11732 3164 11788 3332
rect 16548 3276 16604 3332
rect 30996 3276 31052 3332
rect 14298 3220 14308 3276
rect 14364 3220 16604 3276
rect 20346 3220 20356 3276
rect 20412 3220 21476 3276
rect 21532 3220 23716 3276
rect 23772 3220 23782 3276
rect 28522 3220 28532 3276
rect 28588 3220 29316 3276
rect 29372 3220 29382 3276
rect 29614 3220 29652 3276
rect 29708 3220 29718 3276
rect 30986 3220 30996 3276
rect 31052 3220 31062 3276
rect 4806 3108 4816 3164
rect 4872 3108 4920 3164
rect 4976 3108 5024 3164
rect 5080 3108 5090 3164
rect 7018 3108 7028 3164
rect 7084 3108 7476 3164
rect 7532 3108 7542 3164
rect 7690 3108 7700 3164
rect 7756 3108 7766 3164
rect 8820 3108 9044 3164
rect 9100 3108 11788 3164
rect 12730 3108 12740 3164
rect 12796 3108 13188 3164
rect 13244 3108 13254 3164
rect 13358 3108 13368 3164
rect 13424 3108 13472 3164
rect 13528 3108 13576 3164
rect 13632 3108 13642 3164
rect 19394 3108 19404 3164
rect 19460 3108 20132 3164
rect 20188 3108 20580 3164
rect 20636 3108 20646 3164
rect 21910 3108 21920 3164
rect 21976 3108 22024 3164
rect 22080 3108 22128 3164
rect 22184 3108 22194 3164
rect 26506 3108 26516 3164
rect 26572 3108 28196 3164
rect 28252 3108 28262 3164
rect 28858 3108 28868 3164
rect 28924 3108 29428 3164
rect 29484 3108 29494 3164
rect 30462 3108 30472 3164
rect 30528 3108 30576 3164
rect 30632 3108 30680 3164
rect 30736 3108 30746 3164
rect 1082 2996 1092 3052
rect 1148 2996 2100 3052
rect 2156 2996 3556 3052
rect 3612 2996 3622 3052
rect 8586 2996 8596 3052
rect 8652 2996 9156 3052
rect 9212 2996 9222 3052
rect 12954 2996 12964 3052
rect 13020 2996 14756 3052
rect 14812 2996 16884 3052
rect 16940 2996 16950 3052
rect 26618 2996 26628 3052
rect 26684 2996 26852 3052
rect 26908 2996 26918 3052
rect 27402 2996 27412 3052
rect 27468 2996 31444 3052
rect 31500 2996 31510 3052
rect 2874 2884 2884 2940
rect 2940 2884 7084 2940
rect 7140 2884 7150 2940
rect 7466 2884 7476 2940
rect 7532 2884 8036 2940
rect 8092 2884 8372 2940
rect 8428 2884 8438 2940
rect 10938 2884 10948 2940
rect 11004 2884 12292 2940
rect 12348 2884 12740 2940
rect 12796 2884 13356 2940
rect 13412 2884 13422 2940
rect 14522 2884 14532 2940
rect 14588 2884 16324 2940
rect 16380 2884 17556 2940
rect 17612 2884 18116 2940
rect 18172 2884 18182 2940
rect 26338 2884 26348 2940
rect 26404 2884 27524 2940
rect 27580 2884 34468 2940
rect 34524 2884 34534 2940
rect 7476 2828 7532 2884
rect 6234 2772 6244 2828
rect 6300 2772 7532 2828
rect 8474 2772 8484 2828
rect 8540 2772 9268 2828
rect 9324 2772 12964 2828
rect 13020 2772 13030 2828
rect 15978 2772 15988 2828
rect 16044 2772 16996 2828
rect 17052 2772 20020 2828
rect 20076 2772 20692 2828
rect 20748 2772 21588 2828
rect 21644 2772 21654 2828
rect 22250 2772 22260 2828
rect 22316 2772 23492 2828
rect 23548 2772 23558 2828
rect 25554 2772 25564 2828
rect 25620 2772 27412 2828
rect 27468 2772 27478 2828
rect 30874 2772 30884 2828
rect 30940 2772 31108 2828
rect 31164 2772 31174 2828
rect 5842 2660 5852 2716
rect 5908 2660 6468 2716
rect 6524 2660 6692 2716
rect 6748 2660 8036 2716
rect 8092 2660 8102 2716
rect 12506 2660 12516 2716
rect 12572 2660 13076 2716
rect 13132 2660 13580 2716
rect 13636 2660 14084 2716
rect 14140 2660 18452 2716
rect 18508 2660 19012 2716
rect 19068 2660 19078 2716
rect 23594 2660 23604 2716
rect 23660 2660 23940 2716
rect 23996 2660 24006 2716
rect 25666 2660 25676 2716
rect 25732 2660 28532 2716
rect 28588 2660 28598 2716
rect 29530 2660 29540 2716
rect 29596 2660 29876 2716
rect 29932 2660 29942 2716
rect 33226 2660 33236 2716
rect 33292 2660 33460 2716
rect 33516 2660 33796 2716
rect 33852 2660 33862 2716
rect 35200 2604 36000 2632
rect 7578 2548 7588 2604
rect 7644 2548 7812 2604
rect 7868 2548 11396 2604
rect 11452 2548 11462 2604
rect 13178 2548 13188 2604
rect 13244 2548 13972 2604
rect 14028 2548 14420 2604
rect 14476 2548 14486 2604
rect 16146 2548 16156 2604
rect 16212 2548 18788 2604
rect 18844 2548 18854 2604
rect 21858 2548 21868 2604
rect 21924 2548 23492 2604
rect 23548 2548 23558 2604
rect 23706 2548 23716 2604
rect 23772 2548 24332 2604
rect 24388 2548 24398 2604
rect 25106 2548 25116 2604
rect 25172 2548 25844 2604
rect 25900 2548 25910 2604
rect 26394 2548 26404 2604
rect 26460 2548 27188 2604
rect 27244 2548 27254 2604
rect 31891 2548 36000 2604
rect 31891 2492 31947 2548
rect 35200 2520 36000 2548
rect 3546 2436 3556 2492
rect 3612 2436 5348 2492
rect 5404 2436 8484 2492
rect 8540 2436 8550 2492
rect 12366 2436 12404 2492
rect 12460 2436 12470 2492
rect 18106 2436 18116 2492
rect 18172 2436 19068 2492
rect 19124 2436 19964 2492
rect 20020 2436 20030 2492
rect 23594 2436 23604 2492
rect 23660 2436 26740 2492
rect 26796 2436 28308 2492
rect 28364 2436 28374 2492
rect 29978 2436 29988 2492
rect 30044 2436 31947 2492
rect 9082 2324 9092 2380
rect 9148 2324 9196 2380
rect 9252 2324 9300 2380
rect 9356 2324 9366 2380
rect 12058 2324 12068 2380
rect 12124 2324 14588 2380
rect 14644 2324 14654 2380
rect 17634 2324 17644 2380
rect 17700 2324 17748 2380
rect 17804 2324 17852 2380
rect 17908 2324 17918 2380
rect 18834 2324 18844 2380
rect 18900 2324 19404 2380
rect 19460 2324 19470 2380
rect 20570 2324 20580 2380
rect 20636 2324 21644 2380
rect 21700 2324 21710 2380
rect 23482 2324 23492 2380
rect 23548 2324 24556 2380
rect 24612 2324 25956 2380
rect 26012 2324 26022 2380
rect 26186 2324 26196 2380
rect 26252 2324 26300 2380
rect 26356 2324 26404 2380
rect 26460 2324 26470 2380
rect 7690 2212 7700 2268
rect 7756 2212 8260 2268
rect 8316 2212 8596 2268
rect 8652 2212 8662 2268
rect 10154 2212 10164 2268
rect 10220 2212 10724 2268
rect 10780 2212 20804 2268
rect 20860 2212 23380 2268
rect 23436 2212 23446 2268
rect 23762 2212 23772 2268
rect 23828 2212 24892 2268
rect 24948 2212 25396 2268
rect 25452 2212 28084 2268
rect 28140 2212 28150 2268
rect 5450 2100 5460 2156
rect 5516 2100 5526 2156
rect 6906 2100 6916 2156
rect 6972 2100 7812 2156
rect 7868 2100 7878 2156
rect 13290 2100 13300 2156
rect 13356 2100 15316 2156
rect 15372 2100 15382 2156
rect 16874 2100 16884 2156
rect 16940 2100 17724 2156
rect 17780 2100 17790 2156
rect 18050 2100 18060 2156
rect 18172 2100 18182 2156
rect 18442 2100 18452 2156
rect 18564 2100 18574 2156
rect 19674 2100 19684 2156
rect 19740 2100 23268 2156
rect 23324 2100 24164 2156
rect 24220 2100 24230 2156
rect 28914 2100 28924 2156
rect 28980 2100 29764 2156
rect 29820 2100 34468 2156
rect 34524 2100 34534 2156
rect 3882 1876 3892 1932
rect 3948 1876 4732 1932
rect 4788 1876 5180 1932
rect 5236 1876 5246 1932
rect 5460 1820 5516 2100
rect 7634 1988 7644 2044
rect 7700 1988 8988 2044
rect 9044 1988 9054 2044
rect 17602 1988 17612 2044
rect 17668 1988 18340 2044
rect 18396 1988 18406 2044
rect 19684 1932 19740 2100
rect 21298 1988 21308 2044
rect 21364 1988 22372 2044
rect 22428 1988 22438 2044
rect 22596 1988 22708 2044
rect 22764 1988 22774 2044
rect 23986 1988 23996 2044
rect 24052 1988 24948 2044
rect 25004 1988 25014 2044
rect 26851 1988 27860 2044
rect 27916 1988 29148 2044
rect 29204 1988 29214 2044
rect 22596 1932 22652 1988
rect 26851 1932 26907 1988
rect 8586 1876 8596 1932
rect 8652 1876 12964 1932
rect 13020 1876 13030 1932
rect 13346 1876 13356 1932
rect 13412 1876 14364 1932
rect 14420 1876 19740 1932
rect 20178 1876 20188 1932
rect 20244 1876 21868 1932
rect 21924 1876 22652 1932
rect 22810 1876 22820 1932
rect 22876 1876 23268 1932
rect 23324 1876 23334 1932
rect 25946 1876 25956 1932
rect 26012 1876 26740 1932
rect 26796 1876 26907 1932
rect 27402 1876 27412 1932
rect 27468 1876 27748 1932
rect 27804 1876 28532 1932
rect 28588 1876 28598 1932
rect 4554 1764 4564 1820
rect 4620 1764 6244 1820
rect 6300 1764 6310 1820
rect 15530 1764 15540 1820
rect 15596 1764 20356 1820
rect 20412 1764 21084 1820
rect 21140 1764 21150 1820
rect 22530 1764 22540 1820
rect 22596 1764 25060 1820
rect 25116 1764 26572 1820
rect 26628 1764 26638 1820
rect 5170 1652 5180 1708
rect 5236 1652 5628 1708
rect 5684 1652 9324 1708
rect 9380 1652 9390 1708
rect 11218 1652 11228 1708
rect 11284 1652 13076 1708
rect 13132 1652 13142 1708
rect 15362 1652 15372 1708
rect 15428 1652 15876 1708
rect 15932 1652 15942 1708
rect 17714 1652 17724 1708
rect 17780 1652 18844 1708
rect 18900 1652 19180 1708
rect 19236 1652 19572 1708
rect 19628 1652 19638 1708
rect 19730 1652 19740 1708
rect 19796 1652 22260 1708
rect 22316 1652 22326 1708
rect 24938 1652 24948 1708
rect 25004 1652 28812 1708
rect 28868 1652 30884 1708
rect 30940 1652 30950 1708
rect 31891 1652 33460 1708
rect 33516 1652 33526 1708
rect 4806 1540 4816 1596
rect 4872 1540 4920 1596
rect 4976 1540 5024 1596
rect 5080 1540 5090 1596
rect 12898 1540 12908 1596
rect 12964 1540 13020 1652
rect 31891 1596 31947 1652
rect 13358 1540 13368 1596
rect 13424 1540 13472 1596
rect 13528 1540 13576 1596
rect 13632 1540 13642 1596
rect 19786 1540 19796 1596
rect 19852 1540 20300 1596
rect 20356 1540 20366 1596
rect 21910 1540 21920 1596
rect 21976 1540 22024 1596
rect 22080 1540 22128 1596
rect 22184 1540 22194 1596
rect 25722 1540 25732 1596
rect 25788 1540 26852 1596
rect 26908 1540 26918 1596
rect 30462 1540 30472 1596
rect 30528 1540 30576 1596
rect 30632 1540 30680 1596
rect 30736 1540 30746 1596
rect 30884 1540 31500 1596
rect 31556 1540 31947 1596
rect 30884 1484 30940 1540
rect 20178 1428 20188 1484
rect 20244 1428 20412 1484
rect 20468 1428 20478 1484
rect 21634 1428 21644 1484
rect 21700 1428 22988 1484
rect 23044 1428 23436 1484
rect 23492 1428 23940 1484
rect 23996 1428 24006 1484
rect 28914 1428 28924 1484
rect 28980 1428 29372 1484
rect 29428 1428 30940 1484
rect 19898 1316 19908 1372
rect 19964 1316 20076 1372
rect 20132 1316 20142 1372
rect 20682 1316 20692 1372
rect 20804 1316 20814 1372
rect 21410 1316 21420 1372
rect 21532 1316 21542 1372
rect 33506 1316 33516 1372
rect 33572 1316 34692 1372
rect 34748 1316 34758 1372
rect 17714 1204 17724 1260
rect 17780 1204 18004 1260
rect 18060 1204 18070 1260
rect 19618 1204 19628 1260
rect 19684 1204 20020 1260
rect 20076 1204 23660 1260
rect 23716 1204 24108 1260
rect 24164 1204 24174 1260
rect 24770 1204 24780 1260
rect 24836 1204 25228 1260
rect 25284 1204 25294 1260
rect 26842 1204 26852 1260
rect 26964 1204 26974 1260
rect 27066 1204 27076 1260
rect 27188 1204 27198 1260
rect 28130 1204 28140 1260
rect 28196 1204 30716 1260
rect 30772 1204 30782 1260
rect 32750 1204 32788 1260
rect 32844 1204 32854 1260
rect 19394 1092 19404 1148
rect 19460 1092 19908 1148
rect 19964 1092 19974 1148
rect 22082 1092 22092 1148
rect 22148 1092 23492 1148
rect 23548 1092 26348 1148
rect 26404 1092 26414 1148
rect 26851 1092 31892 1148
rect 31948 1092 32004 1148
rect 32060 1092 32070 1148
rect 32218 1092 32228 1148
rect 32284 1092 33124 1148
rect 33180 1092 33190 1148
rect 26851 1036 26907 1092
rect 17938 980 17948 1036
rect 18004 980 26907 1036
rect 29474 980 29484 1036
rect 29540 980 29876 1036
rect 29932 980 29942 1036
rect 30706 980 30716 1036
rect 30772 980 33684 1036
rect 33740 980 33852 1036
rect 33908 980 33918 1036
rect 35200 924 36000 952
rect 18162 868 18172 924
rect 18228 868 30100 924
rect 30156 868 36000 924
rect 35200 840 36000 868
rect 9082 756 9092 812
rect 9148 756 9196 812
rect 9252 756 9300 812
rect 9356 756 9366 812
rect 17634 756 17644 812
rect 17700 756 17748 812
rect 17804 756 17852 812
rect 17908 756 17918 812
rect 26186 756 26196 812
rect 26252 756 26300 812
rect 26356 756 26404 812
rect 26460 756 26470 812
rect 17490 644 17500 700
rect 17556 644 34468 700
rect 34524 644 34534 700
rect 18386 532 18396 588
rect 18452 532 29988 588
rect 30044 532 30054 588
<< via3 >>
rect 32004 13076 32060 13132
rect 4816 12516 4872 12572
rect 4920 12516 4976 12572
rect 5024 12516 5080 12572
rect 13368 12516 13424 12572
rect 13472 12516 13528 12572
rect 13576 12516 13632 12572
rect 21920 12516 21976 12572
rect 22024 12516 22080 12572
rect 22128 12516 22184 12572
rect 30472 12516 30528 12572
rect 30576 12516 30632 12572
rect 30680 12516 30736 12572
rect 21476 12404 21532 12460
rect 9940 12068 9996 12124
rect 8372 11732 8428 11788
rect 9092 11732 9148 11788
rect 9196 11732 9252 11788
rect 9300 11732 9356 11788
rect 17644 11732 17700 11788
rect 17748 11732 17804 11788
rect 17852 11732 17908 11788
rect 19796 11732 19852 11788
rect 26196 11732 26252 11788
rect 26300 11732 26356 11788
rect 26404 11732 26460 11788
rect 12068 11620 12124 11676
rect 12068 11396 12124 11452
rect 32788 11284 32844 11340
rect 4816 10948 4872 11004
rect 4920 10948 4976 11004
rect 5024 10948 5080 11004
rect 10948 10948 11004 11004
rect 13368 10948 13424 11004
rect 13472 10948 13528 11004
rect 13576 10948 13632 11004
rect 21920 10948 21976 11004
rect 22024 10948 22080 11004
rect 22128 10948 22184 11004
rect 30472 10948 30528 11004
rect 30576 10948 30632 11004
rect 30680 10948 30736 11004
rect 20020 10836 20076 10892
rect 3332 10388 3388 10444
rect 9092 10164 9148 10220
rect 9196 10164 9252 10220
rect 9300 10164 9356 10220
rect 9940 10164 9996 10220
rect 5908 10052 5964 10108
rect 7140 10052 7196 10108
rect 17644 10164 17700 10220
rect 17748 10164 17804 10220
rect 17852 10164 17908 10220
rect 26196 10164 26252 10220
rect 26300 10164 26356 10220
rect 26404 10164 26460 10220
rect 17444 9828 17500 9884
rect 18452 9828 18508 9884
rect 31892 9828 31948 9884
rect 7140 9716 7196 9772
rect 19460 9604 19516 9660
rect 33684 9604 33740 9660
rect 4816 9380 4872 9436
rect 4920 9380 4976 9436
rect 5024 9380 5080 9436
rect 13368 9380 13424 9436
rect 13472 9380 13528 9436
rect 13576 9380 13632 9436
rect 21700 9380 21756 9436
rect 21920 9380 21976 9436
rect 22024 9380 22080 9436
rect 22128 9380 22184 9436
rect 30472 9380 30528 9436
rect 30576 9380 30632 9436
rect 30680 9380 30736 9436
rect 26852 9268 26908 9324
rect 17444 9156 17500 9212
rect 18004 9156 18060 9212
rect 18452 9156 18508 9212
rect 21700 9156 21756 9212
rect 23716 9156 23772 9212
rect 6580 9044 6636 9100
rect 3332 8932 3388 8988
rect 5908 8932 5964 8988
rect 11732 8820 11788 8876
rect 19684 8820 19740 8876
rect 24388 8708 24444 8764
rect 9092 8596 9148 8652
rect 9196 8596 9252 8652
rect 9300 8596 9356 8652
rect 17644 8596 17700 8652
rect 17748 8596 17804 8652
rect 17852 8596 17908 8652
rect 18004 8596 18060 8652
rect 26196 8596 26252 8652
rect 26300 8596 26356 8652
rect 26404 8596 26460 8652
rect 8484 8484 8540 8540
rect 13188 8372 13244 8428
rect 29876 8372 29932 8428
rect 8372 8260 8428 8316
rect 10948 8260 11004 8316
rect 29316 8260 29372 8316
rect 7364 8148 7420 8204
rect 8036 8148 8092 8204
rect 33684 8148 33740 8204
rect 28980 8036 29036 8092
rect 4816 7812 4872 7868
rect 4920 7812 4976 7868
rect 5024 7812 5080 7868
rect 13368 7812 13424 7868
rect 13472 7812 13528 7868
rect 13576 7812 13632 7868
rect 21920 7812 21976 7868
rect 22024 7812 22080 7868
rect 22128 7812 22184 7868
rect 30472 7812 30528 7868
rect 30576 7812 30632 7868
rect 30680 7812 30736 7868
rect 33796 7812 33852 7868
rect 8484 7476 8540 7532
rect 13188 7476 13244 7532
rect 9940 7140 9996 7196
rect 13188 7140 13244 7196
rect 9092 7028 9148 7084
rect 9196 7028 9252 7084
rect 9300 7028 9356 7084
rect 17644 7028 17700 7084
rect 17748 7028 17804 7084
rect 17852 7028 17908 7084
rect 26196 7028 26252 7084
rect 26300 7028 26356 7084
rect 26404 7028 26460 7084
rect 13076 6804 13132 6860
rect 14084 6692 14140 6748
rect 23492 6692 23548 6748
rect 19460 6580 19516 6636
rect 24388 6580 24444 6636
rect 34356 6580 34412 6636
rect 11732 6468 11788 6524
rect 19684 6468 19740 6524
rect 4816 6244 4872 6300
rect 4920 6244 4976 6300
rect 5024 6244 5080 6300
rect 13368 6244 13424 6300
rect 13472 6244 13528 6300
rect 13576 6244 13632 6300
rect 21920 6244 21976 6300
rect 22024 6244 22080 6300
rect 22128 6244 22184 6300
rect 30472 6244 30528 6300
rect 30576 6244 30632 6300
rect 30680 6244 30736 6300
rect 7140 6132 7196 6188
rect 34356 6020 34412 6076
rect 9940 5684 9996 5740
rect 7140 5572 7196 5628
rect 9092 5460 9148 5516
rect 9196 5460 9252 5516
rect 9300 5460 9356 5516
rect 9604 5460 9660 5516
rect 17644 5460 17700 5516
rect 17748 5460 17804 5516
rect 17852 5460 17908 5516
rect 23716 5460 23772 5516
rect 26196 5460 26252 5516
rect 26300 5460 26356 5516
rect 26404 5460 26460 5516
rect 8708 5236 8764 5292
rect 29092 5124 29148 5180
rect 8484 5012 8540 5068
rect 12180 5012 12236 5068
rect 28980 4900 29036 4956
rect 29316 4900 29372 4956
rect 10388 4788 10444 4844
rect 14084 4788 14140 4844
rect 27076 4788 27132 4844
rect 4816 4676 4872 4732
rect 4920 4676 4976 4732
rect 5024 4676 5080 4732
rect 8596 4676 8652 4732
rect 11956 4676 12012 4732
rect 13368 4676 13424 4732
rect 13472 4676 13528 4732
rect 13576 4676 13632 4732
rect 21920 4676 21976 4732
rect 22024 4676 22080 4732
rect 22128 4676 22184 4732
rect 30472 4676 30528 4732
rect 30576 4676 30632 4732
rect 30680 4676 30736 4732
rect 19796 4564 19852 4620
rect 20692 4564 20748 4620
rect 7364 4452 7420 4508
rect 9604 4452 9660 4508
rect 9940 4452 9996 4508
rect 13076 4452 13132 4508
rect 14084 4452 14140 4508
rect 10276 4340 10332 4396
rect 12404 4340 12460 4396
rect 20356 4340 20412 4396
rect 29092 4228 29148 4284
rect 12740 4004 12796 4060
rect 13188 4116 13244 4172
rect 7140 3892 7196 3948
rect 9092 3892 9148 3948
rect 9196 3892 9252 3948
rect 9300 3892 9356 3948
rect 13188 3892 13244 3948
rect 17644 3892 17700 3948
rect 17748 3892 17804 3948
rect 17852 3892 17908 3948
rect 26196 3892 26252 3948
rect 26300 3892 26356 3948
rect 26404 3892 26460 3948
rect 8372 3780 8428 3836
rect 8596 3780 8652 3836
rect 29652 3780 29708 3836
rect 8036 3668 8092 3724
rect 11732 3668 11788 3724
rect 8036 3444 8092 3500
rect 8708 3444 8764 3500
rect 10276 3444 10332 3500
rect 9940 3332 9996 3388
rect 11732 3332 11788 3388
rect 11956 3332 12012 3388
rect 12180 3332 12236 3388
rect 13076 3332 13132 3388
rect 20356 3220 20412 3276
rect 29652 3220 29708 3276
rect 4816 3108 4872 3164
rect 4920 3108 4976 3164
rect 5024 3108 5080 3164
rect 12740 3108 12796 3164
rect 13368 3108 13424 3164
rect 13472 3108 13528 3164
rect 13576 3108 13632 3164
rect 21920 3108 21976 3164
rect 22024 3108 22080 3164
rect 22128 3108 22184 3164
rect 30472 3108 30528 3164
rect 30576 3108 30632 3164
rect 30680 3108 30736 3164
rect 8036 2884 8092 2940
rect 8484 2772 8540 2828
rect 8484 2436 8540 2492
rect 12404 2436 12460 2492
rect 9092 2324 9148 2380
rect 9196 2324 9252 2380
rect 9300 2324 9356 2380
rect 17644 2324 17700 2380
rect 17748 2324 17804 2380
rect 17852 2324 17908 2380
rect 26196 2324 26252 2380
rect 26300 2324 26356 2380
rect 26404 2324 26460 2380
rect 18116 2100 18172 2156
rect 18452 2100 18508 2156
rect 18340 1988 18396 2044
rect 12964 1876 13020 1932
rect 13076 1652 13132 1708
rect 4816 1540 4872 1596
rect 4920 1540 4976 1596
rect 5024 1540 5080 1596
rect 13368 1540 13424 1596
rect 13472 1540 13528 1596
rect 13576 1540 13632 1596
rect 19796 1540 19852 1596
rect 21920 1540 21976 1596
rect 22024 1540 22080 1596
rect 22128 1540 22184 1596
rect 30472 1540 30528 1596
rect 30576 1540 30632 1596
rect 30680 1540 30736 1596
rect 19908 1316 19964 1372
rect 20692 1316 20748 1372
rect 21476 1316 21532 1372
rect 18004 1204 18060 1260
rect 20020 1204 20076 1260
rect 26852 1204 26908 1260
rect 27076 1204 27132 1260
rect 32788 1204 32844 1260
rect 19908 1092 19964 1148
rect 23492 1092 23548 1148
rect 32004 1092 32060 1148
rect 29876 980 29932 1036
rect 9092 756 9148 812
rect 9196 756 9252 812
rect 9300 756 9356 812
rect 17644 756 17700 812
rect 17748 756 17804 812
rect 17852 756 17908 812
rect 26196 756 26252 812
rect 26300 756 26356 812
rect 26404 756 26460 812
<< metal4 >>
rect 32004 13132 32060 13142
rect 4788 12572 5108 12604
rect 4788 12516 4816 12572
rect 4872 12516 4920 12572
rect 4976 12516 5024 12572
rect 5080 12516 5108 12572
rect 4788 11794 5108 12516
rect 4788 11738 4816 11794
rect 4872 11738 4920 11794
rect 4976 11738 5024 11794
rect 5080 11738 5108 11794
rect 4788 11690 5108 11738
rect 4788 11634 4816 11690
rect 4872 11634 4920 11690
rect 4976 11634 5024 11690
rect 5080 11634 5108 11690
rect 4788 11586 5108 11634
rect 4788 11530 4816 11586
rect 4872 11530 4920 11586
rect 4976 11530 5024 11586
rect 5080 11530 5108 11586
rect 4788 11004 5108 11530
rect 4788 10948 4816 11004
rect 4872 10948 4920 11004
rect 4976 10948 5024 11004
rect 5080 10948 5108 11004
rect 3332 10444 3388 10454
rect 3332 8988 3388 10388
rect 3332 8922 3388 8932
rect 4788 9436 5108 10948
rect 8372 11788 8428 11798
rect 4788 9380 4816 9436
rect 4872 9380 4920 9436
rect 4976 9380 5024 9436
rect 5080 9380 5108 9436
rect 4788 8686 5108 9380
rect 5908 10108 5964 10118
rect 5908 8988 5964 10052
rect 7140 10108 7196 10118
rect 7140 9772 7196 10052
rect 6580 9748 6636 9758
rect 7140 9706 7196 9716
rect 6580 9100 6636 9692
rect 6580 9034 6636 9044
rect 5908 8922 5964 8932
rect 4788 8630 4816 8686
rect 4872 8630 4920 8686
rect 4976 8630 5024 8686
rect 5080 8630 5108 8686
rect 4788 8582 5108 8630
rect 4788 8526 4816 8582
rect 4872 8526 4920 8582
rect 4976 8526 5024 8582
rect 5080 8526 5108 8582
rect 4788 8478 5108 8526
rect 4788 8422 4816 8478
rect 4872 8422 4920 8478
rect 4976 8422 5024 8478
rect 5080 8422 5108 8478
rect 4788 7868 5108 8422
rect 8372 8316 8428 11732
rect 9064 11788 9384 12604
rect 13340 12572 13660 12604
rect 13340 12516 13368 12572
rect 13424 12516 13472 12572
rect 13528 12516 13576 12572
rect 13632 12516 13660 12572
rect 9064 11732 9092 11788
rect 9148 11732 9196 11788
rect 9252 11732 9300 11788
rect 9356 11732 9384 11788
rect 9064 10240 9384 11732
rect 9064 10164 9092 10240
rect 9148 10164 9196 10240
rect 9252 10164 9300 10240
rect 9356 10164 9384 10240
rect 9064 10136 9384 10164
rect 9064 10080 9092 10136
rect 9148 10080 9196 10136
rect 9252 10080 9300 10136
rect 9356 10080 9384 10136
rect 9064 10032 9384 10080
rect 9064 9976 9092 10032
rect 9148 9976 9196 10032
rect 9252 9976 9300 10032
rect 9356 9976 9384 10032
rect 9064 8652 9384 9976
rect 9064 8596 9092 8652
rect 9148 8596 9196 8652
rect 9252 8596 9300 8652
rect 9356 8596 9384 8652
rect 8372 8250 8428 8260
rect 8484 8540 8540 8550
rect 4788 7812 4816 7868
rect 4872 7812 4920 7868
rect 4976 7812 5024 7868
rect 5080 7812 5108 7868
rect 4788 6300 5108 7812
rect 4788 6244 4816 6300
rect 4872 6244 4920 6300
rect 4976 6244 5024 6300
rect 5080 6244 5108 6300
rect 4788 5578 5108 6244
rect 7364 8204 7420 8214
rect 4788 5522 4816 5578
rect 4872 5522 4920 5578
rect 4976 5522 5024 5578
rect 5080 5522 5108 5578
rect 4788 5474 5108 5522
rect 4788 5418 4816 5474
rect 4872 5418 4920 5474
rect 4976 5418 5024 5474
rect 5080 5418 5108 5474
rect 4788 5370 5108 5418
rect 4788 5314 4816 5370
rect 4872 5314 4920 5370
rect 4976 5314 5024 5370
rect 5080 5314 5108 5370
rect 4788 4732 5108 5314
rect 4788 4676 4816 4732
rect 4872 4676 4920 4732
rect 4976 4676 5024 4732
rect 5080 4676 5108 4732
rect 4788 3164 5108 4676
rect 7140 6188 7196 6198
rect 7140 5628 7196 6132
rect 7140 3948 7196 5572
rect 7364 4508 7420 8148
rect 7364 4442 7420 4452
rect 8036 8204 8092 8214
rect 7140 3882 7196 3892
rect 8036 3724 8092 8148
rect 8484 7532 8540 8484
rect 8484 7466 8540 7476
rect 9064 7132 9384 8596
rect 9064 6972 9092 7132
rect 9148 6972 9196 7132
rect 9252 6972 9300 7132
rect 9356 6972 9384 7132
rect 9940 12124 9996 12134
rect 9940 10220 9996 12068
rect 13340 11794 13660 12516
rect 13340 11738 13368 11794
rect 13424 11738 13472 11794
rect 13528 11738 13576 11794
rect 13632 11738 13660 11794
rect 13340 11690 13660 11738
rect 12068 11676 12124 11686
rect 12068 11452 12124 11620
rect 9940 7196 9996 10164
rect 10948 11004 11004 11014
rect 10948 8316 11004 10948
rect 12068 9748 12124 11396
rect 12068 9682 12124 9692
rect 13340 11634 13368 11690
rect 13424 11634 13472 11690
rect 13528 11634 13576 11690
rect 13632 11634 13660 11690
rect 13340 11586 13660 11634
rect 13340 11530 13368 11586
rect 13424 11530 13472 11586
rect 13528 11530 13576 11586
rect 13632 11530 13660 11586
rect 13340 11004 13660 11530
rect 13340 10948 13368 11004
rect 13424 10948 13472 11004
rect 13528 10948 13576 11004
rect 13632 10948 13660 11004
rect 13340 9436 13660 10948
rect 17616 11788 17936 12604
rect 21892 12572 22212 12604
rect 21892 12516 21920 12572
rect 21976 12516 22024 12572
rect 22080 12516 22128 12572
rect 22184 12516 22212 12572
rect 21476 12460 21532 12470
rect 17616 11732 17644 11788
rect 17700 11732 17748 11788
rect 17804 11732 17852 11788
rect 17908 11732 17936 11788
rect 17616 10240 17936 11732
rect 17616 10164 17644 10240
rect 17700 10164 17748 10240
rect 17804 10164 17852 10240
rect 17908 10164 17936 10240
rect 17616 10136 17936 10164
rect 17616 10080 17644 10136
rect 17700 10080 17748 10136
rect 17804 10080 17852 10136
rect 17908 10080 17936 10136
rect 17616 10032 17936 10080
rect 17616 9976 17644 10032
rect 17700 9976 17748 10032
rect 17804 9976 17852 10032
rect 17908 9976 17936 10032
rect 13340 9380 13368 9436
rect 13424 9380 13472 9436
rect 13528 9380 13576 9436
rect 13632 9380 13660 9436
rect 10948 8250 11004 8260
rect 11732 8876 11788 8886
rect 9940 7130 9996 7140
rect 9064 6924 9384 6972
rect 9064 6868 9092 6924
rect 9148 6868 9196 6924
rect 9252 6868 9300 6924
rect 9356 6868 9384 6924
rect 9064 5516 9384 6868
rect 11732 6524 11788 8820
rect 13340 8686 13660 9380
rect 17444 9884 17500 9894
rect 17444 9212 17500 9828
rect 17444 9146 17500 9156
rect 13340 8630 13368 8686
rect 13424 8630 13472 8686
rect 13528 8630 13576 8686
rect 13632 8630 13660 8686
rect 13340 8582 13660 8630
rect 13340 8526 13368 8582
rect 13424 8526 13472 8582
rect 13528 8526 13576 8582
rect 13632 8526 13660 8582
rect 13340 8478 13660 8526
rect 13188 8428 13244 8438
rect 13188 7532 13244 8372
rect 13188 7466 13244 7476
rect 13340 8422 13368 8478
rect 13424 8422 13472 8478
rect 13528 8422 13576 8478
rect 13632 8422 13660 8478
rect 13340 7868 13660 8422
rect 13340 7812 13368 7868
rect 13424 7812 13472 7868
rect 13528 7812 13576 7868
rect 13632 7812 13660 7868
rect 13188 7196 13244 7206
rect 11732 6458 11788 6468
rect 13076 6860 13132 6870
rect 9940 5740 9996 5750
rect 9064 5460 9092 5516
rect 9148 5460 9196 5516
rect 9252 5460 9300 5516
rect 9356 5460 9384 5516
rect 8708 5292 8764 5302
rect 8484 5068 8540 5078
rect 8036 3658 8092 3668
rect 8372 3836 8428 3846
rect 4788 3108 4816 3164
rect 4872 3108 4920 3164
rect 4976 3108 5024 3164
rect 5080 3108 5108 3164
rect 4788 2470 5108 3108
rect 8036 3500 8092 3510
rect 8036 2940 8092 3444
rect 8372 3448 8428 3780
rect 8372 3382 8428 3392
rect 8036 2874 8092 2884
rect 4788 2414 4816 2470
rect 4872 2414 4920 2470
rect 4976 2414 5024 2470
rect 5080 2414 5108 2470
rect 8484 2828 8540 5012
rect 8596 4732 8652 4742
rect 8596 3836 8652 4676
rect 8596 3770 8652 3780
rect 8708 3500 8764 5236
rect 8708 3434 8764 3444
rect 9064 4024 9384 5460
rect 9604 5516 9660 5526
rect 9604 4508 9660 5460
rect 9604 4442 9660 4452
rect 9940 4508 9996 5684
rect 12180 5068 12236 5078
rect 9940 4442 9996 4452
rect 10388 4844 10444 4854
rect 10276 4396 10332 4406
rect 9064 3968 9092 4024
rect 9148 3968 9196 4024
rect 9252 3968 9300 4024
rect 9356 3968 9384 4024
rect 9064 3948 9384 3968
rect 9064 3864 9092 3948
rect 9148 3864 9196 3948
rect 9252 3864 9300 3948
rect 9356 3864 9384 3948
rect 9064 3816 9384 3864
rect 9064 3760 9092 3816
rect 9148 3760 9196 3816
rect 9252 3760 9300 3816
rect 9356 3760 9384 3816
rect 8484 2492 8540 2772
rect 8484 2426 8540 2436
rect 4788 2366 5108 2414
rect 4788 2310 4816 2366
rect 4872 2310 4920 2366
rect 4976 2310 5024 2366
rect 5080 2310 5108 2366
rect 4788 2262 5108 2310
rect 4788 2206 4816 2262
rect 4872 2206 4920 2262
rect 4976 2206 5024 2262
rect 5080 2206 5108 2262
rect 4788 1596 5108 2206
rect 4788 1540 4816 1596
rect 4872 1540 4920 1596
rect 4976 1540 5024 1596
rect 5080 1540 5108 1596
rect 4788 724 5108 1540
rect 9064 2380 9384 3760
rect 9940 4340 10276 4348
rect 9940 4292 10332 4340
rect 9940 3388 9996 4292
rect 10388 3628 10444 4788
rect 11956 4732 12012 4742
rect 10276 3572 10444 3628
rect 11732 3724 11788 3734
rect 10276 3500 10332 3572
rect 10276 3434 10332 3444
rect 9940 3322 9996 3332
rect 11732 3388 11788 3668
rect 11732 3322 11788 3332
rect 11956 3448 12012 4676
rect 11956 3388 12012 3392
rect 11956 3322 12012 3332
rect 12180 3388 12236 5012
rect 13076 4508 13132 6804
rect 12180 3322 12236 3332
rect 12404 4396 12460 4406
rect 13076 4348 13132 4452
rect 12404 2492 12460 4340
rect 12964 4292 13132 4348
rect 12740 4060 12796 4070
rect 12740 3164 12796 4004
rect 12740 3098 12796 3108
rect 12404 2426 12460 2436
rect 9064 2324 9092 2380
rect 9148 2324 9196 2380
rect 9252 2324 9300 2380
rect 9356 2324 9384 2380
rect 9064 812 9384 2324
rect 12964 1932 13020 4292
rect 13188 4172 13244 7140
rect 13188 4106 13244 4116
rect 13340 6300 13660 7812
rect 17616 8652 17936 9976
rect 19796 11788 19852 11798
rect 18452 9884 18508 9894
rect 17616 8596 17644 8652
rect 17700 8596 17748 8652
rect 17804 8596 17852 8652
rect 17908 8596 17936 8652
rect 17616 7132 17936 8596
rect 18004 9212 18060 9222
rect 18004 8652 18060 9156
rect 18004 8586 18060 8596
rect 18452 9212 18508 9828
rect 17616 6972 17644 7132
rect 17700 6972 17748 7132
rect 17804 6972 17852 7132
rect 17908 6972 17936 7132
rect 17616 6924 17936 6972
rect 17616 6868 17644 6924
rect 17700 6868 17748 6924
rect 17804 6868 17852 6924
rect 17908 6868 17936 6924
rect 13340 6244 13368 6300
rect 13424 6244 13472 6300
rect 13528 6244 13576 6300
rect 13632 6244 13660 6300
rect 13340 5578 13660 6244
rect 13340 5522 13368 5578
rect 13424 5522 13472 5578
rect 13528 5522 13576 5578
rect 13632 5522 13660 5578
rect 13340 5474 13660 5522
rect 13340 5418 13368 5474
rect 13424 5418 13472 5474
rect 13528 5418 13576 5474
rect 13632 5418 13660 5474
rect 13340 5370 13660 5418
rect 13340 5314 13368 5370
rect 13424 5314 13472 5370
rect 13528 5314 13576 5370
rect 13632 5314 13660 5370
rect 13340 4732 13660 5314
rect 13340 4676 13368 4732
rect 13424 4676 13472 4732
rect 13528 4676 13576 4732
rect 13632 4676 13660 4732
rect 13188 3948 13244 3958
rect 13188 3808 13244 3892
rect 12964 1866 13020 1876
rect 13076 3752 13244 3808
rect 13076 3388 13132 3752
rect 13076 1708 13132 3332
rect 13076 1642 13132 1652
rect 13340 3164 13660 4676
rect 14084 6748 14140 6758
rect 14084 4844 14140 6692
rect 14084 4508 14140 4788
rect 14084 4442 14140 4452
rect 17616 5516 17936 6868
rect 17616 5460 17644 5516
rect 17700 5460 17748 5516
rect 17804 5460 17852 5516
rect 17908 5460 17936 5516
rect 13340 3108 13368 3164
rect 13424 3108 13472 3164
rect 13528 3108 13576 3164
rect 13632 3108 13660 3164
rect 13340 2470 13660 3108
rect 13340 2414 13368 2470
rect 13424 2414 13472 2470
rect 13528 2414 13576 2470
rect 13632 2414 13660 2470
rect 13340 2366 13660 2414
rect 13340 2310 13368 2366
rect 13424 2310 13472 2366
rect 13528 2310 13576 2366
rect 13632 2310 13660 2366
rect 13340 2262 13660 2310
rect 13340 2206 13368 2262
rect 13424 2206 13472 2262
rect 13528 2206 13576 2262
rect 13632 2206 13660 2262
rect 9064 756 9092 812
rect 9148 756 9196 812
rect 9252 756 9300 812
rect 9356 756 9384 812
rect 9064 724 9384 756
rect 13340 1596 13660 2206
rect 13340 1540 13368 1596
rect 13424 1540 13472 1596
rect 13528 1540 13576 1596
rect 13632 1540 13660 1596
rect 13340 724 13660 1540
rect 17616 4024 17936 5460
rect 17616 3968 17644 4024
rect 17700 3968 17748 4024
rect 17804 3968 17852 4024
rect 17908 3968 17936 4024
rect 17616 3948 17936 3968
rect 17616 3864 17644 3948
rect 17700 3864 17748 3948
rect 17804 3864 17852 3948
rect 17908 3864 17936 3948
rect 17616 3816 17936 3864
rect 17616 3760 17644 3816
rect 17700 3760 17748 3816
rect 17804 3760 17852 3816
rect 17908 3760 17936 3816
rect 17616 2380 17936 3760
rect 17616 2324 17644 2380
rect 17700 2324 17748 2380
rect 17804 2324 17852 2380
rect 17908 2324 17936 2380
rect 17616 812 17936 2324
rect 18116 6688 18172 6698
rect 18116 2156 18172 6632
rect 18116 2090 18172 2100
rect 18452 2156 18508 9156
rect 19460 9660 19516 9670
rect 19460 6636 19516 9604
rect 19460 6570 19516 6580
rect 19684 8876 19740 8886
rect 19684 6524 19740 8820
rect 19684 6458 19740 6468
rect 18452 2090 18508 2100
rect 19796 4620 19852 11732
rect 18340 2044 18396 2054
rect 18340 1942 18396 1952
rect 19796 1596 19852 4564
rect 19796 1530 19852 1540
rect 20020 10892 20076 10902
rect 19908 1468 19964 1478
rect 19908 1372 19964 1412
rect 19908 1306 19964 1316
rect 18004 1288 18060 1298
rect 18004 1194 18060 1204
rect 20020 1260 20076 10836
rect 20692 4620 20748 4630
rect 20356 4396 20412 4406
rect 20356 3276 20412 4340
rect 20356 3210 20412 3220
rect 20692 1372 20748 4564
rect 20692 1306 20748 1316
rect 21476 1372 21532 12404
rect 21892 11794 22212 12516
rect 21892 11738 21920 11794
rect 21976 11738 22024 11794
rect 22080 11738 22128 11794
rect 22184 11738 22212 11794
rect 21892 11690 22212 11738
rect 21892 11634 21920 11690
rect 21976 11634 22024 11690
rect 22080 11634 22128 11690
rect 22184 11634 22212 11690
rect 21892 11586 22212 11634
rect 21892 11530 21920 11586
rect 21976 11530 22024 11586
rect 22080 11530 22128 11586
rect 22184 11530 22212 11586
rect 21892 11004 22212 11530
rect 21892 10948 21920 11004
rect 21976 10948 22024 11004
rect 22080 10948 22128 11004
rect 22184 10948 22212 11004
rect 21700 9436 21756 9446
rect 21700 9212 21756 9380
rect 21700 9146 21756 9156
rect 21892 9436 22212 10948
rect 21892 9380 21920 9436
rect 21976 9380 22024 9436
rect 22080 9380 22128 9436
rect 22184 9380 22212 9436
rect 21476 1306 21532 1316
rect 21892 8686 22212 9380
rect 26168 11788 26488 12604
rect 26168 11732 26196 11788
rect 26252 11732 26300 11788
rect 26356 11732 26404 11788
rect 26460 11732 26488 11788
rect 26168 10240 26488 11732
rect 26168 10164 26196 10240
rect 26252 10164 26300 10240
rect 26356 10164 26404 10240
rect 26460 10164 26488 10240
rect 26168 10136 26488 10164
rect 26168 10080 26196 10136
rect 26252 10080 26300 10136
rect 26356 10080 26404 10136
rect 26460 10080 26488 10136
rect 26168 10032 26488 10080
rect 26168 9976 26196 10032
rect 26252 9976 26300 10032
rect 26356 9976 26404 10032
rect 26460 9976 26488 10032
rect 21892 8630 21920 8686
rect 21976 8630 22024 8686
rect 22080 8630 22128 8686
rect 22184 8630 22212 8686
rect 21892 8582 22212 8630
rect 21892 8526 21920 8582
rect 21976 8526 22024 8582
rect 22080 8526 22128 8582
rect 22184 8526 22212 8582
rect 21892 8478 22212 8526
rect 21892 8422 21920 8478
rect 21976 8422 22024 8478
rect 22080 8422 22128 8478
rect 22184 8422 22212 8478
rect 21892 7868 22212 8422
rect 21892 7812 21920 7868
rect 21976 7812 22024 7868
rect 22080 7812 22128 7868
rect 22184 7812 22212 7868
rect 21892 6300 22212 7812
rect 23716 9212 23772 9222
rect 21892 6244 21920 6300
rect 21976 6244 22024 6300
rect 22080 6244 22128 6300
rect 22184 6244 22212 6300
rect 21892 5578 22212 6244
rect 21892 5522 21920 5578
rect 21976 5522 22024 5578
rect 22080 5522 22128 5578
rect 22184 5522 22212 5578
rect 21892 5474 22212 5522
rect 21892 5418 21920 5474
rect 21976 5418 22024 5474
rect 22080 5418 22128 5474
rect 22184 5418 22212 5474
rect 21892 5370 22212 5418
rect 21892 5314 21920 5370
rect 21976 5314 22024 5370
rect 22080 5314 22128 5370
rect 22184 5314 22212 5370
rect 21892 4732 22212 5314
rect 21892 4676 21920 4732
rect 21976 4676 22024 4732
rect 22080 4676 22128 4732
rect 22184 4676 22212 4732
rect 21892 3164 22212 4676
rect 21892 3108 21920 3164
rect 21976 3108 22024 3164
rect 22080 3108 22128 3164
rect 22184 3108 22212 3164
rect 21892 2470 22212 3108
rect 21892 2414 21920 2470
rect 21976 2414 22024 2470
rect 22080 2414 22128 2470
rect 22184 2414 22212 2470
rect 21892 2366 22212 2414
rect 21892 2310 21920 2366
rect 21976 2310 22024 2366
rect 22080 2310 22128 2366
rect 22184 2310 22212 2366
rect 21892 2262 22212 2310
rect 21892 2206 21920 2262
rect 21976 2206 22024 2262
rect 22080 2206 22128 2262
rect 22184 2206 22212 2262
rect 21892 1596 22212 2206
rect 21892 1540 21920 1596
rect 21976 1540 22024 1596
rect 22080 1540 22128 1596
rect 22184 1540 22212 1596
rect 20020 1194 20076 1204
rect 19908 1148 19964 1158
rect 19908 1042 19964 1052
rect 17616 756 17644 812
rect 17700 756 17748 812
rect 17804 756 17852 812
rect 17908 756 17936 812
rect 17616 724 17936 756
rect 21892 724 22212 1540
rect 23492 6748 23548 6758
rect 23492 1148 23548 6692
rect 23716 5516 23772 9156
rect 24388 8764 24444 8774
rect 24388 6636 24444 8708
rect 24388 6570 24444 6580
rect 26168 8652 26488 9976
rect 30444 12572 30764 12604
rect 30444 12516 30472 12572
rect 30528 12516 30576 12572
rect 30632 12516 30680 12572
rect 30736 12516 30764 12572
rect 30444 11794 30764 12516
rect 30444 11738 30472 11794
rect 30528 11738 30576 11794
rect 30632 11738 30680 11794
rect 30736 11738 30764 11794
rect 30444 11690 30764 11738
rect 30444 11634 30472 11690
rect 30528 11634 30576 11690
rect 30632 11634 30680 11690
rect 30736 11634 30764 11690
rect 30444 11586 30764 11634
rect 30444 11530 30472 11586
rect 30528 11530 30576 11586
rect 30632 11530 30680 11586
rect 30736 11530 30764 11586
rect 30444 11004 30764 11530
rect 30444 10948 30472 11004
rect 30528 10948 30576 11004
rect 30632 10948 30680 11004
rect 30736 10948 30764 11004
rect 30444 9436 30764 10948
rect 30444 9380 30472 9436
rect 30528 9380 30576 9436
rect 30632 9380 30680 9436
rect 30736 9380 30764 9436
rect 26168 8596 26196 8652
rect 26252 8596 26300 8652
rect 26356 8596 26404 8652
rect 26460 8596 26488 8652
rect 26168 7132 26488 8596
rect 26168 6972 26196 7132
rect 26252 6972 26300 7132
rect 26356 6972 26404 7132
rect 26460 6972 26488 7132
rect 26168 6924 26488 6972
rect 26168 6868 26196 6924
rect 26252 6868 26300 6924
rect 26356 6868 26404 6924
rect 26460 6868 26488 6924
rect 23716 5450 23772 5460
rect 26168 5516 26488 6868
rect 26168 5460 26196 5516
rect 26252 5460 26300 5516
rect 26356 5460 26404 5516
rect 26460 5460 26488 5516
rect 23492 1082 23548 1092
rect 26168 4024 26488 5460
rect 26168 3968 26196 4024
rect 26252 3968 26300 4024
rect 26356 3968 26404 4024
rect 26460 3968 26488 4024
rect 26168 3948 26488 3968
rect 26168 3864 26196 3948
rect 26252 3864 26300 3948
rect 26356 3864 26404 3948
rect 26460 3864 26488 3948
rect 26168 3816 26488 3864
rect 26168 3760 26196 3816
rect 26252 3760 26300 3816
rect 26356 3760 26404 3816
rect 26460 3760 26488 3816
rect 26168 2380 26488 3760
rect 26168 2324 26196 2380
rect 26252 2324 26300 2380
rect 26356 2324 26404 2380
rect 26460 2324 26488 2380
rect 26168 812 26488 2324
rect 26852 9324 26908 9334
rect 26852 1260 26908 9268
rect 30444 8686 30764 9380
rect 30444 8630 30472 8686
rect 30528 8630 30576 8686
rect 30632 8630 30680 8686
rect 30736 8630 30764 8686
rect 30444 8582 30764 8630
rect 30444 8526 30472 8582
rect 30528 8526 30576 8582
rect 30632 8526 30680 8582
rect 30736 8526 30764 8582
rect 30444 8478 30764 8526
rect 29876 8428 29932 8438
rect 29316 8316 29372 8326
rect 28980 8092 29036 8102
rect 28980 4956 29036 8036
rect 28980 4890 29036 4900
rect 29092 5180 29148 5190
rect 26852 1194 26908 1204
rect 27076 4844 27132 4854
rect 27076 1260 27132 4788
rect 29092 4284 29148 5124
rect 29316 4956 29372 8260
rect 29316 4890 29372 4900
rect 29092 4218 29148 4228
rect 29652 3836 29708 3846
rect 29652 3276 29708 3780
rect 29652 3210 29708 3220
rect 27076 1194 27132 1204
rect 29876 1036 29932 8372
rect 29876 970 29932 980
rect 30444 8422 30472 8478
rect 30528 8422 30576 8478
rect 30632 8422 30680 8478
rect 30736 8422 30764 8478
rect 30444 7868 30764 8422
rect 30444 7812 30472 7868
rect 30528 7812 30576 7868
rect 30632 7812 30680 7868
rect 30736 7812 30764 7868
rect 30444 6300 30764 7812
rect 30444 6244 30472 6300
rect 30528 6244 30576 6300
rect 30632 6244 30680 6300
rect 30736 6244 30764 6300
rect 30444 5578 30764 6244
rect 30444 5522 30472 5578
rect 30528 5522 30576 5578
rect 30632 5522 30680 5578
rect 30736 5522 30764 5578
rect 30444 5474 30764 5522
rect 30444 5418 30472 5474
rect 30528 5418 30576 5474
rect 30632 5418 30680 5474
rect 30736 5418 30764 5474
rect 30444 5370 30764 5418
rect 30444 5314 30472 5370
rect 30528 5314 30576 5370
rect 30632 5314 30680 5370
rect 30736 5314 30764 5370
rect 30444 4732 30764 5314
rect 30444 4676 30472 4732
rect 30528 4676 30576 4732
rect 30632 4676 30680 4732
rect 30736 4676 30764 4732
rect 30444 3164 30764 4676
rect 30444 3108 30472 3164
rect 30528 3108 30576 3164
rect 30632 3108 30680 3164
rect 30736 3108 30764 3164
rect 30444 2470 30764 3108
rect 30444 2414 30472 2470
rect 30528 2414 30576 2470
rect 30632 2414 30680 2470
rect 30736 2414 30764 2470
rect 30444 2366 30764 2414
rect 30444 2310 30472 2366
rect 30528 2310 30576 2366
rect 30632 2310 30680 2366
rect 30736 2310 30764 2366
rect 30444 2262 30764 2310
rect 30444 2206 30472 2262
rect 30528 2206 30576 2262
rect 30632 2206 30680 2262
rect 30736 2206 30764 2262
rect 30444 1596 30764 2206
rect 31892 9884 31948 9894
rect 31892 2008 31948 9828
rect 31892 1942 31948 1952
rect 30444 1540 30472 1596
rect 30528 1540 30576 1596
rect 30632 1540 30680 1596
rect 30736 1540 30764 1596
rect 26168 756 26196 812
rect 26252 756 26300 812
rect 26356 756 26404 812
rect 26460 756 26488 812
rect 26168 724 26488 756
rect 30444 724 30764 1540
rect 32004 1148 32060 13076
rect 32788 11340 32844 11350
rect 32788 1288 32844 11284
rect 33684 9660 33740 9670
rect 33684 8204 33740 9604
rect 33684 1468 33740 8148
rect 33684 1402 33740 1412
rect 33796 7868 33852 7878
rect 32788 1156 32844 1204
rect 32004 1082 32060 1092
rect 33796 1108 33852 7812
rect 34356 6688 34412 6698
rect 34356 6076 34412 6580
rect 34356 6010 34412 6020
rect 33796 1042 33852 1052
<< via4 >>
rect 4816 11738 4872 11794
rect 4920 11738 4976 11794
rect 5024 11738 5080 11794
rect 4816 11634 4872 11690
rect 4920 11634 4976 11690
rect 5024 11634 5080 11690
rect 4816 11530 4872 11586
rect 4920 11530 4976 11586
rect 5024 11530 5080 11586
rect 6580 9692 6636 9748
rect 4816 8630 4872 8686
rect 4920 8630 4976 8686
rect 5024 8630 5080 8686
rect 4816 8526 4872 8582
rect 4920 8526 4976 8582
rect 5024 8526 5080 8582
rect 4816 8422 4872 8478
rect 4920 8422 4976 8478
rect 5024 8422 5080 8478
rect 9092 10220 9148 10240
rect 9092 10184 9148 10220
rect 9196 10220 9252 10240
rect 9196 10184 9252 10220
rect 9300 10220 9356 10240
rect 9300 10184 9356 10220
rect 9092 10080 9148 10136
rect 9196 10080 9252 10136
rect 9300 10080 9356 10136
rect 9092 9976 9148 10032
rect 9196 9976 9252 10032
rect 9300 9976 9356 10032
rect 4816 5522 4872 5578
rect 4920 5522 4976 5578
rect 5024 5522 5080 5578
rect 4816 5418 4872 5474
rect 4920 5418 4976 5474
rect 5024 5418 5080 5474
rect 4816 5314 4872 5370
rect 4920 5314 4976 5370
rect 5024 5314 5080 5370
rect 9092 7084 9148 7132
rect 9092 7076 9148 7084
rect 9092 6972 9148 7028
rect 9196 7084 9252 7132
rect 9196 7076 9252 7084
rect 9196 6972 9252 7028
rect 9300 7084 9356 7132
rect 9300 7076 9356 7084
rect 9300 6972 9356 7028
rect 13368 11738 13424 11794
rect 13472 11738 13528 11794
rect 13576 11738 13632 11794
rect 12068 9692 12124 9748
rect 13368 11634 13424 11690
rect 13472 11634 13528 11690
rect 13576 11634 13632 11690
rect 13368 11530 13424 11586
rect 13472 11530 13528 11586
rect 13576 11530 13632 11586
rect 17644 10220 17700 10240
rect 17644 10184 17700 10220
rect 17748 10220 17804 10240
rect 17748 10184 17804 10220
rect 17852 10220 17908 10240
rect 17852 10184 17908 10220
rect 17644 10080 17700 10136
rect 17748 10080 17804 10136
rect 17852 10080 17908 10136
rect 17644 9976 17700 10032
rect 17748 9976 17804 10032
rect 17852 9976 17908 10032
rect 9092 6868 9148 6924
rect 9196 6868 9252 6924
rect 9300 6868 9356 6924
rect 13368 8630 13424 8686
rect 13472 8630 13528 8686
rect 13576 8630 13632 8686
rect 13368 8526 13424 8582
rect 13472 8526 13528 8582
rect 13576 8526 13632 8582
rect 13368 8422 13424 8478
rect 13472 8422 13528 8478
rect 13576 8422 13632 8478
rect 8372 3392 8428 3448
rect 4816 2414 4872 2470
rect 4920 2414 4976 2470
rect 5024 2414 5080 2470
rect 9092 3968 9148 4024
rect 9196 3968 9252 4024
rect 9300 3968 9356 4024
rect 9092 3892 9148 3920
rect 9092 3864 9148 3892
rect 9196 3892 9252 3920
rect 9196 3864 9252 3892
rect 9300 3892 9356 3920
rect 9300 3864 9356 3892
rect 9092 3760 9148 3816
rect 9196 3760 9252 3816
rect 9300 3760 9356 3816
rect 4816 2310 4872 2366
rect 4920 2310 4976 2366
rect 5024 2310 5080 2366
rect 4816 2206 4872 2262
rect 4920 2206 4976 2262
rect 5024 2206 5080 2262
rect 11956 3392 12012 3448
rect 17644 7084 17700 7132
rect 17644 7076 17700 7084
rect 17644 6972 17700 7028
rect 17748 7084 17804 7132
rect 17748 7076 17804 7084
rect 17748 6972 17804 7028
rect 17852 7084 17908 7132
rect 17852 7076 17908 7084
rect 17852 6972 17908 7028
rect 17644 6868 17700 6924
rect 17748 6868 17804 6924
rect 17852 6868 17908 6924
rect 13368 5522 13424 5578
rect 13472 5522 13528 5578
rect 13576 5522 13632 5578
rect 13368 5418 13424 5474
rect 13472 5418 13528 5474
rect 13576 5418 13632 5474
rect 13368 5314 13424 5370
rect 13472 5314 13528 5370
rect 13576 5314 13632 5370
rect 13368 2414 13424 2470
rect 13472 2414 13528 2470
rect 13576 2414 13632 2470
rect 13368 2310 13424 2366
rect 13472 2310 13528 2366
rect 13576 2310 13632 2366
rect 13368 2206 13424 2262
rect 13472 2206 13528 2262
rect 13576 2206 13632 2262
rect 17644 3968 17700 4024
rect 17748 3968 17804 4024
rect 17852 3968 17908 4024
rect 17644 3892 17700 3920
rect 17644 3864 17700 3892
rect 17748 3892 17804 3920
rect 17748 3864 17804 3892
rect 17852 3892 17908 3920
rect 17852 3864 17908 3892
rect 17644 3760 17700 3816
rect 17748 3760 17804 3816
rect 17852 3760 17908 3816
rect 18116 6632 18172 6688
rect 18340 1988 18396 2008
rect 18340 1952 18396 1988
rect 19908 1412 19964 1468
rect 18004 1260 18060 1288
rect 18004 1232 18060 1260
rect 21920 11738 21976 11794
rect 22024 11738 22080 11794
rect 22128 11738 22184 11794
rect 21920 11634 21976 11690
rect 22024 11634 22080 11690
rect 22128 11634 22184 11690
rect 21920 11530 21976 11586
rect 22024 11530 22080 11586
rect 22128 11530 22184 11586
rect 26196 10220 26252 10240
rect 26196 10184 26252 10220
rect 26300 10220 26356 10240
rect 26300 10184 26356 10220
rect 26404 10220 26460 10240
rect 26404 10184 26460 10220
rect 26196 10080 26252 10136
rect 26300 10080 26356 10136
rect 26404 10080 26460 10136
rect 26196 9976 26252 10032
rect 26300 9976 26356 10032
rect 26404 9976 26460 10032
rect 21920 8630 21976 8686
rect 22024 8630 22080 8686
rect 22128 8630 22184 8686
rect 21920 8526 21976 8582
rect 22024 8526 22080 8582
rect 22128 8526 22184 8582
rect 21920 8422 21976 8478
rect 22024 8422 22080 8478
rect 22128 8422 22184 8478
rect 21920 5522 21976 5578
rect 22024 5522 22080 5578
rect 22128 5522 22184 5578
rect 21920 5418 21976 5474
rect 22024 5418 22080 5474
rect 22128 5418 22184 5474
rect 21920 5314 21976 5370
rect 22024 5314 22080 5370
rect 22128 5314 22184 5370
rect 21920 2414 21976 2470
rect 22024 2414 22080 2470
rect 22128 2414 22184 2470
rect 21920 2310 21976 2366
rect 22024 2310 22080 2366
rect 22128 2310 22184 2366
rect 21920 2206 21976 2262
rect 22024 2206 22080 2262
rect 22128 2206 22184 2262
rect 19908 1092 19964 1108
rect 19908 1052 19964 1092
rect 30472 11738 30528 11794
rect 30576 11738 30632 11794
rect 30680 11738 30736 11794
rect 30472 11634 30528 11690
rect 30576 11634 30632 11690
rect 30680 11634 30736 11690
rect 30472 11530 30528 11586
rect 30576 11530 30632 11586
rect 30680 11530 30736 11586
rect 26196 7084 26252 7132
rect 26196 7076 26252 7084
rect 26196 6972 26252 7028
rect 26300 7084 26356 7132
rect 26300 7076 26356 7084
rect 26300 6972 26356 7028
rect 26404 7084 26460 7132
rect 26404 7076 26460 7084
rect 26404 6972 26460 7028
rect 26196 6868 26252 6924
rect 26300 6868 26356 6924
rect 26404 6868 26460 6924
rect 26196 3968 26252 4024
rect 26300 3968 26356 4024
rect 26404 3968 26460 4024
rect 26196 3892 26252 3920
rect 26196 3864 26252 3892
rect 26300 3892 26356 3920
rect 26300 3864 26356 3892
rect 26404 3892 26460 3920
rect 26404 3864 26460 3892
rect 26196 3760 26252 3816
rect 26300 3760 26356 3816
rect 26404 3760 26460 3816
rect 30472 8630 30528 8686
rect 30576 8630 30632 8686
rect 30680 8630 30736 8686
rect 30472 8526 30528 8582
rect 30576 8526 30632 8582
rect 30680 8526 30736 8582
rect 30472 8422 30528 8478
rect 30576 8422 30632 8478
rect 30680 8422 30736 8478
rect 30472 5522 30528 5578
rect 30576 5522 30632 5578
rect 30680 5522 30736 5578
rect 30472 5418 30528 5474
rect 30576 5418 30632 5474
rect 30680 5418 30736 5474
rect 30472 5314 30528 5370
rect 30576 5314 30632 5370
rect 30680 5314 30736 5370
rect 30472 2414 30528 2470
rect 30576 2414 30632 2470
rect 30680 2414 30736 2470
rect 30472 2310 30528 2366
rect 30576 2310 30632 2366
rect 30680 2310 30736 2366
rect 30472 2206 30528 2262
rect 30576 2206 30632 2262
rect 30680 2206 30736 2262
rect 31892 1952 31948 2008
rect 33684 1412 33740 1468
rect 32788 1260 32844 1288
rect 32788 1232 32844 1260
rect 34356 6636 34412 6688
rect 34356 6632 34412 6636
rect 33796 1052 33852 1108
<< metal5 >>
rect 612 11794 34892 11822
rect 612 11738 4816 11794
rect 4872 11738 4920 11794
rect 4976 11738 5024 11794
rect 5080 11738 13368 11794
rect 13424 11738 13472 11794
rect 13528 11738 13576 11794
rect 13632 11738 21920 11794
rect 21976 11738 22024 11794
rect 22080 11738 22128 11794
rect 22184 11738 30472 11794
rect 30528 11738 30576 11794
rect 30632 11738 30680 11794
rect 30736 11738 34892 11794
rect 612 11690 34892 11738
rect 612 11634 4816 11690
rect 4872 11634 4920 11690
rect 4976 11634 5024 11690
rect 5080 11634 13368 11690
rect 13424 11634 13472 11690
rect 13528 11634 13576 11690
rect 13632 11634 21920 11690
rect 21976 11634 22024 11690
rect 22080 11634 22128 11690
rect 22184 11634 30472 11690
rect 30528 11634 30576 11690
rect 30632 11634 30680 11690
rect 30736 11634 34892 11690
rect 612 11586 34892 11634
rect 612 11530 4816 11586
rect 4872 11530 4920 11586
rect 4976 11530 5024 11586
rect 5080 11530 13368 11586
rect 13424 11530 13472 11586
rect 13528 11530 13576 11586
rect 13632 11530 21920 11586
rect 21976 11530 22024 11586
rect 22080 11530 22128 11586
rect 22184 11530 30472 11586
rect 30528 11530 30576 11586
rect 30632 11530 30680 11586
rect 30736 11530 34892 11586
rect 612 11502 34892 11530
rect 612 10240 34892 10268
rect 612 10184 9092 10240
rect 9148 10184 9196 10240
rect 9252 10184 9300 10240
rect 9356 10184 17644 10240
rect 17700 10184 17748 10240
rect 17804 10184 17852 10240
rect 17908 10184 26196 10240
rect 26252 10184 26300 10240
rect 26356 10184 26404 10240
rect 26460 10184 34892 10240
rect 612 10136 34892 10184
rect 612 10080 9092 10136
rect 9148 10080 9196 10136
rect 9252 10080 9300 10136
rect 9356 10080 17644 10136
rect 17700 10080 17748 10136
rect 17804 10080 17852 10136
rect 17908 10080 26196 10136
rect 26252 10080 26300 10136
rect 26356 10080 26404 10136
rect 26460 10080 34892 10136
rect 612 10032 34892 10080
rect 612 9976 9092 10032
rect 9148 9976 9196 10032
rect 9252 9976 9300 10032
rect 9356 9976 17644 10032
rect 17700 9976 17748 10032
rect 17804 9976 17852 10032
rect 17908 9976 26196 10032
rect 26252 9976 26300 10032
rect 26356 9976 26404 10032
rect 26460 9976 34892 10032
rect 612 9948 34892 9976
rect 6564 9748 12140 9764
rect 6564 9692 6580 9748
rect 6636 9692 12068 9748
rect 12124 9692 12140 9748
rect 6564 9676 12140 9692
rect 612 8686 34892 8714
rect 612 8630 4816 8686
rect 4872 8630 4920 8686
rect 4976 8630 5024 8686
rect 5080 8630 13368 8686
rect 13424 8630 13472 8686
rect 13528 8630 13576 8686
rect 13632 8630 21920 8686
rect 21976 8630 22024 8686
rect 22080 8630 22128 8686
rect 22184 8630 30472 8686
rect 30528 8630 30576 8686
rect 30632 8630 30680 8686
rect 30736 8630 34892 8686
rect 612 8582 34892 8630
rect 612 8526 4816 8582
rect 4872 8526 4920 8582
rect 4976 8526 5024 8582
rect 5080 8526 13368 8582
rect 13424 8526 13472 8582
rect 13528 8526 13576 8582
rect 13632 8526 21920 8582
rect 21976 8526 22024 8582
rect 22080 8526 22128 8582
rect 22184 8526 30472 8582
rect 30528 8526 30576 8582
rect 30632 8526 30680 8582
rect 30736 8526 34892 8582
rect 612 8478 34892 8526
rect 612 8422 4816 8478
rect 4872 8422 4920 8478
rect 4976 8422 5024 8478
rect 5080 8422 13368 8478
rect 13424 8422 13472 8478
rect 13528 8422 13576 8478
rect 13632 8422 21920 8478
rect 21976 8422 22024 8478
rect 22080 8422 22128 8478
rect 22184 8422 30472 8478
rect 30528 8422 30576 8478
rect 30632 8422 30680 8478
rect 30736 8422 34892 8478
rect 612 8394 34892 8422
rect 612 7132 34892 7160
rect 612 7076 9092 7132
rect 9148 7076 9196 7132
rect 9252 7076 9300 7132
rect 9356 7076 17644 7132
rect 17700 7076 17748 7132
rect 17804 7076 17852 7132
rect 17908 7076 26196 7132
rect 26252 7076 26300 7132
rect 26356 7076 26404 7132
rect 26460 7076 34892 7132
rect 612 7028 34892 7076
rect 612 6972 9092 7028
rect 9148 6972 9196 7028
rect 9252 6972 9300 7028
rect 9356 6972 17644 7028
rect 17700 6972 17748 7028
rect 17804 6972 17852 7028
rect 17908 6972 26196 7028
rect 26252 6972 26300 7028
rect 26356 6972 26404 7028
rect 26460 6972 34892 7028
rect 612 6924 34892 6972
rect 612 6868 9092 6924
rect 9148 6868 9196 6924
rect 9252 6868 9300 6924
rect 9356 6868 17644 6924
rect 17700 6868 17748 6924
rect 17804 6868 17852 6924
rect 17908 6868 26196 6924
rect 26252 6868 26300 6924
rect 26356 6868 26404 6924
rect 26460 6868 34892 6924
rect 612 6840 34892 6868
rect 18100 6688 34428 6704
rect 18100 6632 18116 6688
rect 18172 6632 34356 6688
rect 34412 6632 34428 6688
rect 18100 6616 34428 6632
rect 612 5578 34892 5606
rect 612 5522 4816 5578
rect 4872 5522 4920 5578
rect 4976 5522 5024 5578
rect 5080 5522 13368 5578
rect 13424 5522 13472 5578
rect 13528 5522 13576 5578
rect 13632 5522 21920 5578
rect 21976 5522 22024 5578
rect 22080 5522 22128 5578
rect 22184 5522 30472 5578
rect 30528 5522 30576 5578
rect 30632 5522 30680 5578
rect 30736 5522 34892 5578
rect 612 5474 34892 5522
rect 612 5418 4816 5474
rect 4872 5418 4920 5474
rect 4976 5418 5024 5474
rect 5080 5418 13368 5474
rect 13424 5418 13472 5474
rect 13528 5418 13576 5474
rect 13632 5418 21920 5474
rect 21976 5418 22024 5474
rect 22080 5418 22128 5474
rect 22184 5418 30472 5474
rect 30528 5418 30576 5474
rect 30632 5418 30680 5474
rect 30736 5418 34892 5474
rect 612 5370 34892 5418
rect 612 5314 4816 5370
rect 4872 5314 4920 5370
rect 4976 5314 5024 5370
rect 5080 5314 13368 5370
rect 13424 5314 13472 5370
rect 13528 5314 13576 5370
rect 13632 5314 21920 5370
rect 21976 5314 22024 5370
rect 22080 5314 22128 5370
rect 22184 5314 30472 5370
rect 30528 5314 30576 5370
rect 30632 5314 30680 5370
rect 30736 5314 34892 5370
rect 612 5286 34892 5314
rect 612 4024 34892 4052
rect 612 3968 9092 4024
rect 9148 3968 9196 4024
rect 9252 3968 9300 4024
rect 9356 3968 17644 4024
rect 17700 3968 17748 4024
rect 17804 3968 17852 4024
rect 17908 3968 26196 4024
rect 26252 3968 26300 4024
rect 26356 3968 26404 4024
rect 26460 3968 34892 4024
rect 612 3920 34892 3968
rect 612 3864 9092 3920
rect 9148 3864 9196 3920
rect 9252 3864 9300 3920
rect 9356 3864 17644 3920
rect 17700 3864 17748 3920
rect 17804 3864 17852 3920
rect 17908 3864 26196 3920
rect 26252 3864 26300 3920
rect 26356 3864 26404 3920
rect 26460 3864 34892 3920
rect 612 3816 34892 3864
rect 612 3760 9092 3816
rect 9148 3760 9196 3816
rect 9252 3760 9300 3816
rect 9356 3760 17644 3816
rect 17700 3760 17748 3816
rect 17804 3760 17852 3816
rect 17908 3760 26196 3816
rect 26252 3760 26300 3816
rect 26356 3760 26404 3816
rect 26460 3760 34892 3816
rect 612 3732 34892 3760
rect 8356 3448 12028 3464
rect 8356 3392 8372 3448
rect 8428 3392 11956 3448
rect 12012 3392 12028 3448
rect 8356 3376 12028 3392
rect 612 2470 34892 2498
rect 612 2414 4816 2470
rect 4872 2414 4920 2470
rect 4976 2414 5024 2470
rect 5080 2414 13368 2470
rect 13424 2414 13472 2470
rect 13528 2414 13576 2470
rect 13632 2414 21920 2470
rect 21976 2414 22024 2470
rect 22080 2414 22128 2470
rect 22184 2414 30472 2470
rect 30528 2414 30576 2470
rect 30632 2414 30680 2470
rect 30736 2414 34892 2470
rect 612 2366 34892 2414
rect 612 2310 4816 2366
rect 4872 2310 4920 2366
rect 4976 2310 5024 2366
rect 5080 2310 13368 2366
rect 13424 2310 13472 2366
rect 13528 2310 13576 2366
rect 13632 2310 21920 2366
rect 21976 2310 22024 2366
rect 22080 2310 22128 2366
rect 22184 2310 30472 2366
rect 30528 2310 30576 2366
rect 30632 2310 30680 2366
rect 30736 2310 34892 2366
rect 612 2262 34892 2310
rect 612 2206 4816 2262
rect 4872 2206 4920 2262
rect 4976 2206 5024 2262
rect 5080 2206 13368 2262
rect 13424 2206 13472 2262
rect 13528 2206 13576 2262
rect 13632 2206 21920 2262
rect 21976 2206 22024 2262
rect 22080 2206 22128 2262
rect 22184 2206 30472 2262
rect 30528 2206 30576 2262
rect 30632 2206 30680 2262
rect 30736 2206 34892 2262
rect 612 2178 34892 2206
rect 18324 2008 31964 2024
rect 18324 1952 18340 2008
rect 18396 1952 31892 2008
rect 31948 1952 31964 2008
rect 18324 1936 31964 1952
rect 19892 1468 33756 1484
rect 19892 1412 19908 1468
rect 19964 1412 33684 1468
rect 33740 1412 33756 1468
rect 19892 1396 33756 1412
rect 17988 1288 32860 1304
rect 17988 1232 18004 1288
rect 18060 1232 32788 1288
rect 32844 1232 32860 1288
rect 17988 1216 32860 1232
rect 19892 1108 33868 1124
rect 19892 1052 19908 1108
rect 19964 1052 33796 1108
rect 33852 1052 33868 1108
rect 19892 1036 33868 1052
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__A1 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 20048 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__I0
timestamp 1654395037
transform 1 0 30240 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__I1
timestamp 1654395037
transform -1 0 19264 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__I
timestamp 1654395037
transform -1 0 18592 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__I
timestamp 1654395037
transform 1 0 22064 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__A2
timestamp 1654395037
transform 1 0 18816 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__A3
timestamp 1654395037
transform 1 0 20048 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__A2
timestamp 1654395037
transform 1 0 23520 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__B
timestamp 1654395037
transform 1 0 33152 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__A1
timestamp 1654395037
transform -1 0 27552 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__A2
timestamp 1654395037
transform 1 0 24304 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__A2
timestamp 1654395037
transform 1 0 24304 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__A1
timestamp 1654395037
transform 1 0 10640 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__285__I
timestamp 1654395037
transform 1 0 9744 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__294__A1
timestamp 1654395037
transform 1 0 11200 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__295__I
timestamp 1654395037
transform -1 0 12992 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__312__A2
timestamp 1654395037
transform 1 0 18816 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__312__B
timestamp 1654395037
transform 1 0 16688 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__330__A1
timestamp 1654395037
transform -1 0 6944 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__A1
timestamp 1654395037
transform -1 0 20832 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__B
timestamp 1654395037
transform -1 0 22400 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__341__A1
timestamp 1654395037
transform -1 0 21056 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__344__A2
timestamp 1654395037
transform -1 0 21280 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__345__A1
timestamp 1654395037
transform -1 0 28672 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__A1
timestamp 1654395037
transform 1 0 34384 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__I1
timestamp 1654395037
transform -1 0 8512 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__S
timestamp 1654395037
transform 1 0 6944 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__A1
timestamp 1654395037
transform -1 0 26432 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__I
timestamp 1654395037
transform -1 0 28448 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__A1
timestamp 1654395037
transform 1 0 27104 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__A1
timestamp 1654395037
transform -1 0 24864 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__365__A2
timestamp 1654395037
transform 1 0 26880 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__A1
timestamp 1654395037
transform 1 0 25984 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__376__A2
timestamp 1654395037
transform 1 0 9744 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__378__I
timestamp 1654395037
transform 1 0 19712 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__379__A1
timestamp 1654395037
transform 1 0 12208 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__390__A1
timestamp 1654395037
transform -1 0 12656 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__A1
timestamp 1654395037
transform 1 0 18368 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__398__A2
timestamp 1654395037
transform -1 0 22736 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__406__A1
timestamp 1654395037
transform 1 0 17472 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__406__A2
timestamp 1654395037
transform -1 0 14672 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__406__A3
timestamp 1654395037
transform 1 0 17696 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__A1
timestamp 1654395037
transform 1 0 17024 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__A2
timestamp 1654395037
transform 1 0 22960 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__B
timestamp 1654395037
transform 1 0 17136 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__410__A2
timestamp 1654395037
transform 1 0 3024 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__412__A3
timestamp 1654395037
transform 1 0 11312 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__416__A2
timestamp 1654395037
transform -1 0 1456 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__417__A2
timestamp 1654395037
transform 1 0 3920 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__421__A1
timestamp 1654395037
transform -1 0 1792 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__422__A2
timestamp 1654395037
transform -1 0 2352 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__423__A1
timestamp 1654395037
transform 1 0 1904 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__425__A2
timestamp 1654395037
transform -1 0 6944 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__435__A1
timestamp 1654395037
transform 1 0 24304 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__435__C
timestamp 1654395037
transform 1 0 26992 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__436__A1
timestamp 1654395037
transform 1 0 33040 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__439__A1
timestamp 1654395037
transform -1 0 25312 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__440__A1
timestamp 1654395037
transform 1 0 34048 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__A1
timestamp 1654395037
transform -1 0 30352 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__442__A1
timestamp 1654395037
transform -1 0 22176 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__445__CLKN
timestamp 1654395037
transform -1 0 19712 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__445__SETN
timestamp 1654395037
transform 1 0 19040 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__446__CLKN
timestamp 1654395037
transform -1 0 23744 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__446__SETN
timestamp 1654395037
transform 1 0 23744 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__CLKN
timestamp 1654395037
transform -1 0 24192 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__447__SETN
timestamp 1654395037
transform 1 0 24192 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__CLK
timestamp 1654395037
transform -1 0 23072 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__448__RN
timestamp 1654395037
transform 1 0 26656 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__449__CLK
timestamp 1654395037
transform -1 0 25088 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__449__RN
timestamp 1654395037
transform 1 0 30016 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__CLK
timestamp 1654395037
transform 1 0 22624 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__450__SETN
timestamp 1654395037
transform 1 0 15792 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__CLK
timestamp 1654395037
transform 1 0 11760 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__451__RN
timestamp 1654395037
transform 1 0 8176 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__452__CLK
timestamp 1654395037
transform -1 0 28896 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__453__CLK
timestamp 1654395037
transform 1 0 23968 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__454__CLK
timestamp 1654395037
transform 1 0 20160 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__CLK
timestamp 1654395037
transform -1 0 19936 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__SETN
timestamp 1654395037
transform 1 0 19264 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__456__CLK
timestamp 1654395037
transform 1 0 21616 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__456__RN
timestamp 1654395037
transform 1 0 16352 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__CLKN
timestamp 1654395037
transform -1 0 4928 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__457__RN
timestamp 1654395037
transform 1 0 4704 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__CLKN
timestamp 1654395037
transform 1 0 5376 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__458__SETN
timestamp 1654395037
transform 1 0 5600 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__459__CLKN
timestamp 1654395037
transform 1 0 4928 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__459__RN
timestamp 1654395037
transform 1 0 5152 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__CLKN
timestamp 1654395037
transform 1 0 16912 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__460__SETN
timestamp 1654395037
transform 1 0 9520 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__461__CLKN
timestamp 1654395037
transform -1 0 23520 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__461__RN
timestamp 1654395037
transform 1 0 20160 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__462__CLKN
timestamp 1654395037
transform 1 0 19376 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__462__SETN
timestamp 1654395037
transform 1 0 14560 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__463__CLKN
timestamp 1654395037
transform -1 0 13216 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__463__RN
timestamp 1654395037
transform 1 0 9296 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__CLK
timestamp 1654395037
transform 1 0 3472 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__464__RN
timestamp 1654395037
transform 1 0 3696 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__CLK
timestamp 1654395037
transform 1 0 3248 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__465__SETN
timestamp 1654395037
transform 1 0 4816 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__466__CLK
timestamp 1654395037
transform 1 0 12880 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__466__RN
timestamp 1654395037
transform 1 0 6384 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__467__CLK
timestamp 1654395037
transform 1 0 17696 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__467__SETN
timestamp 1654395037
transform 1 0 18816 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__468__CLK
timestamp 1654395037
transform -1 0 19264 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__468__RN
timestamp 1654395037
transform 1 0 18144 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__469__CLK
timestamp 1654395037
transform 1 0 18816 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__469__RN
timestamp 1654395037
transform 1 0 23072 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__470__CLK
timestamp 1654395037
transform -1 0 22624 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__470__RN
timestamp 1654395037
transform 1 0 22624 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__CLK
timestamp 1654395037
transform -1 0 26656 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__471__SETN
timestamp 1654395037
transform 1 0 25984 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__472__CLK
timestamp 1654395037
transform -1 0 21728 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__472__RN
timestamp 1654395037
transform 1 0 21728 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__473__CLK
timestamp 1654395037
transform -1 0 20384 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__473__RN
timestamp 1654395037
transform 1 0 20384 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__474__CLK
timestamp 1654395037
transform 1 0 29568 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__474__SETN
timestamp 1654395037
transform 1 0 29344 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__475__CLK
timestamp 1654395037
transform 1 0 25088 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__475__RN
timestamp 1654395037
transform 1 0 24528 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__476__CLK
timestamp 1654395037
transform 1 0 12992 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__477__CLK
timestamp 1654395037
transform -1 0 30800 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__477__D
timestamp 1654395037
transform 1 0 34272 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__478__CLK
timestamp 1654395037
transform 1 0 24864 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__478__D
timestamp 1654395037
transform 1 0 26656 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__479__CLK
timestamp 1654395037
transform -1 0 28224 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__480__CLK
timestamp 1654395037
transform 1 0 25424 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__480__SETN
timestamp 1654395037
transform 1 0 18592 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__CLK
timestamp 1654395037
transform 1 0 23744 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__481__RN
timestamp 1654395037
transform 1 0 17024 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__482__CLKN
timestamp 1654395037
transform 1 0 13104 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__482__RN
timestamp 1654395037
transform 1 0 9520 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__483__CLKN
timestamp 1654395037
transform 1 0 6832 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__483__SETN
timestamp 1654395037
transform 1 0 7056 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__CLKN
timestamp 1654395037
transform 1 0 4144 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__RN
timestamp 1654395037
transform 1 0 6272 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__485__CLKN
timestamp 1654395037
transform 1 0 18816 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__485__SETN
timestamp 1654395037
transform 1 0 14336 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__486__CLKN
timestamp 1654395037
transform 1 0 3248 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__486__RN
timestamp 1654395037
transform 1 0 1904 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__487__CLKN
timestamp 1654395037
transform 1 0 6384 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__487__SETN
timestamp 1654395037
transform 1 0 6496 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__488__CLKN
timestamp 1654395037
transform 1 0 2576 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__488__RN
timestamp 1654395037
transform 1 0 2800 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__489__CLK
timestamp 1654395037
transform 1 0 3472 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__489__RN
timestamp 1654395037
transform 1 0 3696 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__490__CLK
timestamp 1654395037
transform 1 0 1344 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__490__SETN
timestamp 1654395037
transform 1 0 2128 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__491__CLK
timestamp 1654395037
transform 1 0 1456 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__491__RN
timestamp 1654395037
transform 1 0 1680 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__492__CLK
timestamp 1654395037
transform 1 0 18816 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__492__SETN
timestamp 1654395037
transform 1 0 14560 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__493__CLK
timestamp 1654395037
transform 1 0 33488 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__493__SETN
timestamp 1654395037
transform 1 0 23184 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__494__CLK
timestamp 1654395037
transform -1 0 33936 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__494__RN
timestamp 1654395037
transform 1 0 33712 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__495__CLK
timestamp 1654395037
transform 1 0 18592 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__495__RN
timestamp 1654395037
transform 1 0 31472 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__496__RN
timestamp 1654395037
transform 1 0 21840 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__497__SETN
timestamp 1654395037
transform 1 0 28896 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__498__RN
timestamp 1654395037
transform 1 0 20384 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__499__RN
timestamp 1654395037
transform 1 0 19936 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__500__SETN
timestamp 1654395037
transform 1 0 19488 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__501__RN
timestamp 1654395037
transform 1 0 29120 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1654395037
transform -1 0 18256 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1654395037
transform -1 0 18032 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1654395037
transform -1 0 21504 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1654395037
transform -1 0 17696 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1654395037
transform -1 0 1904 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1654395037
transform -1 0 19488 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1654395037
transform -1 0 20160 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1654395037
transform -1 0 17808 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1654395037
transform -1 0 18480 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1654395037
transform -1 0 17584 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1654395037
transform -1 0 18144 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output12_I
timestamp 1654395037
transform -1 0 6608 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 896 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_34 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 4480 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 4928 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 5824 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_50
timestamp 1654395037
transform 1 0 6272 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 6496 0 1 784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55
timestamp 1654395037
transform 1 0 6832 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67
timestamp 1654395037
transform 1 0 8176 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99
timestamp 1654395037
transform 1 0 11760 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_103
timestamp 1654395037
transform 1 0 12208 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105
timestamp 1654395037
transform 1 0 12432 0 1 784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_112
timestamp 1654395037
transform 1 0 13216 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_144
timestamp 1654395037
transform 1 0 16800 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_148
timestamp 1654395037
transform 1 0 17248 0 1 784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_161
timestamp 1654395037
transform 1 0 18704 0 1 784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_254
timestamp 1654395037
transform 1 0 29120 0 1 784
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_91
timestamp 1654395037
transform 1 0 10864 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_93
timestamp 1654395037
transform 1 0 11088 0 -1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_109
timestamp 1654395037
transform 1 0 12880 0 -1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_126
timestamp 1654395037
transform 1 0 14784 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_128
timestamp 1654395037
transform 1 0 15008 0 -1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_140
timestamp 1654395037
transform 1 0 16352 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_148
timestamp 1654395037
transform 1 0 17248 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_210
timestamp 1654395037
transform 1 0 24192 0 -1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_213
timestamp 1654395037
transform 1 0 24528 0 -1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_260
timestamp 1654395037
transform 1 0 29792 0 -1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_2
timestamp 1654395037
transform 1 0 896 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_10
timestamp 1654395037
transform 1 0 1792 0 1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_109
timestamp 1654395037
transform 1 0 12880 0 1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_215
timestamp 1654395037
transform 1 0 24752 0 1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_220
timestamp 1654395037
transform 1 0 25312 0 1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_259
timestamp 1654395037
transform 1 0 29680 0 1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_266
timestamp 1654395037
transform 1 0 30464 0 1 2352
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_2
timestamp 1654395037
transform 1 0 896 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_6
timestamp 1654395037
transform 1 0 1344 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_8
timestamp 1654395037
transform 1 0 1568 0 -1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_15
timestamp 1654395037
transform 1 0 2352 0 -1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_22
timestamp 1654395037
transform 1 0 3136 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_24
timestamp 1654395037
transform 1 0 3360 0 -1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_53
timestamp 1654395037
transform 1 0 6608 0 -1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_139
timestamp 1654395037
transform 1 0 16240 0 -1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_200
timestamp 1654395037
transform 1 0 23072 0 -1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_213
timestamp 1654395037
transform 1 0 24528 0 -1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_2
timestamp 1654395037
transform 1 0 896 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_159
timestamp 1654395037
transform 1 0 18480 0 1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_192
timestamp 1654395037
transform 1 0 22176 0 1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_266
timestamp 1654395037
transform 1 0 30464 0 1 3920
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_36
timestamp 1654395037
transform 1 0 4704 0 -1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_78
timestamp 1654395037
transform 1 0 9408 0 -1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_106
timestamp 1654395037
transform 1 0 12544 0 -1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_216
timestamp 1654395037
transform 1 0 24864 0 -1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_249
timestamp 1654395037
transform 1 0 28560 0 -1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_302
timestamp 1654395037
transform 1 0 34496 0 -1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_2
timestamp 1654395037
transform 1 0 896 0 1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_45
timestamp 1654395037
transform 1 0 5712 0 1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_115
timestamp 1654395037
transform 1 0 13552 0 1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_223
timestamp 1654395037
transform 1 0 25648 0 1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_266
timestamp 1654395037
transform 1 0 30464 0 1 5488
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_2
timestamp 1654395037
transform 1 0 896 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_7_6
timestamp 1654395037
transform 1 0 1344 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_8
timestamp 1654395037
transform 1 0 1568 0 -1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_15
timestamp 1654395037
transform 1 0 2352 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_164
timestamp 1654395037
transform 1 0 19040 0 -1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_213
timestamp 1654395037
transform 1 0 24528 0 -1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_250
timestamp 1654395037
transform 1 0 28672 0 -1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_2
timestamp 1654395037
transform 1 0 896 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_10
timestamp 1654395037
transform 1 0 1792 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_8_14
timestamp 1654395037
transform 1 0 2240 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_50
timestamp 1654395037
transform 1 0 6272 0 1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_98
timestamp 1654395037
transform 1 0 11648 0 1 7056
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_109
timestamp 1654395037
transform 1 0 12880 0 -1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_134
timestamp 1654395037
transform 1 0 15680 0 -1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_10_2
timestamp 1654395037
transform 1 0 896 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_4
timestamp 1654395037
transform 1 0 1120 0 1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1654395037
transform 1 0 12432 0 1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_164
timestamp 1654395037
transform 1 0 19040 0 1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_198
timestamp 1654395037
transform 1 0 22848 0 1 8624
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_100
timestamp 1654395037
transform 1 0 11872 0 -1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_109
timestamp 1654395037
transform 1 0 12880 0 -1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_201
timestamp 1654395037
transform 1 0 23184 0 -1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_292
timestamp 1654395037
transform 1 0 33376 0 -1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_81
timestamp 1654395037
transform 1 0 9744 0 1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_162
timestamp 1654395037
transform 1 0 18816 0 1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_266
timestamp 1654395037
transform 1 0 30464 0 1 10192
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_2
timestamp 1654395037
transform 1 0 896 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_16
timestamp 1654395037
transform 1 0 2464 0 -1 11760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_65
timestamp 1654395037
transform 1 0 7952 0 -1 11760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_179
timestamp 1654395037
transform 1 0 20720 0 -1 11760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_266
timestamp 1654395037
transform 1 0 30464 0 -1 11760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_2
timestamp 1654395037
transform 1 0 896 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_14_6
timestamp 1654395037
transform 1 0 1344 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_8
timestamp 1654395037
transform 1 0 1568 0 1 11760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_197
timestamp 1654395037
transform 1 0 22736 0 1 11760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_264
timestamp 1654395037
transform 1 0 30240 0 1 11760
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 672 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1654395037
transform -1 0 34832 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1654395037
transform 1 0 672 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1654395037
transform -1 0 34832 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1654395037
transform 1 0 672 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1654395037
transform -1 0 34832 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1654395037
transform 1 0 672 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1654395037
transform -1 0 34832 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1654395037
transform 1 0 672 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1654395037
transform -1 0 34832 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1654395037
transform 1 0 672 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1654395037
transform -1 0 34832 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1654395037
transform 1 0 672 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1654395037
transform -1 0 34832 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1654395037
transform 1 0 672 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1654395037
transform -1 0 34832 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1654395037
transform 1 0 672 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1654395037
transform -1 0 34832 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1654395037
transform 1 0 672 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1654395037
transform -1 0 34832 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1654395037
transform 1 0 672 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1654395037
transform -1 0 34832 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1654395037
transform 1 0 672 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1654395037
transform -1 0 34832 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1654395037
transform 1 0 672 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1654395037
transform -1 0 34832 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1654395037
transform 1 0 672 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1654395037
transform -1 0 34832 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1654395037
transform 1 0 672 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1654395037
transform -1 0 34832 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_30
timestamp 1654395037
transform 1 0 6608 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_31
timestamp 1654395037
transform 1 0 12544 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_32
timestamp 1654395037
transform 1 0 18480 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_33
timestamp 1654395037
transform 1 0 24416 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_34
timestamp 1654395037
transform 1 0 30352 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_35
timestamp 1654395037
transform 1 0 12656 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_36
timestamp 1654395037
transform 1 0 24640 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_37
timestamp 1654395037
transform 1 0 6608 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_38
timestamp 1654395037
transform 1 0 18592 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_39
timestamp 1654395037
transform 1 0 30576 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_40
timestamp 1654395037
transform 1 0 12656 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_41
timestamp 1654395037
transform 1 0 24640 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_42
timestamp 1654395037
transform 1 0 6608 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_43
timestamp 1654395037
transform 1 0 18592 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_44
timestamp 1654395037
transform 1 0 30576 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_45
timestamp 1654395037
transform 1 0 12656 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_46
timestamp 1654395037
transform 1 0 24640 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_47
timestamp 1654395037
transform 1 0 6608 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_48
timestamp 1654395037
transform 1 0 18592 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_49
timestamp 1654395037
transform 1 0 30576 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_50
timestamp 1654395037
transform 1 0 12656 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_51
timestamp 1654395037
transform 1 0 24640 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_52
timestamp 1654395037
transform 1 0 6608 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_53
timestamp 1654395037
transform 1 0 18592 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_54
timestamp 1654395037
transform 1 0 30576 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_55
timestamp 1654395037
transform 1 0 12656 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_56
timestamp 1654395037
transform 1 0 24640 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_57
timestamp 1654395037
transform 1 0 6608 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_58
timestamp 1654395037
transform 1 0 18592 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_59
timestamp 1654395037
transform 1 0 30576 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_60
timestamp 1654395037
transform 1 0 12656 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_61
timestamp 1654395037
transform 1 0 24640 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_62
timestamp 1654395037
transform 1 0 6608 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_63
timestamp 1654395037
transform 1 0 18592 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_64
timestamp 1654395037
transform 1 0 30576 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_65
timestamp 1654395037
transform 1 0 12656 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_66
timestamp 1654395037
transform 1 0 24640 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_67
timestamp 1654395037
transform 1 0 6608 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_68
timestamp 1654395037
transform 1 0 12544 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_69
timestamp 1654395037
transform 1 0 18480 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_70
timestamp 1654395037
transform 1 0 24416 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_71
timestamp 1654395037
transform 1 0 30352 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _220_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 21504 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _221_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 19040 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _222_
timestamp 1654395037
transform 1 0 29008 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _223_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 27776 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _224_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 28560 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _225_
timestamp 1654395037
transform 1 0 22288 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _226_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 22400 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _227_
timestamp 1654395037
transform -1 0 18368 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _228_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 17584 0 -1 5488
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _229_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 18928 0 -1 5488
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _230_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 19264 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _231_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 20832 0 1 11760
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _232_
timestamp 1654395037
transform 1 0 19152 0 1 11760
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _233_
timestamp 1654395037
transform -1 0 18144 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _234_
timestamp 1654395037
transform -1 0 33152 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _235_
timestamp 1654395037
transform -1 0 19600 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _236_
timestamp 1654395037
transform -1 0 20048 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _237_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 20272 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _238_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 17696 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _239_
timestamp 1654395037
transform 1 0 22064 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _240_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 19152 0 1 8624
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _241_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 20608 0 1 8624
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _242_
timestamp 1654395037
transform 1 0 21168 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _243_
timestamp 1654395037
transform 1 0 19040 0 -1 11760
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _244_
timestamp 1654395037
transform -1 0 19040 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _245_
timestamp 1654395037
transform 1 0 29232 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _246_
timestamp 1654395037
transform -1 0 33712 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _247_
timestamp 1654395037
transform -1 0 34048 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _248_
timestamp 1654395037
transform 1 0 4928 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _249_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 6832 0 1 8624
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _250_
timestamp 1654395037
transform -1 0 17472 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _251_
timestamp 1654395037
transform -1 0 16800 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _252_
timestamp 1654395037
transform 1 0 16800 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _253_
timestamp 1654395037
transform 1 0 15232 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _254_
timestamp 1654395037
transform 1 0 27328 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _255_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 30464 0 1 3920
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _256_
timestamp 1654395037
transform 1 0 28224 0 1 3920
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _257_
timestamp 1654395037
transform 1 0 29792 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _258_
timestamp 1654395037
transform 1 0 21056 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _259_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 22400 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _260_
timestamp 1654395037
transform -1 0 17248 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _261_
timestamp 1654395037
transform -1 0 27664 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _262_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 30464 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _263_
timestamp 1654395037
transform 1 0 22960 0 -1 7056
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _264_
timestamp 1654395037
transform 1 0 26208 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _265_
timestamp 1654395037
transform 1 0 22960 0 1 5488
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _266_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 23520 0 -1 5488
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _267_
timestamp 1654395037
transform -1 0 18480 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _268_
timestamp 1654395037
transform 1 0 17136 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _269_
timestamp 1654395037
transform -1 0 5712 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _270_
timestamp 1654395037
transform 1 0 7728 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _271_
timestamp 1654395037
transform 1 0 21504 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _272_
timestamp 1654395037
transform -1 0 26208 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _273_
timestamp 1654395037
transform 1 0 11984 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _274_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 13664 0 1 3920
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _275_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 11984 0 -1 2352
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _276_
timestamp 1654395037
transform 1 0 5936 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _277_
timestamp 1654395037
transform -1 0 14560 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _278_
timestamp 1654395037
transform -1 0 10416 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _279_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 7840 0 -1 3920
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _280_
timestamp 1654395037
transform 1 0 24864 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _281_
timestamp 1654395037
transform -1 0 16688 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _282_
timestamp 1654395037
transform -1 0 10304 0 -1 3920
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _283_
timestamp 1654395037
transform 1 0 7728 0 1 3920
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _284_
timestamp 1654395037
transform -1 0 2352 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _285_
timestamp 1654395037
transform -1 0 9296 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _286_
timestamp 1654395037
transform 1 0 6944 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _287_
timestamp 1654395037
transform 1 0 5824 0 -1 2352
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _288_
timestamp 1654395037
transform -1 0 8288 0 -1 2352
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _289_
timestamp 1654395037
transform 1 0 6832 0 1 2352
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _290_
timestamp 1654395037
transform -1 0 3136 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _291_
timestamp 1654395037
transform 1 0 5712 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _292_
timestamp 1654395037
transform -1 0 11088 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _293_
timestamp 1654395037
transform -1 0 6608 0 1 3920
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _294_
timestamp 1654395037
transform -1 0 11424 0 -1 5488
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _295_
timestamp 1654395037
transform -1 0 12656 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _296_
timestamp 1654395037
transform 1 0 4928 0 1 3920
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _297_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 7504 0 -1 5488
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _298_
timestamp 1654395037
transform -1 0 6496 0 -1 5488
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _299_
timestamp 1654395037
transform 1 0 8288 0 -1 2352
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _300_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 13664 0 1 3920
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _301_
timestamp 1654395037
transform 1 0 13440 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _302_
timestamp 1654395037
transform -1 0 12544 0 1 3920
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _303_
timestamp 1654395037
transform 1 0 12992 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _304_
timestamp 1654395037
transform -1 0 24528 0 -1 3920
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _305_
timestamp 1654395037
transform 1 0 22960 0 -1 2352
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _306_
timestamp 1654395037
transform 1 0 22064 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _307_
timestamp 1654395037
transform -1 0 20496 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _308_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 20384 0 -1 2352
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _309_
timestamp 1654395037
transform -1 0 14560 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _310_
timestamp 1654395037
transform 1 0 12992 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _311_
timestamp 1654395037
transform -1 0 14224 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _312_
timestamp 1654395037
transform 1 0 15120 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _313_
timestamp 1654395037
transform -1 0 15344 0 -1 3920
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _314_
timestamp 1654395037
transform 1 0 15344 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _315_
timestamp 1654395037
transform -1 0 19376 0 1 2352
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _316_
timestamp 1654395037
transform -1 0 16352 0 -1 2352
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _317_
timestamp 1654395037
transform 1 0 10304 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _318_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 12208 0 -1 3920
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _319_
timestamp 1654395037
transform -1 0 10640 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _320_
timestamp 1654395037
transform 1 0 4368 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _321_
timestamp 1654395037
transform -1 0 9072 0 1 2352
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _322_
timestamp 1654395037
transform 1 0 5040 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _323_
timestamp 1654395037
transform -1 0 11760 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _324_
timestamp 1654395037
transform -1 0 7728 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _325_
timestamp 1654395037
transform 1 0 7728 0 -1 8624
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _326_
timestamp 1654395037
transform 1 0 8960 0 -1 3920
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _327_
timestamp 1654395037
transform 1 0 3920 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _328_
timestamp 1654395037
transform 1 0 6832 0 1 5488
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _329_
timestamp 1654395037
transform 1 0 5040 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _330_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 6496 0 -1 5488
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _331_
timestamp 1654395037
transform 1 0 9744 0 -1 5488
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _332_
timestamp 1654395037
transform 1 0 8512 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _333_
timestamp 1654395037
transform -1 0 2352 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _334_
timestamp 1654395037
transform -1 0 9744 0 1 5488
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _335_
timestamp 1654395037
transform 1 0 8848 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _336_
timestamp 1654395037
transform 1 0 7168 0 -1 8624
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _337_
timestamp 1654395037
transform -1 0 9184 0 1 5488
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _338_
timestamp 1654395037
transform -1 0 6608 0 1 5488
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _339_
timestamp 1654395037
transform -1 0 29120 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _340_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 28112 0 -1 3920
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _341_
timestamp 1654395037
transform -1 0 30128 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _342_
timestamp 1654395037
transform 1 0 30800 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _343_
timestamp 1654395037
transform 1 0 25424 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _344_
timestamp 1654395037
transform 1 0 28112 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _345_
timestamp 1654395037
transform 1 0 26880 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _346_
timestamp 1654395037
transform 1 0 26880 0 -1 3920
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _347_
timestamp 1654395037
transform -1 0 26768 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _348_
timestamp 1654395037
transform -1 0 28112 0 1 2352
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _349_
timestamp 1654395037
transform -1 0 25984 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _350_
timestamp 1654395037
transform 1 0 12768 0 1 11760
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _351_
timestamp 1654395037
transform 1 0 11200 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _352_
timestamp 1654395037
transform -1 0 30576 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _353_
timestamp 1654395037
transform -1 0 25424 0 1 5488
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _354_
timestamp 1654395037
transform -1 0 22064 0 -1 7056
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _355_
timestamp 1654395037
transform -1 0 20720 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _356_
timestamp 1654395037
transform -1 0 14784 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _357_
timestamp 1654395037
transform 1 0 9072 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _358_
timestamp 1654395037
transform 1 0 9744 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _359_
timestamp 1654395037
transform -1 0 30464 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _360_
timestamp 1654395037
transform -1 0 18592 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _361_
timestamp 1654395037
transform 1 0 25872 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _362_
timestamp 1654395037
transform 1 0 24864 0 -1 10192
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _363_
timestamp 1654395037
transform -1 0 27216 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _364_
timestamp 1654395037
transform 1 0 23296 0 -1 10192
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _365_
timestamp 1654395037
transform 1 0 26208 0 -1 10192
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _366_
timestamp 1654395037
transform -1 0 22624 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _367_
timestamp 1654395037
transform 1 0 17248 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _368_
timestamp 1654395037
transform -1 0 12432 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _369_
timestamp 1654395037
transform -1 0 11648 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _370_
timestamp 1654395037
transform -1 0 12656 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _371_
timestamp 1654395037
transform 1 0 12544 0 1 8624
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _372_
timestamp 1654395037
transform -1 0 8960 0 1 8624
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _373_
timestamp 1654395037
transform 1 0 9856 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _374_
timestamp 1654395037
transform -1 0 11760 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _375_
timestamp 1654395037
transform 1 0 14560 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _376_
timestamp 1654395037
transform -1 0 12432 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _377_
timestamp 1654395037
transform -1 0 11088 0 1 8624
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _378_
timestamp 1654395037
transform 1 0 32368 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _379_
timestamp 1654395037
transform -1 0 12096 0 -1 8624
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _380_
timestamp 1654395037
transform 1 0 9632 0 -1 8624
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _381_
timestamp 1654395037
transform -1 0 11200 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _382_
timestamp 1654395037
transform 1 0 13664 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _383_
timestamp 1654395037
transform 1 0 12432 0 1 7056
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _384_
timestamp 1654395037
transform 1 0 13216 0 -1 8624
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _385_
timestamp 1654395037
transform 1 0 7280 0 1 7056
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _386_
timestamp 1654395037
transform -1 0 6272 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _387_
timestamp 1654395037
transform -1 0 9856 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _388_
timestamp 1654395037
transform 1 0 11984 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _389_
timestamp 1654395037
transform -1 0 9632 0 -1 8624
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _390_
timestamp 1654395037
transform -1 0 13440 0 -1 7056
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _391_
timestamp 1654395037
transform -1 0 11312 0 -1 8624
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _392_
timestamp 1654395037
transform -1 0 10976 0 -1 10192
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _393_
timestamp 1654395037
transform -1 0 9744 0 1 8624
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _394_
timestamp 1654395037
transform 1 0 12096 0 -1 8624
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _395_
timestamp 1654395037
transform -1 0 15904 0 -1 7056
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _396_
timestamp 1654395037
transform 1 0 14784 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _397_
timestamp 1654395037
transform -1 0 14560 0 1 7056
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _398_
timestamp 1654395037
transform 1 0 18256 0 -1 10192
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _399_
timestamp 1654395037
transform -1 0 20272 0 -1 10192
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _400_
timestamp 1654395037
transform 1 0 16128 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _401_
timestamp 1654395037
transform -1 0 11872 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _402_
timestamp 1654395037
transform -1 0 11088 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _403_
timestamp 1654395037
transform -1 0 9744 0 -1 11760
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _404_
timestamp 1654395037
transform -1 0 11760 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _405_
timestamp 1654395037
transform 1 0 14560 0 1 10192
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _406_
timestamp 1654395037
transform 1 0 15120 0 -1 10192
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _407_
timestamp 1654395037
transform -1 0 18256 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _408_
timestamp 1654395037
transform -1 0 17136 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _409_
timestamp 1654395037
transform -1 0 17024 0 1 10192
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _410_
timestamp 1654395037
transform -1 0 11200 0 1 11760
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _411_
timestamp 1654395037
transform -1 0 9744 0 1 10192
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _412_
timestamp 1654395037
transform 1 0 12992 0 -1 10192
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _413_
timestamp 1654395037
transform 1 0 14224 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _414_
timestamp 1654395037
transform 1 0 3472 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _415_
timestamp 1654395037
transform -1 0 3584 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _416_
timestamp 1654395037
transform 1 0 2352 0 1 8624
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _417_
timestamp 1654395037
transform -1 0 5600 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _418_
timestamp 1654395037
transform 1 0 3584 0 1 8624
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _419_
timestamp 1654395037
transform -1 0 6832 0 -1 10192
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _420_
timestamp 1654395037
transform -1 0 6384 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _421_
timestamp 1654395037
transform 1 0 5376 0 1 10192
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _422_
timestamp 1654395037
transform 1 0 4592 0 1 8624
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _423_
timestamp 1654395037
transform -1 0 5600 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _424_
timestamp 1654395037
transform -1 0 2464 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _425_
timestamp 1654395037
transform -1 0 9072 0 -1 10192
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _426_
timestamp 1654395037
transform 1 0 6832 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _427_
timestamp 1654395037
transform 1 0 6832 0 -1 10192
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _428_
timestamp 1654395037
transform 1 0 7392 0 -1 10192
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _429_
timestamp 1654395037
transform 1 0 7728 0 1 10192
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _430_
timestamp 1654395037
transform -1 0 12544 0 -1 5488
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _431_
timestamp 1654395037
transform 1 0 15904 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _432_
timestamp 1654395037
transform 1 0 13664 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _433_
timestamp 1654395037
transform 1 0 12880 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _434_
timestamp 1654395037
transform -1 0 25536 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _435_
timestamp 1654395037
transform -1 0 21392 0 -1 8624
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _436_
timestamp 1654395037
transform -1 0 25760 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _437_
timestamp 1654395037
transform 1 0 22288 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _438_
timestamp 1654395037
transform -1 0 25984 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _439_
timestamp 1654395037
transform -1 0 25872 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _440_
timestamp 1654395037
transform 1 0 27552 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _441_
timestamp 1654395037
transform -1 0 26992 0 -1 8624
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _442_
timestamp 1654395037
transform 1 0 28672 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _443_
timestamp 1654395037
transform 1 0 31024 0 -1 8624
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _444_
timestamp 1654395037
transform 1 0 32816 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1  _445_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 30576 0 1 11760
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1  _446_
timestamp 1654395037
transform 1 0 25984 0 -1 11760
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1  _447_
timestamp 1654395037
transform 1 0 24640 0 1 11760
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _447__15 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 18704 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _448_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 30576 0 1 8624
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _449_
timestamp 1654395037
transform -1 0 24640 0 -1 11760
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _450_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 16016 0 -1 8624
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _451_
timestamp 1654395037
transform 1 0 14672 0 1 11760
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _452_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 23408 0 1 3920
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _453_
timestamp 1654395037
transform 1 0 20272 0 -1 5488
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _454_
timestamp 1654395037
transform 1 0 19712 0 1 5488
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _455_
timestamp 1654395037
transform 1 0 30352 0 -1 3920
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _456_
timestamp 1654395037
transform 1 0 17248 0 -1 3920
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _457_ pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 896 0 -1 2352
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1  _458_
timestamp 1654395037
transform 1 0 1904 0 1 2352
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _459_
timestamp 1654395037
transform 1 0 1120 0 1 3920
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1  _460_
timestamp 1654395037
transform 1 0 13552 0 -1 5488
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _461_
timestamp 1654395037
transform 1 0 20496 0 1 2352
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1  _462_
timestamp 1654395037
transform 1 0 14560 0 1 2352
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _463_
timestamp 1654395037
transform 1 0 9072 0 1 2352
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _464_
timestamp 1654395037
transform 1 0 896 0 -1 5488
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _465_
timestamp 1654395037
transform 1 0 1008 0 1 5488
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _466_
timestamp 1654395037
transform 1 0 8400 0 -1 7056
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _467_
timestamp 1654395037
transform 1 0 30576 0 -1 2352
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _468_
timestamp 1654395037
transform 1 0 30800 0 1 2352
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _469_
timestamp 1654395037
transform 1 0 24864 0 -1 2352
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _470_
timestamp 1654395037
transform 1 0 29568 0 -1 5488
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _471_
timestamp 1654395037
transform 1 0 25760 0 1 5488
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _472_
timestamp 1654395037
transform -1 0 34608 0 1 5488
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _473_
timestamp 1654395037
transform -1 0 34608 0 1 3920
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _474_
timestamp 1654395037
transform -1 0 32816 0 -1 7056
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _475_
timestamp 1654395037
transform -1 0 28672 0 -1 7056
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _476_
timestamp 1654395037
transform 1 0 12880 0 -1 11760
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _477_
timestamp 1654395037
transform 1 0 26880 0 1 7056
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _478_
timestamp 1654395037
transform 1 0 21392 0 -1 8624
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _479_
timestamp 1654395037
transform -1 0 25984 0 1 10192
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _480_
timestamp 1654395037
transform 1 0 18816 0 1 7056
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _481_
timestamp 1654395037
transform -1 0 22736 0 1 10192
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _482_
timestamp 1654395037
transform 1 0 9744 0 1 5488
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1  _483_
timestamp 1654395037
transform 1 0 4368 0 -1 7056
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _484_
timestamp 1654395037
transform 1 0 2464 0 1 7056
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1  _485_
timestamp 1654395037
transform 1 0 14560 0 1 7056
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _486_
timestamp 1654395037
transform -1 0 10640 0 1 11760
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1  _487_
timestamp 1654395037
transform 1 0 9856 0 1 10192
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1  _488_
timestamp 1654395037
transform 1 0 4144 0 -1 11760
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _489_
timestamp 1654395037
transform -1 0 4704 0 -1 8624
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _490_
timestamp 1654395037
transform 1 0 896 0 1 10192
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _491_
timestamp 1654395037
transform 1 0 896 0 -1 10192
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _492_
timestamp 1654395037
transform 1 0 14560 0 1 5488
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _493_
timestamp 1654395037
transform 1 0 22848 0 1 7056
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _494_
timestamp 1654395037
transform 1 0 27216 0 -1 8624
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _495_
timestamp 1654395037
transform -1 0 34608 0 1 7056
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _496_
timestamp 1654395037
transform -1 0 34608 0 1 8624
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _497_
timestamp 1654395037
transform -1 0 32480 0 -1 10192
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _498_
timestamp 1654395037
transform 1 0 22960 0 1 8624
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _499_
timestamp 1654395037
transform 1 0 30800 0 1 10192
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _500_
timestamp 1654395037
transform 1 0 30576 0 -1 11760
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _501_
timestamp 1654395037
transform -1 0 30016 0 1 10192
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1654395037
transform -1 0 30352 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1654395037
transform 1 0 31696 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  input3 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 28672 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  input4 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 33488 0 -1 10192
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  input5 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 2352 0 1 11760
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1654395037
transform -1 0 34608 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1654395037
transform -1 0 33936 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1654395037
transform -1 0 33040 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1654395037
transform 1 0 29904 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1654395037
transform -1 0 34608 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1654395037
transform -1 0 34608 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output12
timestamp 1654395037
transform 1 0 11872 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output13 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 24416 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output14
timestamp 1654395037
transform 1 0 13888 0 1 10192
box -86 -86 758 870
<< labels >>
flabel metal4 s 4788 724 5108 12604 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 13340 724 13660 12604 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 21892 724 22212 12604 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 30444 724 30764 12604 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 612 2178 34892 2498 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 612 5286 34892 5606 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 612 8394 34892 8714 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 612 11502 34892 11822 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 9064 724 9384 12604 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 17616 724 17936 12604 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 26168 724 26488 12604 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 612 3732 34892 4052 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 612 6840 34892 7160 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 612 9948 34892 10268 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal2 s 12824 13200 12936 14000 0 FreeSans 448 90 0 0 core_clk
port 2 nsew signal tristate
flabel metal2 s 7672 13200 7784 14000 0 FreeSans 448 90 0 0 ext_clk
port 3 nsew signal input
flabel metal3 s 35200 840 36000 952 0 FreeSans 448 0 0 0 ext_clk_sel
port 4 nsew signal input
flabel metal3 s 35200 13048 36000 13160 0 FreeSans 448 0 0 0 ext_reset
port 5 nsew signal input
flabel metal2 s 28280 13200 28392 14000 0 FreeSans 448 90 0 0 pll_clk
port 6 nsew signal input
flabel metal2 s 33432 13200 33544 14000 0 FreeSans 448 90 0 0 pll_clk90
port 7 nsew signal input
flabel metal2 s 2520 13200 2632 14000 0 FreeSans 448 90 0 0 resetb
port 8 nsew signal input
flabel metal2 s 23128 13200 23240 14000 0 FreeSans 448 90 0 0 resetb_sync
port 9 nsew signal tristate
flabel metal3 s 35200 7784 36000 7896 0 FreeSans 448 0 0 0 sel2[0]
port 10 nsew signal input
flabel metal3 s 35200 9576 36000 9688 0 FreeSans 448 0 0 0 sel2[1]
port 11 nsew signal input
flabel metal3 s 35200 11256 36000 11368 0 FreeSans 448 0 0 0 sel2[2]
port 12 nsew signal input
flabel metal3 s 35200 2520 36000 2632 0 FreeSans 448 0 0 0 sel[0]
port 13 nsew signal input
flabel metal3 s 35200 4312 36000 4424 0 FreeSans 448 0 0 0 sel[1]
port 14 nsew signal input
flabel metal3 s 35200 5992 36000 6104 0 FreeSans 448 0 0 0 sel[2]
port 15 nsew signal input
flabel metal2 s 17976 13200 18088 14000 0 FreeSans 448 90 0 0 user_clk
port 16 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 36000 14000
<< end >>
