magic
tech gf180mcuC
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 540 216 756
rect 0 324 216 432
rect 108 108 216 324
rect 0 0 216 108
<< properties >>
string FIXED_BBOX 0 -216 324 756
<< end >>
