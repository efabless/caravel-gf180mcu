* NGSPICE file created from mgmt_protect.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__bufz_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__bufz_8 EN I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

.subckt mgmt_protect VDD VSS caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0]
+ la_data_in_core[10] la_data_in_core[11] la_data_in_core[12] la_data_in_core[13]
+ la_data_in_core[14] la_data_in_core[15] la_data_in_core[16] la_data_in_core[17]
+ la_data_in_core[18] la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21]
+ la_data_in_core[22] la_data_in_core[23] la_data_in_core[24] la_data_in_core[25]
+ la_data_in_core[26] la_data_in_core[27] la_data_in_core[28] la_data_in_core[29]
+ la_data_in_core[2] la_data_in_core[30] la_data_in_core[31] la_data_in_core[32] la_data_in_core[33]
+ la_data_in_core[34] la_data_in_core[35] la_data_in_core[36] la_data_in_core[37]
+ la_data_in_core[38] la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41]
+ la_data_in_core[42] la_data_in_core[43] la_data_in_core[44] la_data_in_core[45]
+ la_data_in_core[46] la_data_in_core[47] la_data_in_core[48] la_data_in_core[49]
+ la_data_in_core[4] la_data_in_core[50] la_data_in_core[51] la_data_in_core[52] la_data_in_core[53]
+ la_data_in_core[54] la_data_in_core[55] la_data_in_core[56] la_data_in_core[57]
+ la_data_in_core[58] la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61]
+ la_data_in_core[62] la_data_in_core[63] la_data_in_core[6] la_data_in_core[7] la_data_in_core[8]
+ la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[10] la_data_in_mprj[11] la_data_in_mprj[12]
+ la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15] la_data_in_mprj[16]
+ la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19] la_data_in_mprj[1] la_data_in_mprj[20]
+ la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23] la_data_in_mprj[24]
+ la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27] la_data_in_mprj[28]
+ la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31] la_data_in_mprj[32]
+ la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35] la_data_in_mprj[36]
+ la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39] la_data_in_mprj[3] la_data_in_mprj[40]
+ la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43] la_data_in_mprj[44]
+ la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47] la_data_in_mprj[48]
+ la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51] la_data_in_mprj[52]
+ la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55] la_data_in_mprj[56]
+ la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59] la_data_in_mprj[5] la_data_in_mprj[60]
+ la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63] la_data_in_mprj[6] la_data_in_mprj[7]
+ la_data_in_mprj[8] la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[10] la_data_out_core[11]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[6] la_data_out_core[7] la_data_out_core[8]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[10] la_data_out_mprj[11]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[6] la_data_out_mprj[7] la_data_out_mprj[8]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[10] la_iena_mprj[11] la_iena_mprj[12]
+ la_iena_mprj[13] la_iena_mprj[14] la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17]
+ la_iena_mprj[18] la_iena_mprj[19] la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21]
+ la_iena_mprj[22] la_iena_mprj[23] la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26]
+ la_iena_mprj[27] la_iena_mprj[28] la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30]
+ la_iena_mprj[31] la_iena_mprj[32] la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35]
+ la_iena_mprj[36] la_iena_mprj[37] la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3]
+ la_iena_mprj[40] la_iena_mprj[41] la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44]
+ la_iena_mprj[45] la_iena_mprj[46] la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49]
+ la_iena_mprj[4] la_iena_mprj[50] la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53]
+ la_iena_mprj[54] la_iena_mprj[55] la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58]
+ la_iena_mprj[59] la_iena_mprj[5] la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62]
+ la_iena_mprj[63] la_iena_mprj[6] la_iena_mprj[7] la_iena_mprj[8] la_iena_mprj[9]
+ la_oenb_core[0] la_oenb_core[10] la_oenb_core[11] la_oenb_core[12] la_oenb_core[13]
+ la_oenb_core[14] la_oenb_core[15] la_oenb_core[16] la_oenb_core[17] la_oenb_core[18]
+ la_oenb_core[19] la_oenb_core[1] la_oenb_core[20] la_oenb_core[21] la_oenb_core[22]
+ la_oenb_core[23] la_oenb_core[24] la_oenb_core[25] la_oenb_core[26] la_oenb_core[27]
+ la_oenb_core[28] la_oenb_core[29] la_oenb_core[2] la_oenb_core[30] la_oenb_core[31]
+ la_oenb_core[32] la_oenb_core[33] la_oenb_core[34] la_oenb_core[35] la_oenb_core[36]
+ la_oenb_core[37] la_oenb_core[38] la_oenb_core[39] la_oenb_core[3] la_oenb_core[40]
+ la_oenb_core[41] la_oenb_core[42] la_oenb_core[43] la_oenb_core[44] la_oenb_core[45]
+ la_oenb_core[46] la_oenb_core[47] la_oenb_core[48] la_oenb_core[49] la_oenb_core[4]
+ la_oenb_core[50] la_oenb_core[51] la_oenb_core[52] la_oenb_core[53] la_oenb_core[54]
+ la_oenb_core[55] la_oenb_core[56] la_oenb_core[57] la_oenb_core[58] la_oenb_core[59]
+ la_oenb_core[5] la_oenb_core[60] la_oenb_core[61] la_oenb_core[62] la_oenb_core[63]
+ la_oenb_core[6] la_oenb_core[7] la_oenb_core[8] la_oenb_core[9] la_oenb_mprj[0]
+ la_oenb_mprj[10] la_oenb_mprj[11] la_oenb_mprj[12] la_oenb_mprj[13] la_oenb_mprj[14]
+ la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18] la_oenb_mprj[19]
+ la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22] la_oenb_mprj[23]
+ la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27] la_oenb_mprj[28]
+ la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31] la_oenb_mprj[32]
+ la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36] la_oenb_mprj[37]
+ la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40] la_oenb_mprj[41]
+ la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45] la_oenb_mprj[46]
+ la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4] la_oenb_mprj[50]
+ la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54] la_oenb_mprj[55]
+ la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59] la_oenb_mprj[5]
+ la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63] la_oenb_mprj[6]
+ la_oenb_mprj[7] la_oenb_mprj[8] la_oenb_mprj[9] mprj_ack_i_core mprj_ack_i_user
+ mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11] mprj_adr_o_core[12] mprj_adr_o_core[13]
+ mprj_adr_o_core[14] mprj_adr_o_core[15] mprj_adr_o_core[16] mprj_adr_o_core[17]
+ mprj_adr_o_core[18] mprj_adr_o_core[19] mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21]
+ mprj_adr_o_core[22] mprj_adr_o_core[23] mprj_adr_o_core[24] mprj_adr_o_core[25]
+ mprj_adr_o_core[26] mprj_adr_o_core[27] mprj_adr_o_core[28] mprj_adr_o_core[29]
+ mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31] mprj_adr_o_core[3] mprj_adr_o_core[4]
+ mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7] mprj_adr_o_core[8] mprj_adr_o_core[9]
+ mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11] mprj_adr_o_user[12] mprj_adr_o_user[13]
+ mprj_adr_o_user[14] mprj_adr_o_user[15] mprj_adr_o_user[16] mprj_adr_o_user[17]
+ mprj_adr_o_user[18] mprj_adr_o_user[19] mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21]
+ mprj_adr_o_user[22] mprj_adr_o_user[23] mprj_adr_o_user[24] mprj_adr_o_user[25]
+ mprj_adr_o_user[26] mprj_adr_o_user[27] mprj_adr_o_user[28] mprj_adr_o_user[29]
+ mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31] mprj_adr_o_user[3] mprj_adr_o_user[4]
+ mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7] mprj_adr_o_user[8] mprj_adr_o_user[9]
+ mprj_cyc_o_core mprj_cyc_o_user mprj_dat_i_core[0] mprj_dat_i_core[10] mprj_dat_i_core[11]
+ mprj_dat_i_core[12] mprj_dat_i_core[13] mprj_dat_i_core[14] mprj_dat_i_core[15]
+ mprj_dat_i_core[16] mprj_dat_i_core[17] mprj_dat_i_core[18] mprj_dat_i_core[19]
+ mprj_dat_i_core[1] mprj_dat_i_core[20] mprj_dat_i_core[21] mprj_dat_i_core[22] mprj_dat_i_core[23]
+ mprj_dat_i_core[24] mprj_dat_i_core[25] mprj_dat_i_core[26] mprj_dat_i_core[27]
+ mprj_dat_i_core[28] mprj_dat_i_core[29] mprj_dat_i_core[2] mprj_dat_i_core[30] mprj_dat_i_core[31]
+ mprj_dat_i_core[3] mprj_dat_i_core[4] mprj_dat_i_core[5] mprj_dat_i_core[6] mprj_dat_i_core[7]
+ mprj_dat_i_core[8] mprj_dat_i_core[9] mprj_dat_i_user[0] mprj_dat_i_user[10] mprj_dat_i_user[11]
+ mprj_dat_i_user[12] mprj_dat_i_user[13] mprj_dat_i_user[14] mprj_dat_i_user[15]
+ mprj_dat_i_user[16] mprj_dat_i_user[17] mprj_dat_i_user[18] mprj_dat_i_user[19]
+ mprj_dat_i_user[1] mprj_dat_i_user[20] mprj_dat_i_user[21] mprj_dat_i_user[22] mprj_dat_i_user[23]
+ mprj_dat_i_user[24] mprj_dat_i_user[25] mprj_dat_i_user[26] mprj_dat_i_user[27]
+ mprj_dat_i_user[28] mprj_dat_i_user[29] mprj_dat_i_user[2] mprj_dat_i_user[30] mprj_dat_i_user[31]
+ mprj_dat_i_user[3] mprj_dat_i_user[4] mprj_dat_i_user[5] mprj_dat_i_user[6] mprj_dat_i_user[7]
+ mprj_dat_i_user[8] mprj_dat_i_user[9] mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11]
+ mprj_dat_o_core[12] mprj_dat_o_core[13] mprj_dat_o_core[14] mprj_dat_o_core[15]
+ mprj_dat_o_core[16] mprj_dat_o_core[17] mprj_dat_o_core[18] mprj_dat_o_core[19]
+ mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21] mprj_dat_o_core[22] mprj_dat_o_core[23]
+ mprj_dat_o_core[24] mprj_dat_o_core[25] mprj_dat_o_core[26] mprj_dat_o_core[27]
+ mprj_dat_o_core[28] mprj_dat_o_core[29] mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31]
+ mprj_dat_o_core[3] mprj_dat_o_core[4] mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7]
+ mprj_dat_o_core[8] mprj_dat_o_core[9] mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11]
+ mprj_dat_o_user[12] mprj_dat_o_user[13] mprj_dat_o_user[14] mprj_dat_o_user[15]
+ mprj_dat_o_user[16] mprj_dat_o_user[17] mprj_dat_o_user[18] mprj_dat_o_user[19]
+ mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21] mprj_dat_o_user[22] mprj_dat_o_user[23]
+ mprj_dat_o_user[24] mprj_dat_o_user[25] mprj_dat_o_user[26] mprj_dat_o_user[27]
+ mprj_dat_o_user[28] mprj_dat_o_user[29] mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31]
+ mprj_dat_o_user[3] mprj_dat_o_user[4] mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7]
+ mprj_dat_o_user[8] mprj_dat_o_user[9] mprj_iena_wb mprj_sel_o_core[0] mprj_sel_o_core[1]
+ mprj_sel_o_core[2] mprj_sel_o_core[3] mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2]
+ mprj_sel_o_user[3] mprj_stb_o_core mprj_stb_o_user mprj_we_o_core mprj_we_o_user
+ user_clock user_clock2 user_irq[0] user_irq[1] user_irq[2] user_irq_core[0] user_irq_core[1]
+ user_irq_core[2] user_irq_ena[0] user_irq_ena[1] user_irq_ena[2] user_reset
XTAP_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__164__I mprj_dat_o_core[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_gates\[8\] mprj_dat_i_user[8] mprj_iena_wb user_wb_dat_gates\[8\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_5_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xla_buf\[36\] _011_/ZN la_data_out_mprj[36] la_data_in_core[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_6_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__074__I la_oenb_mprj[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[25\] la_data_out_core[25] la_iena_mprj[25] user_to_mprj_in_gates\[25\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_user_wb_dat_gates\[16\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__159__I mprj_adr_o_core[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__069__I la_oenb_mprj[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[17\]_A2 la_iena_mprj[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_200_ caravel_clk2 user_clock2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_user_to_mprj_in_gates\[1\]_A2 la_iena_mprj[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_062_ la_oenb_mprj[23] _062_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_131_ mprj_adr_o_core[3] mprj_adr_o_user[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[7\]_A1 mprj_dat_i_user[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[29\]_A1 mprj_dat_i_user[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_045_ la_oenb_mprj[6] _045_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__172__I mprj_dat_o_core[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_114_ la_oenb_mprj[50] la_oenb_core[50] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[62\] user_to_mprj_in_gates\[62\]/ZN la_data_in_mprj[62]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
Xuser_wb_dat_gates\[20\] mprj_dat_i_user[20] mprj_iena_wb user_wb_dat_gates\[20\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__082__I la_oenb_mprj[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[50\]_I user_to_mprj_in_gates\[50\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_buffers\[41\]_I user_to_mprj_in_gates\[41\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[30\]_EN _005_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__167__I mprj_dat_o_core[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_028_ la_oenb_mprj[53] _028_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_4_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[32\]_I user_to_mprj_in_gates\[32\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[55\] la_data_out_core[55] la_iena_mprj[55] user_to_mprj_in_gates\[55\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__077__I la_oenb_mprj[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_buffers\[23\]_I user_to_mprj_in_gates\[23\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[63\]_I la_data_out_mprj[63] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_to_mprj_in_buffers\[14\]_I user_to_mprj_in_gates\[14\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_buffers\[25\] user_to_mprj_in_gates\[25\]/ZN la_data_in_mprj[25]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_la_buf\[54\]_I la_data_out_mprj[54] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[50\]_A2 la_iena_mprj[50] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_la_buf\[45\]_I la_data_out_mprj[45] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[36\]_I la_data_out_mprj[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xla_buf\[29\] _004_/ZN la_data_out_mprj[29] la_data_in_core[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XANTENNA__180__I mprj_dat_o_core[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_la_buf\[27\]_I la_data_out_mprj[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[18\] la_data_out_core[18] la_iena_mprj[18] user_to_mprj_in_gates\[18\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__090__I la_oenb_mprj[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_buffers\[28\] user_wb_dat_gates\[28\]/ZN mprj_dat_i_core[28] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_la_buf\[18\]_I la_data_out_mprj[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[40\]_A1 la_data_out_core[40] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__175__I mprj_dat_o_core[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__085__I la_oenb_mprj[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_wb_dat_buffers\[2\] user_wb_dat_gates\[2\]/ZN mprj_dat_i_core[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_0_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[63\]_A1 la_data_out_core[63] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_130_ mprj_adr_o_core[2] mprj_adr_o_user[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_061_ la_oenb_mprj[22] _061_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[7\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_113_ la_oenb_mprj[49] la_oenb_core[49] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_user_wb_dat_gates\[29\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xla_buf\[7\] _046_/ZN la_data_out_mprj[7] la_data_in_core[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_4_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_044_ la_oenb_mprj[5] _044_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
Xla_buf\[11\] _050_/ZN la_data_out_mprj[11] la_data_in_core[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
Xuser_to_mprj_in_buffers\[55\] user_to_mprj_in_gates\[55\]/ZN la_data_in_mprj[55]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_1_1843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_wb_dat_gates\[13\] mprj_dat_i_user[13] mprj_iena_wb user_wb_dat_gates\[13\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_6_1710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_wb_dat_buffers\[10\] user_wb_dat_gates\[10\]/ZN mprj_dat_i_core[10] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_0_1353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xla_buf\[59\] _034_/ZN la_data_out_mprj[59] la_data_in_core[59] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XANTENNA__183__I mprj_dat_o_core[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_027_ la_oenb_mprj[52] _027_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_to_mprj_in_gates\[48\] la_data_out_core[48] la_iena_mprj[48] user_to_mprj_in_gates\[48\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__093__I la_oenb_mprj[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[19\]_A1 mprj_dat_i_user[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__178__I mprj_dat_o_core[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_buffers\[18\] user_to_mprj_in_gates\[18\]/ZN la_data_in_mprj[18]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XTAP_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__088__I la_oenb_mprj[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_wb_ack_gate_A1 mprj_ack_i_user VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[4\]_A1 la_data_out_core[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xla_buf\[41\] _016_/ZN la_data_out_mprj[41] la_data_in_core[41] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XANTENNA_user_to_mprj_in_gates\[40\]_A2 la_iena_mprj[40] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__191__I mprj_dat_o_core[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_to_mprj_in_gates\[30\] la_data_out_core[30] la_iena_mprj[30] user_to_mprj_in_gates\[30\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_user_to_mprj_in_gates\[63\]_A2 la_iena_mprj[63] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_wb_dat_buffers\[8\]_I user_wb_dat_gates\[8\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_060_ la_oenb_mprj[21] _060_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__186__I mprj_dat_o_core[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_189_ mprj_dat_o_core[28] mprj_dat_o_user[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__096__I la_oenb_mprj[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[30\]_A1 la_data_out_core[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_112_ la_oenb_mprj[48] la_oenb_core[48] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_043_ la_oenb_mprj[4] _043_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_user_to_mprj_in_buffers\[9\]_I user_to_mprj_in_gates\[9\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_buffers\[48\] user_to_mprj_in_gates\[48\]/ZN la_data_in_mprj[48]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_user_to_mprj_in_gates\[53\]_A1 la_data_out_core[53] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_irq_buffers\[2\] user_irq_gates\[2\]/ZN user_irq[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_5_1298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_026_ la_oenb_mprj[51] _026_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_4_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[19\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__194__I mprj_sel_o_core[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_009_ la_oenb_mprj[34] _009_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[60\] la_data_out_core[60] la_iena_mprj[60] user_to_mprj_in_gates\[60\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_wb_ack_gate_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[4\]_A2 la_iena_mprj[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__189__I mprj_dat_o_core[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_to_mprj_in_buffers\[30\] user_to_mprj_in_gates\[30\]/ZN la_data_in_mprj[30]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA__099__I la_oenb_mprj[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_irq_gates\[1\]_A1 user_irq_core[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xla_buf\[34\] _009_/ZN la_data_out_mprj[34] la_data_in_core[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
Xuser_wb_dat_gates\[6\] mprj_dat_i_user[6] mprj_iena_wb user_wb_dat_gates\[6\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_6_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[10\]_EN _049_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[23\] la_data_out_core[23] la_iena_mprj[23] user_to_mprj_in_gates\[23\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_3_1341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_188_ mprj_dat_o_core[27] mprj_dat_o_user[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_buffers\[62\]_I user_to_mprj_in_gates\[62\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[1\]_EN _040_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[53\]_I user_to_mprj_in_gates\[53\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[30\]_A2 la_iena_mprj[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_111_ la_oenb_mprj[47] la_oenb_core[47] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_042_ la_oenb_mprj[3] _042_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_user_to_mprj_in_buffers\[44\]_I user_to_mprj_in_gates\[44\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__197__I mprj_stb_o_core VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_user_to_mprj_in_gates\[53\]_A2 la_iena_mprj[53] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[35\]_I user_to_mprj_in_gates\[35\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_buffers\[26\]_I user_to_mprj_in_gates\[26\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_025_ la_oenb_mprj[50] _025_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[17\]_I user_to_mprj_in_gates\[17\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_buffers\[60\] user_to_mprj_in_gates\[60\]/ZN la_data_in_mprj[60]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_1_1653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[57\]_I la_data_out_mprj[57] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[20\]_A1 la_data_out_core[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[48\]_I la_data_out_mprj[48] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_user_to_mprj_in_gates\[43\]_A1 la_data_out_core[43] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[39\]_I la_data_out_mprj[39] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_008_ la_oenb_mprj[33] _008_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_4_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[53\] la_data_out_core[53] la_iena_mprj[53] user_to_mprj_in_gates\[53\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[23\] user_to_mprj_in_gates\[23\]/ZN la_data_in_mprj[23]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_4_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_irq_gates\[1\]_A2 user_irq_ena[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xla_buf\[27\] _002_/ZN la_data_out_mprj[27] la_data_in_core[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_6_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_wb_dat_gates\[29\] mprj_dat_i_user[29] mprj_iena_wb user_wb_dat_gates\[29\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_to_mprj_in_gates\[16\] la_data_out_core[16] la_iena_mprj[16] user_to_mprj_in_gates\[16\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_wb_dat_buffers\[26\] user_wb_dat_gates\[26\]/ZN mprj_dat_i_core[26] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_3_1397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_187_ mprj_dat_o_core[26] mprj_dat_o_user[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_wb_dat_buffers\[0\] user_wb_dat_gates\[0\]/ZN mprj_dat_i_core[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_5_1426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_110_ la_oenb_mprj[46] la_oenb_core[46] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_041_ la_oenb_mprj[2] _041_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_la_buf\[23\]_EN _062_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_wb_dat_buffers\[12\]_I user_wb_dat_gates\[12\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_user_to_mprj_in_gates\[7\]_A1 la_data_out_core[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_024_ la_oenb_mprj[49] _024_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
Xla_buf\[5\] _044_/ZN la_data_out_mprj[5] la_data_in_core[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_3_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__001__I la_oenb_mprj[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[20\]_A2 la_iena_mprj[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_buffers\[53\] user_to_mprj_in_gates\[53\]/ZN la_data_in_mprj[53]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_1_1632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_wb_dat_gates\[11\] mprj_dat_i_user[11] mprj_iena_wb user_wb_dat_gates\[11\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_6_1565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[1\]_I la_data_out_mprj[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xla_buf\[57\] _032_/ZN la_data_out_mprj[57] la_data_in_core[57] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XANTENNA_user_to_mprj_in_gates\[43\]_A2 la_iena_mprj[43] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_007_ la_oenb_mprj[32] _007_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_4_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_to_mprj_in_gates\[46\] la_data_out_core[46] la_iena_mprj[46] user_to_mprj_in_gates\[46\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_3_1727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_to_mprj_in_gates\[8\] la_data_out_core[8] la_iena_mprj[8] user_to_mprj_in_gates\[8\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_6_1373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[10\]_A1 la_data_out_core[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_buffers\[16\] user_to_mprj_in_gates\[16\]/ZN la_data_in_mprj[16]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_4_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_to_mprj_in_gates\[33\]_A1 la_data_out_core[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_buffers\[8\] user_to_mprj_in_gates\[8\]/ZN la_data_in_mprj[8] VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_6_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[56\]_A1 la_data_out_core[56] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_buffers\[19\] user_wb_dat_gates\[19\]/ZN mprj_dat_i_core[19] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_5_1608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_186_ mprj_dat_o_core[25] mprj_dat_o_user[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__004__I la_oenb_mprj[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_040_ la_oenb_mprj[1] _040_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_169_ mprj_dat_o_core[8] mprj_dat_o_user[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_to_mprj_in_gates\[7\]_A2 la_iena_mprj[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_023_ la_oenb_mprj[48] _023_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[46\] user_to_mprj_in_gates\[46\]/ZN la_data_in_mprj[46]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_1_1699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__102__I la_oenb_mprj[38] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_irq_buffers\[0\] user_irq_gates\[0\]/ZN user_irq[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_0_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_006_ la_oenb_mprj[31] _006_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_4_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__012__I la_oenb_mprj[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_la_buf\[13\]_EN _052_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xuser_to_mprj_in_gates\[39\] la_data_out_core[39] la_iena_mprj[39] user_to_mprj_in_gates\[39\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_6_1352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[10\]_A2 la_iena_mprj[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__007__I la_oenb_mprj[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_la_buf\[4\]_EN _043_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[0\]_A1 mprj_dat_i_user[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[33\]_A2 la_iena_mprj[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[22\]_A1 mprj_dat_i_user[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[56\]_A2 la_iena_mprj[56] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__200__I caravel_clk2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_buffers\[56\]_I user_to_mprj_in_gates\[56\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__110__I la_oenb_mprj[46] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_gates\[4\] mprj_dat_i_user[4] mprj_iena_wb user_wb_dat_gates\[4\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_6_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_185_ mprj_dat_o_core[24] mprj_dat_o_user[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xla_buf\[32\] _007_/ZN la_data_out_mprj[32] la_data_in_core[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XANTENNA_user_to_mprj_in_buffers\[47\]_I user_to_mprj_in_gates\[47\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[20\]_I la_data_out_mprj[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__020__I la_oenb_mprj[45] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_to_mprj_in_gates\[21\] la_data_out_core[21] la_iena_mprj[21] user_to_mprj_in_gates\[21\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_user_to_mprj_in_gates\[23\]_A1 la_data_out_core[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_buffers\[31\] user_wb_dat_gates\[31\]/ZN mprj_dat_i_core[31] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_user_to_mprj_in_buffers\[38\]_I user_to_mprj_in_gates\[38\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[11\]_I la_data_out_mprj[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[29\]_I user_to_mprj_in_gates\[29\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__105__I la_oenb_mprj[41] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[46\]_A1 la_data_out_core[46] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__015__I la_oenb_mprj[40] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_168_ mprj_dat_o_core[7] mprj_dat_o_user[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_099_ la_oenb_mprj[35] la_oenb_core[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_022_ la_oenb_mprj[47] _022_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_4_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_to_mprj_in_buffers\[39\] user_to_mprj_in_gates\[39\]/ZN la_data_in_mprj[39]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_1_1689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_005_ la_oenb_mprj[30] _005_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_1364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__113__I la_oenb_mprj[49] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xla_buf\[62\] _037_/ZN la_data_out_mprj[62] la_data_in_core[62] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_2_1751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__023__I la_oenb_mprj[48] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[51\] la_data_out_core[51] la_iena_mprj[51] user_to_mprj_in_gates\[51\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_3_1559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[0\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__108__I la_oenb_mprj[44] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__018__I la_oenb_mprj[43] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_wb_dat_gates\[22\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_buffers\[21\] user_to_mprj_in_gates\[21\]/ZN la_data_in_mprj[21]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_5_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[26\]_EN _001_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_184_ mprj_dat_o_core[23] mprj_dat_o_user[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xla_buf\[25\] _000_/ZN la_data_out_mprj[25] la_data_in_core[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_6_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_buffers\[24\]_I user_wb_dat_gates\[24\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_gates\[27\] mprj_dat_i_user[27] mprj_iena_wb user_wb_dat_gates\[27\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_to_mprj_in_gates\[14\] la_data_out_core[14] la_iena_mprj[14] user_to_mprj_in_gates\[14\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_user_to_mprj_in_gates\[23\]_A2 la_iena_mprj[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_buffers\[24\] user_wb_dat_gates\[24\]/ZN mprj_dat_i_core[24] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_5_1407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_buffers\[15\]_I user_wb_dat_gates\[15\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__121__I la_oenb_mprj[57] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[12\]_A1 mprj_dat_i_user[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[46\]_A2 la_iena_mprj[46] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_098_ la_oenb_mprj[34] la_oenb_core[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_167_ mprj_dat_o_core[6] mprj_dat_o_user[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__031__I la_oenb_mprj[56] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_buffers\[1\]_I user_wb_dat_gates\[1\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[4\]_I la_data_out_mprj[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__116__I la_oenb_mprj[52] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_021_ la_oenb_mprj[46] _021_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_gates\[13\]_A1 la_data_out_core[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__026__I la_oenb_mprj[51] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_gates\[36\]_A1 la_data_out_core[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_user_to_mprj_in_buffers\[2\]_I user_to_mprj_in_gates\[2\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_004_ la_oenb_mprj[29] _004_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
Xla_buf\[3\] _042_/ZN la_data_out_mprj[3] la_data_in_core[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XTAP_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xuser_to_mprj_in_buffers\[51\] user_to_mprj_in_gates\[51\]/ZN la_data_in_mprj[51]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_user_to_mprj_in_gates\[59\]_A1 la_data_out_core[59] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xla_buf\[55\] _030_/ZN la_data_out_mprj[55] la_data_in_core[55] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_2_1763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_to_mprj_in_gates\[44\] la_data_out_core[44] la_iena_mprj[44] user_to_mprj_in_gates\[44\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_wb_dat_buffers\[9\] user_wb_dat_gates\[9\]/ZN mprj_dat_i_core[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_3_1527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_to_mprj_in_gates\[6\] la_data_out_core[6] la_iena_mprj[6] user_to_mprj_in_gates\[6\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_2_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__124__I la_oenb_mprj[60] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[14\] user_to_mprj_in_gates\[14\]/ZN la_data_in_mprj[14]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA__034__I la_oenb_mprj[59] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__119__I la_oenb_mprj[55] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[6\] user_to_mprj_in_gates\[6\]/ZN la_data_in_mprj[6] VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_6_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_183_ mprj_dat_o_core[22] mprj_dat_o_user[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xla_buf\[18\] _057_/ZN la_data_out_mprj[18] la_data_in_core[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_1_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__029__I la_oenb_mprj[54] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_buffers\[17\] user_wb_dat_gates\[17\]/ZN mprj_dat_i_core[17] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_5_1419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_wb_dat_gates\[12\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_097_ la_oenb_mprj[33] la_oenb_core[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_166_ mprj_dat_o_core[5] mprj_dat_o_user[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__132__I mprj_adr_o_core[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_020_ la_oenb_mprj[45] _020_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_user_to_mprj_in_gates\[13\]_A2 la_iena_mprj[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_149_ mprj_adr_o_core[21] mprj_adr_o_user[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__042__I la_oenb_mprj[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[7\]_EN _046_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_wb_dat_gates\[3\]_A1 mprj_dat_i_user[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[36\]_A2 la_iena_mprj[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_003_ la_oenb_mprj[28] _003_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__127__I la_oenb_mprj[63] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[44\] user_to_mprj_in_gates\[44\]/ZN la_data_in_mprj[44]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_user_to_mprj_in_gates\[59\]_A2 la_iena_mprj[59] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__037__I la_oenb_mprj[62] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_user_wb_dat_gates\[25\]_A1 mprj_dat_i_user[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_buffers\[10\]_I user_to_mprj_in_gates\[10\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xla_buf\[48\] _023_/ZN la_data_out_mprj[48] la_data_in_core[48] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_5_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[50\]_I la_data_out_mprj[50] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[26\]_A1 la_data_out_core[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[37\] la_data_out_core[37] la_iena_mprj[37] user_to_mprj_in_gates\[37\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_1_1296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[41\]_I la_data_out_mprj[41] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[59\]_I user_to_mprj_in_gates\[59\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[32\]_I la_data_out_mprj[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__140__I mprj_adr_o_core[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[49\]_A1 la_data_out_core[49] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_la_buf\[23\]_I la_data_out_mprj[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__050__I la_oenb_mprj[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[14\]_I la_data_out_mprj[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_182_ mprj_dat_o_core[21] mprj_dat_o_user[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__135__I mprj_adr_o_core[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__045__I la_oenb_mprj[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_165_ mprj_dat_o_core[4] mprj_dat_o_user[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xuser_wb_dat_gates\[2\] mprj_dat_i_user[2] mprj_iena_wb user_wb_dat_gates\[2\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xla_buf\[30\] _005_/ZN la_data_out_mprj[30] la_data_in_core[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
X_096_ la_oenb_mprj[32] la_oenb_core[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_1475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_148_ mprj_adr_o_core[20] mprj_adr_o_user[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_079_ la_oenb_mprj[15] la_oenb_core[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_user_wb_dat_gates\[3\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_002_ la_oenb_mprj[27] _002_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_4_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__143__I mprj_adr_o_core[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_wb_dat_gates\[25\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_buffers\[37\] user_to_mprj_in_gates\[37\]/ZN la_data_in_mprj[37]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_1_1489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__053__I la_oenb_mprj[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[29\]_EN _004_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_1710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__138__I mprj_adr_o_core[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__048__I la_oenb_mprj[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[26\]_A2 la_iena_mprj[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[49\]_A2 la_iena_mprj[49] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_wb_dat_gates\[15\]_A1 mprj_dat_i_user[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xla_buf\[60\] _035_/ZN la_data_out_mprj[60] la_data_in_core[60] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_5_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_181_ mprj_dat_o_core[20] mprj_dat_o_user[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_irq_gates\[1\] user_irq_core[1] user_irq_ena[1] user_irq_gates\[1\]/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_user_to_mprj_in_gates\[16\]_A1 la_data_out_core[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__151__I mprj_adr_o_core[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[0\]_A1 la_data_out_core[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__061__I la_oenb_mprj[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_buffers\[4\]_I user_wb_dat_gates\[4\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[39\]_A1 la_data_out_core[39] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[7\]_I la_data_out_mprj[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_164_ mprj_dat_o_core[3] mprj_dat_o_user[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_095_ la_oenb_mprj[31] la_oenb_core[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__146__I mprj_adr_o_core[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xla_buf\[23\] _062_/ZN la_data_out_mprj[23] la_data_in_core[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_2_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_wb_dat_gates\[25\] mprj_dat_i_user[25] mprj_iena_wb user_wb_dat_gates\[25\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__056__I la_oenb_mprj[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[12\] la_data_out_core[12] la_iena_mprj[12] user_to_mprj_in_gates\[12\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_wb_dat_buffers\[22\] user_wb_dat_gates\[22\]/ZN mprj_dat_i_core[22] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_0_1852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[5\]_I user_to_mprj_in_gates\[5\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_078_ la_oenb_mprj[14] la_oenb_core[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_147_ mprj_adr_o_core[19] mprj_adr_o_user[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_001_ la_oenb_mprj[26] _001_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_4_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__154__I mprj_adr_o_core[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xla_buf\[1\] _040_/ZN la_data_out_mprj[1] la_data_in_core[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_5_1390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__064__I la_oenb_mprj[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_wb_dat_gates\[15\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xla_buf\[53\] _028_/ZN la_data_out_mprj[53] la_data_in_core[53] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XANTENNA__149__I mprj_adr_o_core[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__059__I la_oenb_mprj[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[42\] la_data_out_core[42] la_iena_mprj[42] user_to_mprj_in_gates\[42\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_wb_dat_buffers\[7\] user_wb_dat_gates\[7\]/ZN mprj_dat_i_core[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XTAP_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[4\] la_data_out_core[4] la_iena_mprj[4] user_to_mprj_in_gates\[4\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_3_1872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_180_ mprj_dat_o_core[19] mprj_dat_o_user[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_user_to_mprj_in_gates\[16\]_A2 la_iena_mprj[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[0\]_A2 la_iena_mprj[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[12\] user_to_mprj_in_gates\[12\]/ZN la_data_in_mprj[12]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_user_wb_dat_gates\[6\]_A1 mprj_dat_i_user[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[39\]_A2 la_iena_mprj[39] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_to_mprj_in_buffers\[4\] user_to_mprj_in_gates\[4\]/ZN la_data_in_mprj[4] VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
X_094_ la_oenb_mprj[30] la_oenb_core[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_163_ mprj_dat_o_core[2] mprj_dat_o_user[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__162__I mprj_dat_o_core[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xla_buf\[16\] _055_/ZN la_data_out_mprj[16] la_data_in_core[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_2_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[28\]_A1 mprj_dat_i_user[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_gates\[18\] mprj_dat_i_user[18] mprj_iena_wb user_wb_dat_gates\[18\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__072__I la_oenb_mprj[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_buffers\[15\] user_wb_dat_gates\[15\]/ZN mprj_dat_i_core[15] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_0_1875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_buffers\[40\]_I user_to_mprj_in_gates\[40\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__157__I mprj_adr_o_core[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_077_ la_oenb_mprj[13] la_oenb_core[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_146_ mprj_adr_o_core[18] mprj_adr_o_user[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_buffers\[31\]_I user_to_mprj_in_gates\[31\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[29\]_A1 la_data_out_core[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__067__I la_oenb_mprj[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[22\]_I user_to_mprj_in_gates\[22\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_la_buf\[62\]_I la_data_out_mprj[62] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_000_ la_oenb_mprj[25] _000_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_4_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[13\]_I user_to_mprj_in_gates\[13\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_la_buf\[53\]_I la_data_out_mprj[53] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_129_ mprj_adr_o_core[1] mprj_adr_o_user[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_la_buf\[44\]_I la_data_out_mprj[44] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[35\]_I la_data_out_mprj[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__170__I mprj_dat_o_core[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[42\] user_to_mprj_in_gates\[42\]/ZN la_data_in_mprj[42]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_1_1277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_la_buf\[26\]_I la_data_out_mprj[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__080__I la_oenb_mprj[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[17\]_I la_data_out_mprj[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__165__I mprj_dat_o_core[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xla_buf\[46\] _021_/ZN la_data_out_mprj[46] la_data_in_core[46] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_5_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[35\] la_data_out_core[35] la_iena_mprj[35] user_to_mprj_in_gates\[35\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__075__I la_oenb_mprj[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[62\]_A1 la_data_out_core[62] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[6\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_162_ mprj_dat_o_core[1] mprj_dat_o_user[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_093_ la_oenb_mprj[29] la_oenb_core[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[28\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_145_ mprj_adr_o_core[17] mprj_adr_o_user[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__173__I mprj_dat_o_core[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_gates\[0\] mprj_dat_i_user[0] mprj_iena_wb user_wb_dat_gates\[0\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_076_ la_oenb_mprj[12] la_oenb_core[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[29\]_A2 la_iena_mprj[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_gates\[30\] mprj_dat_i_user[30] mprj_iena_wb user_wb_dat_gates\[30\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__083__I la_oenb_mprj[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[18\]_A1 mprj_dat_i_user[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__168__I mprj_dat_o_core[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_128_ mprj_adr_o_core[0] mprj_adr_o_user[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_059_ la_oenb_mprj[20] _059_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_1348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__078__I la_oenb_mprj[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[19\]_A1 la_data_out_core[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[3\]_A1 la_data_out_core[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_buffers\[35\] user_to_mprj_in_gates\[35\]/ZN la_data_in_mprj[35]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_2_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xla_buf\[39\] _014_/ZN la_data_out_mprj[39] la_data_in_core[39] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_5_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__181__I mprj_dat_o_core[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_to_mprj_in_gates\[28\] la_data_out_core[28] la_iena_mprj[28] user_to_mprj_in_gates\[28\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_3_1329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__091__I la_oenb_mprj[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_buffers\[7\]_I user_wb_dat_gates\[7\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[62\]_A2 la_iena_mprj[62] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__176__I mprj_dat_o_core[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__086__I la_oenb_mprj[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_161_ mprj_dat_o_core[0] mprj_dat_o_user[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_092_ la_oenb_mprj[28] la_oenb_core[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[8\]_I user_to_mprj_in_gates\[8\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_user_to_mprj_in_gates\[52\]_A1 la_data_out_core[52] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_075_ la_oenb_mprj[11] la_oenb_core[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_144_ mprj_adr_o_core[16] mprj_adr_o_user[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xla_buf\[21\] _060_/ZN la_data_out_mprj[21] la_data_in_core[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_3_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_wb_dat_gates\[23\] mprj_dat_i_user[23] mprj_iena_wb user_wb_dat_gates\[23\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_to_mprj_in_gates\[10\] la_data_out_core[10] la_iena_mprj[10] user_to_mprj_in_gates\[10\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_wb_dat_buffers\[20\] user_wb_dat_gates\[20\]/ZN mprj_dat_i_core[20] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_0_1630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_wb_dat_gates\[18\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__184__I mprj_dat_o_core[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_127_ la_oenb_mprj[63] la_oenb_core[63] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_058_ la_oenb_mprj[19] _058_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_1338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_to_mprj_in_gates\[58\] la_data_out_core[58] la_iena_mprj[58] user_to_mprj_in_gates\[58\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__094__I la_oenb_mprj[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_to_mprj_in_gates\[19\]_A2 la_iena_mprj[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__179__I mprj_dat_o_core[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[3\]_A2 la_iena_mprj[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_buffers\[28\] user_to_mprj_in_gates\[28\]/ZN la_data_in_mprj[28]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_6_1157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__089__I la_oenb_mprj[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_wb_dat_gates\[9\]_A1 mprj_dat_i_user[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_irq_gates\[0\]_A1 user_irq_core[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xla_buf\[51\] _026_/ZN la_data_out_mprj[51] la_data_in_core[51] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XANTENNA__192__I mprj_dat_o_core[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xuser_to_mprj_in_gates\[40\] la_data_out_core[40] la_iena_mprj[40] user_to_mprj_in_gates\[40\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_user_to_mprj_in_buffers\[61\]_I user_to_mprj_in_gates\[61\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_wb_dat_buffers\[5\] user_wb_dat_gates\[5\]/ZN mprj_dat_i_core[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
Xuser_to_mprj_in_gates\[2\] la_data_out_core[2] la_iena_mprj[2] user_to_mprj_in_gates\[2\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_5_1937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[52\]_I user_to_mprj_in_gates\[52\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[0\]_EN _039_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_091_ la_oenb_mprj[27] la_oenb_core[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_160_ mprj_cyc_o_core mprj_cyc_o_user VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__187__I mprj_dat_o_core[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_buffers\[43\]_I user_to_mprj_in_gates\[43\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xuser_to_mprj_in_buffers\[10\] user_to_mprj_in_gates\[10\]/ZN la_data_in_mprj[10]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_user_to_mprj_in_buffers\[34\]_I user_to_mprj_in_gates\[34\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__097__I la_oenb_mprj[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_gates\[52\]_A2 la_iena_mprj[52] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_to_mprj_in_buffers\[25\]_I user_to_mprj_in_gates\[25\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_buffers\[2\] user_to_mprj_in_gates\[2\]/ZN la_data_in_mprj[2] VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
X_074_ la_oenb_mprj[10] la_oenb_core[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_143_ mprj_adr_o_core[15] mprj_adr_o_user[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xla_buf\[14\] _053_/ZN la_data_out_mprj[14] la_data_in_core[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XANTENNA_user_to_mprj_in_buffers\[16\]_I user_to_mprj_in_gates\[16\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_to_mprj_in_buffers\[58\] user_to_mprj_in_gates\[58\]/ZN la_data_in_mprj[58]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
Xuser_wb_dat_gates\[16\] mprj_dat_i_user[16] mprj_iena_wb user_wb_dat_gates\[16\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_la_buf\[56\]_I la_data_out_mprj[56] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_buffers\[13\] user_wb_dat_gates\[13\]/ZN mprj_dat_i_core[13] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_2_1929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[47\]_I la_data_out_mprj[47] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_la_buf\[38\]_I la_data_out_mprj[38] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_126_ la_oenb_mprj[62] la_oenb_core[62] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_057_ la_oenb_mprj[18] _057_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_gates\[42\]_A1 la_data_out_core[42] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[29\]_I la_data_out_mprj[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__195__I mprj_sel_o_core[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_109_ la_oenb_mprj[45] la_oenb_core[45] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_user_wb_dat_gates\[9\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_irq_gates\[0\]_A2 user_irq_ena[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_buffers\[40\] user_to_mprj_in_gates\[40\]/ZN la_data_in_mprj[40]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_1_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xla_buf\[44\] _019_/ZN la_data_out_mprj[44] la_data_in_core[44] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_2_1386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[33\] la_data_out_core[33] la_iena_mprj[33] user_to_mprj_in_gates\[33\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_3_1117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_090_ la_oenb_mprj[26] la_oenb_core[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_buffers\[11\]_I user_wb_dat_gates\[11\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_142_ mprj_adr_o_core[14] mprj_adr_o_user[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_la_buf\[22\]_EN _061_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_073_ la_oenb_mprj[9] la_oenb_core[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_gates\[6\]_A1 la_data_out_core[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__198__I mprj_we_o_core VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xuser_wb_ack_buffer user_wb_ack_gate/ZN mprj_ack_i_core VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_la_buf\[0\]_I la_data_out_mprj[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_125_ la_oenb_mprj[61] la_oenb_core[61] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_056_ la_oenb_mprj[17] _056_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_1329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_to_mprj_in_gates\[42\]_A2 la_iena_mprj[42] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_wb_dat_gates\[31\]_A1 mprj_dat_i_user[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_108_ la_oenb_mprj[44] la_oenb_core[44] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_039_ la_oenb_mprj[0] _039_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
Xuser_to_mprj_in_gates\[63\] la_data_out_core[63] la_iena_mprj[63] user_to_mprj_in_gates\[63\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_6_1671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[32\]_A1 la_data_out_core[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xuser_to_mprj_in_buffers\[33\] user_to_mprj_in_gates\[33\]/ZN la_data_in_mprj[33]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XTAP_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[55\]_A1 la_data_out_core[55] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xla_buf\[37\] _012_/ZN la_data_out_mprj[37] la_data_in_core[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_6_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_wb_dat_gates\[9\] mprj_dat_i_user[9] mprj_iena_wb user_wb_dat_gates\[9\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_1_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[26\] la_data_out_core[26] la_iena_mprj[26] user_to_mprj_in_gates\[26\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_3_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_141_ mprj_adr_o_core[13] mprj_adr_o_user[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_072_ la_oenb_mprj[8] la_oenb_core[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[6\]_A2 la_iena_mprj[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_124_ la_oenb_mprj[60] la_oenb_core[60] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_055_ la_oenb_mprj[16] _055_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_1319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__002__I la_oenb_mprj[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xuser_to_mprj_in_buffers\[63\] user_to_mprj_in_gates\[63\]/ZN la_data_in_mprj[63]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
Xuser_wb_dat_gates\[21\] mprj_dat_i_user[21] mprj_iena_wb user_wb_dat_gates\[21\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_6_1853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[12\]_EN _051_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_wb_dat_gates\[31\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_107_ la_oenb_mprj[43] la_oenb_core[43] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_038_ la_oenb_mprj[63] _038_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[56\] la_data_out_core[56] la_iena_mprj[56] user_to_mprj_in_gates\[56\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_2_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_la_buf\[3\]_EN _042_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_to_mprj_in_gates\[32\]_A2 la_iena_mprj[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[26\] user_to_mprj_in_gates\[26\]/ZN la_data_in_mprj[26]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XTAP_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[21\]_A1 mprj_dat_i_user[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[55\]_A2 la_iena_mprj[55] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_buffers\[55\]_I user_to_mprj_in_gates\[55\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__100__I la_oenb_mprj[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_to_mprj_in_buffers\[46\]_I user_to_mprj_in_gates\[46\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__010__I la_oenb_mprj[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[19\] la_data_out_core[19] la_iena_mprj[19] user_to_mprj_in_gates\[19\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_user_to_mprj_in_buffers\[37\]_I user_to_mprj_in_gates\[37\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_buffers\[29\] user_wb_dat_gates\[29\]/ZN mprj_dat_i_core[29] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_la_buf\[10\]_I la_data_out_mprj[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_gates\[22\]_A1 la_data_out_core[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_buffers\[28\]_I user_to_mprj_in_gates\[28\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__005__I la_oenb_mprj[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_buffers\[19\]_I user_to_mprj_in_gates\[19\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[45\]_A1 la_data_out_core[45] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[59\]_I la_data_out_mprj[59] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_wb_dat_buffers\[3\] user_wb_dat_gates\[3\]/ZN mprj_dat_i_core[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
Xuser_to_mprj_in_gates\[0\] la_data_out_core[0] la_iena_mprj[0] user_to_mprj_in_gates\[0\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_071_ la_oenb_mprj[7] la_oenb_core[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_140_ mprj_adr_o_core[12] mprj_adr_o_user[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xuser_to_mprj_in_buffers\[0\] user_to_mprj_in_gates\[0\]/ZN la_data_in_mprj[0] VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
X_123_ la_oenb_mprj[59] la_oenb_core[59] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xla_buf\[12\] _051_/ZN la_data_out_mprj[12] la_data_in_core[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
X_054_ la_oenb_mprj[15] _054_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
Xla_buf\[8\] _047_/ZN la_data_out_mprj[8] la_data_in_core[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_3_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_to_mprj_in_buffers\[56\] user_to_mprj_in_gates\[56\]/ZN la_data_in_mprj[56]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_1_1910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_wb_dat_gates\[14\] mprj_dat_i_user[14] mprj_iena_wb user_wb_dat_gates\[14\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_wb_dat_buffers\[11\] user_wb_dat_gates\[11\]/ZN mprj_dat_i_core[11] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_6_1898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__103__I la_oenb_mprj[39] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_106_ la_oenb_mprj[42] la_oenb_core[42] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_037_ la_oenb_mprj[62] _037_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__013__I la_oenb_mprj[38] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[49\] la_data_out_core[49] la_iena_mprj[49] user_to_mprj_in_gates\[49\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_1_1762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__008__I la_oenb_mprj[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_buffers\[19\] user_to_mprj_in_gates\[19\]/ZN la_data_in_mprj[19]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XTAP_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[21\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_la_buf\[25\]_EN _000_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[9\]_A1 la_data_out_core[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__201__I caravel_rstn VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_buffers\[14\]_I user_wb_dat_gates\[14\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[22\]_A2 la_iena_mprj[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__111__I la_oenb_mprj[47] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xla_buf\[42\] _017_/ZN la_data_out_mprj[42] la_data_in_core[42] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_6_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__021__I la_oenb_mprj[46] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_user_wb_dat_gates\[11\]_A1 mprj_dat_i_user[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[45\]_A2 la_iena_mprj[45] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[31\] la_data_out_core[31] la_iena_mprj[31] user_to_mprj_in_gates\[31\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_buffers\[0\]_I user_wb_dat_gates\[0\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[3\]_I la_data_out_mprj[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_070_ la_oenb_mprj[6] la_oenb_core[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__106__I la_oenb_mprj[42] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_199_ caravel_clk user_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__016__I la_oenb_mprj[41] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[12\]_A1 la_data_out_core[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_buffers\[1\]_I user_to_mprj_in_gates\[1\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_122_ la_oenb_mprj[58] la_oenb_core[58] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_053_ la_oenb_mprj[14] _053_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_user_to_mprj_in_gates\[35\]_A1 la_data_out_core[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xuser_to_mprj_in_buffers\[49\] user_to_mprj_in_gates\[49\]/ZN la_data_in_mprj[49]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_6_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[58\]_A1 la_data_out_core[58] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_105_ la_oenb_mprj[41] la_oenb_core[41] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_036_ la_oenb_mprj[61] _036_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__114__I la_oenb_mprj[50] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__024__I la_oenb_mprj[49] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_019_ la_oenb_mprj[44] _019_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_4_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[61\] la_data_out_core[61] la_iena_mprj[61] user_to_mprj_in_gates\[61\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__109__I la_oenb_mprj[45] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[9\]_A2 la_iena_mprj[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[31\] user_to_mprj_in_gates\[31\]/ZN la_data_in_mprj[31]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA__019__I la_oenb_mprj[44] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xla_buf\[35\] _010_/ZN la_data_out_mprj[35] la_data_in_core[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
Xuser_wb_dat_gates\[7\] mprj_dat_i_user[7] mprj_iena_wb user_wb_dat_gates\[7\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_5_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[11\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[24\] la_data_out_core[24] la_iena_mprj[24] user_to_mprj_in_gates\[24\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__122__I la_oenb_mprj[58] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_198_ mprj_we_o_core mprj_we_o_user VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__032__I la_oenb_mprj[57] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[12\]_A2 la_iena_mprj[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[6\]_EN _045_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__117__I la_oenb_mprj[53] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_121_ la_oenb_mprj[57] la_oenb_core[57] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_user_wb_dat_gates\[2\]_A1 mprj_dat_i_user[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_052_ la_oenb_mprj[13] _052_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_user_to_mprj_in_gates\[35\]_A2 la_iena_mprj[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__027__I la_oenb_mprj[52] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[58\]_A2 la_iena_mprj[58] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[24\]_A1 mprj_dat_i_user[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_104_ la_oenb_mprj[40] la_oenb_core[40] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_035_ la_oenb_mprj[60] _035_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_1119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[61\] user_to_mprj_in_gates\[61\]/ZN la_data_in_mprj[61]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_1_1720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_la_buf\[40\]_I la_data_out_mprj[40] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_gates\[25\]_A1 la_data_out_core[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[31\]_I la_data_out_mprj[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_buffers\[58\]_I user_to_mprj_in_gates\[58\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__130__I mprj_adr_o_core[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_018_ la_oenb_mprj[43] _018_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_la_buf\[22\]_I la_data_out_mprj[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_buffers\[49\]_I user_to_mprj_in_gates\[49\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__040__I la_oenb_mprj[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_user_to_mprj_in_gates\[48\]_A1 la_data_out_core[48] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[54\] la_data_out_core[54] la_iena_mprj[54] user_to_mprj_in_gates\[54\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_1_1561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_la_buf\[13\]_I la_data_out_mprj[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__125__I la_oenb_mprj[61] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_to_mprj_in_buffers\[24\] user_to_mprj_in_gates\[24\]/ZN la_data_in_mprj[24]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA__035__I la_oenb_mprj[60] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xla_buf\[28\] _003_/ZN la_data_out_mprj[28] la_data_in_core[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_2_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[17\] la_data_out_core[17] la_iena_mprj[17] user_to_mprj_in_gates\[17\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_wb_dat_buffers\[27\] user_wb_dat_gates\[27\]/ZN mprj_dat_i_core[27] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_3_748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_197_ mprj_stb_o_core mprj_stb_o_user VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xuser_wb_dat_buffers\[1\] user_wb_dat_gates\[1\]/ZN mprj_dat_i_core[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_3_1261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_120_ la_oenb_mprj[56] la_oenb_core[56] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_051_ la_oenb_mprj[12] _051_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA_user_wb_dat_gates\[2\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__133__I mprj_adr_o_core[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__043__I la_oenb_mprj[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[24\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__128__I mprj_adr_o_core[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_103_ la_oenb_mprj[39] la_oenb_core[39] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_034_ la_oenb_mprj[59] _034_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
Xla_buf\[10\] _049_/ZN la_data_out_mprj[10] la_data_in_core[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
Xla_buf\[6\] _045_/ZN la_data_out_mprj[6] la_data_in_core[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_3_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[54\] user_to_mprj_in_gates\[54\]/ZN la_data_in_mprj[54]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_1_1732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_wb_dat_gates\[12\] mprj_dat_i_user[12] mprj_iena_wb user_wb_dat_gates\[12\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__038__I la_oenb_mprj[63] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[25\]_A2 la_iena_mprj[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xla_buf\[58\] _033_/ZN la_data_out_mprj[58] la_data_in_core[58] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XTAP_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_017_ la_oenb_mprj[42] _017_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_buffers\[26\]_I user_wb_dat_gates\[26\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_wb_dat_gates\[14\]_A1 mprj_dat_i_user[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[48\]_A2 la_iena_mprj[48] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[47\] la_data_out_core[47] la_iena_mprj[47] user_to_mprj_in_gates\[47\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_to_mprj_in_gates\[9\] la_data_out_core[9] la_iena_mprj[9] user_to_mprj_in_gates\[9\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_2_1304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__141__I mprj_adr_o_core[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[17\] user_to_mprj_in_gates\[17\]/ZN la_data_in_mprj[17]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_user_to_mprj_in_gates\[15\]_A1 la_data_out_core[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__051__I la_oenb_mprj[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_wb_dat_buffers\[3\]_I user_wb_dat_gates\[3\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[6\]_I la_data_out_mprj[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_to_mprj_in_buffers\[9\] user_to_mprj_in_gates\[9\]/ZN la_data_in_mprj[9] VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_user_to_mprj_in_gates\[38\]_A1 la_data_out_core[38] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__136__I mprj_adr_o_core[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__046__I la_oenb_mprj[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[4\]_I user_to_mprj_in_gates\[4\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xla_buf\[40\] _015_/ZN la_data_out_mprj[40] la_data_in_core[40] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
X_196_ mprj_sel_o_core[3] mprj_sel_o_user[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_050_ la_oenb_mprj[11] _050_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_179_ mprj_dat_o_core[18] mprj_dat_o_user[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_1593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_102_ la_oenb_mprj[38] la_oenb_core[38] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__144__I mprj_adr_o_core[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_033_ la_oenb_mprj[58] _033_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_1_1766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[47\] user_to_mprj_in_gates\[47\]/ZN la_data_in_mprj[47]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA__054__I la_oenb_mprj[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_irq_buffers\[1\] user_irq_gates\[1\]/ZN user_irq[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_5_1198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__139__I mprj_adr_o_core[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_016_ la_oenb_mprj[41] _016_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_4_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[14\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__049__I la_oenb_mprj[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[15\]_A2 la_iena_mprj[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[9\]_EN _048_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_wb_dat_gates\[5\]_A1 mprj_dat_i_user[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[38\]_A2 la_iena_mprj[38] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__152__I mprj_adr_o_core[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__062__I la_oenb_mprj[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[27\]_A1 mprj_dat_i_user[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__147__I mprj_adr_o_core[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_gates\[5\] mprj_dat_i_user[5] mprj_iena_wb user_wb_dat_gates\[5\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_195_ mprj_sel_o_core[2] mprj_sel_o_user[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xla_buf\[33\] _008_/ZN la_data_out_mprj[33] la_data_in_core[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_1_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__057__I la_oenb_mprj[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_buffers\[30\]_I user_to_mprj_in_gates\[30\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[22\] la_data_out_core[22] la_iena_mprj[22] user_to_mprj_in_gates\[22\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_user_to_mprj_in_buffers\[21\]_I user_to_mprj_in_gates\[21\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[28\]_A1 la_data_out_core[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[61\]_I la_data_out_mprj[61] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[12\]_I user_to_mprj_in_gates\[12\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_178_ mprj_dat_o_core[17] mprj_dat_o_user[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_la_buf\[52\]_I la_data_out_mprj[52] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_la_buf\[43\]_I la_data_out_mprj[43] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_101_ la_oenb_mprj[37] la_oenb_core[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__160__I mprj_cyc_o_core VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[34\]_I la_data_out_mprj[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_032_ la_oenb_mprj[57] _032_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_5_1892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[25\]_I la_data_out_mprj[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__070__I la_oenb_mprj[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[16\]_I la_data_out_mprj[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_015_ la_oenb_mprj[40] _015_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__155__I mprj_adr_o_core[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__065__I la_oenb_mprj[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xla_buf\[63\] _038_/ZN la_data_out_mprj[63] la_data_in_core[63] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
Xuser_wb_ack_gate mprj_ack_i_user mprj_iena_wb user_wb_ack_gate/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_5_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[52\] la_data_out_core[52] la_iena_mprj[52] user_to_mprj_in_gates\[52\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_user_to_mprj_in_gates\[61\]_A1 la_data_out_core[61] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[5\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[22\] user_to_mprj_in_gates\[22\]/ZN la_data_in_mprj[22]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_3_1456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[27\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__163__I mprj_dat_o_core[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xla_buf\[26\] _001_/ZN la_data_out_mprj[26] la_data_in_core[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
X_194_ mprj_sel_o_core[1] mprj_sel_o_user[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_wb_dat_gates\[28\] mprj_dat_i_user[28] mprj_iena_wb user_wb_dat_gates\[28\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_to_mprj_in_gates\[15\] la_data_out_core[15] la_iena_mprj[15] user_to_mprj_in_gates\[15\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__073__I la_oenb_mprj[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_buffers\[25\] user_wb_dat_gates\[25\]/ZN mprj_dat_i_core[25] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_user_to_mprj_in_gates\[28\]_A2 la_iena_mprj[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__158__I mprj_adr_o_core[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_177_ mprj_dat_o_core[16] mprj_dat_o_user[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__068__I la_oenb_mprj[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_wb_dat_gates\[17\]_A1 mprj_dat_i_user[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_100_ la_oenb_mprj[36] la_oenb_core[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_031_ la_oenb_mprj[56] _031_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_4_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_1724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[18\]_A1 la_data_out_core[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_wb_dat_buffers\[29\]_I user_wb_dat_gates\[29\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_gates\[2\]_A1 la_data_out_core[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__171__I mprj_dat_o_core[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xla_buf\[4\] _043_/ZN la_data_out_mprj[4] la_data_in_core[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
X_014_ la_oenb_mprj[39] _014_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[52\] user_to_mprj_in_gates\[52\]/ZN la_data_in_mprj[52]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
Xuser_wb_dat_gates\[10\] mprj_dat_i_user[10] mprj_iena_wb user_wb_dat_gates\[10\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_1_1598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__081__I la_oenb_mprj[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_buffers\[6\]_I user_wb_dat_gates\[6\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[9\]_I la_data_out_mprj[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__166__I mprj_dat_o_core[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xla_buf\[56\] _031_/ZN la_data_out_mprj[56] la_data_in_core[56] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_5_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__076__I la_oenb_mprj[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[45\] la_data_out_core[45] la_iena_mprj[45] user_to_mprj_in_gates\[45\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_user_to_mprj_in_gates\[61\]_A2 la_iena_mprj[61] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[7\] la_data_out_core[7] la_iena_mprj[7] user_to_mprj_in_gates\[7\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_6_1284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[7\]_I user_to_mprj_in_gates\[7\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_buffers\[15\] user_to_mprj_in_gates\[15\]/ZN la_data_in_mprj[15]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_1_1192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[7\] user_to_mprj_in_gates\[7\]/ZN la_data_in_mprj[7] VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
X_193_ mprj_sel_o_core[0] mprj_sel_o_user[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_user_to_mprj_in_gates\[51\]_A1 la_data_out_core[51] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xla_buf\[19\] _058_/ZN la_data_out_mprj[19] la_data_in_core[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_1_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_wb_dat_buffers\[18\] user_wb_dat_gates\[18\]/ZN mprj_dat_i_core[18] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_3_1243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__174__I mprj_dat_o_core[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_176_ mprj_dat_o_core[15] mprj_dat_o_user[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_user_wb_dat_gates\[17\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__084__I la_oenb_mprj[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_030_ la_oenb_mprj[55] _030_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__169__I mprj_dat_o_core[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_159_ mprj_adr_o_core[31] mprj_adr_o_user[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_user_to_mprj_in_gates\[18\]_A2 la_iena_mprj[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__079__I la_oenb_mprj[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[2\]_A2 la_iena_mprj[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_wb_dat_gates\[8\]_A1 mprj_dat_i_user[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_013_ la_oenb_mprj[38] _013_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_to_mprj_in_buffers\[45\] user_to_mprj_in_gates\[45\]/ZN la_data_in_mprj[45]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_2_1308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__182__I mprj_dat_o_core[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xla_buf\[49\] _024_/ZN la_data_out_mprj[49] la_data_in_core[49] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_5_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[60\]_I user_to_mprj_in_gates\[60\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[38\] la_data_out_core[38] la_iena_mprj[38] user_to_mprj_in_gates\[38\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__092__I la_oenb_mprj[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_buffers\[51\]_I user_to_mprj_in_gates\[51\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_buffers\[42\]_I user_to_mprj_in_gates\[42\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__177__I mprj_dat_o_core[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__087__I la_oenb_mprj[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_buffers\[33\]_I user_to_mprj_in_gates\[33\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[24\]_I user_to_mprj_in_gates\[24\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_192_ mprj_dat_o_core[31] mprj_dat_o_user[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_user_to_mprj_in_gates\[51\]_A2 la_iena_mprj[51] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_buffers\[15\]_I user_to_mprj_in_gates\[15\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[55\]_I la_data_out_mprj[55] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_la_buf\[46\]_I la_data_out_mprj[46] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[37\]_I la_data_out_mprj[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xla_buf\[31\] _006_/ZN la_data_out_mprj[31] la_data_in_core[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XANTENNA__190__I mprj_dat_o_core[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_175_ mprj_dat_o_core[14] mprj_dat_o_user[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xuser_wb_dat_gates\[3\] mprj_dat_i_user[3] mprj_iena_wb user_wb_dat_gates\[3\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_6_1818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[28\]_I la_data_out_mprj[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[20\] la_data_out_core[20] la_iena_mprj[20] user_to_mprj_in_gates\[20\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_wb_dat_buffers\[30\] user_wb_dat_gates\[30\]/ZN mprj_dat_i_core[30] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_5_1306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[41\]_A1 la_data_out_core[41] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[19\]_I la_data_out_mprj[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__185__I mprj_dat_o_core[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_089_ la_oenb_mprj[25] la_oenb_core[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_158_ mprj_adr_o_core[30] mprj_adr_o_user[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__095__I la_oenb_mprj[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_user_wb_dat_gates\[8\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_012_ la_oenb_mprj[37] _012_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_4_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[38\] user_to_mprj_in_gates\[38\]/ZN la_data_in_mprj[38]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_6_1434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__193__I mprj_sel_o_core[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xla_buf\[61\] _036_/ZN la_data_out_mprj[61] la_data_in_core[61] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_5_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[50\] la_data_out_core[50] la_iena_mprj[50] user_to_mprj_in_gates\[50\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_1_1172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_buffers\[10\]_I user_wb_dat_gates\[10\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_191_ mprj_dat_o_core[30] mprj_dat_o_user[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xuser_irq_gates\[2\] user_irq_core[2] user_irq_ena[2] user_irq_gates\[2\]/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_4_1702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__188__I mprj_dat_o_core[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[20\] user_to_mprj_in_gates\[20\]/ZN la_data_in_mprj[20]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_user_to_mprj_in_gates\[5\]_A1 la_data_out_core[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__098__I la_oenb_mprj[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_174_ mprj_dat_o_core[13] mprj_dat_o_user[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xla_buf\[24\] _063_/ZN la_data_out_mprj[24] la_data_in_core[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_2_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_wb_dat_gates\[26\] mprj_dat_i_user[26] mprj_iena_wb user_wb_dat_gates\[26\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_to_mprj_in_gates\[13\] la_data_out_core[13] la_iena_mprj[13] user_to_mprj_in_gates\[13\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_wb_dat_buffers\[23\] user_wb_dat_gates\[23\]/ZN mprj_dat_i_core[23] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_5_1329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_gates\[41\]_A2 la_iena_mprj[41] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_157_ mprj_adr_o_core[29] mprj_adr_o_user[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_088_ la_oenb_mprj[24] la_oenb_core[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_user_wb_dat_gates\[30\]_A1 mprj_dat_i_user[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_user_wb_dat_buffers\[9\]_I user_wb_dat_gates\[9\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_011_ la_oenb_mprj[36] _011_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_3_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__196__I mprj_sel_o_core[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[31\]_A1 la_data_out_core[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[54\]_A1 la_data_out_core[54] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xla_buf\[2\] _041_/ZN la_data_out_mprj[2] la_data_in_core[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_0_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_to_mprj_in_buffers\[50\] user_to_mprj_in_gates\[50\]/ZN la_data_in_mprj[50]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_6_1276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xla_buf\[54\] _029_/ZN la_data_out_mprj[54] la_data_in_core[54] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_5_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_wb_dat_buffers\[8\] user_wb_dat_gates\[8\]/ZN mprj_dat_i_core[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
Xuser_to_mprj_in_gates\[43\] la_data_out_core[43] la_iena_mprj[43] user_to_mprj_in_gates\[43\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_to_mprj_in_gates\[5\] la_data_out_core[5] la_iena_mprj[5] user_to_mprj_in_gates\[5\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_6_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_190_ mprj_dat_o_core[29] mprj_dat_o_user[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[13\] user_to_mprj_in_gates\[13\]/ZN la_data_in_mprj[13]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_user_to_mprj_in_gates\[5\]_A2 la_iena_mprj[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_173_ mprj_dat_o_core[12] mprj_dat_o_user[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xuser_to_mprj_in_buffers\[5\] user_to_mprj_in_gates\[5\]/ZN la_data_in_mprj[5] VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_2_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xla_buf\[17\] _056_/ZN la_data_out_mprj[17] la_data_in_core[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_6_1809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__199__I caravel_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_gates\[19\] mprj_dat_i_user[19] mprj_iena_wb user_wb_dat_gates\[19\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_5_1308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_wb_dat_buffers\[16\] user_wb_dat_gates\[16\]/ZN mprj_dat_i_core[16] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_3_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_irq_gates\[2\]_A1 user_irq_core[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[11\]_EN _050_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_087_ la_oenb_mprj[23] la_oenb_core[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_156_ mprj_adr_o_core[28] mprj_adr_o_user[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[30\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_010_ la_oenb_mprj[35] _010_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_4_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[2\]_EN _041_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_139_ mprj_adr_o_core[11] mprj_adr_o_user[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_user_to_mprj_in_gates\[31\]_A2 la_iena_mprj[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[54\]_I user_to_mprj_in_gates\[54\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[20\]_A1 mprj_dat_i_user[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_to_mprj_in_gates\[54\]_A2 la_iena_mprj[54] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_buffers\[45\]_I user_to_mprj_in_gates\[45\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__000__I la_oenb_mprj[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_buffers\[43\] user_to_mprj_in_gates\[43\]/ZN la_data_in_mprj[43]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_user_to_mprj_in_buffers\[36\]_I user_to_mprj_in_gates\[36\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_to_mprj_in_buffers\[27\]_I user_to_mprj_in_gates\[27\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[21\]_A1 la_data_out_core[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xla_buf\[47\] _022_/ZN la_data_out_mprj[47] la_data_in_core[47] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_5_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[18\]_I user_to_mprj_in_gates\[18\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[58\]_I la_data_out_mprj[58] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[36\] la_data_out_core[36] la_iena_mprj[36] user_to_mprj_in_gates\[36\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_6_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_user_to_mprj_in_gates\[44\]_A1 la_data_out_core[44] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[49\]_I la_data_out_mprj[49] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_172_ mprj_dat_o_core[11] mprj_dat_o_user[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_irq_gates\[2\]_A2 user_irq_ena[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xuser_wb_dat_gates\[1\] mprj_dat_i_user[1] mprj_iena_wb user_wb_dat_gates\[1\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_086_ la_oenb_mprj[22] la_oenb_core[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_155_ mprj_adr_o_core[27] mprj_adr_o_user[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__003__I la_oenb_mprj[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_wb_dat_gates\[31\] mprj_dat_i_user[31] mprj_iena_wb user_wb_dat_gates\[31\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_1784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_069_ la_oenb_mprj[5] la_oenb_core[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_138_ mprj_adr_o_core[10] mprj_adr_o_user[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_wb_dat_buffers\[31\]_I user_wb_dat_gates\[31\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_wb_dat_gates\[20\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[24\]_EN _063_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[36\] user_to_mprj_in_gates\[36\]/ZN la_data_in_mprj[36]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_user_to_mprj_in_gates\[8\]_A1 la_data_out_core[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_wb_dat_buffers\[13\]_I user_wb_dat_gates\[13\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__101__I la_oenb_mprj[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[21\]_A2 la_iena_mprj[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__011__I la_oenb_mprj[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[29\] la_data_out_core[29] la_iena_mprj[29] user_to_mprj_in_gates\[29\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_user_wb_dat_gates\[10\]_A1 mprj_dat_i_user[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[44\]_A2 la_iena_mprj[44] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[2\]_I la_data_out_mprj[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__006__I la_oenb_mprj[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[11\]_A1 la_data_out_core[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[0\]_I user_to_mprj_in_gates\[0\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_171_ mprj_dat_o_core[10] mprj_dat_o_user[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xuser_irq_gates\[0\] user_irq_core[0] user_irq_ena[0] user_irq_gates\[0\]/ZN VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_2_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[34\]_A1 la_data_out_core[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_to_mprj_in_gates\[57\]_A1 la_data_out_core[57] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_085_ la_oenb_mprj[21] la_oenb_core[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_154_ mprj_adr_o_core[26] mprj_adr_o_user[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xla_buf\[22\] _061_/ZN la_data_out_mprj[22] la_data_in_core[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_0_1218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_wb_dat_gates\[24\] mprj_dat_i_user[24] mprj_iena_wb user_wb_dat_gates\[24\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_to_mprj_in_gates\[11\] la_data_out_core[11] la_iena_mprj[11] user_to_mprj_in_gates\[11\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_wb_dat_buffers\[21\] user_wb_dat_gates\[21\]/ZN mprj_dat_i_core[21] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_0_1774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__104__I la_oenb_mprj[40] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_137_ mprj_adr_o_core[9] mprj_adr_o_user[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_068_ la_oenb_mprj[4] la_oenb_core[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__014__I la_oenb_mprj[39] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[59\] la_data_out_core[59] la_iena_mprj[59] user_to_mprj_in_gates\[59\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_1560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__009__I la_oenb_mprj[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_to_mprj_in_buffers\[29\] user_to_mprj_in_gates\[29\]/ZN la_data_in_mprj[29]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_6_1224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_user_to_mprj_in_gates\[8\]_A2 la_iena_mprj[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xla_buf\[0\] _039_/ZN la_data_out_mprj[0] la_data_in_core[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_5_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_wb_dat_gates\[10\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__112__I la_oenb_mprj[48] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xla_buf\[52\] _027_/ZN la_data_out_mprj[52] la_data_in_core[52] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_5_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__022__I la_oenb_mprj[47] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[41\] la_data_out_core[41] la_iena_mprj[41] user_to_mprj_in_gates\[41\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_wb_dat_buffers\[6\] user_wb_dat_gates\[6\]/ZN mprj_dat_i_core[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XTAP_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[11\]_A2 la_iena_mprj[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[3\] la_data_out_core[3] la_iena_mprj[3] user_to_mprj_in_gates\[3\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_170_ mprj_dat_o_core[9] mprj_dat_o_user[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__107__I la_oenb_mprj[43] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_la_buf\[5\]_EN _044_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[1\]_A1 mprj_dat_i_user[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_buffers\[11\] user_to_mprj_in_gates\[11\]/ZN la_data_in_mprj[11]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA__017__I la_oenb_mprj[42] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[34\]_A2 la_iena_mprj[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_wb_dat_gates\[23\]_A1 mprj_dat_i_user[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_153_ mprj_adr_o_core[25] mprj_adr_o_user[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xuser_to_mprj_in_buffers\[3\] user_to_mprj_in_gates\[3\]/ZN la_data_in_mprj[3] VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_user_to_mprj_in_gates\[57\]_A2 la_iena_mprj[57] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_084_ la_oenb_mprj[20] la_oenb_core[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xla_buf\[15\] _054_/ZN la_data_out_mprj[15] la_data_in_core[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_3_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_to_mprj_in_buffers\[59\] user_to_mprj_in_gates\[59\]/ZN la_data_in_mprj[59]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
Xuser_wb_dat_gates\[17\] mprj_dat_i_user[17] mprj_iena_wb user_wb_dat_gates\[17\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xuser_wb_dat_buffers\[14\] user_wb_dat_gates\[14\]/ZN mprj_dat_i_core[14] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_0_1731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[57\]_I user_to_mprj_in_gates\[57\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[30\]_I la_data_out_mprj[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__120__I la_oenb_mprj[56] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_gates\[24\]_A1 la_data_out_core[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_136_ mprj_adr_o_core[8] mprj_adr_o_user[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_067_ la_oenb_mprj[3] la_oenb_core[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_user_to_mprj_in_buffers\[48\]_I user_to_mprj_in_gates\[48\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[21\]_I la_data_out_mprj[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__030__I la_oenb_mprj[55] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_buffers\[39\]_I user_to_mprj_in_gates\[39\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[12\]_I la_data_out_mprj[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[47\]_A1 la_data_out_core[47] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__115__I la_oenb_mprj[51] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_119_ la_oenb_mprj[55] la_oenb_core[55] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__025__I la_oenb_mprj[50] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[41\] user_to_mprj_in_gates\[41\]/ZN la_data_in_mprj[41]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_2_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xla_buf\[45\] _020_/ZN la_data_out_mprj[45] la_data_in_core[45] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_5_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[34\] la_data_out_core[34] la_iena_mprj[34] user_to_mprj_in_gates\[34\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__123__I la_oenb_mprj[59] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[1\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__033__I la_oenb_mprj[58] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__118__I la_oenb_mprj[54] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_wb_dat_gates\[23\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_083_ la_oenb_mprj[19] la_oenb_core[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_152_ mprj_adr_o_core[24] mprj_adr_o_user[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__028__I la_oenb_mprj[53] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_la_buf\[27\]_EN _002_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_user_to_mprj_in_gates\[24\]_A2 la_iena_mprj[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_066_ la_oenb_mprj[2] la_oenb_core[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_135_ mprj_adr_o_core[7] mprj_adr_o_user[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_to_mprj_in_gates\[47\]_A2 la_iena_mprj[47] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_wb_dat_buffers\[16\]_I user_wb_dat_gates\[16\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_wb_dat_gates\[13\]_A1 mprj_dat_i_user[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__131__I mprj_adr_o_core[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_118_ la_oenb_mprj[54] la_oenb_core[54] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_049_ la_oenb_mprj[10] _049_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_1259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__041__I la_oenb_mprj[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_buffers\[2\]_I user_wb_dat_gates\[2\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[14\]_A1 la_data_out_core[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[5\]_I la_data_out_mprj[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__126__I la_oenb_mprj[62] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_1134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_buffers\[34\] user_to_mprj_in_gates\[34\]/ZN la_data_in_mprj[34]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_user_to_mprj_in_gates\[37\]_A1 la_data_out_core[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__036__I la_oenb_mprj[61] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[3\]_I user_to_mprj_in_gates\[3\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xla_buf\[38\] _013_/ZN la_data_out_mprj[38] la_data_in_core[38] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_5_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_to_mprj_in_gates\[27\] la_data_out_core[27] la_iena_mprj[27] user_to_mprj_in_gates\[27\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_082_ la_oenb_mprj[18] la_oenb_core[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__134__I mprj_adr_o_core[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_151_ mprj_adr_o_core[23] mprj_adr_o_user[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__044__I la_oenb_mprj[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__129__I mprj_adr_o_core[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_065_ la_oenb_mprj[1] la_oenb_core[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_134_ mprj_adr_o_core[6] mprj_adr_o_user[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xla_buf\[20\] _059_/ZN la_data_out_mprj[20] la_data_in_core[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_6_1408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__039__I la_oenb_mprj[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_wb_dat_gates\[22\] mprj_dat_i_user[22] mprj_iena_wb user_wb_dat_gates\[22\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_user_wb_dat_gates\[13\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_117_ la_oenb_mprj[53] la_oenb_core[53] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_048_ la_oenb_mprj[9] _048_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_1216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_to_mprj_in_gates\[57\] la_data_out_core[57] la_iena_mprj[57] user_to_mprj_in_gates\[57\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_1_1894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[14\]_A2 la_iena_mprj[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__142__I mprj_adr_o_core[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_la_buf\[8\]_EN _047_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[4\]_A1 mprj_dat_i_user[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xuser_to_mprj_in_buffers\[27\] user_to_mprj_in_gates\[27\]/ZN la_data_in_mprj[27]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA_user_to_mprj_in_gates\[37\]_A2 la_iena_mprj[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__052__I la_oenb_mprj[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__137__I mprj_adr_o_core[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_wb_dat_gates\[26\]_A1 mprj_dat_i_user[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__047__I la_oenb_mprj[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[20\]_I user_to_mprj_in_gates\[20\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[60\]_I la_data_out_mprj[60] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_buffers\[11\]_I user_to_mprj_in_gates\[11\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[27\]_A1 la_data_out_core[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xla_buf\[50\] _025_/ZN la_data_out_mprj[50] la_data_in_core[50] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_2_1296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[51\]_I la_data_out_mprj[51] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_wb_dat_buffers\[4\] user_wb_dat_gates\[4\]/ZN mprj_dat_i_core[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_0_1937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_la_buf\[42\]_I la_data_out_mprj[42] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xuser_to_mprj_in_gates\[1\] la_data_out_core[1] la_iena_mprj[1] user_to_mprj_in_gates\[1\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_5_1804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_150_ mprj_adr_o_core[22] mprj_adr_o_user[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_081_ la_oenb_mprj[17] la_oenb_core[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_la_buf\[33\]_I la_data_out_mprj[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__150__I mprj_adr_o_core[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[24\]_I la_data_out_mprj[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__060__I la_oenb_mprj[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[15\]_I la_data_out_mprj[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_133_ mprj_adr_o_core[5] mprj_adr_o_user[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xuser_to_mprj_in_buffers\[1\] user_to_mprj_in_gates\[1\]/ZN la_data_in_mprj[1] VDD
+ VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XANTENNA__145__I mprj_adr_o_core[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_064_ la_oenb_mprj[0] la_oenb_core[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xla_buf\[9\] _048_/ZN la_data_out_mprj[9] la_data_in_core[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
Xla_buf\[13\] _052_/ZN la_data_out_mprj[13] la_data_in_core[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_4_1166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_to_mprj_in_buffers\[57\] user_to_mprj_in_gates\[57\]/ZN la_data_in_mprj[57]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
Xuser_wb_dat_gates\[15\] mprj_dat_i_user[15] mprj_iena_wb user_wb_dat_gates\[15\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__055__I la_oenb_mprj[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xuser_wb_dat_buffers\[12\] user_wb_dat_gates\[12\]/ZN mprj_dat_i_core[12] VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_5_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_116_ la_oenb_mprj[52] la_oenb_core[52] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_047_ la_oenb_mprj[8] _047_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_1784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_user_to_mprj_in_gates\[60\]_A1 la_data_out_core[60] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[4\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_gates\[26\]_A2 mprj_iena_wb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__153__I mprj_adr_o_core[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__063__I la_oenb_mprj[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__148__I mprj_adr_o_core[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[27\]_A2 la_iena_mprj[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xla_buf\[43\] _018_/ZN la_data_out_mprj[43] la_data_in_core[43] VDD VSS gf180mcu_fd_sc_mcu7t5v0__bufz_8
XFILLER_5_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__058__I la_oenb_mprj[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xuser_to_mprj_in_gates\[32\] la_data_out_core[32] la_iena_mprj[32] user_to_mprj_in_gates\[32\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_user_wb_dat_gates\[16\]_A1 mprj_dat_i_user[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_080_ la_oenb_mprj[16] la_oenb_core[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_buffers\[28\]_I user_wb_dat_gates\[28\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[17\]_A1 la_data_out_core[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_user_to_mprj_in_gates\[1\]_A1 la_data_out_core[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_201_ caravel_rstn user_reset VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_132_ mprj_adr_o_core[4] mprj_adr_o_user[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_063_ la_oenb_mprj[24] _063_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__161__I mprj_dat_o_core[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__071__I la_oenb_mprj[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_wb_dat_buffers\[5\]_I user_wb_dat_gates\[5\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_la_buf\[8\]_I la_data_out_mprj[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__156__I mprj_adr_o_core[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_046_ la_oenb_mprj[7] _046_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_115_ la_oenb_mprj[51] la_oenb_core[51] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__066__I la_oenb_mprj[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[60\]_A2 la_iena_mprj[60] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_buffers\[6\]_I user_to_mprj_in_gates\[6\]/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_029_ la_oenb_mprj[54] _029_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_6_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xuser_to_mprj_in_gates\[62\] la_data_out_core[62] la_iena_mprj[62] user_to_mprj_in_gates\[62\]/ZN
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_1_1671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xuser_to_mprj_in_buffers\[32\] user_to_mprj_in_gates\[32\]/ZN la_data_in_mprj[32]
+ VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XTAP_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_user_to_mprj_in_gates\[50\]_A1 la_data_out_core[50] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

