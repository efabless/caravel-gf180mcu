magic
tech gf180mcuC
magscale 1 5
timestamp 1655473269
<< checkpaint >>
rect -2518 -1622 302510 301502
<< obsm1 >>
rect 672 1387 299507 298342
<< metal2 >>
rect 5488 299760 5600 300480
rect 16576 299760 16688 300480
rect 27664 299760 27776 300480
rect 38808 299760 38920 300480
rect 49896 299760 50008 300480
rect 61040 299760 61152 300480
rect 72128 299760 72240 300480
rect 83272 299760 83384 300480
rect 94360 299760 94472 300480
rect 105504 299760 105616 300480
rect 116592 299760 116704 300480
rect 127680 299760 127792 300480
rect 138824 299760 138936 300480
rect 149912 299760 150024 300480
rect 161056 299760 161168 300480
rect 172144 299760 172256 300480
rect 183288 299760 183400 300480
rect 194376 299760 194488 300480
rect 205520 299760 205632 300480
rect 216608 299760 216720 300480
rect 227696 299760 227808 300480
rect 238840 299760 238952 300480
rect 249928 299760 250040 300480
rect 261072 299760 261184 300480
rect 272160 299760 272272 300480
rect 283304 299760 283416 300480
rect 294392 299760 294504 300480
rect 392 -480 504 240
rect 1344 -480 1456 240
rect 2352 -480 2464 240
rect 3360 -480 3472 240
rect 4312 -480 4424 240
rect 5320 -480 5432 240
rect 6328 -480 6440 240
rect 7336 -480 7448 240
rect 8288 -480 8400 240
rect 9296 -480 9408 240
rect 10304 -480 10416 240
rect 11312 -480 11424 240
rect 12264 -480 12376 240
rect 13272 -480 13384 240
rect 14280 -480 14392 240
rect 15288 -480 15400 240
rect 16240 -480 16352 240
rect 17248 -480 17360 240
rect 18256 -480 18368 240
rect 19264 -480 19376 240
rect 20216 -480 20328 240
rect 21224 -480 21336 240
rect 22232 -480 22344 240
rect 23240 -480 23352 240
rect 24192 -480 24304 240
rect 25200 -480 25312 240
rect 26208 -480 26320 240
rect 27216 -480 27328 240
rect 28168 -480 28280 240
rect 29176 -480 29288 240
rect 30184 -480 30296 240
rect 31136 -480 31248 240
rect 32144 -480 32256 240
rect 33152 -480 33264 240
rect 34160 -480 34272 240
rect 35112 -480 35224 240
rect 36120 -480 36232 240
rect 37128 -480 37240 240
rect 38136 -480 38248 240
rect 39088 -480 39200 240
rect 40096 -480 40208 240
rect 41104 -480 41216 240
rect 42112 -480 42224 240
rect 43064 -480 43176 240
rect 44072 -480 44184 240
rect 45080 -480 45192 240
rect 46088 -480 46200 240
rect 47040 -480 47152 240
rect 48048 -480 48160 240
rect 49056 -480 49168 240
rect 50064 -480 50176 240
rect 51016 -480 51128 240
rect 52024 -480 52136 240
rect 53032 -480 53144 240
rect 54040 -480 54152 240
rect 54992 -480 55104 240
rect 56000 -480 56112 240
rect 57008 -480 57120 240
rect 58016 -480 58128 240
rect 58968 -480 59080 240
rect 59976 -480 60088 240
rect 60984 -480 61096 240
rect 61936 -480 62048 240
rect 62944 -480 63056 240
rect 63952 -480 64064 240
rect 64960 -480 65072 240
rect 65912 -480 66024 240
rect 66920 -480 67032 240
rect 67928 -480 68040 240
rect 68936 -480 69048 240
rect 69888 -480 70000 240
rect 70896 -480 71008 240
rect 71904 -480 72016 240
rect 72912 -480 73024 240
rect 73864 -480 73976 240
rect 74872 -480 74984 240
rect 75880 -480 75992 240
rect 76888 -480 77000 240
rect 77840 -480 77952 240
rect 78848 -480 78960 240
rect 79856 -480 79968 240
rect 80864 -480 80976 240
rect 81816 -480 81928 240
rect 82824 -480 82936 240
rect 83832 -480 83944 240
rect 84840 -480 84952 240
rect 85792 -480 85904 240
rect 86800 -480 86912 240
rect 87808 -480 87920 240
rect 88816 -480 88928 240
rect 89768 -480 89880 240
rect 90776 -480 90888 240
rect 91784 -480 91896 240
rect 92736 -480 92848 240
rect 93744 -480 93856 240
rect 94752 -480 94864 240
rect 95760 -480 95872 240
rect 96712 -480 96824 240
rect 97720 -480 97832 240
rect 98728 -480 98840 240
rect 99736 -480 99848 240
rect 100688 -480 100800 240
rect 101696 -480 101808 240
rect 102704 -480 102816 240
rect 103712 -480 103824 240
rect 104664 -480 104776 240
rect 105672 -480 105784 240
rect 106680 -480 106792 240
rect 107688 -480 107800 240
rect 108640 -480 108752 240
rect 109648 -480 109760 240
rect 110656 -480 110768 240
rect 111664 -480 111776 240
rect 112616 -480 112728 240
rect 113624 -480 113736 240
rect 114632 -480 114744 240
rect 115640 -480 115752 240
rect 116592 -480 116704 240
rect 117600 -480 117712 240
rect 118608 -480 118720 240
rect 119616 -480 119728 240
rect 120568 -480 120680 240
rect 121576 -480 121688 240
rect 122584 -480 122696 240
rect 123536 -480 123648 240
rect 124544 -480 124656 240
rect 125552 -480 125664 240
rect 126560 -480 126672 240
rect 127512 -480 127624 240
rect 128520 -480 128632 240
rect 129528 -480 129640 240
rect 130536 -480 130648 240
rect 131488 -480 131600 240
rect 132496 -480 132608 240
rect 133504 -480 133616 240
rect 134512 -480 134624 240
rect 135464 -480 135576 240
rect 136472 -480 136584 240
rect 137480 -480 137592 240
rect 138488 -480 138600 240
rect 139440 -480 139552 240
rect 140448 -480 140560 240
rect 141456 -480 141568 240
rect 142464 -480 142576 240
rect 143416 -480 143528 240
rect 144424 -480 144536 240
rect 145432 -480 145544 240
rect 146440 -480 146552 240
rect 147392 -480 147504 240
rect 148400 -480 148512 240
rect 149408 -480 149520 240
rect 150416 -480 150528 240
rect 151368 -480 151480 240
rect 152376 -480 152488 240
rect 153384 -480 153496 240
rect 154336 -480 154448 240
rect 155344 -480 155456 240
rect 156352 -480 156464 240
rect 157360 -480 157472 240
rect 158312 -480 158424 240
rect 159320 -480 159432 240
rect 160328 -480 160440 240
rect 161336 -480 161448 240
rect 162288 -480 162400 240
rect 163296 -480 163408 240
rect 164304 -480 164416 240
rect 165312 -480 165424 240
rect 166264 -480 166376 240
rect 167272 -480 167384 240
rect 168280 -480 168392 240
rect 169288 -480 169400 240
rect 170240 -480 170352 240
rect 171248 -480 171360 240
rect 172256 -480 172368 240
rect 173264 -480 173376 240
rect 174216 -480 174328 240
rect 175224 -480 175336 240
rect 176232 -480 176344 240
rect 177240 -480 177352 240
rect 178192 -480 178304 240
rect 179200 -480 179312 240
rect 180208 -480 180320 240
rect 181160 -480 181272 240
rect 182168 -480 182280 240
rect 183176 -480 183288 240
rect 184184 -480 184296 240
rect 185136 -480 185248 240
rect 186144 -480 186256 240
rect 187152 -480 187264 240
rect 188160 -480 188272 240
rect 189112 -480 189224 240
rect 190120 -480 190232 240
rect 191128 -480 191240 240
rect 192136 -480 192248 240
rect 193088 -480 193200 240
rect 194096 -480 194208 240
rect 195104 -480 195216 240
rect 196112 -480 196224 240
rect 197064 -480 197176 240
rect 198072 -480 198184 240
rect 199080 -480 199192 240
rect 200088 -480 200200 240
rect 201040 -480 201152 240
rect 202048 -480 202160 240
rect 203056 -480 203168 240
rect 204064 -480 204176 240
rect 205016 -480 205128 240
rect 206024 -480 206136 240
rect 207032 -480 207144 240
rect 208040 -480 208152 240
rect 208992 -480 209104 240
rect 210000 -480 210112 240
rect 211008 -480 211120 240
rect 211960 -480 212072 240
rect 212968 -480 213080 240
rect 213976 -480 214088 240
rect 214984 -480 215096 240
rect 215936 -480 216048 240
rect 216944 -480 217056 240
rect 217952 -480 218064 240
rect 218960 -480 219072 240
rect 219912 -480 220024 240
rect 220920 -480 221032 240
rect 221928 -480 222040 240
rect 222936 -480 223048 240
rect 223888 -480 224000 240
rect 224896 -480 225008 240
rect 225904 -480 226016 240
rect 226912 -480 227024 240
rect 227864 -480 227976 240
rect 228872 -480 228984 240
rect 229880 -480 229992 240
rect 230888 -480 231000 240
rect 231840 -480 231952 240
rect 232848 -480 232960 240
rect 233856 -480 233968 240
rect 234864 -480 234976 240
rect 235816 -480 235928 240
rect 236824 -480 236936 240
rect 237832 -480 237944 240
rect 238840 -480 238952 240
rect 239792 -480 239904 240
rect 240800 -480 240912 240
rect 241808 -480 241920 240
rect 242760 -480 242872 240
rect 243768 -480 243880 240
rect 244776 -480 244888 240
rect 245784 -480 245896 240
rect 246736 -480 246848 240
rect 247744 -480 247856 240
rect 248752 -480 248864 240
rect 249760 -480 249872 240
rect 250712 -480 250824 240
rect 251720 -480 251832 240
rect 252728 -480 252840 240
rect 253736 -480 253848 240
rect 254688 -480 254800 240
rect 255696 -480 255808 240
rect 256704 -480 256816 240
rect 257712 -480 257824 240
rect 258664 -480 258776 240
rect 259672 -480 259784 240
rect 260680 -480 260792 240
rect 261688 -480 261800 240
rect 262640 -480 262752 240
rect 263648 -480 263760 240
rect 264656 -480 264768 240
rect 265664 -480 265776 240
rect 266616 -480 266728 240
rect 267624 -480 267736 240
rect 268632 -480 268744 240
rect 269640 -480 269752 240
rect 270592 -480 270704 240
rect 271600 -480 271712 240
rect 272608 -480 272720 240
rect 273560 -480 273672 240
rect 274568 -480 274680 240
rect 275576 -480 275688 240
rect 276584 -480 276696 240
rect 277536 -480 277648 240
rect 278544 -480 278656 240
rect 279552 -480 279664 240
rect 280560 -480 280672 240
rect 281512 -480 281624 240
rect 282520 -480 282632 240
rect 283528 -480 283640 240
rect 284536 -480 284648 240
rect 285488 -480 285600 240
rect 286496 -480 286608 240
rect 287504 -480 287616 240
rect 288512 -480 288624 240
rect 289464 -480 289576 240
rect 290472 -480 290584 240
rect 291480 -480 291592 240
rect 292488 -480 292600 240
rect 293440 -480 293552 240
rect 294448 -480 294560 240
rect 295456 -480 295568 240
rect 296464 -480 296576 240
rect 297416 -480 297528 240
rect 298424 -480 298536 240
rect 299432 -480 299544 240
<< obsm2 >>
rect 826 299730 5458 299838
rect 5630 299730 16546 299838
rect 16718 299730 27634 299838
rect 27806 299730 38778 299838
rect 38950 299730 49866 299838
rect 50038 299730 61010 299838
rect 61182 299730 72098 299838
rect 72270 299730 83242 299838
rect 83414 299730 94330 299838
rect 94502 299730 105474 299838
rect 105646 299730 116562 299838
rect 116734 299730 127650 299838
rect 127822 299730 138794 299838
rect 138966 299730 149882 299838
rect 150054 299730 161026 299838
rect 161198 299730 172114 299838
rect 172286 299730 183258 299838
rect 183430 299730 194346 299838
rect 194518 299730 205490 299838
rect 205662 299730 216578 299838
rect 216750 299730 227666 299838
rect 227838 299730 238810 299838
rect 238982 299730 249898 299838
rect 250070 299730 261042 299838
rect 261214 299730 272130 299838
rect 272302 299730 283274 299838
rect 283446 299730 294362 299838
rect 294534 299730 299502 299838
rect 826 270 299502 299730
rect 826 210 1314 270
rect 1486 210 2322 270
rect 2494 210 3330 270
rect 3502 210 4282 270
rect 4454 210 5290 270
rect 5462 210 6298 270
rect 6470 210 7306 270
rect 7478 210 8258 270
rect 8430 210 9266 270
rect 9438 210 10274 270
rect 10446 210 11282 270
rect 11454 210 12234 270
rect 12406 210 13242 270
rect 13414 210 14250 270
rect 14422 210 15258 270
rect 15430 210 16210 270
rect 16382 210 17218 270
rect 17390 210 18226 270
rect 18398 210 19234 270
rect 19406 210 20186 270
rect 20358 210 21194 270
rect 21366 210 22202 270
rect 22374 210 23210 270
rect 23382 210 24162 270
rect 24334 210 25170 270
rect 25342 210 26178 270
rect 26350 210 27186 270
rect 27358 210 28138 270
rect 28310 210 29146 270
rect 29318 210 30154 270
rect 30326 210 31106 270
rect 31278 210 32114 270
rect 32286 210 33122 270
rect 33294 210 34130 270
rect 34302 210 35082 270
rect 35254 210 36090 270
rect 36262 210 37098 270
rect 37270 210 38106 270
rect 38278 210 39058 270
rect 39230 210 40066 270
rect 40238 210 41074 270
rect 41246 210 42082 270
rect 42254 210 43034 270
rect 43206 210 44042 270
rect 44214 210 45050 270
rect 45222 210 46058 270
rect 46230 210 47010 270
rect 47182 210 48018 270
rect 48190 210 49026 270
rect 49198 210 50034 270
rect 50206 210 50986 270
rect 51158 210 51994 270
rect 52166 210 53002 270
rect 53174 210 54010 270
rect 54182 210 54962 270
rect 55134 210 55970 270
rect 56142 210 56978 270
rect 57150 210 57986 270
rect 58158 210 58938 270
rect 59110 210 59946 270
rect 60118 210 60954 270
rect 61126 210 61906 270
rect 62078 210 62914 270
rect 63086 210 63922 270
rect 64094 210 64930 270
rect 65102 210 65882 270
rect 66054 210 66890 270
rect 67062 210 67898 270
rect 68070 210 68906 270
rect 69078 210 69858 270
rect 70030 210 70866 270
rect 71038 210 71874 270
rect 72046 210 72882 270
rect 73054 210 73834 270
rect 74006 210 74842 270
rect 75014 210 75850 270
rect 76022 210 76858 270
rect 77030 210 77810 270
rect 77982 210 78818 270
rect 78990 210 79826 270
rect 79998 210 80834 270
rect 81006 210 81786 270
rect 81958 210 82794 270
rect 82966 210 83802 270
rect 83974 210 84810 270
rect 84982 210 85762 270
rect 85934 210 86770 270
rect 86942 210 87778 270
rect 87950 210 88786 270
rect 88958 210 89738 270
rect 89910 210 90746 270
rect 90918 210 91754 270
rect 91926 210 92706 270
rect 92878 210 93714 270
rect 93886 210 94722 270
rect 94894 210 95730 270
rect 95902 210 96682 270
rect 96854 210 97690 270
rect 97862 210 98698 270
rect 98870 210 99706 270
rect 99878 210 100658 270
rect 100830 210 101666 270
rect 101838 210 102674 270
rect 102846 210 103682 270
rect 103854 210 104634 270
rect 104806 210 105642 270
rect 105814 210 106650 270
rect 106822 210 107658 270
rect 107830 210 108610 270
rect 108782 210 109618 270
rect 109790 210 110626 270
rect 110798 210 111634 270
rect 111806 210 112586 270
rect 112758 210 113594 270
rect 113766 210 114602 270
rect 114774 210 115610 270
rect 115782 210 116562 270
rect 116734 210 117570 270
rect 117742 210 118578 270
rect 118750 210 119586 270
rect 119758 210 120538 270
rect 120710 210 121546 270
rect 121718 210 122554 270
rect 122726 210 123506 270
rect 123678 210 124514 270
rect 124686 210 125522 270
rect 125694 210 126530 270
rect 126702 210 127482 270
rect 127654 210 128490 270
rect 128662 210 129498 270
rect 129670 210 130506 270
rect 130678 210 131458 270
rect 131630 210 132466 270
rect 132638 210 133474 270
rect 133646 210 134482 270
rect 134654 210 135434 270
rect 135606 210 136442 270
rect 136614 210 137450 270
rect 137622 210 138458 270
rect 138630 210 139410 270
rect 139582 210 140418 270
rect 140590 210 141426 270
rect 141598 210 142434 270
rect 142606 210 143386 270
rect 143558 210 144394 270
rect 144566 210 145402 270
rect 145574 210 146410 270
rect 146582 210 147362 270
rect 147534 210 148370 270
rect 148542 210 149378 270
rect 149550 210 150386 270
rect 150558 210 151338 270
rect 151510 210 152346 270
rect 152518 210 153354 270
rect 153526 210 154306 270
rect 154478 210 155314 270
rect 155486 210 156322 270
rect 156494 210 157330 270
rect 157502 210 158282 270
rect 158454 210 159290 270
rect 159462 210 160298 270
rect 160470 210 161306 270
rect 161478 210 162258 270
rect 162430 210 163266 270
rect 163438 210 164274 270
rect 164446 210 165282 270
rect 165454 210 166234 270
rect 166406 210 167242 270
rect 167414 210 168250 270
rect 168422 210 169258 270
rect 169430 210 170210 270
rect 170382 210 171218 270
rect 171390 210 172226 270
rect 172398 210 173234 270
rect 173406 210 174186 270
rect 174358 210 175194 270
rect 175366 210 176202 270
rect 176374 210 177210 270
rect 177382 210 178162 270
rect 178334 210 179170 270
rect 179342 210 180178 270
rect 180350 210 181130 270
rect 181302 210 182138 270
rect 182310 210 183146 270
rect 183318 210 184154 270
rect 184326 210 185106 270
rect 185278 210 186114 270
rect 186286 210 187122 270
rect 187294 210 188130 270
rect 188302 210 189082 270
rect 189254 210 190090 270
rect 190262 210 191098 270
rect 191270 210 192106 270
rect 192278 210 193058 270
rect 193230 210 194066 270
rect 194238 210 195074 270
rect 195246 210 196082 270
rect 196254 210 197034 270
rect 197206 210 198042 270
rect 198214 210 199050 270
rect 199222 210 200058 270
rect 200230 210 201010 270
rect 201182 210 202018 270
rect 202190 210 203026 270
rect 203198 210 204034 270
rect 204206 210 204986 270
rect 205158 210 205994 270
rect 206166 210 207002 270
rect 207174 210 208010 270
rect 208182 210 208962 270
rect 209134 210 209970 270
rect 210142 210 210978 270
rect 211150 210 211930 270
rect 212102 210 212938 270
rect 213110 210 213946 270
rect 214118 210 214954 270
rect 215126 210 215906 270
rect 216078 210 216914 270
rect 217086 210 217922 270
rect 218094 210 218930 270
rect 219102 210 219882 270
rect 220054 210 220890 270
rect 221062 210 221898 270
rect 222070 210 222906 270
rect 223078 210 223858 270
rect 224030 210 224866 270
rect 225038 210 225874 270
rect 226046 210 226882 270
rect 227054 210 227834 270
rect 228006 210 228842 270
rect 229014 210 229850 270
rect 230022 210 230858 270
rect 231030 210 231810 270
rect 231982 210 232818 270
rect 232990 210 233826 270
rect 233998 210 234834 270
rect 235006 210 235786 270
rect 235958 210 236794 270
rect 236966 210 237802 270
rect 237974 210 238810 270
rect 238982 210 239762 270
rect 239934 210 240770 270
rect 240942 210 241778 270
rect 241950 210 242730 270
rect 242902 210 243738 270
rect 243910 210 244746 270
rect 244918 210 245754 270
rect 245926 210 246706 270
rect 246878 210 247714 270
rect 247886 210 248722 270
rect 248894 210 249730 270
rect 249902 210 250682 270
rect 250854 210 251690 270
rect 251862 210 252698 270
rect 252870 210 253706 270
rect 253878 210 254658 270
rect 254830 210 255666 270
rect 255838 210 256674 270
rect 256846 210 257682 270
rect 257854 210 258634 270
rect 258806 210 259642 270
rect 259814 210 260650 270
rect 260822 210 261658 270
rect 261830 210 262610 270
rect 262782 210 263618 270
rect 263790 210 264626 270
rect 264798 210 265634 270
rect 265806 210 266586 270
rect 266758 210 267594 270
rect 267766 210 268602 270
rect 268774 210 269610 270
rect 269782 210 270562 270
rect 270734 210 271570 270
rect 271742 210 272578 270
rect 272750 210 273530 270
rect 273702 210 274538 270
rect 274710 210 275546 270
rect 275718 210 276554 270
rect 276726 210 277506 270
rect 277678 210 278514 270
rect 278686 210 279522 270
rect 279694 210 280530 270
rect 280702 210 281482 270
rect 281654 210 282490 270
rect 282662 210 283498 270
rect 283670 210 284506 270
rect 284678 210 285458 270
rect 285630 210 286466 270
rect 286638 210 287474 270
rect 287646 210 288482 270
rect 288654 210 289434 270
rect 289606 210 290442 270
rect 290614 210 291450 270
rect 291622 210 292458 270
rect 292630 210 293410 270
rect 293582 210 294418 270
rect 294590 210 295426 270
rect 295598 210 296434 270
rect 296606 210 297386 270
rect 297558 210 298394 270
rect 298566 210 299402 270
<< metal3 >>
rect 299760 296576 300480 296688
rect -480 296352 240 296464
rect 299760 289912 300480 290024
rect -480 289184 240 289296
rect 299760 283248 300480 283360
rect -480 282072 240 282184
rect 299760 276584 300480 276696
rect -480 274904 240 275016
rect 299760 269920 300480 270032
rect -480 267792 240 267904
rect 299760 263256 300480 263368
rect -480 260624 240 260736
rect 299760 256592 300480 256704
rect -480 253512 240 253624
rect 299760 249928 300480 250040
rect -480 246344 240 246456
rect 299760 243264 300480 243376
rect -480 239232 240 239344
rect 299760 236600 300480 236712
rect -480 232064 240 232176
rect 299760 229936 300480 230048
rect -480 224896 240 225008
rect 299760 223272 300480 223384
rect -480 217784 240 217896
rect 299760 216608 300480 216720
rect -480 210616 240 210728
rect 299760 209944 300480 210056
rect -480 203504 240 203616
rect 299760 203280 300480 203392
rect 299760 196616 300480 196728
rect -480 196336 240 196448
rect 299760 189952 300480 190064
rect -480 189224 240 189336
rect 299760 183288 300480 183400
rect -480 182056 240 182168
rect 299760 176624 300480 176736
rect -480 174944 240 175056
rect 299760 169960 300480 170072
rect -480 167776 240 167888
rect 299760 163296 300480 163408
rect -480 160664 240 160776
rect 299760 156632 300480 156744
rect -480 153496 240 153608
rect 299760 149912 300480 150024
rect -480 146328 240 146440
rect 299760 143248 300480 143360
rect -480 139216 240 139328
rect 299760 136584 300480 136696
rect -480 132048 240 132160
rect 299760 129920 300480 130032
rect -480 124936 240 125048
rect 299760 123256 300480 123368
rect -480 117768 240 117880
rect 299760 116592 300480 116704
rect -480 110656 240 110768
rect 299760 109928 300480 110040
rect -480 103488 240 103600
rect 299760 103264 300480 103376
rect 299760 96600 300480 96712
rect -480 96376 240 96488
rect 299760 89936 300480 90048
rect -480 89208 240 89320
rect 299760 83272 300480 83384
rect -480 82096 240 82208
rect 299760 76608 300480 76720
rect -480 74928 240 75040
rect 299760 69944 300480 70056
rect -480 67760 240 67872
rect 299760 63280 300480 63392
rect -480 60648 240 60760
rect 299760 56616 300480 56728
rect -480 53480 240 53592
rect 299760 49952 300480 50064
rect -480 46368 240 46480
rect 299760 43288 300480 43400
rect -480 39200 240 39312
rect 299760 36624 300480 36736
rect -480 32088 240 32200
rect 299760 29960 300480 30072
rect -480 24920 240 25032
rect 299760 23296 300480 23408
rect -480 17808 240 17920
rect 299760 16632 300480 16744
rect -480 10640 240 10752
rect 299760 9968 300480 10080
rect -480 3528 240 3640
rect 299760 3304 300480 3416
<< obsm3 >>
rect 240 296718 299838 298158
rect 240 296546 299730 296718
rect 240 296494 299838 296546
rect 270 296322 299838 296494
rect 240 290054 299838 296322
rect 240 289882 299730 290054
rect 240 289326 299838 289882
rect 270 289154 299838 289326
rect 240 283390 299838 289154
rect 240 283218 299730 283390
rect 240 282214 299838 283218
rect 270 282042 299838 282214
rect 240 276726 299838 282042
rect 240 276554 299730 276726
rect 240 275046 299838 276554
rect 270 274874 299838 275046
rect 240 270062 299838 274874
rect 240 269890 299730 270062
rect 240 267934 299838 269890
rect 270 267762 299838 267934
rect 240 263398 299838 267762
rect 240 263226 299730 263398
rect 240 260766 299838 263226
rect 270 260594 299838 260766
rect 240 256734 299838 260594
rect 240 256562 299730 256734
rect 240 253654 299838 256562
rect 270 253482 299838 253654
rect 240 250070 299838 253482
rect 240 249898 299730 250070
rect 240 246486 299838 249898
rect 270 246314 299838 246486
rect 240 243406 299838 246314
rect 240 243234 299730 243406
rect 240 239374 299838 243234
rect 270 239202 299838 239374
rect 240 236742 299838 239202
rect 240 236570 299730 236742
rect 240 232206 299838 236570
rect 270 232034 299838 232206
rect 240 230078 299838 232034
rect 240 229906 299730 230078
rect 240 225038 299838 229906
rect 270 224866 299838 225038
rect 240 223414 299838 224866
rect 240 223242 299730 223414
rect 240 217926 299838 223242
rect 270 217754 299838 217926
rect 240 216750 299838 217754
rect 240 216578 299730 216750
rect 240 210758 299838 216578
rect 270 210586 299838 210758
rect 240 210086 299838 210586
rect 240 209914 299730 210086
rect 240 203646 299838 209914
rect 270 203474 299838 203646
rect 240 203422 299838 203474
rect 240 203250 299730 203422
rect 240 196758 299838 203250
rect 240 196586 299730 196758
rect 240 196478 299838 196586
rect 270 196306 299838 196478
rect 240 190094 299838 196306
rect 240 189922 299730 190094
rect 240 189366 299838 189922
rect 270 189194 299838 189366
rect 240 183430 299838 189194
rect 240 183258 299730 183430
rect 240 182198 299838 183258
rect 270 182026 299838 182198
rect 240 176766 299838 182026
rect 240 176594 299730 176766
rect 240 175086 299838 176594
rect 270 174914 299838 175086
rect 240 170102 299838 174914
rect 240 169930 299730 170102
rect 240 167918 299838 169930
rect 270 167746 299838 167918
rect 240 163438 299838 167746
rect 240 163266 299730 163438
rect 240 160806 299838 163266
rect 270 160634 299838 160806
rect 240 156774 299838 160634
rect 240 156602 299730 156774
rect 240 153638 299838 156602
rect 270 153466 299838 153638
rect 240 150054 299838 153466
rect 240 149882 299730 150054
rect 240 146470 299838 149882
rect 270 146298 299838 146470
rect 240 143390 299838 146298
rect 240 143218 299730 143390
rect 240 139358 299838 143218
rect 270 139186 299838 139358
rect 240 136726 299838 139186
rect 240 136554 299730 136726
rect 240 132190 299838 136554
rect 270 132018 299838 132190
rect 240 130062 299838 132018
rect 240 129890 299730 130062
rect 240 125078 299838 129890
rect 270 124906 299838 125078
rect 240 123398 299838 124906
rect 240 123226 299730 123398
rect 240 117910 299838 123226
rect 270 117738 299838 117910
rect 240 116734 299838 117738
rect 240 116562 299730 116734
rect 240 110798 299838 116562
rect 270 110626 299838 110798
rect 240 110070 299838 110626
rect 240 109898 299730 110070
rect 240 103630 299838 109898
rect 270 103458 299838 103630
rect 240 103406 299838 103458
rect 240 103234 299730 103406
rect 240 96742 299838 103234
rect 240 96570 299730 96742
rect 240 96518 299838 96570
rect 270 96346 299838 96518
rect 240 90078 299838 96346
rect 240 89906 299730 90078
rect 240 89350 299838 89906
rect 270 89178 299838 89350
rect 240 83414 299838 89178
rect 240 83242 299730 83414
rect 240 82238 299838 83242
rect 270 82066 299838 82238
rect 240 76750 299838 82066
rect 240 76578 299730 76750
rect 240 75070 299838 76578
rect 270 74898 299838 75070
rect 240 70086 299838 74898
rect 240 69914 299730 70086
rect 240 67902 299838 69914
rect 270 67730 299838 67902
rect 240 63422 299838 67730
rect 240 63250 299730 63422
rect 240 60790 299838 63250
rect 270 60618 299838 60790
rect 240 56758 299838 60618
rect 240 56586 299730 56758
rect 240 53622 299838 56586
rect 270 53450 299838 53622
rect 240 50094 299838 53450
rect 240 49922 299730 50094
rect 240 46510 299838 49922
rect 270 46338 299838 46510
rect 240 43430 299838 46338
rect 240 43258 299730 43430
rect 240 39342 299838 43258
rect 270 39170 299838 39342
rect 240 36766 299838 39170
rect 240 36594 299730 36766
rect 240 32230 299838 36594
rect 270 32058 299838 32230
rect 240 30102 299838 32058
rect 240 29930 299730 30102
rect 240 25062 299838 29930
rect 270 24890 299838 25062
rect 240 23438 299838 24890
rect 240 23266 299730 23438
rect 240 17950 299838 23266
rect 270 17778 299838 17950
rect 240 16774 299838 17778
rect 240 16602 299730 16774
rect 240 10782 299838 16602
rect 270 10610 299838 10782
rect 240 10110 299838 10610
rect 240 9938 299730 10110
rect 240 3670 299838 9938
rect 270 3498 299838 3670
rect 240 3446 299838 3498
rect 240 3402 299730 3446
<< metal4 >>
rect -1518 -622 -1208 300502
rect -1038 -142 -728 300022
rect 1017 -622 1327 300502
rect 10017 -622 10327 300502
rect 19017 -622 19327 300502
rect 28017 -622 28327 300502
rect 37017 -622 37327 300502
rect 46017 -622 46327 300502
rect 55017 -622 55327 300502
rect 64017 -622 64327 300502
rect 73017 -622 73327 300502
rect 82017 -622 82327 300502
rect 91017 -622 91327 300502
rect 100017 -622 100327 300502
rect 109017 -622 109327 300502
rect 118017 -622 118327 300502
rect 127017 -622 127327 300502
rect 136017 -622 136327 300502
rect 145017 -622 145327 300502
rect 154017 -622 154327 300502
rect 163017 -622 163327 300502
rect 172017 -622 172327 300502
rect 181017 -622 181327 300502
rect 190017 -622 190327 300502
rect 199017 -622 199327 300502
rect 208017 -622 208327 300502
rect 217017 -622 217327 300502
rect 226017 -622 226327 300502
rect 235017 -622 235327 300502
rect 244017 -622 244327 300502
rect 253017 -622 253327 300502
rect 262017 -622 262327 300502
rect 271017 -622 271327 300502
rect 280017 -622 280327 300502
rect 289017 -622 289327 300502
rect 298017 -622 298327 300502
rect 300720 -142 301030 300022
rect 301200 -622 301510 300502
<< metal5 >>
rect -1518 300192 301510 300502
rect -1038 299712 301030 300022
rect -1518 289913 301510 290223
rect -1518 280913 301510 281223
rect -1518 271913 301510 272223
rect -1518 262913 301510 263223
rect -1518 253913 301510 254223
rect -1518 244913 301510 245223
rect -1518 235913 301510 236223
rect -1518 226913 301510 227223
rect -1518 217913 301510 218223
rect -1518 208913 301510 209223
rect -1518 199913 301510 200223
rect -1518 190913 301510 191223
rect -1518 181913 301510 182223
rect -1518 172913 301510 173223
rect -1518 163913 301510 164223
rect -1518 154913 301510 155223
rect -1518 145913 301510 146223
rect -1518 136913 301510 137223
rect -1518 127913 301510 128223
rect -1518 118913 301510 119223
rect -1518 109913 301510 110223
rect -1518 100913 301510 101223
rect -1518 91913 301510 92223
rect -1518 82913 301510 83223
rect -1518 73913 301510 74223
rect -1518 64913 301510 65223
rect -1518 55913 301510 56223
rect -1518 46913 301510 47223
rect -1518 37913 301510 38223
rect -1518 28913 301510 29223
rect -1518 19913 301510 20223
rect -1518 10913 301510 11223
rect -1518 1913 301510 2223
rect -1038 -142 301030 168
rect -1518 -622 301510 -312
<< labels >>
rlabel metal3 s 299760 3304 300480 3416 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 299760 203280 300480 203392 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 299760 223272 300480 223384 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 299760 243264 300480 243376 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 299760 263256 300480 263368 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 299760 283248 300480 283360 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 294392 299760 294504 300480 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 261072 299760 261184 300480 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 227696 299760 227808 300480 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 194376 299760 194488 300480 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 161056 299760 161168 300480 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 299760 23296 300480 23408 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 127680 299760 127792 300480 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 94360 299760 94472 300480 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 61040 299760 61152 300480 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 27664 299760 27776 300480 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s -480 296352 240 296464 4 io_in[24]
port 17 nsew signal input
rlabel metal3 s -480 274904 240 275016 4 io_in[25]
port 18 nsew signal input
rlabel metal3 s -480 253512 240 253624 4 io_in[26]
port 19 nsew signal input
rlabel metal3 s -480 232064 240 232176 4 io_in[27]
port 20 nsew signal input
rlabel metal3 s -480 210616 240 210728 4 io_in[28]
port 21 nsew signal input
rlabel metal3 s -480 189224 240 189336 4 io_in[29]
port 22 nsew signal input
rlabel metal3 s 299760 43288 300480 43400 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s -480 167776 240 167888 4 io_in[30]
port 24 nsew signal input
rlabel metal3 s -480 146328 240 146440 4 io_in[31]
port 25 nsew signal input
rlabel metal3 s -480 124936 240 125048 4 io_in[32]
port 26 nsew signal input
rlabel metal3 s -480 103488 240 103600 4 io_in[33]
port 27 nsew signal input
rlabel metal3 s -480 82096 240 82208 4 io_in[34]
port 28 nsew signal input
rlabel metal3 s -480 60648 240 60760 4 io_in[35]
port 29 nsew signal input
rlabel metal3 s -480 39200 240 39312 4 io_in[36]
port 30 nsew signal input
rlabel metal3 s -480 17808 240 17920 4 io_in[37]
port 31 nsew signal input
rlabel metal3 s 299760 63280 300480 63392 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 299760 83272 300480 83384 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 299760 103264 300480 103376 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 299760 123256 300480 123368 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 299760 143248 300480 143360 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 299760 163296 300480 163408 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 299760 183288 300480 183400 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 299760 16632 300480 16744 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 299760 216608 300480 216720 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 299760 236600 300480 236712 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 299760 256592 300480 256704 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 299760 276584 300480 276696 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 299760 296576 300480 296688 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 272160 299760 272272 300480 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 238840 299760 238952 300480 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 205520 299760 205632 300480 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 172144 299760 172256 300480 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 138824 299760 138936 300480 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 299760 36624 300480 36736 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 105504 299760 105616 300480 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 72128 299760 72240 300480 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 38808 299760 38920 300480 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 5488 299760 5600 300480 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s -480 282072 240 282184 4 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s -480 260624 240 260736 4 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s -480 239232 240 239344 4 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s -480 217784 240 217896 4 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s -480 196336 240 196448 4 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s -480 174944 240 175056 4 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 299760 56616 300480 56728 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s -480 153496 240 153608 4 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s -480 132048 240 132160 4 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s -480 110656 240 110768 4 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s -480 89208 240 89320 4 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s -480 67760 240 67872 4 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s -480 46368 240 46480 4 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s -480 24920 240 25032 4 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s -480 3528 240 3640 4 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 299760 76608 300480 76720 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 299760 96600 300480 96712 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 299760 116592 300480 116704 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 299760 136584 300480 136696 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 299760 156632 300480 156744 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 299760 176624 300480 176736 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 299760 196616 300480 196728 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 299760 9968 300480 10080 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 299760 209944 300480 210056 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 299760 229936 300480 230048 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 299760 249928 300480 250040 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 299760 269920 300480 270032 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 299760 289912 300480 290024 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 283304 299760 283416 300480 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 249928 299760 250040 300480 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 216608 299760 216720 300480 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 183288 299760 183400 300480 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 149912 299760 150024 300480 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 299760 29960 300480 30072 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 116592 299760 116704 300480 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 83272 299760 83384 300480 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 49896 299760 50008 300480 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 16576 299760 16688 300480 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s -480 289184 240 289296 4 io_out[24]
port 93 nsew signal output
rlabel metal3 s -480 267792 240 267904 4 io_out[25]
port 94 nsew signal output
rlabel metal3 s -480 246344 240 246456 4 io_out[26]
port 95 nsew signal output
rlabel metal3 s -480 224896 240 225008 4 io_out[27]
port 96 nsew signal output
rlabel metal3 s -480 203504 240 203616 4 io_out[28]
port 97 nsew signal output
rlabel metal3 s -480 182056 240 182168 4 io_out[29]
port 98 nsew signal output
rlabel metal3 s 299760 49952 300480 50064 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s -480 160664 240 160776 4 io_out[30]
port 100 nsew signal output
rlabel metal3 s -480 139216 240 139328 4 io_out[31]
port 101 nsew signal output
rlabel metal3 s -480 117768 240 117880 4 io_out[32]
port 102 nsew signal output
rlabel metal3 s -480 96376 240 96488 4 io_out[33]
port 103 nsew signal output
rlabel metal3 s -480 74928 240 75040 4 io_out[34]
port 104 nsew signal output
rlabel metal3 s -480 53480 240 53592 4 io_out[35]
port 105 nsew signal output
rlabel metal3 s -480 32088 240 32200 4 io_out[36]
port 106 nsew signal output
rlabel metal3 s -480 10640 240 10752 4 io_out[37]
port 107 nsew signal output
rlabel metal3 s 299760 69944 300480 70056 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 299760 89936 300480 90048 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 299760 109928 300480 110040 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 299760 129920 300480 130032 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 299760 149912 300480 150024 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 299760 169960 300480 170072 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 299760 189952 300480 190064 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 105672 -480 105784 240 8 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 135464 -480 135576 240 8 la_data_in[10]
port 116 nsew signal input
rlabel metal2 s 138488 -480 138600 240 8 la_data_in[11]
port 117 nsew signal input
rlabel metal2 s 141456 -480 141568 240 8 la_data_in[12]
port 118 nsew signal input
rlabel metal2 s 144424 -480 144536 240 8 la_data_in[13]
port 119 nsew signal input
rlabel metal2 s 147392 -480 147504 240 8 la_data_in[14]
port 120 nsew signal input
rlabel metal2 s 150416 -480 150528 240 8 la_data_in[15]
port 121 nsew signal input
rlabel metal2 s 153384 -480 153496 240 8 la_data_in[16]
port 122 nsew signal input
rlabel metal2 s 156352 -480 156464 240 8 la_data_in[17]
port 123 nsew signal input
rlabel metal2 s 159320 -480 159432 240 8 la_data_in[18]
port 124 nsew signal input
rlabel metal2 s 162288 -480 162400 240 8 la_data_in[19]
port 125 nsew signal input
rlabel metal2 s 108640 -480 108752 240 8 la_data_in[1]
port 126 nsew signal input
rlabel metal2 s 165312 -480 165424 240 8 la_data_in[20]
port 127 nsew signal input
rlabel metal2 s 168280 -480 168392 240 8 la_data_in[21]
port 128 nsew signal input
rlabel metal2 s 171248 -480 171360 240 8 la_data_in[22]
port 129 nsew signal input
rlabel metal2 s 174216 -480 174328 240 8 la_data_in[23]
port 130 nsew signal input
rlabel metal2 s 177240 -480 177352 240 8 la_data_in[24]
port 131 nsew signal input
rlabel metal2 s 180208 -480 180320 240 8 la_data_in[25]
port 132 nsew signal input
rlabel metal2 s 183176 -480 183288 240 8 la_data_in[26]
port 133 nsew signal input
rlabel metal2 s 186144 -480 186256 240 8 la_data_in[27]
port 134 nsew signal input
rlabel metal2 s 189112 -480 189224 240 8 la_data_in[28]
port 135 nsew signal input
rlabel metal2 s 192136 -480 192248 240 8 la_data_in[29]
port 136 nsew signal input
rlabel metal2 s 111664 -480 111776 240 8 la_data_in[2]
port 137 nsew signal input
rlabel metal2 s 195104 -480 195216 240 8 la_data_in[30]
port 138 nsew signal input
rlabel metal2 s 198072 -480 198184 240 8 la_data_in[31]
port 139 nsew signal input
rlabel metal2 s 201040 -480 201152 240 8 la_data_in[32]
port 140 nsew signal input
rlabel metal2 s 204064 -480 204176 240 8 la_data_in[33]
port 141 nsew signal input
rlabel metal2 s 207032 -480 207144 240 8 la_data_in[34]
port 142 nsew signal input
rlabel metal2 s 210000 -480 210112 240 8 la_data_in[35]
port 143 nsew signal input
rlabel metal2 s 212968 -480 213080 240 8 la_data_in[36]
port 144 nsew signal input
rlabel metal2 s 215936 -480 216048 240 8 la_data_in[37]
port 145 nsew signal input
rlabel metal2 s 218960 -480 219072 240 8 la_data_in[38]
port 146 nsew signal input
rlabel metal2 s 221928 -480 222040 240 8 la_data_in[39]
port 147 nsew signal input
rlabel metal2 s 114632 -480 114744 240 8 la_data_in[3]
port 148 nsew signal input
rlabel metal2 s 224896 -480 225008 240 8 la_data_in[40]
port 149 nsew signal input
rlabel metal2 s 227864 -480 227976 240 8 la_data_in[41]
port 150 nsew signal input
rlabel metal2 s 230888 -480 231000 240 8 la_data_in[42]
port 151 nsew signal input
rlabel metal2 s 233856 -480 233968 240 8 la_data_in[43]
port 152 nsew signal input
rlabel metal2 s 236824 -480 236936 240 8 la_data_in[44]
port 153 nsew signal input
rlabel metal2 s 239792 -480 239904 240 8 la_data_in[45]
port 154 nsew signal input
rlabel metal2 s 242760 -480 242872 240 8 la_data_in[46]
port 155 nsew signal input
rlabel metal2 s 245784 -480 245896 240 8 la_data_in[47]
port 156 nsew signal input
rlabel metal2 s 248752 -480 248864 240 8 la_data_in[48]
port 157 nsew signal input
rlabel metal2 s 251720 -480 251832 240 8 la_data_in[49]
port 158 nsew signal input
rlabel metal2 s 117600 -480 117712 240 8 la_data_in[4]
port 159 nsew signal input
rlabel metal2 s 254688 -480 254800 240 8 la_data_in[50]
port 160 nsew signal input
rlabel metal2 s 257712 -480 257824 240 8 la_data_in[51]
port 161 nsew signal input
rlabel metal2 s 260680 -480 260792 240 8 la_data_in[52]
port 162 nsew signal input
rlabel metal2 s 263648 -480 263760 240 8 la_data_in[53]
port 163 nsew signal input
rlabel metal2 s 266616 -480 266728 240 8 la_data_in[54]
port 164 nsew signal input
rlabel metal2 s 269640 -480 269752 240 8 la_data_in[55]
port 165 nsew signal input
rlabel metal2 s 272608 -480 272720 240 8 la_data_in[56]
port 166 nsew signal input
rlabel metal2 s 275576 -480 275688 240 8 la_data_in[57]
port 167 nsew signal input
rlabel metal2 s 278544 -480 278656 240 8 la_data_in[58]
port 168 nsew signal input
rlabel metal2 s 281512 -480 281624 240 8 la_data_in[59]
port 169 nsew signal input
rlabel metal2 s 120568 -480 120680 240 8 la_data_in[5]
port 170 nsew signal input
rlabel metal2 s 284536 -480 284648 240 8 la_data_in[60]
port 171 nsew signal input
rlabel metal2 s 287504 -480 287616 240 8 la_data_in[61]
port 172 nsew signal input
rlabel metal2 s 290472 -480 290584 240 8 la_data_in[62]
port 173 nsew signal input
rlabel metal2 s 293440 -480 293552 240 8 la_data_in[63]
port 174 nsew signal input
rlabel metal2 s 123536 -480 123648 240 8 la_data_in[6]
port 175 nsew signal input
rlabel metal2 s 126560 -480 126672 240 8 la_data_in[7]
port 176 nsew signal input
rlabel metal2 s 129528 -480 129640 240 8 la_data_in[8]
port 177 nsew signal input
rlabel metal2 s 132496 -480 132608 240 8 la_data_in[9]
port 178 nsew signal input
rlabel metal2 s 106680 -480 106792 240 8 la_data_out[0]
port 179 nsew signal output
rlabel metal2 s 136472 -480 136584 240 8 la_data_out[10]
port 180 nsew signal output
rlabel metal2 s 139440 -480 139552 240 8 la_data_out[11]
port 181 nsew signal output
rlabel metal2 s 142464 -480 142576 240 8 la_data_out[12]
port 182 nsew signal output
rlabel metal2 s 145432 -480 145544 240 8 la_data_out[13]
port 183 nsew signal output
rlabel metal2 s 148400 -480 148512 240 8 la_data_out[14]
port 184 nsew signal output
rlabel metal2 s 151368 -480 151480 240 8 la_data_out[15]
port 185 nsew signal output
rlabel metal2 s 154336 -480 154448 240 8 la_data_out[16]
port 186 nsew signal output
rlabel metal2 s 157360 -480 157472 240 8 la_data_out[17]
port 187 nsew signal output
rlabel metal2 s 160328 -480 160440 240 8 la_data_out[18]
port 188 nsew signal output
rlabel metal2 s 163296 -480 163408 240 8 la_data_out[19]
port 189 nsew signal output
rlabel metal2 s 109648 -480 109760 240 8 la_data_out[1]
port 190 nsew signal output
rlabel metal2 s 166264 -480 166376 240 8 la_data_out[20]
port 191 nsew signal output
rlabel metal2 s 169288 -480 169400 240 8 la_data_out[21]
port 192 nsew signal output
rlabel metal2 s 172256 -480 172368 240 8 la_data_out[22]
port 193 nsew signal output
rlabel metal2 s 175224 -480 175336 240 8 la_data_out[23]
port 194 nsew signal output
rlabel metal2 s 178192 -480 178304 240 8 la_data_out[24]
port 195 nsew signal output
rlabel metal2 s 181160 -480 181272 240 8 la_data_out[25]
port 196 nsew signal output
rlabel metal2 s 184184 -480 184296 240 8 la_data_out[26]
port 197 nsew signal output
rlabel metal2 s 187152 -480 187264 240 8 la_data_out[27]
port 198 nsew signal output
rlabel metal2 s 190120 -480 190232 240 8 la_data_out[28]
port 199 nsew signal output
rlabel metal2 s 193088 -480 193200 240 8 la_data_out[29]
port 200 nsew signal output
rlabel metal2 s 112616 -480 112728 240 8 la_data_out[2]
port 201 nsew signal output
rlabel metal2 s 196112 -480 196224 240 8 la_data_out[30]
port 202 nsew signal output
rlabel metal2 s 199080 -480 199192 240 8 la_data_out[31]
port 203 nsew signal output
rlabel metal2 s 202048 -480 202160 240 8 la_data_out[32]
port 204 nsew signal output
rlabel metal2 s 205016 -480 205128 240 8 la_data_out[33]
port 205 nsew signal output
rlabel metal2 s 208040 -480 208152 240 8 la_data_out[34]
port 206 nsew signal output
rlabel metal2 s 211008 -480 211120 240 8 la_data_out[35]
port 207 nsew signal output
rlabel metal2 s 213976 -480 214088 240 8 la_data_out[36]
port 208 nsew signal output
rlabel metal2 s 216944 -480 217056 240 8 la_data_out[37]
port 209 nsew signal output
rlabel metal2 s 219912 -480 220024 240 8 la_data_out[38]
port 210 nsew signal output
rlabel metal2 s 222936 -480 223048 240 8 la_data_out[39]
port 211 nsew signal output
rlabel metal2 s 115640 -480 115752 240 8 la_data_out[3]
port 212 nsew signal output
rlabel metal2 s 225904 -480 226016 240 8 la_data_out[40]
port 213 nsew signal output
rlabel metal2 s 228872 -480 228984 240 8 la_data_out[41]
port 214 nsew signal output
rlabel metal2 s 231840 -480 231952 240 8 la_data_out[42]
port 215 nsew signal output
rlabel metal2 s 234864 -480 234976 240 8 la_data_out[43]
port 216 nsew signal output
rlabel metal2 s 237832 -480 237944 240 8 la_data_out[44]
port 217 nsew signal output
rlabel metal2 s 240800 -480 240912 240 8 la_data_out[45]
port 218 nsew signal output
rlabel metal2 s 243768 -480 243880 240 8 la_data_out[46]
port 219 nsew signal output
rlabel metal2 s 246736 -480 246848 240 8 la_data_out[47]
port 220 nsew signal output
rlabel metal2 s 249760 -480 249872 240 8 la_data_out[48]
port 221 nsew signal output
rlabel metal2 s 252728 -480 252840 240 8 la_data_out[49]
port 222 nsew signal output
rlabel metal2 s 118608 -480 118720 240 8 la_data_out[4]
port 223 nsew signal output
rlabel metal2 s 255696 -480 255808 240 8 la_data_out[50]
port 224 nsew signal output
rlabel metal2 s 258664 -480 258776 240 8 la_data_out[51]
port 225 nsew signal output
rlabel metal2 s 261688 -480 261800 240 8 la_data_out[52]
port 226 nsew signal output
rlabel metal2 s 264656 -480 264768 240 8 la_data_out[53]
port 227 nsew signal output
rlabel metal2 s 267624 -480 267736 240 8 la_data_out[54]
port 228 nsew signal output
rlabel metal2 s 270592 -480 270704 240 8 la_data_out[55]
port 229 nsew signal output
rlabel metal2 s 273560 -480 273672 240 8 la_data_out[56]
port 230 nsew signal output
rlabel metal2 s 276584 -480 276696 240 8 la_data_out[57]
port 231 nsew signal output
rlabel metal2 s 279552 -480 279664 240 8 la_data_out[58]
port 232 nsew signal output
rlabel metal2 s 282520 -480 282632 240 8 la_data_out[59]
port 233 nsew signal output
rlabel metal2 s 121576 -480 121688 240 8 la_data_out[5]
port 234 nsew signal output
rlabel metal2 s 285488 -480 285600 240 8 la_data_out[60]
port 235 nsew signal output
rlabel metal2 s 288512 -480 288624 240 8 la_data_out[61]
port 236 nsew signal output
rlabel metal2 s 291480 -480 291592 240 8 la_data_out[62]
port 237 nsew signal output
rlabel metal2 s 294448 -480 294560 240 8 la_data_out[63]
port 238 nsew signal output
rlabel metal2 s 124544 -480 124656 240 8 la_data_out[6]
port 239 nsew signal output
rlabel metal2 s 127512 -480 127624 240 8 la_data_out[7]
port 240 nsew signal output
rlabel metal2 s 130536 -480 130648 240 8 la_data_out[8]
port 241 nsew signal output
rlabel metal2 s 133504 -480 133616 240 8 la_data_out[9]
port 242 nsew signal output
rlabel metal2 s 107688 -480 107800 240 8 la_oenb[0]
port 243 nsew signal input
rlabel metal2 s 137480 -480 137592 240 8 la_oenb[10]
port 244 nsew signal input
rlabel metal2 s 140448 -480 140560 240 8 la_oenb[11]
port 245 nsew signal input
rlabel metal2 s 143416 -480 143528 240 8 la_oenb[12]
port 246 nsew signal input
rlabel metal2 s 146440 -480 146552 240 8 la_oenb[13]
port 247 nsew signal input
rlabel metal2 s 149408 -480 149520 240 8 la_oenb[14]
port 248 nsew signal input
rlabel metal2 s 152376 -480 152488 240 8 la_oenb[15]
port 249 nsew signal input
rlabel metal2 s 155344 -480 155456 240 8 la_oenb[16]
port 250 nsew signal input
rlabel metal2 s 158312 -480 158424 240 8 la_oenb[17]
port 251 nsew signal input
rlabel metal2 s 161336 -480 161448 240 8 la_oenb[18]
port 252 nsew signal input
rlabel metal2 s 164304 -480 164416 240 8 la_oenb[19]
port 253 nsew signal input
rlabel metal2 s 110656 -480 110768 240 8 la_oenb[1]
port 254 nsew signal input
rlabel metal2 s 167272 -480 167384 240 8 la_oenb[20]
port 255 nsew signal input
rlabel metal2 s 170240 -480 170352 240 8 la_oenb[21]
port 256 nsew signal input
rlabel metal2 s 173264 -480 173376 240 8 la_oenb[22]
port 257 nsew signal input
rlabel metal2 s 176232 -480 176344 240 8 la_oenb[23]
port 258 nsew signal input
rlabel metal2 s 179200 -480 179312 240 8 la_oenb[24]
port 259 nsew signal input
rlabel metal2 s 182168 -480 182280 240 8 la_oenb[25]
port 260 nsew signal input
rlabel metal2 s 185136 -480 185248 240 8 la_oenb[26]
port 261 nsew signal input
rlabel metal2 s 188160 -480 188272 240 8 la_oenb[27]
port 262 nsew signal input
rlabel metal2 s 191128 -480 191240 240 8 la_oenb[28]
port 263 nsew signal input
rlabel metal2 s 194096 -480 194208 240 8 la_oenb[29]
port 264 nsew signal input
rlabel metal2 s 113624 -480 113736 240 8 la_oenb[2]
port 265 nsew signal input
rlabel metal2 s 197064 -480 197176 240 8 la_oenb[30]
port 266 nsew signal input
rlabel metal2 s 200088 -480 200200 240 8 la_oenb[31]
port 267 nsew signal input
rlabel metal2 s 203056 -480 203168 240 8 la_oenb[32]
port 268 nsew signal input
rlabel metal2 s 206024 -480 206136 240 8 la_oenb[33]
port 269 nsew signal input
rlabel metal2 s 208992 -480 209104 240 8 la_oenb[34]
port 270 nsew signal input
rlabel metal2 s 211960 -480 212072 240 8 la_oenb[35]
port 271 nsew signal input
rlabel metal2 s 214984 -480 215096 240 8 la_oenb[36]
port 272 nsew signal input
rlabel metal2 s 217952 -480 218064 240 8 la_oenb[37]
port 273 nsew signal input
rlabel metal2 s 220920 -480 221032 240 8 la_oenb[38]
port 274 nsew signal input
rlabel metal2 s 223888 -480 224000 240 8 la_oenb[39]
port 275 nsew signal input
rlabel metal2 s 116592 -480 116704 240 8 la_oenb[3]
port 276 nsew signal input
rlabel metal2 s 226912 -480 227024 240 8 la_oenb[40]
port 277 nsew signal input
rlabel metal2 s 229880 -480 229992 240 8 la_oenb[41]
port 278 nsew signal input
rlabel metal2 s 232848 -480 232960 240 8 la_oenb[42]
port 279 nsew signal input
rlabel metal2 s 235816 -480 235928 240 8 la_oenb[43]
port 280 nsew signal input
rlabel metal2 s 238840 -480 238952 240 8 la_oenb[44]
port 281 nsew signal input
rlabel metal2 s 241808 -480 241920 240 8 la_oenb[45]
port 282 nsew signal input
rlabel metal2 s 244776 -480 244888 240 8 la_oenb[46]
port 283 nsew signal input
rlabel metal2 s 247744 -480 247856 240 8 la_oenb[47]
port 284 nsew signal input
rlabel metal2 s 250712 -480 250824 240 8 la_oenb[48]
port 285 nsew signal input
rlabel metal2 s 253736 -480 253848 240 8 la_oenb[49]
port 286 nsew signal input
rlabel metal2 s 119616 -480 119728 240 8 la_oenb[4]
port 287 nsew signal input
rlabel metal2 s 256704 -480 256816 240 8 la_oenb[50]
port 288 nsew signal input
rlabel metal2 s 259672 -480 259784 240 8 la_oenb[51]
port 289 nsew signal input
rlabel metal2 s 262640 -480 262752 240 8 la_oenb[52]
port 290 nsew signal input
rlabel metal2 s 265664 -480 265776 240 8 la_oenb[53]
port 291 nsew signal input
rlabel metal2 s 268632 -480 268744 240 8 la_oenb[54]
port 292 nsew signal input
rlabel metal2 s 271600 -480 271712 240 8 la_oenb[55]
port 293 nsew signal input
rlabel metal2 s 274568 -480 274680 240 8 la_oenb[56]
port 294 nsew signal input
rlabel metal2 s 277536 -480 277648 240 8 la_oenb[57]
port 295 nsew signal input
rlabel metal2 s 280560 -480 280672 240 8 la_oenb[58]
port 296 nsew signal input
rlabel metal2 s 283528 -480 283640 240 8 la_oenb[59]
port 297 nsew signal input
rlabel metal2 s 122584 -480 122696 240 8 la_oenb[5]
port 298 nsew signal input
rlabel metal2 s 286496 -480 286608 240 8 la_oenb[60]
port 299 nsew signal input
rlabel metal2 s 289464 -480 289576 240 8 la_oenb[61]
port 300 nsew signal input
rlabel metal2 s 292488 -480 292600 240 8 la_oenb[62]
port 301 nsew signal input
rlabel metal2 s 295456 -480 295568 240 8 la_oenb[63]
port 302 nsew signal input
rlabel metal2 s 125552 -480 125664 240 8 la_oenb[6]
port 303 nsew signal input
rlabel metal2 s 128520 -480 128632 240 8 la_oenb[7]
port 304 nsew signal input
rlabel metal2 s 131488 -480 131600 240 8 la_oenb[8]
port 305 nsew signal input
rlabel metal2 s 134512 -480 134624 240 8 la_oenb[9]
port 306 nsew signal input
rlabel metal2 s 296464 -480 296576 240 8 user_clock2
port 307 nsew signal input
rlabel metal2 s 297416 -480 297528 240 8 user_irq[0]
port 308 nsew signal output
rlabel metal2 s 298424 -480 298536 240 8 user_irq[1]
port 309 nsew signal output
rlabel metal2 s 299432 -480 299544 240 8 user_irq[2]
port 310 nsew signal output
rlabel metal4 s -1038 -142 -728 300022 4 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1038 -142 301030 168 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1038 299712 301030 300022 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 300720 -142 301030 300022 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 1017 -622 1327 300502 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 19017 -622 19327 300502 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 37017 -622 37327 300502 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 55017 -622 55327 300502 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 73017 -622 73327 300502 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 91017 -622 91327 300502 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 109017 -622 109327 300502 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 127017 -622 127327 300502 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 145017 -622 145327 300502 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 163017 -622 163327 300502 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 181017 -622 181327 300502 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 199017 -622 199327 300502 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 217017 -622 217327 300502 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 235017 -622 235327 300502 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 253017 -622 253327 300502 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 271017 -622 271327 300502 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 289017 -622 289327 300502 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1518 1913 301510 2223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1518 19913 301510 20223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1518 37913 301510 38223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1518 55913 301510 56223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1518 73913 301510 74223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1518 91913 301510 92223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1518 109913 301510 110223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1518 127913 301510 128223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1518 145913 301510 146223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1518 163913 301510 164223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1518 181913 301510 182223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1518 199913 301510 200223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1518 217913 301510 218223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1518 235913 301510 236223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1518 253913 301510 254223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1518 271913 301510 272223 6 vdd
port 311 nsew power bidirectional
rlabel metal5 s -1518 289913 301510 290223 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s -1518 -622 -1208 300502 4 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 -622 301510 -312 8 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 300192 301510 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 301200 -622 301510 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 10017 -622 10327 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 28017 -622 28327 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 46017 -622 46327 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 64017 -622 64327 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 82017 -622 82327 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 100017 -622 100327 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 118017 -622 118327 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 136017 -622 136327 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 154017 -622 154327 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 172017 -622 172327 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 190017 -622 190327 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 208017 -622 208327 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 226017 -622 226327 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 244017 -622 244327 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 262017 -622 262327 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 280017 -622 280327 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 298017 -622 298327 300502 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 10913 301510 11223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 28913 301510 29223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 46913 301510 47223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 64913 301510 65223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 82913 301510 83223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 100913 301510 101223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 118913 301510 119223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 136913 301510 137223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 154913 301510 155223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 172913 301510 173223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 190913 301510 191223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 208913 301510 209223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 226913 301510 227223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 244913 301510 245223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 262913 301510 263223 6 vss
port 312 nsew ground bidirectional
rlabel metal5 s -1518 280913 301510 281223 6 vss
port 312 nsew ground bidirectional
rlabel metal2 s 392 -480 504 240 8 wb_clk_i
port 313 nsew signal input
rlabel metal2 s 1344 -480 1456 240 8 wb_rst_i
port 314 nsew signal input
rlabel metal2 s 2352 -480 2464 240 8 wbs_ack_o
port 315 nsew signal output
rlabel metal2 s 6328 -480 6440 240 8 wbs_adr_i[0]
port 316 nsew signal input
rlabel metal2 s 40096 -480 40208 240 8 wbs_adr_i[10]
port 317 nsew signal input
rlabel metal2 s 43064 -480 43176 240 8 wbs_adr_i[11]
port 318 nsew signal input
rlabel metal2 s 46088 -480 46200 240 8 wbs_adr_i[12]
port 319 nsew signal input
rlabel metal2 s 49056 -480 49168 240 8 wbs_adr_i[13]
port 320 nsew signal input
rlabel metal2 s 52024 -480 52136 240 8 wbs_adr_i[14]
port 321 nsew signal input
rlabel metal2 s 54992 -480 55104 240 8 wbs_adr_i[15]
port 322 nsew signal input
rlabel metal2 s 58016 -480 58128 240 8 wbs_adr_i[16]
port 323 nsew signal input
rlabel metal2 s 60984 -480 61096 240 8 wbs_adr_i[17]
port 324 nsew signal input
rlabel metal2 s 63952 -480 64064 240 8 wbs_adr_i[18]
port 325 nsew signal input
rlabel metal2 s 66920 -480 67032 240 8 wbs_adr_i[19]
port 326 nsew signal input
rlabel metal2 s 10304 -480 10416 240 8 wbs_adr_i[1]
port 327 nsew signal input
rlabel metal2 s 69888 -480 70000 240 8 wbs_adr_i[20]
port 328 nsew signal input
rlabel metal2 s 72912 -480 73024 240 8 wbs_adr_i[21]
port 329 nsew signal input
rlabel metal2 s 75880 -480 75992 240 8 wbs_adr_i[22]
port 330 nsew signal input
rlabel metal2 s 78848 -480 78960 240 8 wbs_adr_i[23]
port 331 nsew signal input
rlabel metal2 s 81816 -480 81928 240 8 wbs_adr_i[24]
port 332 nsew signal input
rlabel metal2 s 84840 -480 84952 240 8 wbs_adr_i[25]
port 333 nsew signal input
rlabel metal2 s 87808 -480 87920 240 8 wbs_adr_i[26]
port 334 nsew signal input
rlabel metal2 s 90776 -480 90888 240 8 wbs_adr_i[27]
port 335 nsew signal input
rlabel metal2 s 93744 -480 93856 240 8 wbs_adr_i[28]
port 336 nsew signal input
rlabel metal2 s 96712 -480 96824 240 8 wbs_adr_i[29]
port 337 nsew signal input
rlabel metal2 s 14280 -480 14392 240 8 wbs_adr_i[2]
port 338 nsew signal input
rlabel metal2 s 99736 -480 99848 240 8 wbs_adr_i[30]
port 339 nsew signal input
rlabel metal2 s 102704 -480 102816 240 8 wbs_adr_i[31]
port 340 nsew signal input
rlabel metal2 s 18256 -480 18368 240 8 wbs_adr_i[3]
port 341 nsew signal input
rlabel metal2 s 22232 -480 22344 240 8 wbs_adr_i[4]
port 342 nsew signal input
rlabel metal2 s 25200 -480 25312 240 8 wbs_adr_i[5]
port 343 nsew signal input
rlabel metal2 s 28168 -480 28280 240 8 wbs_adr_i[6]
port 344 nsew signal input
rlabel metal2 s 31136 -480 31248 240 8 wbs_adr_i[7]
port 345 nsew signal input
rlabel metal2 s 34160 -480 34272 240 8 wbs_adr_i[8]
port 346 nsew signal input
rlabel metal2 s 37128 -480 37240 240 8 wbs_adr_i[9]
port 347 nsew signal input
rlabel metal2 s 3360 -480 3472 240 8 wbs_cyc_i
port 348 nsew signal input
rlabel metal2 s 7336 -480 7448 240 8 wbs_dat_i[0]
port 349 nsew signal input
rlabel metal2 s 41104 -480 41216 240 8 wbs_dat_i[10]
port 350 nsew signal input
rlabel metal2 s 44072 -480 44184 240 8 wbs_dat_i[11]
port 351 nsew signal input
rlabel metal2 s 47040 -480 47152 240 8 wbs_dat_i[12]
port 352 nsew signal input
rlabel metal2 s 50064 -480 50176 240 8 wbs_dat_i[13]
port 353 nsew signal input
rlabel metal2 s 53032 -480 53144 240 8 wbs_dat_i[14]
port 354 nsew signal input
rlabel metal2 s 56000 -480 56112 240 8 wbs_dat_i[15]
port 355 nsew signal input
rlabel metal2 s 58968 -480 59080 240 8 wbs_dat_i[16]
port 356 nsew signal input
rlabel metal2 s 61936 -480 62048 240 8 wbs_dat_i[17]
port 357 nsew signal input
rlabel metal2 s 64960 -480 65072 240 8 wbs_dat_i[18]
port 358 nsew signal input
rlabel metal2 s 67928 -480 68040 240 8 wbs_dat_i[19]
port 359 nsew signal input
rlabel metal2 s 11312 -480 11424 240 8 wbs_dat_i[1]
port 360 nsew signal input
rlabel metal2 s 70896 -480 71008 240 8 wbs_dat_i[20]
port 361 nsew signal input
rlabel metal2 s 73864 -480 73976 240 8 wbs_dat_i[21]
port 362 nsew signal input
rlabel metal2 s 76888 -480 77000 240 8 wbs_dat_i[22]
port 363 nsew signal input
rlabel metal2 s 79856 -480 79968 240 8 wbs_dat_i[23]
port 364 nsew signal input
rlabel metal2 s 82824 -480 82936 240 8 wbs_dat_i[24]
port 365 nsew signal input
rlabel metal2 s 85792 -480 85904 240 8 wbs_dat_i[25]
port 366 nsew signal input
rlabel metal2 s 88816 -480 88928 240 8 wbs_dat_i[26]
port 367 nsew signal input
rlabel metal2 s 91784 -480 91896 240 8 wbs_dat_i[27]
port 368 nsew signal input
rlabel metal2 s 94752 -480 94864 240 8 wbs_dat_i[28]
port 369 nsew signal input
rlabel metal2 s 97720 -480 97832 240 8 wbs_dat_i[29]
port 370 nsew signal input
rlabel metal2 s 15288 -480 15400 240 8 wbs_dat_i[2]
port 371 nsew signal input
rlabel metal2 s 100688 -480 100800 240 8 wbs_dat_i[30]
port 372 nsew signal input
rlabel metal2 s 103712 -480 103824 240 8 wbs_dat_i[31]
port 373 nsew signal input
rlabel metal2 s 19264 -480 19376 240 8 wbs_dat_i[3]
port 374 nsew signal input
rlabel metal2 s 23240 -480 23352 240 8 wbs_dat_i[4]
port 375 nsew signal input
rlabel metal2 s 26208 -480 26320 240 8 wbs_dat_i[5]
port 376 nsew signal input
rlabel metal2 s 29176 -480 29288 240 8 wbs_dat_i[6]
port 377 nsew signal input
rlabel metal2 s 32144 -480 32256 240 8 wbs_dat_i[7]
port 378 nsew signal input
rlabel metal2 s 35112 -480 35224 240 8 wbs_dat_i[8]
port 379 nsew signal input
rlabel metal2 s 38136 -480 38248 240 8 wbs_dat_i[9]
port 380 nsew signal input
rlabel metal2 s 8288 -480 8400 240 8 wbs_dat_o[0]
port 381 nsew signal output
rlabel metal2 s 42112 -480 42224 240 8 wbs_dat_o[10]
port 382 nsew signal output
rlabel metal2 s 45080 -480 45192 240 8 wbs_dat_o[11]
port 383 nsew signal output
rlabel metal2 s 48048 -480 48160 240 8 wbs_dat_o[12]
port 384 nsew signal output
rlabel metal2 s 51016 -480 51128 240 8 wbs_dat_o[13]
port 385 nsew signal output
rlabel metal2 s 54040 -480 54152 240 8 wbs_dat_o[14]
port 386 nsew signal output
rlabel metal2 s 57008 -480 57120 240 8 wbs_dat_o[15]
port 387 nsew signal output
rlabel metal2 s 59976 -480 60088 240 8 wbs_dat_o[16]
port 388 nsew signal output
rlabel metal2 s 62944 -480 63056 240 8 wbs_dat_o[17]
port 389 nsew signal output
rlabel metal2 s 65912 -480 66024 240 8 wbs_dat_o[18]
port 390 nsew signal output
rlabel metal2 s 68936 -480 69048 240 8 wbs_dat_o[19]
port 391 nsew signal output
rlabel metal2 s 12264 -480 12376 240 8 wbs_dat_o[1]
port 392 nsew signal output
rlabel metal2 s 71904 -480 72016 240 8 wbs_dat_o[20]
port 393 nsew signal output
rlabel metal2 s 74872 -480 74984 240 8 wbs_dat_o[21]
port 394 nsew signal output
rlabel metal2 s 77840 -480 77952 240 8 wbs_dat_o[22]
port 395 nsew signal output
rlabel metal2 s 80864 -480 80976 240 8 wbs_dat_o[23]
port 396 nsew signal output
rlabel metal2 s 83832 -480 83944 240 8 wbs_dat_o[24]
port 397 nsew signal output
rlabel metal2 s 86800 -480 86912 240 8 wbs_dat_o[25]
port 398 nsew signal output
rlabel metal2 s 89768 -480 89880 240 8 wbs_dat_o[26]
port 399 nsew signal output
rlabel metal2 s 92736 -480 92848 240 8 wbs_dat_o[27]
port 400 nsew signal output
rlabel metal2 s 95760 -480 95872 240 8 wbs_dat_o[28]
port 401 nsew signal output
rlabel metal2 s 98728 -480 98840 240 8 wbs_dat_o[29]
port 402 nsew signal output
rlabel metal2 s 16240 -480 16352 240 8 wbs_dat_o[2]
port 403 nsew signal output
rlabel metal2 s 101696 -480 101808 240 8 wbs_dat_o[30]
port 404 nsew signal output
rlabel metal2 s 104664 -480 104776 240 8 wbs_dat_o[31]
port 405 nsew signal output
rlabel metal2 s 20216 -480 20328 240 8 wbs_dat_o[3]
port 406 nsew signal output
rlabel metal2 s 24192 -480 24304 240 8 wbs_dat_o[4]
port 407 nsew signal output
rlabel metal2 s 27216 -480 27328 240 8 wbs_dat_o[5]
port 408 nsew signal output
rlabel metal2 s 30184 -480 30296 240 8 wbs_dat_o[6]
port 409 nsew signal output
rlabel metal2 s 33152 -480 33264 240 8 wbs_dat_o[7]
port 410 nsew signal output
rlabel metal2 s 36120 -480 36232 240 8 wbs_dat_o[8]
port 411 nsew signal output
rlabel metal2 s 39088 -480 39200 240 8 wbs_dat_o[9]
port 412 nsew signal output
rlabel metal2 s 9296 -480 9408 240 8 wbs_sel_i[0]
port 413 nsew signal input
rlabel metal2 s 13272 -480 13384 240 8 wbs_sel_i[1]
port 414 nsew signal input
rlabel metal2 s 17248 -480 17360 240 8 wbs_sel_i[2]
port 415 nsew signal input
rlabel metal2 s 21224 -480 21336 240 8 wbs_sel_i[3]
port 416 nsew signal input
rlabel metal2 s 4312 -480 4424 240 8 wbs_stb_i
port 417 nsew signal input
rlabel metal2 s 5320 -480 5432 240 8 wbs_we_i
port 418 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 300000 300000
string GDS_END 17415220
string GDS_FILE ../gds/user_project_wrapper.gds.gz
string GDS_START 53688
string LEFclass BLOCK
string LEFview TRUE
<< end >>
