* NGSPICE file created from housekeeping.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_4 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_4 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_4 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_4 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 D RN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 D SETN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

.subckt housekeeping VDD VSS debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oe
+ pad_flash_csb pad_flash_csb_oe pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ie
+ pad_flash_io0_oe pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ie pad_flash_io1_oe
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out qspi_enabled reset
+ ser_rx ser_tx serial_clock serial_data_1 serial_data_2 serial_load serial_resetn
+ spi_csb spi_enabled spi_sck spi_sdi spi_sdo spi_sdoenb spimemio_flash_clk spimemio_flash_csb
+ spimemio_flash_io0_di spimemio_flash_io0_do spimemio_flash_io0_oeb spimemio_flash_io1_di
+ spimemio_flash_io1_do spimemio_flash_io1_oeb spimemio_flash_io2_di spimemio_flash_io2_do
+ spimemio_flash_io2_oeb spimemio_flash_io3_di spimemio_flash_io3_do spimemio_flash_io3_oeb
+ trap uart_enabled user_clock wb_ack_o wb_adr_i[0] wb_adr_i[10] wb_adr_i[11] wb_adr_i[12]
+ wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17] wb_adr_i[18] wb_adr_i[19]
+ wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23] wb_adr_i[24] wb_adr_i[25]
+ wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2] wb_adr_i[30] wb_adr_i[31]
+ wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7] wb_adr_i[8] wb_adr_i[9]
+ wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11] wb_dat_i[12] wb_dat_i[13]
+ wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18] wb_dat_i[19] wb_dat_i[1]
+ wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24] wb_dat_i[25] wb_dat_i[26]
+ wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30] wb_dat_i[31] wb_dat_i[3]
+ wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8] wb_dat_i[9] wb_dat_o[0]
+ wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14] wb_dat_o[15] wb_dat_o[16]
+ wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20] wb_dat_o[21] wb_dat_o[22]
+ wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27] wb_dat_o[28] wb_dat_o[29]
+ wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4] wb_dat_o[5] wb_dat_o[6]
+ wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0] wb_sel_i[1] wb_sel_i[2]
+ wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_95_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6914_ hold73/Z _6915_/RN _6914_/CLK hold72/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6845_ _6845_/D _7170_/RN _6845_/CLK _6845_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6776_ _6776_/D _7194_/RN _6776_/CLK _6776_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3988_ _3988_/I0 _6658_/Q _3988_/S _6658_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5727_ _5775_/I0 hold655/Z _5727_/S _5727_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5658_ hold977/Z _5796_/I0 _5664_/S _5658_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4609_ _4601_/Z _5285_/B _4607_/Z _5021_/B _4612_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_184_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5589_ hold556/Z _5781_/I0 hold34/Z _6952_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold340 _5684_/Z _7036_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_117_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold351 _7041_/Q hold351/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold362 _5649_/Z _7005_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold373 _7058_/Q hold373/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold384 _4224_/Z _6752_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_78_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7259_ _7259_/D _7259_/RN _7260_/CLK _7259_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold395 _5778_/Z _7119_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_117_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold1040 _6870_/Q _3799_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1051 _6917_/Q _5550_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1062 _6716_/Q _4174_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1073 _7304_/Q _3490_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_1_0__f__1062_ clkbuf_0__1062_/Z _4297_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_68_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4960_ _4960_/A1 _5055_/A2 _5270_/A1 _4761_/I _4960_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_17_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3911_ hold258/I _3525_/Z _3913_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_60_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4891_ _5315_/A2 _5399_/A1 _5380_/B2 _5260_/A1 _4891_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_189_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6630_ _7162_/RN _6652_/A2 _6630_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_177_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3842_ _3519_/Z _4185_/A2 _3950_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_177_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1202_461 _4073__37/I _6704_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1202_472 net852_131/I _6693_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6561_ _6561_/A1 _7261_/Q _6833_/D _6561_/B2 _6562_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3773_ _3773_/A1 _3773_/A2 _3773_/A3 _3773_/A4 _3773_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_158_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet1202_483 net1202_483/I _6682_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet1202_494 net1202_494/I _6671_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5512_ _5796_/I0 hold561/Z _5512_/S _5512_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6492_ _6492_/A1 _6492_/A2 _6492_/A3 _6492_/A4 _6492_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_121_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5443_ _5443_/A1 _5245_/Z _5444_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_146_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5374_ _5374_/A1 _5374_/A2 _5374_/A3 _5374_/A4 _5374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7113_ _7113_/D _7185_/RN _7113_/CLK _7113_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4325_ _6613_/I1 hold747/Z _4325_/S _4325_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7044_ _7044_/D _7090_/RN _7044_/CLK _7044_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_101_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4256_ _5860_/I0 hold128/Z _4261_/S _4256_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4187_ _4343_/I0 hold509/Z _4187_/S _4187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6828_ _6828_/D _7261_/RN _7279_/CLK _6828_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_11_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6759_ _6759_/D _7255_/RN _6759_/CLK _6759_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_12_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold170 _6954_/Q hold170/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_151_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold181 _6747_/Q hold181/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold192 _5533_/Z _6903_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_120_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout650 fanout656/Z _7162_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout661 _7171_/RN _7146_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_59_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout672 fanout685/Z _7171_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout683 _7019_/RN _7027_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_93_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout694 _7173_/RN _7205_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4110_ _5798_/I0 hold775/Z _4118_/S _4110_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5090_ _5090_/A1 _5090_/A2 _5400_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_4_3_0__1359_ clkbuf_0__1359_/Z _4073__49/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4041_ _3425_/S _7283_/Q _4041_/A3 _4041_/B1 _3409_/Z _6733_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_49_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5992_ _5992_/A1 _5991_/Z _5995_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_18_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4943_ _4759_/Z _4903_/Z _5330_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_178_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4874_ _4641_/Z _4833_/Z _4874_/B _4874_/C _4876_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_20_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6613_ hold841/Z _6613_/I1 _6613_/S _6613_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3825_ _3519_/Z _5510_/A2 _3933_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_178_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6544_ _6711_/Q _6544_/A2 _6544_/B1 _6810_/Q _6546_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3756_ _6685_/Q _3945_/C2 _3941_/A2 _7161_/Q _3757_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6475_ _6475_/I _6476_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3687_ _3687_/A1 _3687_/A2 _3687_/A3 _3686_/Z _3687_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5426_ _5426_/A1 _4369_/Z _5172_/B _5172_/C _5426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xoutput220 _4062_/Z mgmt_gpio_out[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_134_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput231 _6749_/Q mgmt_gpio_out[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput242 _6752_/Q mgmt_gpio_out[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput253 _4079_/I pad_flash_io0_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput264 hold76/I pll_div[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_161_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5357_ _5357_/A1 _5357_/A2 _5357_/A3 _5357_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xoutput275 hold66/I pll_trim[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput286 hold68/I pll_trim[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput297 _6892_/Q pwr_ctrl_out VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ _6567_/I0 _6814_/Q _4312_/S _6814_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5288_ _5288_/A1 _5468_/A2 _5288_/B _5288_/C _5292_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_87_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7027_ _7027_/D _7027_/RN _7027_/CLK _7027_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_114_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4239_ _4238_/Z hold385/Z _4245_/S _4239_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet852_106 net852_106/I _7119_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet852_117 _4073__17/I _7108_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet852_128 net802_64/I _7097_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout480 _4510_/Z _5236_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout491 hold6/Z _5547_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xnet852_139 net902_185/I _7086_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_171_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3610_ _6571_/I0 _6874_/Q _3898_/S _3610_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4590_ _5269_/A1 _4878_/A2 _4635_/A4 _5367_/A2 _4590_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_174_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3541_ _5875_/A1 _3540_/Z _3541_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_127_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold906 _5711_/Z _7060_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_115_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold917 _7156_/Q hold917/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold928 _5743_/Z _7088_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6260_ _6260_/A1 _6260_/A2 _6260_/A3 _6259_/Z _6260_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold939 _7045_/Q hold939/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3472_ _3472_/I0 hold26/Z _3500_/S hold27/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_43_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5211_ _4892_/B _4683_/Z _5211_/B _5211_/C _5396_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_6191_ _7076_/Q _5965_/Z _5980_/Z _6694_/Q _5967_/Z _6720_/Q _6193_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_130_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5142_ _5281_/C _4539_/I _5142_/A3 _5278_/B _4547_/Z _5470_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_96_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5073_ _4699_/Z _5255_/B _5073_/B _5335_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4024_ _4024_/I _6731_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5975_ _7044_/Q _3386_/I _3387_/I _6211_/A2 _5975_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_80_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4926_ _5324_/A1 _4926_/A2 _4926_/B _4929_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_178_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4857_ _5478_/A1 _4833_/Z _5289_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3808_ _4185_/A2 _3617_/Z _5728_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4788_ _5414_/A2 _5218_/B _5125_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6527_ _6554_/A1 _6521_/Z _6526_/Z _6527_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_3739_ _3739_/A1 _3739_/A2 _3739_/A3 _3739_/A4 _3739_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_134_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6458_ _7116_/Q _6240_/Z _6297_/Z _6704_/Q _6459_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_162_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5409_ _5334_/Z _5409_/A2 _5448_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_121_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6389_ _7031_/Q _6552_/A2 _6273_/Z _6975_/Q _6390_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_121_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_184_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ hold325/Z _5832_/I0 _5766_/S _5760_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4711_ _5307_/A3 _5099_/A1 _5099_/A2 _5401_/A2 _4711_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_1290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5691_ hold291/Z _5775_/I0 _5691_/S _5691_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4642_ _5315_/A1 _5315_/A2 _4990_/A1 _5364_/B _5038_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_175_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4573_ _5373_/A2 _5364_/B _5471_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold703 _6994_/Q hold703/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_7_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6312_ _6989_/Q _6533_/A2 _6533_/A3 _6533_/A4 _6318_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold714 _5726_/Z _7074_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3524_ _5611_/A1 _3523_/Z _3957_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold725 _7082_/Q hold725/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7292_ _7292_/D _6646_/Z _7304_/CLK _7292_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold736 _5730_/Z _7077_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold747 _6823_/Q hold747/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold758 _4273_/Z _6786_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold769 _6971_/Q hold769/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6243_ _6484_/A2 _6533_/A4 _6285_/A2 _6302_/A4 _6243_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_170_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3455_ hold14/Z hold38/Z _3460_/S _7289_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6174_ _7067_/Q _5985_/Z _6000_/Z _7133_/Q _6174_/C _6180_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_58_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3386_ _3386_/I _6002_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_5125_ _5317_/A1 _5123_/Z _5125_/A3 _5126_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_29_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5056_ _5403_/A1 _5051_/Z _5056_/B _5056_/C _5057_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_66_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4007_ _3990_/I _4006_/Z _4008_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet802_55 net802_55/I _7170_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet802_66 net802_66/I _7159_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet802_77 _4073__5/I _7148_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_134__1359_ net1152_446/I _4073__3/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xnet802_88 net802_91/I _7137_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_54__1359_ clkbuf_4_14_0__1359_/Z net952_234/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xnet802_99 net802_99/I _7126_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5958_ _3386_/I _3387_/I _6210_/C _6210_/A2 _5958_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_179_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4909_ _4500_/Z _4973_/A4 _3408_/I _4494_/Z _4909_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5889_ _5889_/I0 hold86/Z _5892_/S hold87/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold30 hold30/I hold30/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold41 hold41/I hold41/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_48_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold52 hold52/I hold52/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold63 hold63/I hold63/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold74 hold74/I hold74/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold85 hold85/I hold85/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold96 hold96/I hold96/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_57_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_7__f_wb_clk_i clkbuf_0_wb_clk_i/Z _4067_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_189_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_84_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_5 _7015_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6930_ _6930_/D _7034_/RN _6930_/CLK _6930_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6861_ _6861_/D _6865_/RN _6865_/CLK _6861_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5812_ _5884_/A2 _5839_/A2 _5857_/A4 _5820_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_6792_ _6792_/D _7258_/CLK _6792_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5743_ _5869_/I0 hold927/Z _5748_/S _5743_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5674_ _5674_/A1 _5674_/A2 _5682_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_148_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4625_ _4887_/A1 _4868_/A1 _5373_/A2 _5364_/B _4625_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_117_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold500 _4241_/Z _6760_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold511 _7090_/Q hold511/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4556_ _4528_/Z _4536_/Z _4556_/A3 _4547_/Z _4556_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold522 _5581_/Z _6945_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_117_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold533 _6935_/Q hold533/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold544 _6857_/Q hold544/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3507_ _3904_/A3 _3680_/A3 hold211/I hold221/I _3507_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold555 _5644_/Z _7001_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7275_ _7275_/D _7278_/RN _7279_/CLK _7275_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_171_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold566 _5511_/Z _6889_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4487_ _4687_/A2 _4687_/A3 _5220_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold577 _7026_/Q hold577/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold588 _6851_/Q hold588/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6226_ _6727_/Q _5994_/I _6226_/B _6227_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_44_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold599 _5640_/Z _6997_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3438_ _4056_/I1 _3438_/I1 _3438_/S _7295_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6157_ _7116_/Q _5984_/Z _5997_/Z _7100_/Q _7074_/Q _5980_/Z _6158_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3369_ _7007_/Q _3369_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _5400_/A1 _5108_/A2 _5310_/C _5107_/I _5108_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6088_ _6088_/I _6089_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5039_ _5035_/Z _5036_/Z _5205_/C _5039_/A4 _5040_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_39_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput120 wb_adr_i[3] input120/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput131 wb_dat_i[12] _6591_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput142 wb_dat_i[22] _6597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput153 wb_dat_i[3] _3396_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput164 wb_sel_i[3] _6575_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4410_ _4412_/B _4412_/C _5003_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_172_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5390_ _5390_/A1 _5390_/A2 _5350_/Z _5390_/A4 _5390_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4341_ _4353_/A1 _3560_/Z _4350_/A3 _4343_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_67_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7060_ _7060_/D _7090_/RN _7060_/CLK _7060_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4272_ _5867_/I0 hold743/Z _4273_/S _4272_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6011_ _6011_/A1 _6450_/S _6011_/B1 _6310_/A3 _7241_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_86_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6913_ _6913_/D _6915_/RN _6913_/CLK _6913_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6844_ _6844_/D _6844_/RN _6844_/CLK _6844_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_62_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6775_ _6775_/D _7194_/RN _6775_/CLK _6775_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3987_ _3984_/S _3972_/Z _3987_/A3 _3987_/B _3988_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_10_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5726_ _5855_/I0 hold713/Z _5727_/S _5726_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5657_ hold933/Z _5795_/I0 _5664_/S _5657_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4608_ _5373_/A2 _4449_/B _4853_/A1 _4635_/A4 _5021_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5588_ hold460/Z _5798_/I0 hold34/Z _6951_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold330 _4231_/Z _6755_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold341 _7056_/Q hold341/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4539_ _4539_/I _5281_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xhold352 _5689_/Z _7041_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold363 _7177_/Q hold363/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold374 _5708_/Z _7058_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold385 _6759_/Q hold385/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_131_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold396 _7022_/Q hold396/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7258_ _7258_/D _7258_/RN _7258_/CLK _7258_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_120_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6209_ _7297_/Q _5969_/Z _6227_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_132_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7189_ _7189_/D _7201_/RN _7189_/CLK _7189_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1030 _5840_/Z _7174_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1041 _6871_/Q _3762_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold1052 _7272_/Q _4107_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold1063 _7010_/Q hold233/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1074 _7105_/Q hold479/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_133_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3910_ _6932_/Q _3910_/A2 _3953_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_189_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4890_ _4890_/I _5259_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_189_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3841_ _6695_/Q _4143_/A1 _3868_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_20_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3772_ hold36/I _3912_/A2 _3930_/A2 _7128_/Q _3773_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xnet1202_462 net852_150/I _6703_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6560_ _6561_/B2 _6559_/Z _6561_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xnet1202_473 net852_131/I _6692_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_186_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1202_484 net1202_485/I _6681_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1202_495 net802_84/I _6670_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5511_ _5795_/I0 hold565/Z _5512_/S _5511_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6491_ _7173_/Q _6544_/A2 _6544_/B1 _6963_/Q _6545_/B1 _7019_/Q _6492_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_8_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5442_ _5442_/A1 _5442_/A2 _5442_/A3 _5442_/A4 _5442_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_146_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5373_ _5287_/C _5373_/A2 _5287_/B _5373_/B _5374_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_4324_ _6612_/I1 hold787/Z _4325_/S _4324_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7112_ _7112_/D _7019_/RN _7112_/CLK _7112_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_59_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7043_ _7043_/D _7237_/RN _7043_/CLK _7043_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_87_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4255_ hold54/Z hold94/Z _4261_/S hold95/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4186_ _4103_/I hold537/Z _4187_/S _4186_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6827_ _6827_/D _7261_/RN _7279_/CLK _6833_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_6758_ _6758_/D _7255_/RN _6758_/CLK _6758_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_6_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5709_ hold250/Z _5892_/I0 _5709_/S _5709_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6689_ hold71/Z _6847_/RN _6689_/CLK hold70/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_109_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold160 _6920_/Q hold160/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold171 _6904_/Q hold171/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_176_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold182 _4214_/Z _6747_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_78_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold193 _6878_/Q hold193/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_137_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout640 _7154_/RN _7170_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout651 fanout656/Z _7194_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout662 _7171_/RN _7090_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout673 _6821_/RN _7211_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout684 fanout685/Z _7019_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_86_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout695 fanout714/Z _7173_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_92_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4040_ _4040_/I _6734_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_76_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5991_ _6117_/A2 _5991_/A2 _6021_/A4 _5991_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_92_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4942_ _4939_/Z _4942_/A2 _5062_/B _4948_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_17_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4873_ _4641_/Z _4873_/A2 _4873_/A3 _4681_/Z _4874_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_32_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6612_ hold825/Z _6612_/I1 _6613_/S _6612_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3824_ _3844_/A1 _3653_/Z _3935_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_165_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6543_ _6852_/Q _6543_/A2 _6285_/Z _6693_/Q _6707_/Q _6254_/Z _6546_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3755_ _6951_/Q _5584_/A1 _3956_/A2 _7121_/Q _7145_/Q _3951_/C1 _3757_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3686_ _3686_/A1 _3686_/A2 _3686_/A3 _3686_/A4 _3686_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6474_ _3324_/I _7256_/Q _6474_/B _6475_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_146_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput210 _4056_/Z mgmt_gpio_out[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5425_ _5425_/A1 _5425_/A2 _5425_/A3 _5425_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
Xoutput221 _6739_/Q mgmt_gpio_out[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_145_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput232 hold72/I mgmt_gpio_out[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput243 _4059_/Z mgmt_gpio_out[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput254 _7307_/Z pad_flash_io1_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5356_ _5356_/A1 _5387_/A2 _5356_/B _5356_/C _5357_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xoutput265 _6881_/Q pll_div[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput276 _6680_/Q pll_trim[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput287 _6889_/Q pll_trim[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4307_ _6566_/I0 _6813_/Q _4312_/S _6813_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput298 _3907_/Z reset VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_87_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5287_ _5290_/A2 _5287_/A2 _5287_/B _5287_/C _5487_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_7026_ _7026_/D _7027_/RN _7026_/CLK _7026_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4238_ hold160/Z _5880_/I0 _4242_/S _4238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4169_ _5538_/I1 hold649/Z _4169_/S _4169_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet852_107 net852_147/I _7118_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout470 _5291_/C _5276_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet852_118 net802_62/I _7107_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout481 _4495_/Z _4982_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet852_129 net802_73/I _7096_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout492 hold5/Z hold6/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_46_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3540_ _3653_/A1 hold144/I _3500_/Z _3492_/Z _3540_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_128_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold907 _7086_/Q hold907/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold918 _5819_/Z _7156_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_171_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold929 _6948_/Q hold929/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3471_ _3471_/I _3472_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5210_ _5209_/Z _5208_/Z _5417_/A1 _5210_/A4 _5210_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6190_ _6716_/Q _5997_/Z _6014_/Z _6809_/Q _6193_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_130_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5141_ _5293_/A1 _5290_/A3 _5289_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_36_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5072_ _4500_/Z _4906_/Z _5078_/A2 _5072_/A4 _5072_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_97_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4023_ _4023_/A1 _4022_/Z _4024_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_77_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5974_ _5974_/A1 _5974_/A2 _5974_/A3 _5974_/A4 _5983_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4925_ _5080_/B _5080_/C _5370_/B _4926_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_80_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4856_ _5478_/A1 _4817_/Z _4858_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_165_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3807_ _5629_/A1 _3519_/Z _3923_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4787_ _5220_/B2 _5092_/A1 _4787_/A3 _4491_/B _4787_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_181_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6526_ _6526_/A1 _6526_/A2 _6526_/A3 _6526_/A4 _6526_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3738_ input67/Z _4227_/S _4242_/S input38/Z _5701_/A1 _7055_/Q _3739_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_147_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6457_ _7188_/Q _6532_/A2 _6293_/Z _7156_/Q _6296_/Z _7164_/Q _6465_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3669_ _6953_/Q _5584_/A1 _3959_/B1 _6671_/Q _3673_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5408_ _4761_/I _5245_/Z _5481_/B1 _4908_/Z _5408_/C _5409_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_47_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6388_ _6943_/Q _6551_/A2 _6288_/Z _7121_/Q _6390_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xclkbuf_leaf_77__1359_ net902_187/I _4073__41/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5339_ _5261_/I _5338_/Z _5262_/Z _5339_/A4 _5340_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_47_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7009_ _7009_/D _7259_/RN _7009_/CLK _7009_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_28_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_6__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7279_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_83_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4710_ _4694_/Z _5401_/A2 _5308_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_1291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5690_ hold279/Z _5855_/I0 _5691_/S _5690_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4641_ _5281_/C _4467_/B _4472_/B _3406_/I _4641_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_187_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4572_ _4572_/I _5472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_129_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6311_ _6973_/Q _6402_/A2 _6311_/A3 _6533_/A2 _6327_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold704 _5636_/Z _6994_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3523_ _3904_/A3 hold144/I hold211/I hold221/I _3523_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold715 _7181_/Q hold715/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold726 _5736_/Z _7082_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_155_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7291_ _7291_/D _6645_/Z _7302_/CLK _7291_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold737 _6978_/Q hold737/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold748 _4325_/Z _6823_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6242_ _7110_/Q _6240_/Z _6550_/A2 _7044_/Q _6260_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold759 _6986_/Q hold759/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_131_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3454_ hold4/Z hold14/Z _3460_/S _7290_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3385_ _3385_/I _3385_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6173_ _6173_/I _6174_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5124_ _5414_/A2 _5228_/A3 _5124_/B _5317_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_69_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5055_ _5130_/B2 _5055_/A2 _4367_/Z _5276_/B _5055_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_111_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4006_ _5900_/A1 _5911_/A1 _7225_/Q _7224_/Q _4006_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_2909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet802_56 net802_64/I _7169_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet802_67 net802_67/I _7158_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet802_78 net802_78/I _7147_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet802_89 net802_89/I _7136_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_1__1359_ net1152_451/I net1152_421/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5957_ _3990_/I _5957_/I1 _5957_/S _6476_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4908_ _5324_/A1 _4759_/Z _4494_/Z _4496_/Z _4908_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5888_ _5888_/I0 hold548/Z _5892_/S _5888_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4839_ _4887_/A1 _5364_/A1 _5399_/A2 _5369_/A1 _5369_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_166_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6509_ _6692_/Q _6285_/Z _6299_/Z _6857_/Q _6511_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_106_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold20 hold20/I hold20/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_130_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold31 hold31/I hold31/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold42 hold42/I hold42/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_76_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold53 hold53/I hold53/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold64 hold64/I hold64/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_188_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold75 hold75/I hold75/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_29_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold86 hold86/I hold86/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_63_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold97 hold97/I hold97/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_75_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_6 _6943_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_60__1359_ clkbuf_4_13_0__1359_/Z net902_191/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_140__1359_ net1152_446/I net802_75/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_140_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6860_ _6860_/D _6865_/RN _6865_/CLK _6860_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5811_ _5811_/I0 hold857/Z _5811_/S _5811_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6791_ _6791_/D _7262_/CLK _6791_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5742_ _5859_/I0 hold881/Z _5748_/S _5742_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5673_ hold789/Z _5784_/I0 _5673_/S _5673_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4624_ _5365_/A3 _5281_/C _4752_/A2 _3406_/I _4624_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_129_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold501 _6764_/Q hold501/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_156_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4555_ _5129_/A3 _4715_/A1 _4555_/B _4555_/C _4556_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xhold512 _5745_/Z _7090_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold523 _6726_/Q hold523/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold534 _5570_/Z _6935_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold545 _4360_/Z _6857_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3506_ _5875_/A1 _3505_/Z _3909_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_104_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold556 hold556/I hold556/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_1_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7274_ _7274_/D _7278_/RN _7279_/CLK _7274_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4486_ _4486_/A1 _4877_/A2 _4486_/B1 _4484_/Z _5312_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold567 _6970_/Q hold567/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold578 _5672_/Z _7026_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_131_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6225_ _6800_/Q _5958_/Z _5967_/Z _6721_/Q _6227_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold589 _4351_/Z _6851_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_103_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3437_ _3442_/B _6663_/Q _6664_/Q _3441_/C _3438_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_98_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6156_ _7156_/Q _5960_/Z _5965_/Z _6704_/Q _6006_/Z _7172_/Q _6158_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3368_ _7015_/Q _3368_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ _5107_/I _5309_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6087_ _6364_/C _7243_/Q _6087_/B _6088_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_57_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3299_ _3441_/C _3465_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5038_ _5038_/A1 _4606_/Z _5003_/Z _5038_/B _5205_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XTAP_2706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6989_ _6989_/D fanout658/Z _6989_/CLK _6989_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_53_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet1002_290 _4073__8/I _6935_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_166_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput110 wb_adr_i[23] _4026_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_1_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput121 wb_adr_i[4] input121/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput132 wb_dat_i[13] _6594_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput143 wb_dat_i[23] _6600_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput154 wb_dat_i[4] _3397_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput165 wb_stb_i _4032_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_91_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4340_ _4361_/I1 hold615/Z _4340_/S _4340_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4271_ _5821_/A1 _5510_/A2 _4347_/A3 _5839_/A3 _4273_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6010_ _6010_/A1 _6010_/A2 _6924_/Q _6201_/A3 _6011_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_97_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6912_ _6912_/D _6915_/RN _6912_/CLK _6912_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_70_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6843_ _6843_/D _6844_/RN _6843_/CLK _6843_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_63_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6774_ _6774_/D _7194_/RN _6774_/CLK _6774_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3986_ _7305_/Q _3415_/Z _6658_/Q _3987_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5725_ hold40/Z hold46/Z _5727_/S hold47/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5656_ _5656_/A1 _5674_/A2 _5664_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_163_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4607_ _4607_/A1 _4570_/Z _4606_/Z _4449_/B _4607_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5587_ hold392/Z _5797_/I0 hold34/Z _5587_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold320 _4209_/Z _6741_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold331 _6922_/Q hold331/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_151_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4538_ _5288_/B _4467_/B _4472_/B _4539_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_117_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold342 _5706_/Z _7056_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold353 _6737_/Q hold353/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold364 _5843_/Z _7177_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_132_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold375 _7039_/Q hold375/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7257_ _7257_/D _7257_/RN _7257_/CLK _7257_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4469_ _4459_/Z _4469_/A2 _4690_/B _4690_/C _4786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold386 _4239_/Z _6759_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold397 _5668_/Z _7022_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6208_ _7249_/Q _6208_/I1 _6558_/S _7249_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7188_ _7188_/D _7188_/RN _7188_/CLK _7188_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6139_ _7058_/Q _6139_/A2 _6210_/B _6210_/C _6155_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1020 _5869_/Z _7200_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1031 _7143_/Q _5805_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1042 _6869_/Q _3899_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold1053 _5878_/Z hold3/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1064 _6717_/Q hold492/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1075 _7007_/Q hold232/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3840_ _4185_/A2 _3680_/Z _4143_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_32_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet1202_452 net1202_452/I _6713_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1202_463 net1202_463/I _6702_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3771_ _7070_/Q _3943_/A2 _3945_/B1 _7088_/Q _3773_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xnet1202_474 net1202_474/I _6691_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1202_485 net1202_485/I _6680_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5510_ _5776_/A1 _5510_/A2 _5794_/A3 _5512_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_157_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1202_496 net1202_499/I _6669_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_186_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6490_ _7085_/Q _6290_/Z _6302_/Z _7093_/Q _6490_/C _6492_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_145_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5441_ _5437_/Z _5440_/Z _5441_/B _5463_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_145_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5372_ _5372_/A1 _5139_/Z _5055_/Z _5372_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_99_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7111_ _7111_/D _7215_/RN _7111_/CLK _7111_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4323_ _4332_/A1 _5821_/A3 hold146/Z _5794_/A3 _4325_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_114_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7042_ _7042_/D _7188_/RN _7042_/CLK _7042_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_99_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4254_ hold64/Z hold118/Z _4261_/S _4254_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4185_ _5520_/C _4185_/A2 hold146/Z _5629_/A3 _4187_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_68_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6826_ _6826_/D _7261_/RN _7279_/CLK _6826_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_23_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6757_ _6757_/D _7257_/RN _6757_/CLK _6757_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3969_ _3427_/Z _6663_/Q _6664_/Q _3970_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5708_ hold373/Z _5891_/I0 _5709_/S _5708_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6688_ _6688_/D _7296_/RN _6688_/CLK _6688_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_12_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_opt_3_0__1359_ _4073__24/I clkbuf_opt_3_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_137_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5639_ hold273/Z _5876_/I0 _5646_/S _5639_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold150 hold150/I hold150/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7309_ _7309_/I _7309_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_1070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold161 _5553_/Z _6920_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold172 _5534_/Z _6904_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold183 _6753_/Q hold183/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold194 _5498_/Z _6878_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xfanout630 _5426_/A1 _5097_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout641 _7077_/RN _7154_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_120_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout652 fanout656/Z _7218_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout663 _7171_/RN _7141_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout674 _6821_/RN _7202_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout685 input75/Z fanout685/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_19_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout696 _7149_/RN _7125_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_3001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5990_ _7020_/Q _6211_/A2 _6002_/A2 _6956_/Q _6211_/B1 _6988_/Q _5992_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_91_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4941_ _5464_/A1 _5410_/A1 _5062_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4073__50 net802_99/I _7175_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4872_ _4872_/A1 _5215_/C _5117_/A2 _5215_/B _4874_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_60_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6611_ _6611_/A1 _6611_/A2 _6613_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3823_ _6981_/Q _3901_/A2 _3889_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_177_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6542_ _6542_/A1 _6542_/A2 _6542_/A3 _6542_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_3754_ _7137_/Q _3951_/A2 _3954_/B1 input23/Z _3754_/C _3757_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_119_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6473_ _6466_/Z _6472_/Z _6473_/B1 _6286_/Z _6500_/C _6474_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3685_ _6961_/Q _3957_/A2 _3941_/B1 _7171_/Q _3686_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_146_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5424_ _5489_/A1 _5423_/Z _5427_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_160_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput200 _4050_/Z mgmt_gpio_oeb[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput211 _6758_/Q mgmt_gpio_out[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput222 _6740_/Q mgmt_gpio_out[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput233 _6915_/Q mgmt_gpio_out[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput244 _6754_/Q mgmt_gpio_out[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_142_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5355_ _5437_/A2 _5350_/Z _5352_/Z _5354_/Z _5355_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xoutput255 _4077_/ZN pad_flash_io1_ie VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput266 _6882_/Q pll_div[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput277 hold56/I pll_trim[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4306_ _6565_/I0 _6812_/Q _4312_/S _6812_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput288 _6890_/Q pll_trim[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput299 _4085_/Z ser_rx VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5286_ _5286_/A1 _5374_/A3 _5374_/A2 _5292_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_102_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7025_ _7025_/D _7122_/RN _7025_/CLK _7025_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_87_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4237_ _4236_/Z hold420/Z _4245_/S _4237_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4168_ _5537_/I1 hold635/Z _4169_/S _4168_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_3_5__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7260_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4099_ hold9/Z _6608_/I0 _4117_/S hold10/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6809_ _6809_/D _6847_/RN _6809_/CLK _6809_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_177_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout460 _4700_/Z _5260_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet852_108 net952_234/I _7117_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_119 net852_119/I _7106_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout471 _4990_/A1 _5373_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout482 _4446_/Z _5287_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout493 hold16/Z _5645_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_93_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold908 _5741_/Z _7086_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_183_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold919 _7078_/Q hold919/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_7_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3470_ _6660_/Q _3978_/S _3470_/B hold255/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_155_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5140_ _5293_/A1 _4549_/Z _5147_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_69_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5071_ _4376_/Z _5071_/A2 _5257_/A1 _4699_/Z _5408_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_56_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4022_ _7282_/Q _3409_/Z _4022_/A3 _6730_/Q _4022_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_65_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5973_ _7012_/Q _5971_/Z _5972_/Z _6940_/Q _5974_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4924_ _5259_/A1 _5337_/A2 _5258_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_21_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4855_ _5287_/C _4844_/Z _4855_/B _4855_/C _4858_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_127_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3806_ _5629_/A1 _4350_/A2 _3924_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_178_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4786_ _4786_/A1 _4786_/A2 _4786_/A3 _5137_/B1 _4787_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_165_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6525_ _6694_/Q _6248_/Z _6300_/Z _6720_/Q _6526_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3737_ _6927_/Q _3935_/A2 _3916_/A2 _7153_/Q _3912_/B1 _6886_/Q _3739_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_107_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6456_ _7140_/Q _6253_/Z _6540_/A2 _7204_/Q _6456_/C _6465_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_174_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3668_ _7083_/Q _3923_/C1 _3956_/A2 _7123_/Q _3668_/C _3674_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_109_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5407_ _5406_/Z _5454_/A2 _5419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6387_ _7047_/Q _6550_/A2 _6550_/B1 _6983_/Q _6268_/Z _6951_/Q _6390_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3599_ _7011_/Q _3934_/A2 _5683_/A1 _7043_/Q _7051_/Q _3952_/A2 _3601_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_47_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5338_ _5332_/Z _5334_/Z _5447_/A1 _5338_/A4 _5338_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_87_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5269_ _5269_/A1 _5269_/A2 _4651_/Z _5380_/B2 _5464_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_130_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7008_ _7008_/D _7259_/RN _7008_/CLK _7008_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_75_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_20__1359_ _4073__49/I net902_157/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_100__1359_ clkbuf_4_5_0__1359_/Z net802_78/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_83__1359_ net902_187/I net802_81/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_148_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4640_ _5315_/A1 _5315_/A2 _5468_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_147_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4571_ _4549_/Z _4570_/Z _4572_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_128_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6310_ _6308_/Z _6310_/A2 _6310_/A3 _6450_/S _6310_/B2 _7251_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_3522_ _5629_/A1 _5776_/A1 _3910_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold705 _6958_/Q hold705/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7290_ _7290_/D _6644_/Z _7302_/CLK hold4/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold716 _5847_/Z _7181_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold727 _6855_/Q hold727/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold738 _5618_/Z _6978_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6241_ _3328_/I _6300_/A1 _6300_/A2 _6275_/A4 _6241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold749 _7185_/Q hold749/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3453_ _4041_/B1 _3442_/B _6732_/Q _3460_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_115_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6172_ _6979_/Q _5964_/Z _6014_/Z _6963_/Q _5999_/Z _7035_/Q _6173_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3384_ _6786_/Q _6555_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_58_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5123_ _5456_/A1 _5220_/B2 _5312_/A2 _5137_/B1 _5123_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_112_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5054_ _5370_/B _5258_/A2 _4977_/Z _5248_/A3 _5324_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_38_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4005_ _4005_/A1 _4003_/Z _5945_/A1 _6901_/Q _6743_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_37_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet802_57 net802_73/I _7168_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet802_68 net802_68/I _7157_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet802_79 net802_89/I _7146_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5956_ _5957_/S _5957_/I1 _6310_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4907_ _4759_/Z _4906_/Z _5257_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5887_ hold2/Z hold36/Z _5892_/S hold37/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4838_ _4555_/C _4876_/A2 _4838_/B1 _5276_/B _4841_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_178_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4769_ _5401_/A2 _4764_/Z _5117_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_5_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6508_ _6724_/Q _6240_/Z _6247_/Z _6728_/Q _6511_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_147_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6439_ _6434_/Z _6439_/A2 _6439_/A3 _6439_/A4 _6439_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_122_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold10 hold10/I hold10/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold21 hold21/I hold21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold32 hold32/I hold32/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_102_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold43 hold43/I hold43/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold54 hold54/I hold54/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold65 hold65/I hold65/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold76 hold76/I hold76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold87 hold87/I hold87/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold98 hold98/I hold98/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_90_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet1052_350 _4073__31/I _6867_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_7 user_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5810_ _5891_/I0 hold843/Z _5811_/S _5810_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6790_ _6790_/D _6933_/RN _6790_/CLK _6790_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_76_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5741_ _5867_/I0 hold907/Z _5748_/S _5741_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_188_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5672_ hold577/Z _5837_/I0 _5673_/S _5672_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4623_ _4887_/A1 _4868_/A1 _5376_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_176_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4554_ _5426_/A1 _4836_/A3 _5420_/A4 _4873_/A2 _4554_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold502 _4248_/Z _6764_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold513 _7049_/Q hold513/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold524 _4189_/Z _6726_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3505_ hold144/I hold210/Z _3489_/I _3492_/Z _3505_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold535 _6841_/Q hold535/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7273_ _7273_/D _7278_/RN _7279_/CLK _7273_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold546 _6728_/Q hold546/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4485_ _4381_/Z _4485_/A2 _4486_/B1 _4424_/B _4687_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold557 _6846_/Q hold557/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold568 _5609_/Z _6970_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6224_ _6719_/Q _5960_/Z _5965_/Z _7077_/Q _6006_/Z _6711_/Q _6227_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold579 _7120_/Q hold579/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3436_ _3441_/C _6664_/Q _6663_/Q _3898_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_106_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6155_ _6155_/A1 _6155_/A2 _6155_/A3 _6155_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XTAP_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3367_ _7023_/Q _3367_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5106_ _5106_/A1 _5106_/A2 _5107_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ _6073_/Z _6085_/Z _6392_/B1 _6118_/B _6744_/Q _6087_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_100_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3298_ hold8/Z hold9/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5037_ _5039_/A4 _5036_/Z _5357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_100_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6988_ _6988_/D fanout658/Z _6988_/CLK _6988_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5939_ _5957_/I1 _5939_/A2 _5913_/I _6282_/A2 _7233_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_40_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1002_280 net1052_328/I _6945_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1002_291 net952_206/I _6934_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput100 wb_adr_i[14] _4386_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput111 wb_adr_i[24] _4029_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput122 wb_adr_i[5] _5322_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_76_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput133 wb_dat_i[14] _6597_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput144 wb_dat_i[24] _6579_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput155 wb_dat_i[5] _3398_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput166 wb_we_i _6575_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_91_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4270_ hold293/Z _5784_/I0 _4270_/S _4270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6911_ _6911_/D _6915_/RN _6911_/CLK _6911_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6842_ _6842_/D _6844_/RN _6842_/CLK _6842_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_62_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6773_ hold99/Z _7193_/RN _6773_/CLK hold98/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3985_ _3984_/Z _6659_/Q _3988_/S _6659_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5724_ _5724_/I0 hold480/Z _5727_/S _5724_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5655_ hold234/Z _5811_/I0 _5655_/S _5655_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4606_ _4648_/A2 _4944_/A1 _4648_/A1 _4606_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_5586_ _5586_/I0 _5796_/I0 hold34/Z _5586_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold310 _5799_/Z _7138_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_105_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold321 _6879_/Q hold321/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4537_ _5365_/A3 _3406_/I _5399_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_2_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold332 _5555_/Z _6922_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold343 _7057_/Q hold343/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold354 _4201_/Z _6737_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7256_ _7256_/D _7257_/RN _7257_/CLK _7256_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold365 _7055_/Q hold365/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4468_ _4467_/B _4736_/A1 _4468_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
Xhold376 _5687_/Z _7039_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold387 _6863_/Q hold387/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold398 _6942_/Q hold398/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6207_ _6207_/I _6208_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3419_ _4041_/B1 _6730_/Q _7304_/Q _3421_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7187_ _7187_/D _7211_/RN _7187_/CLK _7187_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4399_ _4402_/B _4395_/B _4026_/B _4026_/C _4399_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6138_ _7108_/Q _5967_/Z _6147_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1010 _5695_/Z _7046_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1021 _7199_/Q _5868_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1032 _5805_/Z _7143_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1043 _6873_/Q _3691_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ _7063_/Q _5985_/Z _6084_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold1054 _6659_/Q _3475_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1065 _6953_/Q hold541/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold1076 _6819_/Q hold1076/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3770_ _7160_/Q _3941_/A2 _5503_/A2 _3904_/A2 _3770_/C _3773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xnet1202_453 net1202_453/I _6712_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1202_464 net852_150/I _6701_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_160_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet1202_475 net802_55/I _6690_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet1202_486 net1202_486/I _6679_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1202_497 net802_84/I _6668_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5440_ _5440_/A1 _5357_/Z _5388_/Z _5440_/A4 _5440_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_173_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5371_ _5371_/A1 _5278_/B _5470_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_59_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7110_ _7110_/D _7215_/RN _7110_/CLK _7110_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4322_ _5859_/I0 hold569/Z _4322_/S _4322_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7041_ _7041_/D _7163_/RN _7041_/CLK _7041_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4253_ _5857_/A1 _3540_/Z _4060_/S _5884_/A3 _4261_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_101_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4184_ hold845/Z _4361_/I1 _4184_/S _4184_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_4__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7257_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_27_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6825_ _6825_/D _6839_/RN _6825_/CLK _6825_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6756_ _6756_/D _7125_/RN _6756_/CLK _6756_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3968_ _3441_/C _3967_/Z _6665_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_10_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5707_ hold343/Z _5881_/I0 _5709_/S _5707_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6687_ hold51/Z _7296_/RN _6687_/CLK hold50/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_148_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3899_ _3898_/Z _3899_/I1 _3899_/S _6869_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5638_ _5638_/A1 _5674_/A2 _5646_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_163_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5569_ _5806_/I0 hold909/Z _5574_/S _5569_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold140 _6684_/Q hold140/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7308_ _7308_/I _7308_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold151 _3493_/Z hold151/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_2_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold162 _6676_/Q hold162/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_132_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold173 _6777_/Q hold173/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold184 _4226_/Z _6753_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold195 _6780_/Q hold195/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7239_ _7239_/D _7240_/RN _4067_/I1 _7239_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_144_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout620 _4441_/B _5365_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout631 _3401_/I _5426_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xfanout642 _6847_/RN _7296_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout653 fanout656/Z _7098_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_59_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout664 _7171_/RN _7155_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout675 fanout677/Z _6821_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_19_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout686 _7219_/RN _7179_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_86_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout697 _7149_/RN _7034_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4940_ _5010_/A1 _5410_/A1 _4942_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_45_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4871_ _4641_/Z _5142_/A3 _5117_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4073__40 net802_96/I _7185_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__51 _4073__51/I _7174_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3822_ _6788_/Q _4274_/A1 _3947_/B1 _6717_/Q _3873_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_21_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6610_ _6610_/A1 _6610_/A2 _6610_/A3 _6610_/A4 _7279_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6541_ _6725_/Q _6240_/Z _6248_/Z _6695_/Q _6542_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_20_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3753_ _3753_/I _3754_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6472_ _6554_/A1 _6472_/A2 _6472_/A3 _6472_/A4 _6472_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3684_ _7155_/Q _3916_/A2 _5528_/S _3683_/Z _3686_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_145_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5423_ _5423_/A1 _5423_/A2 _5377_/Z _5422_/Z _5423_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_134_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput201 _4049_/Z mgmt_gpio_oeb[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput212 _6759_/Q mgmt_gpio_out[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_161_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput223 _6741_/Q mgmt_gpio_out[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5354_ _5354_/A1 _5354_/A2 _5354_/A3 _5354_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xoutput234 _4053_/Z mgmt_gpio_out[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput245 _4058_/Z mgmt_gpio_out[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput256 _4077_/I pad_flash_io1_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput267 _6876_/Q pll_ena VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4305_ _6564_/I0 _6811_/Q _4312_/S _6811_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput278 _6666_/Q pll_trim[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput289 _6684_/Q pll_trim[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5285_ _4598_/Z _5287_/A2 _5285_/B _5374_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_99_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7024_ _7024_/D _7024_/RN _7024_/CLK _7024_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4236_ hold359/Z _5879_/I0 _4242_/S _4236_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4167_ _4350_/A2 _4185_/A2 _4350_/A3 _4169_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_4098_ _6656_/A1 _6657_/A2 _4098_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_36_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6808_ _6808_/D _7262_/CLK _6808_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6739_ _6739_/D _7193_/RN _6739_/CLK _6739_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout450 _6533_/A2 _6275_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_48_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout461 _4699_/Z _5403_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xfanout472 _4551_/Z _4990_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xnet852_109 net802_93/I _7116_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout483 _4421_/Z _5010_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_24_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout494 _5555_/I0 _5837_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_74_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold909 _6934_/Q hold909/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_182_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5070_ _5070_/A1 _5070_/A2 _5334_/A1 _5070_/A4 _5074_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xclkbuf_leaf_43__1359_ clkbuf_4_11_0__1359_/Z _4073__5/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_123__1359_ _4073__49/I net852_146/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_78_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4021_ _4021_/I _6746_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5972_ _5991_/A2 _6210_/C _6015_/A3 _6139_/A2 _5972_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4923_ _4423_/Z _4923_/A2 _4923_/B _5080_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_33_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4854_ _5290_/A1 _5364_/A1 _5478_/A1 _4483_/B _4855_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_20_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3805_ _3519_/Z _5839_/A2 _3912_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4785_ _4808_/A2 _5220_/B2 _5092_/A1 _4491_/B _5124_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_118_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6524_ _6690_/Q _6257_/Z _6536_/B1 _6849_/Q _6526_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3736_ _7217_/Q _3912_/A2 _4194_/A1 input55/Z _3948_/C1 input64/Z _3739_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_109_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3667_ _3667_/I _3668_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6455_ _7084_/Q _6290_/Z _6299_/Z _7058_/Q _6466_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5406_ _5406_/A1 _5404_/Z _5406_/A3 _4799_/Z _5406_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_162_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6386_ _7023_/Q _6549_/A2 _6549_/B1 _7007_/Q _6265_/Z _6999_/Q _6391_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3598_ _7165_/Q _3941_/A2 _3947_/A2 _7101_/Q _7059_/Q _5701_/A1 _3601_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_115_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5337_ _5337_/A1 _5337_/A2 _5337_/B _5337_/C _5449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_88_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5268_ _5368_/A1 _4650_/Z _5172_/C _5268_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_4219_ hold195/Z _5798_/I0 _4227_/S _4219_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7007_ _7007_/D _7125_/RN _7007_/CLK _7007_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_69_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ _5191_/Z _5196_/Z _5390_/A2 _5476_/A2 _5199_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_29_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4570_ _5270_/A1 _5269_/A1 _5364_/B _4570_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_162_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3521_ hold221/I _3492_/Z _3680_/A3 hold211/Z _3521_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_128_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold706 _5596_/Z _6958_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_7_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold717 _7188_/Q hold717/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold728 _4357_/Z _6855_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6240_ _7236_/Q _6533_/A4 _6302_/A4 _6533_/A3 _6240_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold739 _6981_/Q hold739/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3452_ _3451_/Z _7291_/Q _3452_/S _7291_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6171_ _7149_/Q _5987_/Z _6002_/Z _7093_/Q _6003_/Z _7165_/Q _6181_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3383_ _7077_/Q _3866_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5122_ _5456_/A1 _5231_/A2 _5122_/B _5213_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_85_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5053_ _5325_/B _5078_/A2 _5060_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_133_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4004_ _4005_/A1 _4003_/Z _5894_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_38_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet802_58 net802_64/I _7167_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet802_69 _4073__4/I _7156_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5955_ _5954_/Z _7240_/Q _5955_/S _7240_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4906_ _4494_/Z _5259_/A1 _4496_/Z _4407_/Z _4906_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5886_ _5886_/I0 hold663/Z _5892_/S _5886_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4837_ _5278_/C _5164_/A4 _4838_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4768_ _5236_/A1 _4764_/Z _4770_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_146_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6507_ _6726_/Q _6253_/Z _6296_/Z _6714_/Q _6511_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_181_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3719_ _3719_/A1 _3719_/A2 _3719_/A3 _3719_/A4 _3719_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_107_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4699_ _5420_/A3 _4835_/A2 _5420_/A4 _4878_/A4 _4699_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_20_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6438_ _7083_/Q _6290_/Z _6302_/Z _7091_/Q _6438_/C _6439_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_150_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6369_ _6967_/Q _6531_/A2 _6391_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xnet902_190 net952_218/I _7035_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold11 hold11/I hold11/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold22 hold22/I hold22/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_130_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold33 hold33/I hold33/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_75_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold44 hold44/I hold44/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_152_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold55 hold55/I hold55/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold66 hold66/I hold66/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold77 hold77/I hold77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold88 hold88/I hold88/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_91_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold99 hold99/I hold99/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_56_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet1052_340 net1052_346/I _6885_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xnet1052_351 net802_64/I _6866_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_8 hold258/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5740_ _5884_/A2 _5767_/A3 _5857_/A4 _5748_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_176_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5671_ hold482/Z _5782_/I0 _5673_/S _5671_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4622_ _4622_/A1 _5029_/B _5353_/B _4627_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_175_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4553_ _4836_/A4 _5270_/A2 _5370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold503 _6968_/Q hold503/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold514 _5698_/Z _7049_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold525 _7024_/Q hold525/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3504_ hold152/Z _5857_/A3 hold153/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold536 _4336_/Z _6841_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7272_ _7272_/D _7278_/RN _7279_/CLK _7272_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4484_ _4381_/Z _4385_/Z _4387_/Z _4424_/B _4484_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold547 _4192_/Z _6728_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold558 _4343_/Z _6846_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6223_ _6691_/Q _5985_/Z _6014_/Z _6810_/Q _6228_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold569 _6821_/Q hold569/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3435_ _3435_/A1 _3435_/A2 _7298_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_143_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6154_ _7018_/Q _5971_/Z _6005_/Z _7042_/Q _7050_/Q _6019_/Z _6155_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3366_ _7031_/Q _3366_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5105_ _5105_/A1 _5104_/Z _5310_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_97_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6085_ _6078_/Z _6085_/A2 _6085_/A3 _6084_/Z _6085_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_111_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3297_ _7291_/Q _3451_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5036_ _5356_/C _5389_/C _5328_/A1 _5356_/B _5036_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_26_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6987_ _6987_/D _7124_/RN _6987_/CLK _6987_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_80_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5938_ _6484_/A2 _6302_/A3 _5939_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_139_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5869_ _5869_/I0 _5869_/I1 _5874_/S _5869_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1002_270 net802_78/I _6955_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1002_281 net1052_328/I _6944_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1002_292 net1202_485/I _6933_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_166_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput101 wb_adr_i[15] _4386_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_103_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput112 wb_adr_i[25] _3334_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput123 wb_adr_i[6] _4549_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput134 wb_dat_i[15] _6600_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput145 wb_dat_i[25] _6582_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput156 wb_dat_i[6] _3399_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_3__f_wb_clk_i clkbuf_0_wb_clk_i/Z _6865_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_6_0__1359_ clkbuf_0__1359_/Z net952_221/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6910_ hold93/Z _7193_/RN _6910_/CLK hold92/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6841_ _6841_/D _6844_/RN _6841_/CLK _6841_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_51_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6772_ hold97/Z _7224_/RN _6772_/CLK hold96/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3984_ _3983_/Z _6658_/Q _3984_/S _3984_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5723_ _5852_/I0 hold819/Z _5727_/S _5723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5654_ hold233/Z _5681_/I1 _5655_/S _7010_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4605_ _4638_/A2 _4648_/B _5356_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_175_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5585_ hold929/Z _5795_/I0 hold34/Z _5585_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold300 _4126_/Z _6680_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold311 _6754_/Q hold311/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4536_ _5414_/A2 _5295_/A2 _4472_/B _5399_/A1 _4536_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold322 _5499_/Z _6879_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold333 _7102_/Q hold333/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold344 _5707_/Z _7057_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_132_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold355 _7176_/Q hold355/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_117_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7255_ _7255_/D _7255_/RN _7257_/CLK _7255_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold366 _5705_/Z _7055_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4467_ _4467_/A1 _4555_/B _4467_/B _4690_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_131_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold377 _6921_/Q hold377/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold388 _3480_/Z _3481_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6206_ _6529_/S _7248_/Q _6206_/B _6207_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold399 _5578_/Z _6942_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3418_ _3417_/Z _7305_/Q _3988_/S _7305_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7186_ _7186_/D _7211_/RN _7186_/CLK _7186_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4398_ _5002_/A3 _5002_/A4 _5165_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_86_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6137_ _7246_/Q _6136_/Z _6558_/S _7246_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold1000 _5721_/Z _7069_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3349_ _7161_/Q _3349_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1011 _7068_/Q _5720_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1022 _5868_/Z _7199_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1033 _6989_/Q _5631_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1044 _6868_/Q _3965_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_85_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6068_ _7145_/Q _6068_/A2 _6210_/B _6164_/A2 _6076_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_133_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold1055 _3475_/Z _3476_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1066 _6892_/Q _5516_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold1077 _7282_/Q _3466_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5019_ _5191_/A3 _5019_/A2 _5390_/A1 _5019_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XTAP_2516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet1202_454 net1202_487/I _6711_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_186_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1202_465 _4073__41/I _6700_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_157_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1202_476 net1202_481/I _6689_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1202_487 net1202_487/I _6678_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_158_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1202_498 net802_90/I _6667_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5370_ _5370_/A1 _5172_/B _5370_/B _5370_/C _5371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_4321_ _5867_/I0 hold571/Z _4322_/S _4321_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7040_ _7040_/D _7098_/RN _7040_/CLK _7040_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4252_ _5890_/I0 hold228/Z _4252_/S _4252_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4183_ hold827/Z _4360_/I1 _4184_/S _4183_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6824_ _6824_/D _6839_/RN _6824_/CLK _6824_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_24_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6755_ _6755_/D _7257_/RN _6755_/CLK _6755_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3967_ _3427_/Z _6663_/Q _6664_/Q _3967_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_32_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5706_ hold341/Z _5724_/I0 _5709_/S _5706_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6686_ _6686_/D _7296_/RN _6686_/CLK _6686_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3898_ _6565_/I0 _6868_/Q _3898_/S _3898_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_177_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5637_ _5775_/I0 hold653/Z _5637_/S _5637_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5568_ _5778_/I0 hold631/Z _5574_/S _5568_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold130 _7114_/Q hold130/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7307_ _7307_/I _7307_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold141 _4131_/Z _6684_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_137_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4519_ _5170_/A2 _5269_/A2 _5328_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold152 hold152/I hold152/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_5499_ hold321/Z _5538_/I1 hold29/Z _5499_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold163 _4122_/Z _6676_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold174 _4263_/Z _6777_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold185 _7130_/Q hold185/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7238_ _7238_/D _7238_/RN _7260_/CLK _7238_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_120_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold196 _4266_/Z _6780_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_137_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout610 _4422_/Z _5290_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout621 _4715_/A1 _4835_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_104_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout632 input95/Z _3401_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout643 _7297_/RN _6847_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_58_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout654 fanout655/Z _7215_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_7169_ _7169_/D _7218_/RN _7169_/CLK _7169_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
Xfanout665 _7024_/RN _7002_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout676 fanout677/Z _7207_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_59_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout687 _7177_/RN _7219_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout698 fanout714/Z _7149_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_100_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4073__30 _4073__46/I _7195_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4870_ _5293_/B _4844_/Z _5215_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_2880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__41 _4073__41/I _7184_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3821_ _4185_/A2 _3653_/Z _3947_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_60_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6540_ _6867_/Q _6540_/A2 _6293_/Z _6719_/Q _6540_/C _6547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3752_ _6975_/Q _3923_/A2 _3959_/B1 _6669_/Q _5656_/A1 _7015_/Q _3753_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xclkbuf_leaf_66__1359_ clkbuf_4_13_0__1359_/Z net952_238/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_146__1359_ net1152_451/I net1202_491/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_159_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6471_ _6946_/Q _6245_/Z _6273_/Z _6978_/Q _7124_/Q _6288_/Z _6472_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3683_ _7250_/Q _6898_/Q _6900_/Q _3683_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5422_ _5034_/B _4866_/Z _5422_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
Xoutput202 _3376_/ZN mgmt_gpio_oeb[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput213 _4068_/Z mgmt_gpio_out[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput224 _6742_/Q mgmt_gpio_out[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5353_ _5353_/A1 _5387_/A2 _5353_/B _5354_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xoutput235 _4054_/Z mgmt_gpio_out[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_126_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput246 _4057_/Z mgmt_gpio_out[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput257 _6886_/Q pll90_sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput268 _6883_/Q pll_sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4304_ _6829_/Q _6563_/A2 _4312_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xoutput279 _6667_/Q pll_trim[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5284_ _5284_/A1 _5369_/B _5284_/A3 _5277_/I _5286_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_4_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7023_ _7023_/D _7125_/RN _7023_/CLK _7023_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_101_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4235_ _4234_/Z hold369/Z _4245_/S _4235_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4166_ _5538_/I1 hold899/Z _4166_/S _4166_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4097_ _4097_/A1 _4415_/B _6828_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6807_ _6807_/D _7262_/CLK _6807_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4999_ _4999_/A1 _4999_/A2 _4998_/Z _5341_/B _5000_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_6738_ _6738_/D _6771_/RN _6738_/CLK _6738_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_177_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6669_ _6669_/D fanout659/Z _6669_/CLK _6669_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_137_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout440 _5884_/A3 _5848_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_59_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout451 _6233_/ZN _6533_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout462 _5478_/A2 _5287_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xfanout473 _4546_/Z _5146_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_150_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout484 _5083_/B _5080_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_19_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout495 _5555_/I0 _5681_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4020_ _4014_/Z _4020_/A2 _5951_/B _4003_/Z _4021_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_49_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5971_ _5991_/A2 _6021_/A4 _6211_/B1 _6139_/A2 _5971_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4922_ _4373_/Z _4385_/Z _4922_/A3 _4922_/A4 _4923_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_127_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4853_ _4853_/A1 _4873_/A3 _5228_/A3 _3406_/I _4853_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_20_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3804_ _6842_/Q _3930_/B1 _3884_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4784_ _4960_/A1 _3402_/I _3403_/I _3404_/I _4784_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_147_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6523_ _6866_/Q _6540_/A2 _6290_/Z _6708_/Q _6526_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3735_ _7113_/Q _3917_/A2 _5674_/A1 _7031_/Q _3735_/C _3760_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_147_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6454_ _7100_/Q _6250_/Z _6302_/Z _7092_/Q _6292_/Z _7148_/Q _6466_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_134_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3666_ _6929_/Q _3935_/A2 _5656_/A1 _7017_/Q _3667_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_106_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5405_ _5454_/A1 _4791_/Z _5126_/I _5406_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6385_ _6385_/A1 _6385_/A2 _6385_/A3 _6384_/Z _6385_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3597_ hold56/I _3546_/Z _3945_/C2 hold70/I _3913_/A2 input19/Z _3601_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_115_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5336_ _5412_/A1 _5412_/A3 _5338_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5267_ _4898_/C _5428_/A4 _4893_/Z _5267_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_130_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7006_ _7006_/D _7258_/RN _7006_/CLK _7006_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4218_ _4217_/Z hold201/Z _4228_/S _4218_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5198_ _5309_/B2 _5205_/A1 _5351_/C _5205_/B1 _5198_/C _5476_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4149_ _3507_/Z _5731_/A2 _5794_/A3 _4157_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_28_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet952_250 net952_250/I _6975_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3520_ _5884_/A1 _3519_/Z _3520_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_116_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold707 _7213_/Q hold707/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_157_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold718 _5855_/Z _7188_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold729 _7146_/Q hold729/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_170_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3451_ _3451_/I0 _4056_/I1 _6730_/Q _3451_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3382_ _6785_/Q _6528_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_6170_ _6971_/Q _5979_/Z _5981_/Z _6939_/Q _5996_/Z _7085_/Q _6181_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_124_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5121_ _5121_/A1 _4876_/C _5457_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_85_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5052_ _4936_/I _5051_/Z _5064_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4003_ _5954_/A3 _7225_/Q _7226_/Q _7223_/Q _4003_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_38_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet802_59 net802_67/I _7166_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5954_ _7223_/Q _5954_/A2 _5954_/A3 _5951_/B _5954_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_52_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4905_ _4944_/A1 _4495_/Z _5263_/A2 _5324_/A1 _4905_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_178_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5885_ _5885_/I0 _5885_/I1 _5892_/S _5885_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4836_ _5420_/A3 _4549_/Z _4836_/A3 _4836_/A4 _4836_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_14_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4767_ _5226_/A1 _4764_/Z _5118_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6506_ _6820_/Q _6531_/A2 _6552_/A2 _6847_/Q _6512_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3718_ input16/Z _3913_/A2 _3945_/B1 _7090_/Q _3719_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_135_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4698_ _5097_/A1 _4704_/A2 _4698_/B _5094_/B _4714_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_161_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6437_ _6437_/I _6438_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3649_ _3648_/Z _3649_/I1 _3899_/S _6874_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6368_ _7145_/Q _6292_/Z _6383_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_1_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet902_180 _4073__27/I _7045_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet902_191 net902_191/I _7034_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5319_ _5392_/B _4801_/Z _5319_/A3 _5319_/A4 _5319_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_142_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6299_ _5946_/S _6299_/A2 _6452_/A4 _6302_/A4 _6299_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold12 hold12/I hold12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_88_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold23 hold23/I hold23/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold34 hold34/I hold34/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_60_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold45 hold45/I hold45/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold56 hold56/I hold56/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_29_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold67 hold67/I hold67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold78 hold78/I hold78/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold89 hold89/I hold89/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_17_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1052_330 net902_179/I _6895_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xnet1052_341 net1052_346/I _6884_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_9 _4108_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_2__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7269_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5670_ hold525/Z _5781_/I0 _5673_/S _5670_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4621_ _4367_/Z _4555_/B _5291_/C _5353_/A1 _5353_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_30_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4552_ _4549_/Z _5373_/A2 _5011_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_144_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold504 _5607_/Z _6968_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold515 _6961_/Q hold515/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3503_ _3680_/A3 _3500_/Z _3503_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7271_ _7271_/D _7278_/RN _7279_/CLK _7271_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold526 _5670_/Z _7024_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4483_ _4489_/A1 _4692_/B _4483_/B _4687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xhold537 _6724_/Q hold537/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold548 _7217_/Q hold548/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6222_ _6823_/Q _5964_/Z _5999_/Z _6848_/Q _6729_/Q _6000_/Z _6228_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold559 _6893_/Q hold559/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3434_ _3442_/B _3409_/Z _3434_/B _3435_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_100_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6153_ _6946_/Q _5972_/Z _6021_/Z _7002_/Q _6155_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3365_ _7039_/Q _3365_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5104_ _5104_/A1 _5139_/A3 _5094_/B _5104_/A4 _5104_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6084_ _6084_/A1 _6084_/A2 _6084_/A3 _6084_/A4 _6084_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_39_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3296_ _7294_/Q _4084_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5035_ _5035_/A1 _5032_/Z _5204_/C _5035_/A4 _5035_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_73_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6986_ _6986_/D _7124_/RN _6986_/CLK _6986_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_40_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5937_ _6279_/A3 _7233_/Q _6302_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_40_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5868_ _5877_/I0 _5868_/I1 _5874_/S _5868_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4819_ _5290_/A1 _4624_/Z _4673_/Z _4483_/B _4819_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5799_ _5871_/I0 hold309/Z hold12/Z _5799_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet1002_260 _4073__42/I _6965_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1002_271 net952_228/I _6954_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_166_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1002_282 net1052_328/I _6943_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1002_293 net802_83/I _6932_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput102 wb_adr_i[16] _4391_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_1_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput113 wb_adr_i[26] _4031_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput124 wb_adr_i[7] input124/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput135 wb_dat_i[16] _6579_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput146 wb_dat_i[26] _6585_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput157 wb_dat_i[7] _3400_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6840_ _6840_/D _6933_/RN _6840_/CLK _6840_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_22_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6771_ _6771_/D _6771_/RN _6771_/CLK _6771_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3983_ _6659_/Q _3972_/Z _3983_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5722_ _5860_/I0 hold120/Z _5727_/S _5722_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5653_ hold307/Z _5827_/I0 _5655_/S _5653_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4604_ _4449_/B _4604_/A2 _4604_/A3 _4604_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_5584_ _5584_/A1 _5674_/A2 hold34/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_7_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold301 _7201_/Q hold301/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4535_ _5414_/A2 _4534_/Z _5323_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold312 _4228_/Z _6754_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_172_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold323 _6742_/Q hold323/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold334 _5759_/Z _7102_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold345 _7107_/Q hold345/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7254_ _7254_/D _7257_/RN _7257_/CLK _7254_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold356 _5842_/Z _7176_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4466_ _5270_/A2 _4367_/Z _4363_/Z _4690_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xhold367 _6782_/Q hold367/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold378 _5554_/Z _6921_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_132_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6205_ _6193_/Z _6204_/Z _6528_/B1 _6118_/B _6555_/C _6206_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold389 _3508_/Z hold389/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3417_ _3416_/Z _7304_/Q _3984_/S _3417_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7185_ _7185_/D _7185_/RN _7185_/CLK _7185_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4397_ _5002_/A3 _5002_/A4 _4397_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_98_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6136_ _6136_/I0 _7245_/Q _6529_/S _6136_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3348_ _7169_/Q _3348_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1001 _7175_/Q _5841_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1012 _5720_/Z _7068_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1023 _7214_/Q _5885_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1034 _5631_/Z _6989_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6067_ _6067_/A1 _5991_/Z _6072_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold1045 _6875_/Q _3611_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_86_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1056 _7303_/Q _3498_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1067 _6952_/Q hold556/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5018_ _5389_/B _5439_/B2 _5018_/B _5390_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold1078 _6947_/Q _5583_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_2506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6969_ _6969_/D _7122_/RN _6969_/CLK _6969_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_13_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold890 _5601_/Z _6963_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_174_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet1202_455 net1202_487/I _6710_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1202_466 net802_91/I _6699_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1202_477 net1202_481/I _6688_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1202_488 net1202_489/I _6677_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1202_499 net1202_499/I _6666_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_185_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4320_ _5848_/A3 _3535_/Z hold389/Z _5620_/A4 _4322_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_172_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4251_ _5889_/I0 hold104/Z _4252_/S _4251_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4182_ _4182_/A1 _6611_/A2 _4184_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_79_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_106__1359_ clkbuf_4_5_0__1359_/Z net802_87/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_68_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_89__1359_ clkbuf_4_7_0__1359_/Z net952_208/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_55_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6823_ _6823_/D _6839_/RN _6823_/CLK _6823_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6754_ _6754_/D _7124_/RN _6754_/CLK _6754_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_189_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3966_ _3966_/I _6868_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5705_ hold365/Z _5852_/I0 _5709_/S _5705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6685_ _6685_/D _7296_/RN _6685_/CLK _6685_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_31_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3897_ _3897_/A1 _3897_/A2 _3855_/Z _3896_/Z _6565_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_177_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5636_ _5855_/I0 hold703/Z _5637_/S _5636_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5567_ _5795_/I0 hold745/Z _5574_/S _5567_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold120 _7070_/Q hold120/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold131 _5772_/Z _7114_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4518_ _4835_/A2 _3403_/I _5269_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_2_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold142 _6860_/Q hold142/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_5498_ hold193/Z _5537_/I1 hold29/Z _5498_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold153 hold153/I hold153/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold164 _6766_/Q hold164/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold175 _6899_/Q hold175/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7237_ _7237_/D _7237_/RN _7257_/CLK _7237_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
Xhold186 _5790_/Z _7130_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4449_ _4501_/A1 _5201_/A1 _4449_/B _4451_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xhold197 _6751_/Q hold197/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xfanout600 _4643_/A4 _4635_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_59_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout611 _5201_/A1 _5464_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout622 _3404_/ZN _4715_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout633 _6907_/RN _6894_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout644 _6933_/RN _6839_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_7168_ _7168_/D fanout677/Z _7168_/CLK _7168_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_101_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout655 fanout656/Z fanout655/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout666 _7024_/RN _7238_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6119_ _7155_/Q _5960_/Z _6133_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout677 fanout685/Z fanout677/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_86_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout688 _7193_/RN _7177_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7099_ _7099_/D _7211_/RN _7099_/CLK _7099_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_74_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout699 _7257_/RN _7255_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_3004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4073__20 net802_68/I _7205_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4073__31 _4073__31/I _7194_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__42 _4073__42/I _7183_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3820_ _5510_/A2 _3578_/Z _4274_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_178_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3751_ _3751_/A1 _3751_/A2 _3732_/Z _3751_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_174_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6470_ _7050_/Q _6550_/A2 _6251_/Z _6986_/Q _6550_/C1 _6954_/Q _6472_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_119_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3682_ _7001_/Q _5638_/A1 _3912_/B1 _6888_/Q _3686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_118_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5421_ _5420_/Z _5421_/A2 _5421_/A3 _5421_/A4 _5489_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_145_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput203 _3375_/ZN mgmt_gpio_oeb[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput214 _4067_/Z mgmt_gpio_out[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5352_ _5191_/Z _5352_/A2 _5285_/B _5020_/Z _5352_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xoutput225 hold82/I mgmt_gpio_out[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput236 hold90/I mgmt_gpio_out[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput247 _4075_/Z pad_flash_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput258 _6887_/Q pll90_sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4303_ hold877/Z _6613_/I1 _4303_/S _4303_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput269 _6884_/Q pll_sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5283_ _5278_/C _4554_/Z _5283_/B _5471_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_142_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7022_ _7022_/D _7122_/RN _7022_/CLK _7022_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_87_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4234_ hold132/Z _5860_/I0 _4242_/S _4234_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4165_ _4103_/I hold965/Z _4166_/S _4165_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4096_ _4097_/A1 _4096_/A2 _6829_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_169_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6806_ _6806_/D _7258_/CLK _6806_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4998_ _5340_/A1 _4998_/A2 _5262_/A2 _5343_/A2 _4998_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_11_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3949_ _3949_/A1 _3949_/A2 _3949_/A3 _3949_/A4 _3949_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6737_ _6737_/D _6771_/RN _6737_/CLK _6737_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_17_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6668_ _6668_/D fanout659/Z _6668_/CLK _6668_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_104_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5619_ _5784_/I0 hold973/Z _5619_/S _5619_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6599_ _6599_/I0 _7276_/Q _6602_/S _7276_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout430 _6168_/C _6118_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_132_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout441 hold11/Z _5884_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout452 _4784_/Z _5228_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_63_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout463 _4683_/Z _5478_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_171_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout474 _4532_/ZN _5364_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout485 _4313_/Z _6601_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xfanout496 _5855_/I0 _5891_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_72__1359_ clkbuf_4_14_0__1359_/Z net802_52/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5970_ _7102_/Q _5967_/Z _5969_/Z _7118_/Q _5974_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4921_ _4920_/Z _4890_/I _4926_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_61_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4852_ _4852_/A1 _5106_/A2 _4852_/A3 _4855_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3803_ _4353_/A1 _3680_/Z _3930_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_127_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4783_ _4836_/A4 _4530_/I _5137_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_165_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6522_ _6696_/Q _6532_/A2 _6302_/Z _6712_/Q _6526_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_159_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3734_ _3734_/I _3735_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6453_ _7066_/Q _6257_/Z _6536_/B1 _7042_/Q _6300_/Z _7108_/Q _6466_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3665_ _7009_/Q _3934_/A2 _3954_/A2 _6993_/Q _3674_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_106_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5404_ _5404_/A1 _5314_/Z _5404_/A3 _5404_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_118_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6384_ _6384_/A1 _6384_/A2 _6380_/Z _6383_/Z _6384_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3596_ _3592_/Z _3596_/A2 _3596_/A3 _3596_/A4 _3596_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5335_ _4908_/Z _5245_/Z _5481_/B1 _4905_/Z _5335_/C _5447_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_114_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5266_ _5265_/Z _5341_/B _4994_/Z _5266_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_142_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7005_ _7005_/D _7098_/RN _7005_/CLK _7005_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4217_ hold189/Z _5797_/I0 _4227_/S _4217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5197_ _5346_/A2 _5349_/A1 _5276_/C _5205_/A1 _5197_/C _5390_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4148_ hold661/Z _4361_/I1 _4148_/S _4148_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4079_ _4079_/I _4079_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet952_240 net952_250/I _6985_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet952_251 net952_251/I _6974_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_109_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_1__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7258_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_182_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold708 _5883_/Z _7213_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_7_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold719 _7205_/Q hold719/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3450_ _3450_/A1 _3450_/A2 _7292_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_6_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3381_ _6931_/Q _6500_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_171_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5120_ _5118_/Z _5238_/A1 _5127_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5051_ _4698_/B _5343_/A1 _5051_/S _5051_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_112_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4002_ _7225_/Q _7226_/Q _5954_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_37_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5953_ _5953_/I0 _7239_/Q _5955_/S _7239_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4904_ _5263_/A2 _4903_/Z _5255_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5884_ _5884_/A1 _5884_/A2 _5884_/A3 _5892_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_33_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4835_ _4555_/C _4835_/A2 _5129_/A3 _5420_/A2 _5368_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_178_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4766_ _4766_/A1 _4766_/A2 _4762_/Z _4765_/Z _4770_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_140_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6505_ _6853_/Q _6550_/A2 _6297_/Z _7076_/Q _6512_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3717_ _6928_/Q _3935_/A2 _3943_/A2 _7072_/Q _6895_/Q _5528_/S _3719_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_174_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4697_ _4467_/B _4463_/Z _5302_/B _5099_/A2 _4697_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_106_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6436_ _7147_/Q _6292_/Z _6300_/Z _7107_/Q _6437_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_20_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3648_ _6570_/I0 _6873_/Q _3898_/S _3648_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6367_ _7253_/Q _6367_/I1 _6450_/S _7253_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3579_ _5517_/A2 _3578_/Z _3959_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xnet902_170 net902_170/I _7055_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_181 net902_181/I _7044_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_192 net952_216/I _7033_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5318_ _5318_/A1 _5314_/Z _5316_/Z _5318_/A4 _5320_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_88_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6298_ _7158_/Q _6296_/Z _6297_/Z _6698_/Q _6298_/C _6307_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_130_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold13 hold13/I hold13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold24 hold24/I hold24/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_29_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5249_ _5410_/A1 _5245_/Z _5250_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_29_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold35 hold35/I hold35/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_57_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold46 hold46/I hold46/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold57 hold57/I hold57/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold68 hold68/I hold68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_29_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold79 hold79/I hold79/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_188_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1052_320 net852_136/I _6905_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_331 net1152_427/I _6894_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xnet1052_342 net1052_346/I _6883_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_131_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4620_ _4557_/Z _4604_/Z _5353_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4551_ _4930_/A1 _3404_/I _5129_/A4 _3402_/I _4551_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_156_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3502_ hold144/Z hold211/Z _3904_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold505 _7054_/Q hold505/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7270_ _7270_/D _7278_/RN _7279_/CLK hold62/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold516 _5599_/Z _6961_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4482_ _4381_/Z _4485_/A2 _4390_/Z _5170_/A3 _4486_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold527 _6944_/Q hold527/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_7_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold538 _4186_/Z _6724_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6221_ _6725_/Q _5984_/Z _5997_/Z _6717_/Q _6695_/Q _5980_/Z _6228_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold549 _5888_/Z _7217_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3433_ _3427_/Z _3433_/A2 _3433_/B _3435_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_103_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6152_ _6152_/A1 _6152_/A2 _6152_/A3 _6152_/A4 _6152_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3364_ _7047_/Q _3364_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ _5103_/A1 _5101_/Z _5103_/A3 _5308_/A2 _5108_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6083_ _6975_/Q _5964_/Z _5999_/Z _7031_/Q _6084_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3295_ _7283_/Q _4022_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ _5190_/A2 _4604_/Z _5003_/Z _5034_/B _5204_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_38_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6985_ _6985_/D _7122_/RN _6985_/CLK _6985_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5936_ _5957_/I1 _7233_/Q _7232_/Q _5936_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_5867_ _5867_/I0 _5867_/I1 _5874_/S _5867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4818_ _4624_/Z _5142_/A3 _5313_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5798_ _5798_/I0 hold581/Z hold12/Z _7137_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet1002_261 net952_245/I _6964_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1002_272 net802_78/I _6953_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_182_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet1002_283 net1052_328/I _6942_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4749_ _5401_/A2 _5230_/B _5313_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_175_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet1002_294 net902_194/I _6931_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6419_ _6500_/C _7254_/Q _6419_/B _6420_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_150_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput103 wb_adr_i[17] _4391_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_130_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput114 wb_adr_i[27] _4027_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput125 wb_adr_i[8] _4388_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput136 wb_dat_i[17] _6582_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput147 wb_dat_i[27] _6588_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput158 wb_dat_i[8] _6579_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_173_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3982_ _3981_/Z _6660_/Q _3988_/S _6660_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6770_ hold95/Z _6771_/RN _6770_/CLK hold94/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_189_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5721_ _5886_/I0 hold999/Z _5727_/S _5721_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5652_ _5652_/I0 _5781_/I0 _5655_/S _5652_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4603_ _4580_/B _4604_/A3 _5351_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5583_ _5583_/I0 hold6/Z _5583_/S hold7/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_129__1359_ net1152_446/I net1202_489/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_49__1359_ clkbuf_4_11_0__1359_/Z _4073__45/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4534_ _4782_/A1 _4736_/A3 _4736_/A1 _4752_/A2 _4534_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_7_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold302 _5870_/Z _7201_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold313 _6688_/Q hold313/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold324 _4211_/Z _6742_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold335 _6735_/Q hold335/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold346 _5764_/Z _7107_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4465_ _5315_/A1 _4481_/A2 _4473_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_116_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7253_ _7253_/D _7253_/RN _7257_/CLK _7253_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold357 _6896_/Q hold357/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_132_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold368 _4268_/Z _6782_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6204_ _6198_/Z _6201_/Z _6204_/A3 _6204_/A4 _6204_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold379 _7118_/Q hold379/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3416_ _7305_/Q _3415_/Z _3416_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7184_ _7184_/D fanout677/Z _7184_/CLK _7184_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4396_ _5385_/A1 _4385_/Z _4922_/A3 _4424_/B _5002_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6135_ _6127_/Z _6134_/Z _6447_/B1 _6118_/B _6136_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3347_ _7177_/Q _3732_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1002 _5841_/Z _7175_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1013 _7158_/Q _5822_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1024 _5885_/Z _7214_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6066_ _7023_/Q _6164_/A2 _6164_/B1 _6991_/Q _6067_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold1035 _7160_/Q _5824_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1046 _6731_/Q _4023_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_73_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold1057 _6662_/Q _3483_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_5017_ _5017_/A1 _5197_/C _5019_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_3219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold1068 _6731_/Q _3312_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1079 _6983_/Q _5624_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_2507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6968_ _6968_/D _7260_/RN _6968_/CLK _6968_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_53_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5919_ _6002_/A3 _6015_/A3 _5984_/A1 _5957_/I1 _5919_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6899_ _6899_/D _7238_/RN _6899_/CLK _6899_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xhold880 _5828_/Z _7164_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold891 _7018_/Q hold891/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_67_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet1202_456 net902_189/I _6709_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1202_467 net952_245/I _6698_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1202_478 net1202_481/I _6687_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1202_489 net1202_489/I _6676_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_157_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4250_ _5834_/I0 hold164/Z _4252_/S _4250_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4181_ _4361_/I1 hold871/Z _4181_/S _4181_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6822_ _6822_/D _6847_/RN _6822_/CLK _6822_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6753_ _6753_/D _6854_/RN _6753_/CLK _6753_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3965_ _6564_/I0 _3965_/A2 _3965_/B1 _3899_/S _3966_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_32_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5704_ hold505/Z _5869_/I0 _5709_/S _5704_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3896_ _3860_/Z _3869_/Z _3885_/Z _3895_/Z _3896_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6684_ _6684_/D _7296_/RN _6684_/CLK _6684_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_5635_ _5818_/I0 hold765/Z _5637_/S _5635_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5566_ _5875_/A3 _5776_/A1 hold389/Z _5620_/A4 _5574_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_145_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold110 _6887_/Q hold110/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold121 _5722_/Z _7070_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7305_ _7305_/D _6657_/Z _4072_/B2 _7305_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
Xhold132 _6918_/Q hold132/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_132_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4517_ _5165_/A4 _5003_/A2 _4491_/B _4517_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_5497_ hold153/I hold28/Z _5647_/A2 _5620_/A4 hold29/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_117_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold143 _3496_/Z _3497_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold154 _5648_/S _5655_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold165 _4250_/Z _6766_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold176 _5526_/Z _6899_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7236_ _7236_/D _7075_/RN _4067_/I1 _7236_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_104_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4448_ _3401_/I _5288_/C _4369_/Z _4522_/A2 _4451_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold187 _6781_/Q hold187/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_120_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout601 _4643_/A4 _5278_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xhold198 _4222_/Z _6751_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout612 _5076_/A1 _5201_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_144_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout623 _3403_/ZN _5129_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_144_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout634 _6907_/RN _6854_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_58_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7167_ _7167_/D _7218_/RN _7167_/CLK _7167_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_99_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4379_ _4853_/A1 _5201_/A1 _4604_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xfanout645 _7297_/RN _6933_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout656 fanout685/Z fanout656/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout667 _7024_/RN _7122_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6118_ _7057_/Q _5924_/Z _6118_/B _6127_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout678 _7163_/RN _7258_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_7098_ _7098_/D _7098_/RN _7098_/CLK _7098_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout689 _6915_/RN _7193_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_86_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6049_ _6942_/Q _5972_/Z _6021_/Z _6998_/Q _6049_/C _6053_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_3027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_112__1359_ clkbuf_4_4_0__1359_/Z net802_90/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_95__1359_ clkbuf_4_5_0__1359_/Z net1152_425/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_136_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073__10 _4073__7/I _7215_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4073__21 net802_68/I _7204_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4073__32 _4073__32/I _7193_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__43 net802_82/I _7182_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3750_ _7007_/Q _3934_/A2 _5638_/A1 _6999_/Q _3916_/B1 _6881_/Q _3751_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_13_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3681_ _5510_/A2 _3680_/Z _3912_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_186_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5420_ _5420_/A1 _5420_/A2 _5420_/A3 _5420_/A4 _5420_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_185_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput204 _3374_/ZN mgmt_gpio_oeb[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5351_ _5356_/A1 _5387_/A2 _5356_/B _5351_/C _5352_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_57_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput215 _4066_/Z mgmt_gpio_out[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput226 hold74/I mgmt_gpio_out[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_182_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput237 _4055_/Z mgmt_gpio_out[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput248 _4094_/ZN pad_flash_clk_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4302_ hold941/Z _6612_/I1 _4303_/S _4302_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput259 _6888_/Q pll90_sel[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5282_ _5281_/C _4467_/B _5399_/A2 _5478_/A2 _5283_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7021_ _7021_/D _7155_/RN _7021_/CLK _7021_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4233_ _4232_/Z hold207/Z _4245_/S _4233_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4164_ _5520_/C _5821_/A2 _5517_/A3 _5517_/A1 _4166_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_110_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4095_ _4097_/A1 _4900_/B _6831_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_70_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6805_ _6805_/D _7258_/CLK _6805_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4997_ _5146_/A1 _5329_/A2 _4997_/B _4997_/C _4999_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_168_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6736_ _6736_/D _6771_/RN _6736_/CLK _6736_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3948_ input43/Z _4210_/S _4194_/A1 input52/Z _3948_/C1 input61/Z _3949_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_139_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6667_ _6667_/D _6892_/RN _6667_/CLK _6667_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3879_ _7087_/Q _3945_/B1 _3952_/A2 _7045_/Q _3950_/C1 _6844_/Q _3880_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_176_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5618_ _5681_/I1 hold737/Z _5619_/S _5618_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6598_ _6598_/A1 _6601_/A2 _6598_/B _6599_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_3_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5549_ hold64/Z hold116/Z _5556_/S _5549_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_0__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7262_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_133_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1102_400 net1102_400/I _6774_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7219_ _7219_/D _7219_/RN _7219_/CLK _7219_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout420 _6261_/Z _6544_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_87_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout431 _4817_/Z _5142_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_48_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout442 hold10/Z hold11/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout453 _4784_/Z _5164_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout464 _4675_/Z _5380_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_150_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout475 _4532_/ZN _5414_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout486 _5811_/I0 _5784_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_19_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout497 _5555_/I0 _5855_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_171_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4920_ _5130_/B2 _4960_/A1 _4367_/Z _4920_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_80_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4851_ _5287_/C _4833_/Z _4852_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3802_ _4332_/A1 _3540_/Z _3925_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_21_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4782_ _4782_/A1 _5236_/A1 _5302_/B _5099_/A1 _5213_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6521_ _6521_/A1 _6521_/A2 _6521_/A3 _6521_/A4 _6521_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_158_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3733_ _7193_/Q _3909_/A2 _5683_/A1 _7039_/Q _3952_/A2 _7047_/Q _3734_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_146_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6452_ _7074_/Q _6452_/A2 _6452_/A3 _6452_/A4 _6456_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3664_ input17/Z _3913_/A2 _5674_/A1 _7033_/Q _3674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5403_ _5403_/A1 _5403_/A2 _5456_/A2 _5403_/B2 _5403_/C _5404_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_174_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3595_ _6995_/Q _3954_/A2 _3927_/A2 _6705_/Q _3596_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6383_ _6383_/A1 _6383_/A2 _6383_/A3 _6383_/A4 _6383_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_155_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5334_ _5334_/A1 _5334_/A2 _5334_/A3 _5334_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_86_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5265_ _5265_/A1 _4991_/C _5392_/B _5265_/A4 _5265_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_134_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7004_ _7004_/D _7090_/RN _7004_/CLK _7004_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4216_ _4215_/Z hold315/Z _4228_/S _4216_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5196_ _5347_/A1 _5437_/A1 _5195_/Z _5347_/A3 _5196_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_56_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4147_ hold671/Z _5822_/I0 _4148_/S _4147_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4078_ _4081_/A1 input86/Z _4079_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_36_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6719_ _6719_/D _6847_/RN _6719_/CLK _6719_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_11_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet952_230 _4073__12/I _6995_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet952_241 net952_241/I _6984_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold709 _6704_/Q hold709/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_156_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3380_ _6930_/Q _6473_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_124_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5050_ _5343_/A2 _5389_/A2 _5078_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_46_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4001_ _4001_/I _6836_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5952_ _6746_/Q _3324_/I _5952_/A3 _5952_/B _5955_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_18_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4903_ _4903_/A1 _4407_/Z _4495_/Z _5259_/A1 _4903_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_179_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5883_ _5892_/I0 hold707/Z _5883_/S _5883_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4834_ _4834_/A1 _4834_/A2 _4846_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_33_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4765_ _4765_/A1 _4774_/A3 _5478_/B1 _5226_/C _4765_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_147_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6504_ _6789_/Q _6551_/A2 _6543_/A2 _6851_/Q _6512_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3716_ _7130_/Q _3930_/A2 _3925_/A2 input7/Z hold153/I _3904_/A2 _3719_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_4696_ _5099_/A2 _4695_/Z _4704_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_107_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6435_ _7187_/Q _6532_/A2 _6299_/Z _7057_/Q _6993_/Q _6237_/Z _6439_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3647_ _3647_/A1 _3625_/Z _3646_/Z _3647_/A4 _6570_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_161_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6366_ _6366_/I _6367_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_160 net802_54/I _7065_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3578_ _3653_/A1 _3904_/A3 hold144/I _3500_/Z _3578_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xnet902_171 _4073__41/I _7054_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_182 net802_60/I _7043_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_193 net952_225/I _7032_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5317_ _5317_/A1 _5454_/A1 _5318_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_143_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6297_ _6300_/A2 _6484_/A3 _6300_/A4 _5942_/S _6297_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold14 hold14/I hold14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_5248_ _5246_/Z _5248_/A2 _5248_/A3 _5056_/C _5248_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold25 hold25/I hold25/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_130_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold36 hold36/I hold36/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_29_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold47 hold47/I hold47/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_102_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold58 hold58/I hold58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold69 hold69/I hold69/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_96_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5179_ _5240_/B _5343_/A2 _5179_/B _5242_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_60_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1052_310 net1052_312/I _6915_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_43_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1052_321 net852_136/I _6904_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_332 net1202_491/I _6893_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xnet1052_343 net1202_453/I _6882_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_61_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4550_ _5269_/A1 _5269_/A2 _5368_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3501_ _3499_/I _3305_/I _4113_/S _3501_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold506 _5704_/Z _7054_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4481_ _4481_/A1 _4481_/A2 _4486_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold517 _6845_/Q hold517/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold528 _5580_/Z _6944_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold539 _6977_/Q hold539/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6220_ _6217_/Z _6220_/A2 _6220_/A3 _6220_/A4 _6220_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_116_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3432_ _3432_/I _7299_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6151_ _7148_/Q _5987_/Z _6015_/Z _7010_/Q _6152_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3363_ _7055_/Q _3363_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _5367_/A2 _5142_/A3 _5103_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_44_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3294_ _7300_/Q _4081_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_6082_ _7169_/Q _6006_/Z _6014_/Z hold88/I _6084_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ _5035_/A4 _5032_/Z _5388_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_26_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6984_ _6984_/D _7122_/RN _6984_/CLK _6984_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_80_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5935_ _6282_/A2 _6279_/A3 _6300_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_22_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5866_ _5875_/A1 _3507_/Z _5866_/A3 _5874_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_90_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4817_ _5420_/A3 _5369_/A1 _3402_/I _5269_/A2 _4817_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_178_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5797_ _5797_/I0 hold428/Z hold12/Z _5797_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet1002_262 net902_187/I _6963_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1002_273 net952_241/I _6952_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4748_ _5236_/A1 _5478_/A3 _5099_/A1 _5226_/C _4748_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xclkbuf_4_11_0__1359_ clkbuf_0__1359_/Z clkbuf_4_11_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet1002_284 net1202_463/I _6941_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1002_295 net902_191/I _6930_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4679_ _4670_/Z _5451_/C _4685_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_174_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6418_ _6411_/Z _6417_/Z _6418_/B1 _6286_/Z _6529_/S _6419_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_116_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6349_ _7200_/Q _6540_/A2 _6532_/A2 _7184_/Q _6296_/Z _7160_/Q _6356_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_88_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput104 wb_adr_i[18] _4391_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xclkbuf_0__1359_ _4072_/ZN clkbuf_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput115 wb_adr_i[28] _4027_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput126 wb_adr_i[9] _4388_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput137 wb_dat_i[18] _6585_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput148 wb_dat_i[28] _6591_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput159 wb_dat_i[9] _6582_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_3981_ _3981_/A1 _3981_/A2 _3981_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5720_ _5867_/I0 _5720_/I1 _5727_/S _5720_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5651_ hold232/Z _5879_/I0 _5655_/S _7007_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4602_ _5399_/A1 _5399_/A2 _5290_/A2 _5364_/B _5285_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_148_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5582_ hold168/Z _5645_/I1 _5583_/S _5582_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4533_ _4736_/A3 _4690_/C _4713_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold303 _6671_/Q hold303/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_156_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold314 _4135_/Z _6688_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold325 _7103_/Q hold325/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7252_ _7252_/D _7257_/RN _7257_/CLK _7252_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4464_ _5420_/A4 _4873_/A2 _4460_/B _4752_/A2 _4464_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold336 _4197_/Z _6735_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold347 _7106_/Q hold347/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold358 _5523_/Z _6896_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6203_ _6724_/Q _5984_/Z _6000_/Z _6728_/Q _6710_/Q _6006_/Z _6204_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_104_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold369 _6757_/Q hold369/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_131_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3415_ _7304_/Q _7303_/Q _3415_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_7183_ _7183_/D _7207_/RN _7183_/CLK _7183_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4395_ _4580_/C _4489_/A1 _4395_/B _5002_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_98_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6134_ _6134_/A1 _6134_/A2 _6134_/A3 _6133_/Z _6134_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3346_ _7185_/Q _3346_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold1003 _7167_/Q _5832_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold1014 _5822_/Z _7158_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ _7243_/Q _6065_/I1 _6558_/S _7243_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1025 _7191_/Q _5859_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1036 _5824_/Z _7160_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_85_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold1047 _7298_/Q _3433_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1058 _6897_/Q _5524_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_5016_ _5438_/C _5373_/A2 _4586_/Z _5003_/Z _5016_/B2 _5197_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_27_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold1069 _7139_/Q hold600/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_39_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _6967_/D _6967_/RN _6967_/CLK _6967_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_158_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5918_ _5957_/I1 _5917_/Z _5913_/I _6021_/A2 _7228_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6898_ _6898_/D _7122_/RN _6898_/CLK _6898_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_167_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5849_ _5876_/I0 hold454/Z _5856_/S _5849_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold870 _5664_/Z _7019_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_122_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold881 _7087_/Q hold881/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold892 _5663_/Z _7018_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_107_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_55__1359_ clkbuf_4_15_0__1359_/Z net902_170/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_60_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1202_457 net902_189/I _6708_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1202_468 net1202_468/I _6697_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_160_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1202_479 net1202_483/I _6686_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_185_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4180_ _4180_/I0 hold134/Z _4181_/S _4180_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6821_ _6821_/D _6821_/RN _6821_/CLK _6821_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_91_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6752_ _6752_/D _7247_/RN _6752_/CLK _6752_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3964_ _3898_/S _3899_/S _3965_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_50_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5703_ hold416/Z _5877_/I0 _5709_/S _5703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6683_ _6683_/D _7296_/RN _6683_/CLK _6683_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3895_ _3895_/A1 _3889_/Z _3895_/A3 _3894_/Z _3895_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_148_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5634_ _5808_/I0 hold681/Z _5637_/S _5634_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5565_ _5811_/I0 hold645/Z _5565_/S _5565_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold100 _6912_/Q hold100/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7304_ _7304_/D _6656_/Z _7304_/CLK _7304_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold111 _5508_/Z _6887_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4516_ _5003_/A2 _4561_/A2 _5389_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_176_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold122 _7186_/Q hold122/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_160_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5496_ _5538_/I1 hold156/Z _5496_/S _5496_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold133 _5551_/Z _6918_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold144 hold144/I hold144/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold155 _5652_/Z _7008_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7235_ _7235_/D _7237_/RN _7257_/CLK _7235_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold166 _7002_/Q hold166/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4447_ _5055_/A2 _4501_/A1 _5270_/A1 _4501_/B _4504_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold177 _6905_/Q hold177/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold188 _4267_/Z _6781_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold199 _6750_/Q hold199/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xfanout602 _4563_/Z _4643_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_59_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout613 _4455_/A2 _5270_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7166_ _7166_/D _6786_/RN _7166_/CLK _7166_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xfanout624 _3403_/ZN _4930_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout635 _6886_/RN _6882_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_98_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4378_ _4652_/A4 _5201_/A1 _4648_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_98_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout646 _7077_/RN _7297_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout657 _7146_/RN _6892_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6117_ hold46/I _6117_/A2 _6210_/C _6117_/A4 _6128_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xfanout668 _7171_/RN _7024_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3329_ _3329_/I _5942_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XTAP_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout679 _7163_/RN _7247_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_7097_ _7097_/D _7194_/RN _7097_/CLK _7097_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XTAP_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6048_ _5925_/Z _6048_/A2 _6048_/B _6048_/C _6049_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_3006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__11 _4073__7/I _7214_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__22 _4073__46/I _7203_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__33 net802_53/I _7192_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4073__44 _4073__4/I _7181_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3680_ hold221/I _3492_/Z _3680_/A3 _3500_/Z _3680_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_118_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5350_ _5350_/A1 _5350_/A2 _5350_/A3 _5350_/A4 _5350_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xoutput205 _3373_/ZN mgmt_gpio_oeb[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_127_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput216 _6735_/Q mgmt_gpio_out[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput227 hold92/I mgmt_gpio_out[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4301_ _4301_/A1 _5647_/A2 _4303_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
Xoutput238 _4048_/Z mgmt_gpio_out[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput249 _4074_/Z pad_flash_csb VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5281_ _5288_/A1 _5281_/A2 _5281_/B _5281_/C _5369_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_7020_ _7020_/D _7260_/RN _7020_/CLK _7020_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_141_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4232_ _4232_/I0 hold54/Z _4242_/S _4232_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4163_ hold849/Z _5832_/I0 _4163_/S _4163_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4094_ _4094_/I _4094_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6804_ _6804_/D _7262_/CLK _6804_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4996_ _5083_/C _4997_/C _5329_/A2 _4422_/Z _5341_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_149_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6735_ _6735_/D _6771_/RN _6735_/CLK _6735_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3947_ _7094_/Q _3947_/A2 _3947_/B1 _6716_/Q _3949_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_51_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6666_ _6666_/D _6892_/RN _6666_/CLK _6666_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_165_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3878_ _6904_/Q _5532_/A1 _3935_/B1 _6850_/Q _3885_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_137_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5617_ _5782_/I0 hold539/Z _5619_/S _5617_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6597_ _6600_/A1 _6597_/A2 _6597_/B1 _3316_/I _6597_/C1 _6597_/C2 _6598_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5548_ hold258/Z _3542_/Z _4064_/S _5875_/A3 _5556_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_173_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5479_ _5479_/A1 _5479_/A2 _5479_/A3 _5479_/A4 _5479_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7218_ hold87/Z _7218_/RN _7218_/CLK hold86/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout410 _5731_/A2 _5767_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet1102_401 net1152_431/I _6773_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout421 _6245_/Z _6551_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_132_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout432 _5072_/A4 _4973_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout443 _6452_/A2 _6484_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_63_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout454 _5095_/B1 _5226_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7149_ _7149_/D _7149_/RN _7149_/CLK _7149_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_63_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout465 _4666_/Z _5475_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout476 _4672_/A2 _4530_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_86_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout487 _5865_/I0 _5811_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout498 hold16/Z _5555_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_100_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4850_ _5287_/C _5142_/A3 _5106_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3801_ _4332_/A1 _3653_/Z _3928_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4781_ _4781_/A1 _5121_/A1 _5456_/B _5122_/B _4790_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_1990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6520_ _6710_/Q _6544_/A2 _6292_/Z _6722_/Q _6521_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3732_ _3732_/A1 _5857_/A3 _5839_/A3 _3732_/A4 _3732_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_174_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6451_ _7212_/Q _6256_/Z _6464_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3663_ _3663_/A1 _3663_/A2 _3663_/A3 _3663_/A4 _3663_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_9_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5402_ _5480_/A1 _5480_/A2 _5406_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_103_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6382_ _7039_/Q _6275_/Z _6300_/Z _7105_/Q _6383_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3594_ _6963_/Q _3957_/A2 _3927_/C2 input33/Z _5575_/A1 _6947_/Q _3596_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_86_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5333_ _4761_/I _5481_/B1 _5334_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_173_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5264_ _5264_/A1 _5412_/A3 _5264_/A3 _5263_/Z _5265_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_173_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7003_ _7003_/D _7027_/RN _7003_/CLK _7003_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_130_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4215_ hold297/Z _5850_/I0 _4225_/S _4215_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5195_ _5350_/A1 _5350_/A3 _5195_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_68_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4146_ _4146_/A1 _5647_/A2 _4148_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_4077_ _4077_/I _4077_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4979_ _4419_/Z _4973_/Z _4979_/B _4979_/C _4986_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_138_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6718_ _6718_/D _6847_/RN _6718_/CLK _6718_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xnet952_220 _4073__27/I _7005_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet952_231 _4073__37/I _6994_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet952_242 net952_247/I _6983_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6649_ _6650_/A1 _6650_/A2 _6649_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_109_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4000_ _6597_/C1 _4097_/A1 _6831_/Q _4001_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_19_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_9_0__1359_ clkbuf_0__1359_/Z _4073__46/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_77_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5951_ _7225_/Q _7226_/Q _5951_/A3 _5951_/B _5952_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_65_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4902_ _3408_/I _4494_/Z _5248_/A3 _4902_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_33_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5882_ _5891_/I0 hold679/Z _5883_/S _5882_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4833_ _5290_/A1 _4530_/I _4878_/A2 _4483_/B _4833_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4764_ _4765_/A1 _5315_/A4 _4764_/A3 _4692_/C _4764_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_159_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6503_ _7258_/Q _6503_/I1 _6558_/S _7258_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3715_ _3715_/A1 _3715_/A2 _3715_/A3 _3715_/A4 _3715_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4695_ _4736_/A3 _4467_/B _4736_/A1 _4695_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_146_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6434_ _6434_/A1 _6434_/A2 _6434_/A3 _6434_/A4 _6434_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3646_ _3646_/A1 _3630_/Z _3646_/A3 _3645_/Z _3646_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_161_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6365_ _3324_/I _7252_/Q _6365_/B _6366_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3577_ _3512_/Z _5731_/A2 _3947_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_115_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet902_161 net952_209/I _7064_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_172 net902_197/I _7053_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5316_ _5316_/A1 _5316_/A2 _5315_/Z _4772_/Z _5316_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xnet902_183 _4073__37/I _7042_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet902_194 net902_194/I _7031_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6296_ _3328_/I _6296_/A2 _6484_/A2 _6484_/A3 _6296_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_114_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5247_ _5246_/Z _5248_/A3 _5056_/C _4496_/Z _5247_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold15 hold15/I hold15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold26 hold26/I hold26/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold37 hold37/I hold37/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold48 hold48/I hold48/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_69_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5178_ _5180_/A3 _5180_/A2 _5211_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold59 hold59/I hold59/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_29_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4129_ _6612_/I1 hold809/Z _4136_/S _4129_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1052_311 net1052_312/I _6914_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_322 net852_136/I _6903_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_333 net1202_485/I _6892_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_169_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1052_344 net1052_346/I _6881_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3500_ _3500_/I0 _3500_/I1 _3500_/S _3500_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_7_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4480_ _4463_/Z _4468_/Z _4786_/A2 _4786_/A3 _4808_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold507 _7202_/Q hold507/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold518 _4342_/Z _6845_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold529 _6867_/Q hold529/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3431_ _6734_/Q _3434_/B _7299_/Q _3432_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_98_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6150_ _7092_/Q _6002_/Z _6003_/Z _7164_/Q _6152_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_125_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3362_ _7063_/Q _3362_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5101_ _5303_/A1 _5460_/A1 _5101_/A3 _5303_/A2 _5101_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_140_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6081_ _7113_/Q _5984_/Z _5997_/Z _7097_/Q _7071_/Q _5980_/Z _6084_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3293_ _7301_/Q _3428_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5032_ _4397_/Z _4411_/Z _5328_/A1 _5387_/A1 _5032_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6983_ hold61/Z _7124_/RN _6983_/CLK _6983_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_25_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5934_ _5934_/I _7232_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5865_ _5865_/I0 hold685/Z _5865_/S _5865_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4816_ _5369_/A1 _4673_/Z _5132_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_22_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5796_ _5796_/I0 hold935/Z hold12/Z _5796_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1002_252 _4073__42/I _6973_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4747_ _4747_/A1 _4747_/A2 _5231_/C _4751_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xnet1002_263 net902_175/I _6962_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1002_274 net952_228/I _6951_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1002_285 net1202_499/I _6940_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1002_296 net952_227/I _6929_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4678_ _4997_/C _4673_/Z _5380_/B2 _5451_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_6417_ _6554_/A1 _6417_/A2 _6417_/A3 _6417_/A4 _6417_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3629_ _7124_/Q _3956_/A2 _3927_/B1 _7066_/Q _3630_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_123_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6348_ _7136_/Q _6253_/Z _6293_/Z _7152_/Q _6348_/C _6356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_88_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6279_ _6282_/A4 _6285_/A2 _6279_/A3 _7237_/Q _6279_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xinput105 wb_adr_i[19] _4391_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput116 wb_adr_i[29] _4031_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput127 wb_cyc_i _4032_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput138 wb_dat_i[19] _6588_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput149 wb_dat_i[29] _6594_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_15__1359_ net1152_430/I net802_64/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_21_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_78__1359_ net952_221/I net852_119/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_98_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3980_ _3978_/S _3972_/Z _6659_/Q _3981_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XPHY_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5650_ hold371/Z _5806_/I0 _5655_/S _5650_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4601_ _4601_/A1 _4595_/Z _4599_/Z _4600_/Z _4601_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_176_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5581_ hold521/Z _5818_/I0 _5583_/S _5581_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4532_ _5420_/A2 _3403_/I _3404_/I _5129_/A4 _4532_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_7_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold304 _4114_/Z _6671_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold315 _6748_/Q hold315/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7251_ _7251_/D _7257_/RN _7260_/CLK _7251_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold326 _5760_/Z _7103_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4463_ _4460_/B _4481_/A2 _4463_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
XFILLER_117_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold337 _6883_/Q hold337/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold348 _5763_/Z _7106_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_172_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6202_ _6799_/Q _5958_/Z _5969_/Z _7296_/Q _6726_/Q _5994_/I _6204_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold359 _6919_/Q hold359/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3414_ _3304_/I _3413_/Z _3442_/B _3988_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7182_ _7182_/D _6821_/RN _7182_/CLK _7182_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_125_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4394_ _4427_/A3 _4481_/A1 _4922_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6133_ _6133_/A1 _6133_/A2 _6133_/A3 _6133_/A4 _6133_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3345_ _7193_/Q _3345_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ _6064_/I _6065_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold1004 _5832_/Z _7167_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1015 _7198_/Q _5867_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1026 _5859_/Z _7191_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1037 _7044_/Q _5693_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_5015_ _5013_/Z _5350_/A2 _5017_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold1048 _7295_/Q _3438_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1059 _6882_/Q _5502_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_39_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6966_ _6966_/D _7122_/RN _6966_/CLK _6966_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_41_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5917_ _5991_/A2 _5914_/S _5917_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6897_ _6897_/D _7002_/RN _6897_/CLK _6897_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_107_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _5875_/A1 _3521_/Z _5848_/A3 _5856_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_50_995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5779_ _5833_/I0 hold579/Z _5784_/S _5779_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold860 _4171_/Z _6714_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_66_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold871 _6721_/Q hold871/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold882 _5742_/Z _7087_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold893 _7142_/Q hold893/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_103_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_2__1359_ net1152_451/I net1202_468/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_83_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1202_458 net802_66/I _6707_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_185_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet1202_469 net802_63/I _6696_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6820_ _6820_/D _6821_/RN _6820_/CLK _6820_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3963_ _3915_/Z _3919_/Z _3963_/A3 _3962_/Z _6564_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6751_ _6751_/D _7260_/RN _6751_/CLK _6751_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_90_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5702_ hold414/Z _5876_/I0 _5709_/S _5702_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6682_ _6682_/D _7296_/RN _6682_/CLK _6682_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3894_ _3894_/A1 _3894_/A2 _3894_/A3 _3894_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_149_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5633_ _5852_/I0 hold613/Z _5637_/S _5633_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5564_ _5837_/I0 hold594/Z _5565_/S _5564_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold101 _5544_/Z _6912_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7303_ _7303_/D _6655_/Z _4072_/B2 _7303_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4515_ _5002_/A3 _5002_/A4 _5080_/B _4561_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xhold112 _7040_/Q hold112/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5495_ _5537_/I1 _6876_/Q _5496_/S _5495_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold123 _5853_/Z _7186_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_172_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold134 _6720_/Q hold134/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold145 hold145/I hold145/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_171_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold156 _6877_/Q hold156/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4446_ _5365_/A3 _5281_/C _4467_/B _3406_/I _4446_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7234_ _7234_/D _7237_/RN _7257_/CLK _7234_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold167 _5645_/Z _7002_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold178 _5535_/Z _6905_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold189 _6779_/Q hold189/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xclkbuf_leaf_141__1359_ net1152_446/I net1052_346/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_61__1359_ clkbuf_4_15_0__1359_/Z net1152_416/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xfanout603 _4554_/Z _5290_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7165_ _7165_/D _7205_/RN _7165_/CLK _7165_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_160_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4377_ _3401_/I _4836_/A3 _4456_/B _4456_/C _5076_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xfanout614 _4501_/A1 _4853_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_86_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout625 _5055_/A2 _5420_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout636 _6907_/RN _6886_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout647 fanout685/Z _7077_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6116_ _6116_/A1 _5991_/Z _6132_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout658 _7146_/RN fanout658/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3328_ _3328_/I _5943_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7096_ _7096_/D _7202_/RN _7096_/CLK _7096_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_85_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout669 _7083_/RN _7260_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6047_ _7144_/Q _5987_/Z _6015_/Z _7006_/Q _6047_/C _6048_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_74_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6949_ _6949_/D fanout659/Z _6949_/CLK _6949_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_169_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold690 _5833_/Z _7168_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_150_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__12 _4073__12/I _7213_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__23 _4073__23/I _7202_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4073__34 net802_99/I _7191_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__45 _4073__45/I _7180_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput206 _3372_/ZN mgmt_gpio_oeb[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput217 _6736_/Q mgmt_gpio_out[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4300_ _6571_/I0 _6808_/Q _4300_/S _6808_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput228 _6911_/Q mgmt_gpio_out[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5280_ _5372_/A1 _5055_/Z _5284_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xoutput239 _4047_/Z mgmt_gpio_out[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_126_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4231_ _4230_/Z hold329/Z _4245_/S _4231_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4162_ hold861/Z _5822_/I0 _4163_/S _4162_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4093_ _7299_/Q _6894_/RN _4094_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_67_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6803_ _6803_/D _7262_/CLK _6803_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4995_ _4892_/B _5329_/A2 _5428_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_51_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6734_ _6734_/D _6625_/Z _7304_/CLK _6734_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3946_ _6720_/Q _3946_/A2 _4161_/A1 _6708_/Q _6674_/Q _3546_/Z _3949_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_182_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3877_ _7005_/Q _3934_/A2 _3916_/B1 _6879_/Q _3885_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6665_ _6665_/D _6620_/Z _7302_/CLK _6665_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_20_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5616_ _5808_/I0 hold659/Z _5619_/S _5616_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6596_ _6596_/I0 _7275_/Q _6602_/S _7275_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5547_ _5547_/I0 hold275/Z _5547_/S _5547_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5478_ _5478_/A1 _5478_/A2 _5478_/A3 _5478_/B1 _5230_/B _5479_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_132_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7217_ _7217_/D _7219_/RN _7217_/CLK _7217_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4429_ _5083_/C _5173_/A2 _5340_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xfanout400 _6256_/Z _6535_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xfanout411 _3537_/Z _5731_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_48_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout422 _6484_/A4 _6533_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_59_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout433 _4350_/A3 _5520_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_101_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7148_ _7148_/D _7221_/RN _7148_/CLK _7148_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout444 _6402_/A2 _6452_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout455 _5329_/A2 _5095_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_87_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout466 _4614_/Z _5478_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout477 _5164_/A2 _5315_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7079_ _7079_/D fanout655/Z _7079_/CLK _7079_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_100_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout488 _5547_/I0 _5865_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout499 hold15/Z hold16/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_46_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3800_ _4332_/A1 _3680_/Z _3928_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_60_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4780_ _5095_/B1 _4778_/Z _5122_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_14_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3731_ input14/Z _3913_/A2 _3758_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_147_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3662_ _7131_/Q _3930_/A2 _3901_/A2 _6985_/Q _3663_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6450_ _7256_/Q _6450_/I1 _6450_/S _7256_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5401_ _4694_/Z _5401_/A2 _5401_/B _5401_/C _5480_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_6381_ _7097_/Q _6250_/Z _6290_/Z _7081_/Q _6302_/Z _7089_/Q _6383_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3593_ _6939_/Q _3910_/A2 _3901_/A2 _6987_/Q _3596_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_161_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5332_ _5444_/A2 _5327_/Z _5482_/A1 _5332_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_47_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5263_ _4997_/B _5263_/A2 _5329_/A2 _5263_/A4 _5263_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_130_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4214_ _4213_/Z hold181/Z _4228_/S _4214_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7002_ _7002_/D _7002_/RN _7002_/CLK _7002_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5194_ _4555_/C _5205_/A1 _5194_/B1 _5346_/A2 _5350_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_68_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4145_ hold641/Z _5538_/I1 _4145_/S _4145_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4076_ _7299_/Q input88/Z _4077_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_23_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4978_ _5258_/A2 _4977_/Z _4979_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6717_ _6717_/D _6850_/RN _6717_/CLK _6717_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3929_ _3926_/Z _3929_/A2 _3929_/A3 _3929_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_20_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet952_210 net952_250/I _7015_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet952_221 net952_221/I _7004_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet952_232 net802_89/I _6993_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet952_243 net802_81/I _6982_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6648_ _7224_/RN _6648_/A2 _6648_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_20_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6579_ _6600_/A1 _6579_/A2 _6579_/B1 _3316_/I _3317_/I _6579_/C2 _6580_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_146_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5950_ _5950_/A1 _5950_/A2 _5950_/B1 _6302_/A4 _7237_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_46_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4901_ _5260_/A1 _5329_/A2 _5442_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_3190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5881_ _5881_/I0 hold665/Z _5883_/S _5881_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4832_ _5287_/B _5287_/A2 _5281_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_92_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4763_ _4765_/A1 _5315_/A4 _5226_/C _5403_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_187_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6502_ _6502_/I _6503_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3714_ _7024_/Q _5665_/A1 _3923_/C1 _7082_/Q _3714_/C _3715_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4694_ _5307_/A3 _4778_/A4 _4468_/Z _5099_/A2 _4694_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_174_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6433_ hold46/I _6248_/Z _6297_/Z hold42/I _6433_/C _6434_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3645_ _3638_/Z _3642_/Z _3645_/A3 _3645_/A4 _3645_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_106_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3576_ _5776_/A1 _3844_/A1 _5638_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6364_ _6357_/Z _6363_/Z _6364_/B1 _6286_/Z _6364_/C _6365_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_127_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet902_162 net902_162/I _7063_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_173 net902_197/I _7052_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5315_ _5315_/A1 _5315_/A2 _5478_/A2 _5315_/A4 _5315_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6295_ _6295_/I _6298_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_184 net902_184/I _7041_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet902_195 net802_81/I _7030_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5246_ _5258_/B2 _5343_/A2 _5389_/A2 _5255_/A2 _5246_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_60_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold16 hold16/I hold16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold27 hold27/I hold27/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold38 hold38/I hold38/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_29_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold49 hold49/I hold49/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_68_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5177_ _4414_/Z _4878_/Z _5180_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_28_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4128_ _4350_/A3 _5517_/A2 hold146/Z _5629_/A3 _4136_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4059_ _6753_/Q input77/Z _4059_/S _4059_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1052_312 net1052_312/I _6913_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1052_323 net802_64/I _6902_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_334 net1202_491/I _6891_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xnet1052_345 net1202_490/I _6880_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_118__1359_ net952_221/I _4073__39/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold508 _5871_/Z _7202_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_128_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3430_ _7300_/Q _7283_/Q _3430_/S _7300_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold519 _6984_/Q hold519/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_171_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3361_ _7071_/Q _3361_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5100_ _5100_/A1 _5312_/A2 _5220_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6080_ _6943_/Q _5972_/Z _6021_/Z _6999_/Q _6085_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_151_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3292_ _7303_/Q _3422_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5031_ _5028_/Z _5354_/A1 _5202_/A3 _5035_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6982_ _6982_/D _6967_/RN _6982_/CLK _6982_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_65_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5933_ _5913_/I _5957_/I1 _7232_/Q _5934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5864_ _5891_/I0 hold699/Z _5865_/S _5864_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4815_ _5364_/A1 _4764_/Z _5215_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_179_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5795_ _5795_/I0 hold921/Z hold12/Z _5795_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1002_253 net852_138/I _6972_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4746_ _5226_/A1 _5230_/B _5231_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xnet1002_264 net952_229/I _6961_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_175_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1002_275 net952_228/I _6950_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1002_286 net802_76/I _6939_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1002_297 net952_227/I _6928_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4677_ _4673_/Z _4892_/B _5392_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_147_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6416_ _6944_/Q _6551_/A2 _6531_/A2 _6968_/Q _7032_/Q _6552_/A2 _6417_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_135_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3628_ input27/Z _3954_/B1 _3925_/A2 input9/Z _3630_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6347_ _7038_/Q _6536_/B1 _6300_/Z _7104_/Q _6347_/C _6357_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3559_ _3523_/Z _5731_/A2 _3923_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_131_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6278_ _6276_/Z _6277_/Z _6287_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_131_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput106 wb_adr_i[1] _4547_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput117 wb_adr_i[2] input117/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput128 wb_dat_i[0] _3393_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5229_ _5229_/A1 _5479_/A2 _5234_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_88_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput139 wb_dat_i[1] _3394_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4600_ _5399_/A1 _5399_/A2 _5146_/A1 _5364_/B _4600_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_157_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5580_ hold527/Z _5781_/I0 _5583_/S _5580_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4531_ _5270_/A1 _4530_/I _5214_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold305 _6739_/Q hold305/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7250_ _7250_/D _7260_/RN _7260_/CLK _7250_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold316 _4216_/Z _6748_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4462_ _4736_/A1 _4736_/A3 _4778_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold327 _6685_/Q hold327/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold338 _5504_/Z _6883_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6201_ _6201_/A1 _6201_/A2 _6201_/A3 _6201_/A4 _6201_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold349 _6677_/Q hold349/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3413_ _3412_/Z _3409_/Z _6732_/Q _3413_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_7181_ _7181_/D _7201_/RN _7181_/CLK _7181_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4393_ _4385_/Z _4387_/Z _4390_/Z _4489_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_98_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6132_ _7139_/Q _5994_/I _6132_/B _6133_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3344_ _6926_/Q _6364_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6063_ _6364_/C _7242_/Q _6063_/B _6064_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1005 _6949_/Q _5586_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_39_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1016 _5867_/Z _7198_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1027 _7190_/Q _5858_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1038 _5693_/Z _7044_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_5014_ _4555_/C _5439_/A1 _5349_/A1 _5439_/B2 _5350_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold1049 _6955_/Q _5592_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_27_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _6965_/D fanout655/Z _6965_/CLK _6965_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5916_ _5991_/A2 _5914_/S _6210_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xclkbuf_leaf_21__1359_ _4073__49/I net802_99/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_146_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_101__1359_ clkbuf_4_5_0__1359_/Z net952_235/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6896_ _6896_/D _6967_/RN _6896_/CLK _6896_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_84__1359_ clkbuf_4_13_0__1359_/Z net952_247/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5847_ _5892_/I0 hold715/Z _5847_/S _5847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5778_ _5778_/I0 hold394/Z _5784_/S _5778_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4729_ _4765_/A1 _5307_/A3 _5099_/A2 _5478_/B1 _4729_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_181_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold850 _4163_/Z _6709_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold861 _6708_/Q hold861/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold872 _4181_/Z _6721_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold883 _6853_/Q hold883/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold894 _5804_/Z _7142_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_27_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet1202_459 net852_131/I _6706_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_186_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6750_ _6750_/D _7122_/RN _6750_/CLK _6750_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_17_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3962_ _3938_/Z _3944_/Z _3949_/Z _3961_/Z _3962_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_51_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5701_ _5701_/A1 hold33/Z _5709_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_188_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6681_ hold57/Z _6839_/RN _6681_/CLK hold56/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3893_ _7151_/Q _3916_/A2 _5536_/A1 _6907_/Q _3894_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_177_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5632_ _5797_/I0 hold436/Z _5637_/S _5632_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5563_ _5827_/I0 hold755/Z _5565_/S _5563_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7302_ _7302_/D _6654_/Z _7302_/CLK _7302_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_145_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4514_ _4414_/Z _5010_/A1 _4452_/Z _4810_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
Xhold102 _6885_/Q hold102/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_7_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold113 _5688_/Z _7040_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_5494_ _3508_/Z _5884_/A2 _5848_/A3 hold137/Z _5494_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold124 _7210_/Q hold124/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_117_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold135 _4180_/Z _6720_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_172_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7233_ _7233_/D _7253_/RN _7257_/CLK _7233_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xhold146 hold146/I hold146/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4445_ _4853_/A1 _4449_/B _5309_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold157 _5496_/Z _6877_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold168 _6946_/Q hold168/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold179 _7062_/Q hold179/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7164_ _7164_/D _7201_/RN _7164_/CLK _7164_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout604 _4526_/Z _4997_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout615 _4944_/A1 _4467_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4376_ _3401_/I _4836_/A3 _4456_/B _4456_/C _4376_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xfanout626 _3402_/ZN _5055_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6115_ _7025_/Q _6211_/A2 _6211_/B1 _6993_/Q _6116_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xfanout637 _7077_/RN _6907_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout648 fanout656/Z _6786_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_3327_ _7232_/Q _6279_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
Xfanout659 _7140_/RN fanout659/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7095_ _7095_/D _6856_/RN _7095_/CLK _7095_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XTAP_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6046_ _7160_/Q _6117_/A2 _6164_/A2 _6117_/A4 _6047_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_3008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6948_ _6948_/D fanout659/Z _6948_/CLK _6948_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_169_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6879_ _6879_/D _6882_/RN _6879_/CLK _6879_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold680 _5882_/Z _7212_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold691 _6789_/Q hold691/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_150_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__13 _4073__17/I _7212_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__24 _4073__24/I _7201_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__35 _4073__35/I _7190_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__46 _4073__46/I _7179_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput207 _3371_/ZN mgmt_gpio_oeb[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_154_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput218 _6737_/Q mgmt_gpio_out[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput229 _6912_/Q mgmt_gpio_out[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_154_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4230_ hold116/Z hold64/I _4244_/S _4230_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4161_ _4161_/A1 _5647_/A2 _4163_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_4092_ _4092_/I _4092_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6802_ _6802_/D _7262_/CLK _6802_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4994_ _5083_/C _4997_/C _5146_/A1 _4422_/Z _4994_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_23_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6733_ _6733_/D _6624_/Z _7304_/CLK _6733_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3945_ _7174_/Q _3945_/A2 _3945_/B1 _7086_/Q _6682_/Q _3945_/C2 _3949_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_23_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6664_ _6664_/D _6619_/Z _7302_/CLK _6664_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3876_ _3873_/Z _3876_/A2 _3876_/A3 _3876_/A4 _3876_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_17_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5615_ _5798_/I0 hold463/Z _5619_/S _5615_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6595_ _6595_/A1 _6601_/A2 _6595_/B _6596_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_118_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5546_ hold16/Z hold72/Z _5547_/S hold73/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5477_ _5352_/Z _5390_/Z _5437_/Z _5476_/Z _5477_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_133_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7216_ hold37/Z _7220_/RN _7216_/CLK hold36/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4428_ _4427_/Z _4428_/A2 _4373_/Z _4428_/B2 _5337_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xfanout401 _6251_/Z _6550_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_160_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout412 hold212/I _5517_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_2_3__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _7302_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout423 _6235_/Z _6549_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_132_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout434 _5821_/A1 _4350_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_7147_ _7147_/D _7155_/RN _7147_/CLK _7147_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_113_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4359_ _4359_/A1 _6611_/A2 _4361_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_48_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout445 hold210/Z hold211/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_87_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout456 _4716_/Z _5329_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_171_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout467 _4614_/Z _5290_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_101_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout478 _5093_/A1 _5020_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7078_ _7078_/D _7077_/RN _7078_/CLK _7078_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_74_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout489 _5775_/I0 _5892_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6029_ _7103_/Q _5967_/Z _5969_/Z _7119_/Q _6030_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_100_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3730_ _7071_/Q _3943_/A2 _3945_/B1 _7089_/Q _3757_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_147_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3661_ _7057_/Q _5701_/A1 _3925_/A2 input8/Z _3663_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_173_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5400_ _5400_/A1 _5400_/A2 _5399_/Z _4729_/Z _5401_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6380_ _6380_/A1 _6380_/A2 _6380_/A3 _6380_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_3592_ _3592_/A1 _3592_/A2 _3592_/A3 _3592_/A4 _3592_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_55_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5331_ _5331_/I _5482_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5262_ _5340_/A1 _5262_/A2 _5328_/A2 _5442_/A4 _5262_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_173_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7001_ _7001_/D _7141_/RN _7001_/CLK _7001_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_69_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4213_ hold173/Z _4103_/I _4225_/S _4213_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5193_ _5193_/A1 _5193_/A2 _5437_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_96_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4144_ hold643/Z _5537_/I1 _4145_/S _4144_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4075_ input83/Z _4075_/I1 _7299_/Q _4075_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4977_ _5262_/A2 _5343_/A2 _4982_/A2 _4497_/Z _4977_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_51_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6716_ _6716_/D _6850_/RN _6716_/CLK _6716_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3928_ _6940_/Q _5575_/A1 _3928_/B1 _6789_/Q _3928_/C1 _6822_/Q _3929_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xnet952_211 net802_81/I _7014_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet952_222 net952_226/I _7003_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet952_233 net802_78/I _6992_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6647_ _7224_/RN _6648_/A2 _6647_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
Xnet952_244 net952_244/I _6981_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3859_ _6933_/Q _3910_/A2 _3959_/B1 _6667_/Q _3925_/A2 input35/Z _3860_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_146_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6578_ _6578_/A1 _6578_/A2 _6602_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_30_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5529_ hold33/Z hold65/Z _6901_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_3_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4900_ _5343_/B _5255_/A2 _4900_/B _5341_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_3180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5880_ _5880_/I0 hold124/Z _5883_/S _5880_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4831_ _5214_/A2 _5420_/A1 _5223_/A2 _5276_/B _5276_/A1 _4840_/B1 _4834_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_2490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4762_ _5055_/A2 _5270_/A1 _4761_/I _3401_/I _4762_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6501_ _6500_/C _7257_/Q _6501_/B _6502_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3713_ _3713_/I _3714_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4693_ _5099_/A1 _5099_/A2 _5097_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_146_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6432_ _6432_/A1 _6239_/Z _6433_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_174_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3644_ _7010_/Q _3934_/A2 _3916_/A2 _7156_/Q _3645_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_128_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6363_ _6554_/A1 _6363_/A2 _6363_/A3 _6363_/A4 _6363_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3575_ _7067_/Q _3927_/B1 _3592_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_136_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet902_152 net902_162/I _7073_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5314_ _5314_/A1 _5314_/A2 _5314_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
Xnet902_163 net902_170/I _7062_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6294_ _7142_/Q _6292_/Z _6293_/Z _7150_/Q _6295_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xnet902_174 net952_238/I _7051_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_185 net902_185/I _7040_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_196 _4073__23/I _7029_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5245_ _4421_/Z _4510_/Z _5475_/A4 _5415_/A1 _5245_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_130_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold17 hold17/I hold17/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_102_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold28 hold28/I hold28/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_69_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5176_ _5175_/Z _4313_/Z _5184_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold39 hold39/I hold39/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_57_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4127_ hold6/Z hold56/Z _4127_/S hold57/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4058_ _6755_/Q input67/Z _7302_/Q _4058_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1052_302 _4073__48/I _6923_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_313 net1052_315/I _6912_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1052_324 net902_170/I _6901_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_335 net1202_499/I _6890_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xnet1052_346 net1052_346/I _6879_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold509 _6725_/Q hold509/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_156_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3360_ _6701_/Q _3360_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5030_ _5471_/B2 _5376_/B2 _5002_/Z _5353_/A1 _5202_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6981_ _6981_/D fanout658/Z _6981_/CLK _6981_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_18_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5932_ _5932_/I _7231_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5863_ hold40/Z hold230/Z _5865_/S _5863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4814_ _5414_/A2 _5369_/A1 _4876_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5794_ _3507_/Z _5794_/A2 _5794_/A3 hold12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_178_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _5478_/B1 _5230_/B _4747_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xnet1002_254 net952_226/I _6971_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1002_265 net952_209/I _6960_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1002_276 net1202_463/I _6949_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1002_287 net802_52/I _6938_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet1002_298 net802_98/I _6927_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4676_ _5380_/B2 _5295_/A2 _4472_/B _4524_/Z _4892_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_174_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6415_ _7048_/Q _6550_/A2 _6550_/B1 _6984_/Q _6550_/C1 _6952_/Q _6417_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_179_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3627_ _7002_/Q _5638_/A1 _3959_/B1 hold48/I input32/Z _3927_/C2 _3630_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_179_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6346_ _7096_/Q _6250_/Z _6302_/Z _7088_/Q _6292_/Z _7144_/Q _6357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3558_ _5884_/A2 _5839_/A2 _3916_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_143_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6277_ _6544_/B1 _6549_/C1 _6550_/C1 _6552_/A2 _6277_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3489_ _3489_/I _3653_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
Xclkbuf_leaf_44__1359_ _4073__46/I _4073__9/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_124__1359_ _4073__49/I _4073__27/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_103_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput107 wb_adr_i[20] input107/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput118 wb_adr_i[30] _4035_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5228_ _5287_/C _5478_/A3 _5228_/A3 _5228_/B _5479_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
Xinput129 wb_dat_i[10] _6585_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5159_ _5290_/A1 _5438_/A1 _4641_/Z _4483_/B _5160_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_5_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_189_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4530_ _4530_/I _4860_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_157_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold306 _4205_/Z _6739_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4461_ _4652_/A4 _4481_/A2 _4469_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold317 _7171_/Q hold317/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold328 _4132_/Z _6685_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6200_ _6843_/Q _5971_/Z _5981_/Z _6787_/Q _6005_/Z _6849_/Q _6201_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold339 _7036_/Q hold339/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_171_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3412_ _3451_/I0 _7292_/Q _7293_/Q _3412_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_7180_ _7180_/D _7201_/RN _7180_/CLK _7180_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_171_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4392_ _4385_/Z _4387_/Z _4390_/Z _4392_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_113_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6131_ hold42/I _5965_/Z _5967_/Z _7107_/Q _7171_/Q _6006_/Z _6133_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3343_ _7136_/Q _6051_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ _6053_/Z _6061_/Z _6364_/B1 _6118_/B _6529_/S _6063_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_100_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1006 _5586_/Z _6949_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_97_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold1017 _7079_/Q _5733_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _5347_/A1 _5012_/Z _5347_/A4 _5192_/B _5013_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1028 _5858_/Z _7190_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1039 _6874_/Q _3649_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_38_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6964_ _6964_/D _7090_/RN _6964_/CLK _6964_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_41_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5915_ _5945_/A1 _5957_/I1 _5941_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_179_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6895_ _6895_/D _7247_/RN _6895_/CLK _6895_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_62_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5846_ _5891_/I0 hold733/Z _5847_/S _5846_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5777_ _6612_/I1 hold379/Z _5784_/S _5777_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4728_ _4765_/A1 _5478_/A3 _5099_/A2 _4728_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_175_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4659_ _5281_/C _3408_/I _5295_/A3 _4501_/B _4659_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_163_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold840 _4346_/Z _6848_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold851 _6847_/Q hold851/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_66_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold862 _4162_/Z _6708_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold873 _7166_/Q hold873/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold884 _4354_/Z _6853_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6329_ _6329_/A1 _6329_/A2 _6322_/Z _6328_/Z _6329_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_66_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold895 _7165_/Q hold895/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_153_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_90__1359_ clkbuf_4_7_0__1359_/Z net902_168/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_76_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3961_ _3953_/Z _3958_/Z _3961_/A3 _3961_/A4 _3961_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_16_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5700_ _5784_/I0 hold947/Z _5700_/S _5700_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_177_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6680_ _6680_/D _6839_/RN _6680_/CLK _6680_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3892_ _7111_/Q _3917_/A2 _3950_/B1 _6725_/Q _3894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_177_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5631_ _5796_/I0 _5631_/I1 _5637_/S _5631_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5562_ _5724_/I0 hold475/Z _5565_/S _5562_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7301_ _7301_/D _6653_/Z _7302_/CLK _7301_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4513_ _5010_/A1 _4506_/Z _5180_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_8_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold103 _5506_/Z _6885_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_5493_ _5751_/I0 hold529/Z _5493_/S _5493_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold114 _6686_/Q hold114/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold125 _5880_/Z _7210_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7232_ _7232_/D _7237_/RN _4067_/I1 _7232_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4444_ _5288_/B _4472_/B _4868_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold136 _6864_/Q _3309_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold147 _4173_/Z _4175_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold158 _6783_/Q hold158/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_171_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold169 _5582_/Z _6946_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7163_ _7163_/D _7163_/RN _7163_/CLK _7163_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4375_ _3401_/I _4836_/A3 _5170_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xfanout605 _4526_/Z _4889_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout616 _4903_/A1 _4944_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6114_ _6953_/Q _5958_/Z _5969_/Z _7123_/Q _6133_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout627 _4960_/A1 _5420_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout638 _7077_/RN _6844_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3326_ _7233_/Q _6282_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
X_7094_ _7094_/D _7162_/RN _7094_/CLK _7094_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xfanout649 _7162_/RN _6856_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6045_ _7088_/Q _6002_/Z _6048_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_37_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ hold7/Z _7238_/RN _6947_/CLK _6947_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_179_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6878_ _6878_/D _6882_/RN _6878_/CLK _6878_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_139_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5829_ _5892_/I0 hold895/Z _5829_/S _5829_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold670 _4330_/Z _6837_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold681 _6992_/Q hold681/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_2_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold692 _4278_/Z _6789_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_134_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__14 net802_62/I _7211_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073__25 net802_95/I _7200_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__36 _4073__45/I _7189_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__47 net802_98/I _7178_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput208 _3370_/ZN mgmt_gpio_oeb[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_127_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput219 _6738_/Q mgmt_gpio_out[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_175_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4160_ _5832_/I0 hold617/Z _4160_/S _4160_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4091_ _7300_/Q _6894_/RN _4092_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_56_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6801_ _6801_/D _7262_/CLK _6801_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4993_ _4993_/A1 _4988_/Z _4993_/A3 _4999_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_3944_ _3944_/A1 _3944_/A2 _3944_/A3 _3944_/A4 _3944_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6732_ _6732_/D _6623_/Z _7304_/CLK _6732_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_189_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6663_ _6663_/D _6618_/Z _7302_/CLK _6663_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3875_ _7053_/Q _5701_/A1 _4188_/A1 _6727_/Q _3914_/B1 _6877_/Q _3876_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_165_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5614_ _5806_/I0 hold949/Z _5619_/S _5614_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6594_ _6600_/A1 _6594_/A2 _6594_/B1 _3316_/I _3317_/I _6594_/C2 _6595_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5545_ _5890_/I0 hold224/Z _5547_/S _5545_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5476_ _5476_/A1 _5476_/A2 _5475_/Z _5151_/B _5476_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_7215_ _7215_/D _7215_/RN _7215_/CLK _7215_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4427_ _4374_/Z _4427_/A2 _4427_/A3 _4481_/A1 _4427_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_63_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout402 _6243_/Z _6549_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xfanout413 _3521_/Z _5776_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7146_ _7146_/D _7146_/RN _7146_/CLK _7146_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_48_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4358_ _5832_/I0 hold693/Z _4358_/S _4358_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout424 _5968_/ZN _6211_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_98_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout435 hold11/Z _5821_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_24_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout446 _3497_/I _3680_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_58_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout457 _4703_/Z _5401_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_171_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3309_ _3309_/I _5474_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
Xfanout468 _4586_/Z _5367_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_150_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7077_ _7077_/D _7077_/RN _7077_/CLK _7077_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4289_ _4289_/A1 _6611_/A2 _4291_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
Xfanout479 _5093_/A1 _5359_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_87_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6028_ _7151_/Q _5960_/Z _5965_/Z _6699_/Q _6030_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_2105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3660_ _6937_/Q _3910_/A2 _5575_/A1 _6945_/Q _3663_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_16_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3591_ _7141_/Q _3951_/A2 _3954_/B1 input28/Z _3959_/B1 hold68/I _3592_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_127_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5330_ _4936_/I _5246_/Z _5445_/B2 _5330_/B2 _5330_/C _5331_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_154_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5261_ _5261_/I _5264_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7000_ _7000_/D _7260_/RN _7000_/CLK _7000_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4212_ _4225_/S _4194_/Z _4060_/S _3519_/Z hold33/Z _4228_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_5192_ _4517_/Z _4547_/Z _5192_/B _5192_/C _5193_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_4143_ _4143_/A1 _6611_/A2 _4145_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_110_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4074_ input84/Z input67/Z _7300_/Q _4074_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4976_ _4421_/Z _5263_/A2 _4976_/A3 _5263_/A4 _5337_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_11_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6715_ _6715_/D _7154_/RN _6715_/CLK _6715_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3927_ _6698_/Q _3927_/A2 _3927_/B1 _7060_/Q input4/Z _3927_/C2 _3929_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xnet952_212 net802_91/I _7013_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet952_223 net952_228/I _7002_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3858_ _6699_/Q _3927_/A2 _3902_/A2 _6890_/Q input15/Z _3927_/C2 _3860_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xnet952_234 net952_234/I _6991_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6646_ _7224_/RN _6648_/A2 _6646_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
Xnet952_245 net952_245/I _6980_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3789_ _7006_/Q _3934_/A2 _5528_/S _6897_/Q _3790_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6577_ _6600_/A1 _6607_/A2 _6605_/A2 _3316_/I _6577_/C _6578_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xclkbuf_4_14_0__1359_ clkbuf_0__1359_/Z clkbuf_4_14_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5528_ _6901_/Q hold64/Z _5528_/S hold65/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5459_ _5459_/A1 _5098_/B _5098_/C _5458_/Z _5460_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_105_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7129_ _7129_/D _7221_/RN _7129_/CLK _7129_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_8_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_8__1359_ net1152_430/I net802_67/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_151_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4830_ _5369_/A1 _5367_/A2 _4840_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_2480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4761_ _4761_/I _5071_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3712_ _6992_/Q _3954_/A2 _3954_/B1 input24/Z _3713_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6500_ _6493_/Z _6499_/Z _6500_/B1 _6286_/Z _6500_/C _6501_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_14_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4692_ _4735_/A2 _4764_/A3 _4692_/B _4692_/C _5099_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_14_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3643_ _6688_/Q _3945_/C2 _3941_/A2 _7164_/Q _3645_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6431_ _7131_/Q _6484_/A2 _6533_/A3 hold44/I _6432_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_134_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6362_ _6942_/Q _6551_/A2 _6273_/Z _6974_/Q _7120_/Q _6288_/Z _6363_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3574_ _5776_/A1 _5767_/A3 _3927_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_155_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5313_ _5313_/A1 _5313_/A2 _5313_/A3 _5312_/Z _5314_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xnet902_153 net902_184/I _7072_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_164 net802_82/I _7061_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6293_ _3328_/I _3329_/I _6302_/A3 _6484_/A3 _6293_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xnet902_175 net902_175/I _7050_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_186 net802_93/I _7039_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet902_197 net902_197/I _7028_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5244_ _5324_/A1 _5324_/A2 _5324_/C _5250_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_170_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold18 hold18/I hold18/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold29 hold29/I hold29/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_5175_ _5175_/A1 _5380_/C _5175_/A3 _5175_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_28_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4126_ _5645_/I1 hold299/Z _4127_/S _4126_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ _6756_/Q _4072_/B2 _7301_/Q _4057_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1052_303 net1152_415/I _6922_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_314 net1052_315/I _6911_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_325 net1052_328/I _6900_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_336 net1202_499/I _6889_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xnet1052_347 net1202_453/I _6878_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4959_ _4959_/A1 _4959_/A2 _4957_/Z _4958_/Z _4963_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xclkbuf_leaf_67__1359_ clkbuf_4_13_0__1359_/Z net902_175/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_184_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_147__1359_ net1152_451/I net1152_427/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_138_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6629_ _6844_/RN _6652_/A2 _6629_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_119_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6980_ _6980_/D _7090_/RN _6980_/CLK _6980_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_20_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5931_ _5931_/I0 _6068_/A2 _5931_/S _5932_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5862_ hold20/Z hold80/Z _5865_/S hold81/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4813_ _5173_/A2 _4997_/C _4554_/Z _4877_/A2 _5167_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_22_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5793_ _5892_/I0 hold773/Z _5793_/S _5793_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4744_ _5315_/A4 _3406_/I _4786_/A2 _5099_/A1 _5230_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_159_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1002_255 net902_199/I _6970_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1002_266 net952_208/I _6959_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1002_277 net1202_463/I _6948_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4675_ _4424_/B _4026_/B _4026_/C _4402_/B _4675_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xnet1002_288 net952_235/I _6937_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1002_299 net852_119/I _6926_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6414_ _7008_/Q _6549_/B1 _6273_/Z _6976_/Q _6414_/C _6417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3626_ _7188_/Q _3959_/C1 _3923_/C1 _7084_/Q _3951_/C1 _7148_/Q _3646_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_150_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6345_ _6345_/I _6347_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3557_ _3523_/Z _5692_/A1 _5665_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_1_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6276_ _6549_/A2 _6237_/Z _6549_/B1 _6545_/B1 _6276_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_163_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3488_ _3487_/Z hold219/Z _3500_/S _3488_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_142_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5227_ _5227_/I _5228_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput108 wb_adr_i[21] input108/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput119 wb_adr_i[31] _4035_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5158_ _5293_/A1 _5293_/B _5161_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4109_ hold58/Z _7273_/Q _4117_/S hold59/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_186_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5089_ _4506_/Z _5475_/A4 _5341_/C _5265_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_16_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_130__1359_ net1152_446/I net1202_486/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_50__1359_ clkbuf_4_11_0__1359_/Z net802_96/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_184_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4460_ _5270_/A2 _4367_/Z _4460_/B _4736_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_172_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold307 _7009_/Q hold307/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_7_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold318 _5836_/Z _7171_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold329 _6755_/Q hold329/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3411_ _7293_/Q _7292_/Q _4042_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_172_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4391_ _4391_/A1 _4391_/A2 _4391_/A3 _4391_/A4 _4481_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6130_ _6937_/Q _5981_/Z _5984_/Z hold44/I _6134_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_125_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3342_ _7251_/Q _6310_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6061_ _6057_/Z _6061_/A2 _6061_/A3 _6061_/A4 _6061_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_86_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1007 _7127_/Q _5787_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_5012_ _5350_/A1 _5192_/C _5009_/Z _4576_/C _5012_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1018 _5733_/Z _7079_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold1029 _7174_/Q _5840_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_66_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6963_ _6963_/D _7019_/RN _6963_/CLK _6963_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_81_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5914_ _5957_/I1 _5913_/I _5914_/S _7227_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6894_ _6894_/D _6894_/RN _6894_/CLK _6894_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_146_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5845_ _5890_/I0 hold586/Z _5847_/S _5845_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5776_ _5776_/A1 _5821_/A2 hold11/Z _5784_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_4727_ _4727_/A1 _5223_/C _4727_/A3 _5090_/A1 _4733_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_148_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_2_0__1359_ clkbuf_0__1359_/Z net1152_430/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4658_ _4887_/A1 _5315_/A2 _5172_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_174_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput90 spimemio_flash_io2_oeb input90/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold830 _5827_/Z _7163_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3609_ _7294_/Q _6732_/Q _3899_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold841 _7297_/Q hold841/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold852 _4345_/Z _6847_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4589_ _4715_/A1 _5270_/A2 _4643_/A4 _4589_/A4 _4589_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold863 _6715_/Q hold863/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold874 _5831_/Z _7166_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6328_ _6328_/A1 _6328_/A2 _6328_/A3 _6328_/A4 _6328_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold885 _7152_/Q hold885/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold896 _5829_/Z _7165_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6259_ _6259_/A1 _6259_/A2 _6259_/A3 _6259_/A4 _6259_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_104_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3960_ _7206_/Q _3960_/A2 _3960_/B1 _6718_/Q _3960_/C _3961_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_50_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3891_ _6949_/Q _5584_/A1 _3954_/B1 input21/Z _5575_/A1 _6941_/Q _3894_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_32_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5630_ _5795_/I0 hold959/Z _5637_/S _5630_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5561_ _5834_/I0 hold426/Z _5565_/S _5561_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7300_ _7300_/D _6652_/Z _4075_/I1 _7300_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_145_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4512_ _5010_/A1 _4452_/Z _5043_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5492_ _5885_/I0 hold484/Z _5493_/S _5492_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold104 _6767_/Q hold104/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold115 _4133_/Z _6686_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_145_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold126 _7178_/Q hold126/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_105_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7231_ _7231_/D _7240_/RN _7257_/CLK _7231_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_160_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4443_ _4522_/A2 _4380_/Z _4580_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold137 _3477_/Z hold137/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold148 _4174_/Z _6716_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold159 _4269_/Z _6783_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7162_ hold79/Z _7162_/RN _7162_/CLK hold78/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4374_ _4522_/A2 _4853_/A1 _4884_/A1 _4374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_171_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout606 _4524_/Z _5399_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout617 _4652_/A4 _5281_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6113_ _7245_/Q _6113_/I1 _6558_/S _7245_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3325_ _4009_/B _5950_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
XTAP_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7093_ _7093_/D _7173_/RN _7093_/CLK _7093_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_140_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout628 _3401_/ZN _4960_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout639 _7077_/RN _6850_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_98_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6044_ _6210_/A2 _7054_/Q _6048_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6946_ _6946_/D _7002_/RN _6946_/CLK _6946_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_53_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6877_ _6877_/D _6882_/RN _6877_/CLK _6877_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_167_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5828_ _5891_/I0 hold879/Z _5829_/S _5828_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5759_ hold333/Z _5822_/I0 _5766_/S _5759_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold660 _5616_/Z _6976_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_1_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold671 _6696_/Q hold671/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold682 _5634_/Z _6992_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold693 _6856_/Q hold693/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_1_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4073__15 _4073__23/I _7210_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__26 _4073__42/I _7199_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__37 _4073__37/I _7188_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__48 _4073__48/I _7177_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput209 _4063_/Z mgmt_gpio_out[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_182_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4090_ _4097_/A1 _4686_/B _6827_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_64_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6800_ _6800_/D _6847_/RN _6800_/CLK _6800_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_91_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4992_ _5337_/A2 _5130_/B2 _5368_/A1 _5080_/B _5415_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_56_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6731_ _6731_/D _6622_/Z _7302_/CLK _6731_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3943_ _7068_/Q _3943_/A2 _5728_/A1 _7076_/Q _4182_/A1 _6722_/Q _3944_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_143_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6662_ _6662_/D _6617_/Z _4072_/B2 _6662_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3874_ _6884_/Q _3912_/B1 _3934_/B1 _6846_/Q _6858_/Q _4359_/A1 _3876_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_143_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ _5850_/I0 hold452/Z _5619_/S _5613_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6593_ _6593_/I0 _7274_/Q _6602_/S _7274_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5544_ _5889_/I0 hold100/Z _5547_/S _5544_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5475_ _5438_/C _4604_/Z _5475_/A3 _5475_/A4 _5475_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7214_ _7214_/D _7218_/RN _7214_/CLK _7214_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4426_ _4721_/A1 _4721_/A2 _5083_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xfanout403 _6241_/Z _6550_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xfanout414 _3517_/ZN _5629_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_98_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7145_ _7145_/D _7221_/RN _7145_/CLK _7145_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4357_ _5885_/I0 hold727/Z _4358_/S _4357_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout425 _5968_/ZN _6164_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout436 hold11/Z _5794_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_101_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout447 _3489_/I hold221/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_98_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3308_ _6863_/Q _5431_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout458 _4703_/Z _5415_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7076_ _7076_/D _7077_/RN _7076_/CLK _7076_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4288_ _6571_/I0 _6798_/Q _4288_/S _6798_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout469 _4568_/Z _5438_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_39_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6027_ _6949_/Q _5958_/Z _5994_/I _7135_/Q _6027_/C _6030_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_104_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6929_ _6929_/D _7258_/RN _6929_/CLK _6929_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold490 _6985_/Q hold490/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_78_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3590_ _7019_/Q _5656_/A1 _3925_/A2 input10/Z _5665_/A1 _7027_/Q _3592_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_139_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5260_ _5260_/A1 _4982_/Z _5260_/B _5261_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_5_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4211_ _4210_/Z hold323/Z _4211_/S _4211_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5191_ _4600_/Z _5190_/Z _5191_/A3 _5191_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_4142_ _5832_/I0 hold677/Z _4142_/S _4142_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4975_ _4975_/A1 _4975_/A2 _4975_/A3 _4979_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6714_ _6714_/D _7154_/RN _6714_/CLK _6714_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_149_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3926_ _3926_/A1 _3926_/A2 _3926_/A3 _3926_/A4 _3926_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_177_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet952_202 net952_218/I _7023_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet952_213 net802_91/I _7012_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet952_224 net802_78/I _7001_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6645_ _7224_/RN _6648_/A2 _6645_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3857_ _6838_/Q _3923_/B1 _3960_/B1 _6719_/Q _3860_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xnet952_235 net952_235/I _6990_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xnet952_246 net952_247/I _6979_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6576_ _6832_/Q _6608_/I1 _6606_/A2 _3317_/I _6578_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3788_ _7104_/Q _5758_/A1 _3947_/A2 _7096_/Q _3941_/B1 _7168_/Q _3790_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_164_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5527_ hold215/Z _5877_/I0 _5527_/S _5527_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5458_ _4539_/I _5478_/A2 _5302_/B _5458_/A4 _5458_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_160_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4409_ _4407_/Z _4390_/Z _4485_/A2 _5385_/A1 _4412_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_99_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5389_ _5389_/A1 _5389_/A2 _5389_/B _5389_/C _5390_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_160_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7128_ _7128_/D _7207_/RN _7128_/CLK _7128_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xclkbuf_leaf_107__1359_ clkbuf_4_5_0__1359_/Z net802_84/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_27__1359_ clkbuf_opt_1_0__1359_/Z net1152_431/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7059_ _7059_/D _7188_/RN _7059_/CLK _7059_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_189_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _5324_/A1 _3408_/I _4982_/A2 _4759_/Z _4761_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_1791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3711_ _7016_/Q _5656_/A1 _3924_/A2 _6968_/Q _3927_/A2 _6702_/Q _3715_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_14_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4691_ _4786_/A2 _4692_/B _4692_/C _4691_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_119_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6430_ _7203_/Q _6540_/A2 _6536_/B1 _7041_/Q _6293_/Z _7155_/Q _6434_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_174_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3642_ _3642_/A1 _3642_/A2 _3642_/A3 _3642_/A4 _3642_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_146_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6361_ _7046_/Q _6550_/A2 _6550_/B1 _6982_/Q _6550_/C1 _6950_/Q _6363_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3573_ _3523_/Z _3732_/A4 _3951_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_143_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5312_ _5312_/A1 _5312_/A2 _5376_/B2 _5312_/A4 _5312_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet902_154 net902_170/I _7071_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6292_ _3328_/I _6300_/A1 _6484_/A3 _6299_/A2 _6292_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xnet902_165 net952_245/I _7060_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_176 net952_229/I _7049_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_187 net902_187/I _7038_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_198 net902_199/I _7027_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5243_ _5243_/A1 _4890_/I _5324_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_130_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold19 hold19/I hold19/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_5174_ _5392_/B _4893_/Z _4991_/C _5175_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_69_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4125_ hold40/Z hold66/Z _4127_/S hold67/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4056_ _6757_/Q _4056_/I1 _7302_/Q _4056_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1052_304 _4073__8/I _6921_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1052_315 net1052_315/I _6910_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_326 net1102_394/I _6899_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_337 net1202_483/I _6888_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xnet1052_348 net1202_490/I _6877_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4958_ _5258_/B2 _5248_/A3 _5248_/A2 _4958_/A4 _4958_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_177_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3909_ _7190_/Q _3909_/A2 _3915_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4889_ _4889_/A1 _5478_/B1 _4890_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6628_ _6844_/RN _6652_/A2 _6628_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_138_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6559_ _6833_/D _6830_/Q _6826_/Q _6833_/Q _6559_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_118_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_10__1359_ net1152_430/I net852_131/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_38_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_73__1359_ _4073__46/I net802_97/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5930_ _5924_/Z _6210_/A2 _6201_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_47_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5861_ _5888_/I0 hold281/Z _5865_/S _5861_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4812_ _4812_/A1 _4812_/A2 _5179_/B _4812_/B _5000_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_5792_ _5855_/I0 hold833/Z _5793_/S _5792_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4743_ _4743_/A1 _4740_/Z _4741_/Z _5111_/C _4747_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xnet1002_256 net1152_425/I _6969_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1002_267 net952_206/I _6958_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_175_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet1002_278 net952_228/I _6947_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4674_ _4424_/B _5173_/A2 _5172_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xnet1002_289 net952_209/I _6936_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6413_ _6413_/I _6414_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3625_ _3625_/A1 _3625_/A2 _3625_/A3 _3866_/B _3625_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_162_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6344_ _7062_/Q _6257_/Z _6299_/Z _7054_/Q _6345_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_116_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3556_ _3525_/Z _5692_/A1 _5701_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_142_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6275_ _3328_/I _6296_/A2 _6484_/A2 _6275_/A4 _6275_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_170_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3487_ _6658_/Q _7305_/Q _3984_/S _3487_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5226_ _5226_/A1 _5310_/A2 _5226_/B _5226_/C _5227_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
Xinput109 wb_adr_i[22] _4026_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5157_ _5157_/A1 _5423_/A1 _5161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_99_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4108_ _5797_/I0 hold434/Z _4118_/S _4108_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5088_ _5340_/C _5417_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4039_ _6730_/Q _3464_/Z _6734_/Q _4040_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_25_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold308 _5653_/Z _7009_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold319 _6741_/Q hold319/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3410_ _6732_/Q _3409_/Z _3991_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4390_ _4391_/A1 _4391_/A2 _4391_/A3 _4391_/A4 _4390_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_124_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3341_ _6925_/Q _6336_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_171_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _6974_/Q _5964_/Z _5984_/Z _7112_/Q _6061_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_98_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold1008 _5787_/Z _7127_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_5011_ _5389_/C _5011_/A2 _5002_/Z _5194_/B1 _5350_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1019 _7200_/Q _5869_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_78_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6962_ _6962_/D _7149_/RN _6962_/CLK _6962_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5913_ _5913_/I _5952_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6893_ _6893_/D _6894_/RN _6893_/CLK _6893_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5844_ _5889_/I0 hold126/Z _5847_/S _5844_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5775_ _5775_/I0 hold651/Z _5775_/S _5775_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4726_ _5401_/A2 _5222_/A1 _5090_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_148_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4657_ _4657_/A1 _4654_/Z _4657_/A3 _4656_/Z _4664_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_162_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput80 spi_sck input80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3608_ _3589_/Z _3596_/Z _3607_/Z _6571_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xhold820 _5723_/Z _7071_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xinput91 spimemio_flash_io3_do input91/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold831 _7092_/Q hold831/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4588_ _5146_/A1 _4635_/A4 _5205_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold842 _6613_/Z _7297_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold853 _6799_/Q hold853/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold864 _4172_/Z _6715_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6327_ _7021_/Q _6549_/A2 _6531_/A2 _6965_/Q _6327_/C _6328_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_162_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold875 _7147_/Q hold875/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3539_ _5611_/A1 _3525_/Z _3954_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_107_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold886 _5815_/Z _7152_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_103_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold897 _7112_/Q hold897/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6258_ _7206_/Q _6535_/A2 _6257_/Z _7060_/Q _6259_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_107_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5209_ _5438_/B _4397_/Z _5209_/A3 _5475_/A4 _5209_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6189_ _6690_/Q _5985_/Z _5999_/Z _6847_/Q _6822_/Q _5964_/Z _6193_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_29_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3890_ _7135_/Q _3951_/A2 _3924_/B1 _6821_/Q _3951_/C1 _7143_/Q _3895_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_32_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5560_ _5833_/I0 hold467/Z _5565_/S _5560_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4511_ _4930_/A1 _5343_/B _4715_/A1 _4878_/A4 _4511_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_185_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5491_ _5857_/A1 _5857_/A2 hold212/I _5857_/A4 _5493_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_156_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold105 _4251_/Z _6767_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7230_ _7230_/D _7255_/RN _7257_/CLK _7230_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
Xhold116 _6916_/Q hold116/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4442_ _4380_/Z _4579_/A2 _4607_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold127 _5844_/Z _7178_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold138 _5494_/Z _5496_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_172_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold149 _6861_/Q _3307_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_132_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7161_ _7161_/D _7194_/RN _7161_/CLK _7161_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_125_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4373_ _4501_/B _5288_/C _4369_/Z _4373_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XTAP_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6112_ _6529_/S _6109_/Z _6112_/A3 _6112_/B _6113_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
Xfanout607 _5270_/A2 _5269_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3324_ _3324_/I _5957_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
Xfanout618 _3407_/ZN _4652_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7092_ _7092_/D _7173_/RN _7092_/CLK _7092_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout629 _5097_/B2 _5129_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_101_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6043_ _7022_/Q _6211_/A2 _6211_/B1 _6990_/Q _6051_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ _6945_/D _7002_/RN _6945_/CLK _6945_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_81_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6876_ _6876_/D _6882_/RN _6876_/CLK _6876_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5827_ _5827_/I0 hold829/Z _5829_/S _5827_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5758_ _5758_/A1 hold33/Z _5766_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_148_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4709_ _5459_/A1 _5098_/B _4705_/Z _4709_/A4 _4709_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5689_ hold351/Z _5827_/I0 _5691_/S _5689_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold650 _4169_/Z _6713_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_151_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold661 _6697_/Q hold661/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_78_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold672 _4147_/Z _6696_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold683 _7187_/Q hold683/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold694 _4358_/Z _6856_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_77_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__16 _4073__28/I _7209_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__27 _4073__27/I _7198_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__38 _4073__39/I _7187_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__49 _4073__49/I _7176_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4991_ _5340_/A1 _5370_/B _4991_/B _4991_/C _4993_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_1_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6730_ _6730_/D _6621_/Z _7304_/CLK _6730_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_189_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3942_ _3907_/Z _3942_/A2 _7036_/Q _5683_/A1 _3942_/C1 _6853_/Q _3944_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_189_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6661_ _6661_/D _6616_/Z _4072_/B2 _6661_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3873_ _3873_/A1 _3873_/A2 _3873_/A3 _3873_/A4 _3873_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5612_ _5867_/I0 hold975/Z _5619_/S _5612_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6592_ _6592_/A1 _6601_/A2 _6592_/B _6593_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_20_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5543_ _5888_/I0 hold283/Z _5547_/S _5543_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5474_ _5474_/A1 _5299_/C _5466_/Z _5473_/Z _5474_/C _6864_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_105_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7213_ _7213_/D _7220_/RN _7213_/CLK _7213_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4425_ _4395_/B _4373_/Z _4485_/A2 _4390_/Z _4721_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_172_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7144_ _7144_/D _6967_/RN _7144_/CLK _7144_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xfanout404 _5948_/Z _6544_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_4356_ _5857_/A1 _3560_/Z _5857_/A4 _4358_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
Xfanout415 _3517_/ZN _5839_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout426 _6164_/A2 _6211_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_87_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout437 _5884_/A3 _5857_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_101_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3307_ _3307_/I hold150/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout448 _6282_/A4 _6452_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_113_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7075_ _7075_/D _7075_/RN _7075_/CLK _7075_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout459 _4700_/Z _5478_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4287_ _6570_/I0 _6797_/Q _4288_/S _6797_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6026_ _6026_/A1 _6026_/A2 _6026_/A3 _6026_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_100_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6928_ _6928_/D _7258_/RN _6928_/CLK _6928_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_22_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6859_ _6859_/D _6865_/RN _6865_/CLK _6859_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_167_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold480 _7072_/Q hold480/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold491 _5626_/Z _6985_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_1_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4210_ hold265/Z _5547_/I0 _4210_/S _4210_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5190_ _5201_/A1 _5190_/A2 _5438_/C _5435_/A2 _5190_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_69_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4141_ _5822_/I0 hold657/Z _4142_/S _4141_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4072_ _4117_/S _4072_/A2 _4072_/B1 _4072_/B2 _4072_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_62_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4974_ _5359_/A1 _4973_/Z _4975_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_51_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3925_ input34/Z _3925_/A2 _3925_/B1 _6824_/Q _6839_/Q _3925_/C2 _3926_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6713_ _6713_/D _6882_/RN _6713_/CLK _6713_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xnet952_203 net952_250/I _7022_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6644_ _6644_/A1 _6656_/A2 _6644_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_20_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3856_ _7013_/Q _5656_/A1 _5638_/A1 _6997_/Q _5665_/A1 _7021_/Q _3860_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xnet952_214 net952_218/I _7011_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet952_225 net952_225/I _7000_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet952_236 net952_244/I _6989_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet952_247 net952_247/I _6978_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6575_ _6575_/A1 _6575_/A2 _6606_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3787_ _7192_/Q _3909_/A2 _4202_/S input45/Z _4227_/S _4056_/I1 _3795_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_146_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5526_ hold175/Z _5645_/I1 _5527_/S _5526_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5457_ _5457_/A1 _5457_/A2 _5316_/Z _5457_/A4 _5457_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_161_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4408_ _4719_/A2 _4489_/A1 _4428_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5388_ _5388_/A1 _5202_/Z _5354_/Z _5388_/A4 _5388_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_120_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7127_ _7127_/D fanout655/Z _7127_/CLK _7127_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4339_ _4360_/I1 hold531/Z _4340_/S _4339_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7058_ _7058_/D _7220_/RN _7058_/CLK _7058_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_189_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6009_ _6009_/A1 _6009_/A2 _6009_/A3 _6008_/Z _6010_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_189_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3710_ _6976_/Q _3923_/A2 _3910_/A2 _6936_/Q _3956_/A2 _7122_/Q _3715_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_53_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4690_ _4736_/A1 _4736_/A3 _4690_/B _4690_/C _5099_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_147_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3641_ _6704_/Q _3927_/A2 _3924_/A2 _6970_/Q _3642_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xclkbuf_leaf_33__1359_ _4073__24/I net852_120/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_113__1359_ clkbuf_4_4_0__1359_/Z net952_244/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6360_ _6966_/Q _6531_/A2 _6552_/A2 _7030_/Q _6360_/C _6363_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xclkbuf_leaf_96__1359_ clkbuf_4_5_0__1359_/Z net1102_394/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3572_ _5692_/A1 _5830_/A1 _3952_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5311_ _5308_/Z _5479_/A3 _5318_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_53_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6291_ _7190_/Q _6285_/Z _6290_/Z _7078_/Q _6307_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_114_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet902_155 net802_68/I _7070_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_166 net802_94/I _7059_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_177 net952_225/I _7048_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5242_ _4812_/B _5242_/A2 _5242_/A3 _4810_/B _5242_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_130_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet902_188 _4073__51/I _7037_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_199 net902_199/I _7026_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5173_ _4424_/B _5173_/A2 _5269_/A2 _4997_/C _5173_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4124_ hold20/Z _6678_/Q _4127_/S hold21/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput1 debug_mode input1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_84_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4055_ _6766_/Q input81/Z _4055_/S _4055_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1052_305 net1152_415/I _6920_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1052_316 _4073__32/I _6909_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_327 net1152_425/I _6898_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_338 net1052_346/I _6887_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xnet1052_349 net1202_490/I _6876_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_4957_ _5389_/A2 _5248_/A3 _5248_/A2 _4958_/A4 _4957_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3908_ _5517_/A1 _5517_/A2 _5517_/A3 _3942_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_131_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4888_ _5263_/A2 _5478_/B1 _5445_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_178_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6627_ _6844_/RN _6652_/A2 _6627_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3839_ _5884_/A1 _3680_/Z _3922_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_119_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6558_ _7260_/Q _6558_/I1 _6558_/S _7260_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5509_ _6888_/Q hold40/Z _5509_/S hold41/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6489_ _6489_/I _6490_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5860_ _5860_/I0 hold236/Z _5865_/S _5860_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4811_ _5094_/C _5312_/A2 _5137_/B1 _5220_/B2 _5179_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_179_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5791_ _5890_/I0 hold203/Z _5793_/S _5791_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4742_ _5478_/A3 _4695_/Z _5401_/A2 _5226_/C _5111_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_119_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet1002_257 net952_225/I _6968_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1002_268 net852_146/I _6957_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4673_ _5420_/A3 _5129_/A3 _3404_/I _3402_/I _4673_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_174_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1002_279 net952_228/I _6946_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6412_ _7024_/Q _6549_/A2 _6549_/C1 _7000_/Q _6288_/Z _7122_/Q _6413_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3624_ _7058_/Q _5701_/A1 _5674_/A1 _7034_/Q _3952_/A2 _7050_/Q _3625_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_179_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6343_ hold84/I _6290_/Z _6357_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3555_ _3507_/Z _3732_/A4 _3951_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6274_ _6296_/A2 _6282_/A1 _6302_/A3 _6300_/A4 _6274_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_0_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3486_ _7305_/Q _3984_/S _3987_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_102_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5225_ _4728_/Z _5310_/A2 _5225_/B _5310_/C _5229_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_29_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5156_ _5356_/A1 _5403_/B2 _5156_/B _5423_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_130_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4107_ hold1/Z _4107_/I1 _4117_/S hold2/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5087_ _5087_/A1 _4982_/Z _5340_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_186_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4038_ _4038_/A1 _6561_/B2 _6826_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_72_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5989_ _7142_/Q _5987_/Z _5988_/Z _6980_/Q _6009_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_24_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput190 _3352_/ZN mgmt_gpio_oeb[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_88_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_2_0__1359_ _4073__6/I clkbuf_opt_2_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_189_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold309 _7138_/Q hold309/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_183_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _5010_/A1 _4517_/Z _5435_/A2 _4606_/Z _5192_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold1009 _7046_/Q _5695_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_39_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6961_ _6961_/D _7083_/RN _6961_/CLK _6961_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_81_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5912_ _6743_/Q _4009_/B _5913_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6892_ _6892_/D _6892_/RN _6892_/CLK _6892_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_146_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5843_ _5888_/I0 hold363/Z _5847_/S _5843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5774_ _5855_/I0 hold887/Z _5775_/S _5774_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4725_ _5236_/A1 _5325_/B _4727_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_175_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4656_ _4960_/A1 _4374_/Z _5165_/A4 _5209_/A3 _4656_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_147_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput70 mgmt_gpio_in[7] input70/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3607_ _3601_/Z _3607_/A2 _3606_/Z _3607_/A4 _3607_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xinput81 spi_sdo input81/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold810 _4129_/Z _6682_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold821 _7113_/Q hold821/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4587_ _5269_/A1 _5269_/A2 _4635_/A4 _5367_/A2 _4587_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xinput92 spimemio_flash_io3_oeb input92/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold832 _5747_/Z _7092_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold843 _7148_/Q hold843/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold854 _4290_/Z _6799_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6326_ _7079_/Q _6290_/Z _6302_/Z _7087_/Q _6326_/C _6328_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3538_ _3505_/Z _5767_/A3 _3943_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold865 _7085_/Q hold865/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold876 _5809_/Z _7147_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_153_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold887 _7116_/Q hold887/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold898 _5770_/Z _7112_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_103_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6257_ _6484_/A3 _6282_/A2 _7232_/Q _6452_/A4 _6257_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3469_ _3991_/A1 _3469_/A2 _7280_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_153_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5208_ _5206_/Z _4662_/B _5433_/A1 _5208_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_88_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6188_ _6857_/Q _5924_/Z _6201_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5139_ _4376_/Z _5139_/A2 _5139_/A3 _5276_/B _5139_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_123_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_180_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4510_ _5420_/A2 _3403_/I _3404_/I _5129_/A4 _4510_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_184_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5490_ _5490_/A1 _5299_/C _5466_/Z _5489_/Z _5490_/C _6865_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_7_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold106 _7100_/Q hold106/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4441_ _4960_/A1 _5315_/A1 _4884_/A1 _4441_/B _4579_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_156_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold117 _5549_/Z _6916_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_145_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold128 _6771_/Q hold128/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold139 _5495_/Z _6876_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7160_ _7160_/D _7207_/RN _7160_/CLK _7160_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4372_ _4853_/A1 _4884_/A1 _4759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_153_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6111_ _6529_/S _7244_/Q _6112_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout608 _4454_/Z _5270_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_3323_ _6832_/Q _4096_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7091_ _7091_/D _7211_/RN _7091_/CLK _7091_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout619 _4522_/A2 _5288_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6042_ _7168_/Q _6006_/Z _6053_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6944_ _6944_/D _7238_/RN _6944_/CLK _6944_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_54_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6875_ _6875_/D _6633_/Z _4075_/I1 _6875_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_34_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5826_ hold20/Z hold78/Z _5829_/S hold79/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5757_ _5865_/I0 hold601/Z _5757_/S _5757_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4708_ _4708_/A1 _5312_/A2 _5312_/A1 _5094_/C _4709_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_163_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5688_ hold112/Z hold20/Z _5691_/S _5688_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4639_ _4639_/A1 _5039_/A4 _4638_/Z _4644_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_135_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold640 _4193_/Z _6729_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_151_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold651 _7117_/Q hold651/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold662 _4148_/Z _6697_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold673 _7066_/Q hold673/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold684 _5854_/Z _7187_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6309_ _6554_/A1 _6924_/Q _6310_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold695 _6964_/Q hold695/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7289_ _7289_/D _6643_/Z _7302_/CLK hold14/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_131_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__17 _4073__17/I _7208_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073__28 _4073__28/I _7197_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__39 _4073__39/I _7186_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4990_ _4990_/A1 _4892_/B _4991_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_1_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3941_ _7158_/Q _3941_/A2 _3941_/B1 _7166_/Q _3941_/C _3944_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_95_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3872_ _6675_/Q _3546_/Z _3945_/C2 _6683_/Q _3873_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6660_ _6660_/D _6615_/Z _4072_/B2 _6660_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_177_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5611_ _5611_/A1 _5848_/A3 _5821_/A3 _5857_/A3 _5619_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_83_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6591_ _6600_/A1 _6591_/A2 _6591_/B1 _3316_/I _3317_/I _6591_/C2 _6592_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5542_ _5860_/I0 hold92/Z _5547_/S hold93/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5473_ _5469_/Z _5489_/A2 _5472_/Z _5473_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_117_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7212_ _7212_/D _7220_/RN _7212_/CLK _7212_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4424_ _4374_/Z _4489_/A1 _4424_/B _4721_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_144_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4355_ _5538_/I1 hold997/Z _4355_/S _4355_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7143_ _7143_/D _6821_/RN _7143_/CLK _7143_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xfanout405 _5442_/A2 _5323_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout416 hold151/Z _3904_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout427 _5959_/ZN _6164_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_3306_ _6860_/Q _5185_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout438 _5848_/A3 _5866_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7074_ _7074_/D _7220_/RN _7074_/CLK _7074_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4286_ _6569_/I0 _6796_/Q _4288_/S _6796_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout449 _6299_/A2 _6533_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_101_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6025_ _7053_/Q _5924_/Z _6002_/Z _7087_/Q _6118_/B _6026_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_74_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6927_ _6927_/D _7215_/RN _6927_/CLK _6927_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_70_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6858_ _6858_/D _7154_/RN _6858_/CLK _6858_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_11_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5809_ _5818_/I0 hold875/Z _5811_/S _5809_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6789_ _6789_/D _6839_/RN _6789_/CLK _6789_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_155_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold470 _5531_/Z _6902_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_145_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold481 _5724_/Z _7072_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_78_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold492 hold492/I hold492/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_150_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4140_ _5857_/A1 _5857_/A2 _4347_/A3 _5857_/A4 _4142_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_68_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4071_ _3994_/Z _4117_/S _4072_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_83_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_56__1359_ clkbuf_4_14_0__1359_/Z net902_162/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_136__1359_ net1152_446/I net1102_382/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4973_ _5324_/A1 _5263_/A4 _4718_/B _4973_/A4 _4973_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6712_ _6712_/D _6882_/RN _6712_/CLK _6712_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3924_ _6964_/Q _3924_/A2 _3924_/B1 _6820_/Q _3926_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_20_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet952_204 net952_250/I _7021_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6643_ _6644_/A1 _6656_/A2 _6643_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3855_ _3855_/A1 _3855_/A2 _3855_/A3 _3855_/A4 _3855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xnet952_215 net952_218/I _7010_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet952_226 net952_226/I _6999_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet952_237 net802_91/I _6988_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet952_248 net952_248/I _6977_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3786_ _3786_/A1 _3786_/A2 _3786_/A3 _3786_/A4 _3786_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6574_ _6575_/A2 _6574_/A2 _6605_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5525_ hold217/Z _5818_/I0 _5527_/S _5525_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5456_ _5456_/A1 _5456_/A2 _5456_/B _5457_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_133_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4407_ _4428_/A2 _4395_/B _4407_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_5387_ _5387_/A1 _5387_/A2 _5387_/B _5388_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_87_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7126_ _7126_/D _7215_/RN _7126_/CLK _7126_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4338_ _4353_/A1 _5520_/C _5517_/A3 _5857_/A2 _4340_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7057_ _7057_/D _7163_/RN _7057_/CLK _7057_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4269_ hold158/Z _5645_/I1 _4270_/S _4269_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6008_ _6008_/A1 _6008_/A2 _6008_/A3 _6008_/A4 _6008_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_28_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3640_ _6962_/Q _3957_/A2 _3901_/A2 _6986_/Q _3642_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_140_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3571_ _5830_/A1 _5839_/A2 _3941_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_143_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5310_ _4728_/Z _5310_/A2 _5310_/B _5310_/C _5479_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_155_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6290_ _6484_/A3 _6300_/A4 _6300_/A1 _6299_/A2 _6290_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_154_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet902_156 net802_99/I _7069_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet902_167 _4073__45/I _7058_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_46_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet902_178 net902_194/I _7047_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5241_ _5321_/A1 _5241_/A2 _5451_/B _5242_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_115_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet902_189 net902_189/I _7036_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5172_ _5172_/A1 _5368_/A1 _5172_/B _5172_/C _5380_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_96_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4123_ _5834_/I0 hold349/Z _4127_/S _4123_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 debug_oeb input2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4054_ _6764_/Q input78/Z _4055_/S _4054_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1052_306 net1152_416/I _6919_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1052_317 _4073__32/I _6908_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_328 net1052_328/I _6897_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1052_339 net802_75/I _6886_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4956_ _5020_/A2 _4761_/I _4959_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3907_ _7300_/Q _7283_/Q _6893_/Q _3907_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_20_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ _4887_/A1 _5315_/A2 _5290_/A2 _5380_/B2 _4887_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6626_ _6844_/RN _6652_/A2 _6626_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3838_ _5884_/A1 _3617_/Z _3920_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_165_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6557_ _6557_/I _6558_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3769_ _7038_/Q _5683_/A1 _5674_/A1 _7030_/Q _3912_/B1 _6885_/Q _3773_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_118_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5508_ hold110/Z hold20/Z _5509_/S _5508_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6488_ _7149_/Q _6292_/Z _6300_/Z _7109_/Q _6489_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_10_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5439_ _5439_/A1 _5468_/A1 _5439_/B1 _5439_/B2 _5439_/C _5440_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_160_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7109_ _7109_/D _7253_/RN _7109_/CLK _7109_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_75_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4810_ _4997_/C _5380_/B2 _5478_/A2 _4810_/B _4812_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XTAP_2280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ _5880_/I0 hold185/Z _5793_/S _5790_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4741_ _5236_/A1 _5478_/A3 _4695_/Z _5226_/C _4741_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xnet1002_258 net952_247/I _6967_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4672_ _5269_/A2 _4672_/A2 _5291_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xnet1002_269 net902_181/I _6956_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6411_ _6401_/Z _6408_/Z _6411_/A3 _6411_/A4 _6411_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_135_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3623_ _7108_/Q _5758_/A1 _5683_/A1 _7042_/Q _6930_/Q _3935_/A2 _3625_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_116_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6342_ _7070_/Q _6484_/A2 _6452_/A3 _6452_/A4 _6348_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3554_ _3505_/Z _5839_/A2 _3930_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_115_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3485_ hold256/Z _5620_/A4 _3480_/Z _3484_/Z _3485_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6273_ _6484_/A2 _6300_/A4 _6300_/A1 _6275_/A4 _6273_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5224_ _5224_/A1 _5224_/A2 _5401_/B _5400_/A2 _5225_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_102_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5155_ _5275_/B _5153_/Z _5157_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_29_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4106_ _5796_/I0 hold791/Z _4118_/S _4106_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5086_ _5086_/A1 _5412_/A1 _5412_/A2 _5260_/B _5182_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_56_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4037_ _4036_/I _6826_/Q _6561_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_186_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5988_ _5991_/A2 _6021_/A4 _6002_/A2 _6139_/A2 _5988_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_36_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4939_ _4939_/A1 _5061_/B _4937_/Z _4938_/Z _4939_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_178_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6609_ _6608_/Z _6833_/Q _6830_/Q _4313_/Z _6610_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_166_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput180 _3361_/ZN mgmt_gpio_oeb[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_121_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput191 _3351_/ZN mgmt_gpio_oeb[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_88_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet802_100 net952_239/I _7125_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6960_ _6960_/D _7140_/RN _6960_/CLK _6960_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_47_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5911_ _5911_/A1 _5901_/B _5911_/B _7226_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6891_ _6891_/D _6894_/RN _6891_/CLK _6891_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_59_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5842_ _5842_/I0 hold355/Z _5847_/S _5842_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5773_ hold40/Z hold44/Z _5775_/S hold45/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4724_ _5248_/A3 _4500_/Z _4973_/A4 _5248_/A2 _5325_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_175_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4655_ _5043_/A2 _5043_/B _4657_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold800 _5559_/Z _6925_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3606_ _3606_/A1 _3606_/A2 _3606_/A3 _3606_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xinput60 mgmt_gpio_in[31] input60/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold811 _7017_/Q hold811/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xinput71 mgmt_gpio_in[8] input71/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput82 spi_sdoenb input82/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4586_ _5288_/B _5281_/C _4652_/A1 _4472_/B _4586_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xinput93 trap _3339_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold822 _5771_/Z _7113_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold833 _7132_/Q hold833/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6325_ _6325_/I _6326_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold844 _5810_/Z _7148_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold855 _6998_/Q hold855/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3537_ hold137/Z _3481_/I _3484_/Z hold256/Z _3537_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_66_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold866 _5739_/Z _7085_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold877 _6810_/Q hold877/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold888 _5774_/Z _7116_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold899 _6711_/Q hold899/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6256_ _6282_/A1 _6300_/A4 _6296_/A2 _6533_/A3 _6256_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3468_ _7295_/Q hold8/Z _3469_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_130_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5207_ _4662_/B _5433_/A1 _5362_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6187_ _6187_/A1 _5991_/Z _6192_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3399_ _3399_/I _6598_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5138_ _5138_/A1 _5278_/B _5148_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_85_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5069_ _4761_/I _5078_/A2 _5070_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_72_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4440_ _4436_/B _4648_/A1 _4440_/B _4604_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold107 _5756_/Z _7100_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold118 _6769_/Q hold118/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold129 _4256_/Z _6771_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_160_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4371_ _4836_/A3 _4456_/B _4456_/C _3407_/I _4497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_113_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6110_ _6201_/A3 _6928_/Q _6112_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3322_ _5951_/B _4005_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7090_ _7090_/D _7090_/RN _7090_/CLK _7090_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_140_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout609 _4422_/Z _5173_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _7242_/Q _6041_/I1 _6450_/S _7242_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6943_ _6943_/D _7238_/RN _6943_/CLK _6943_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_183_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6874_ _6874_/D _6632_/Z _4075_/I1 _6874_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_5825_ _5834_/I0 hold242/Z _5829_/S _5825_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5756_ hold16/Z hold106/Z _5757_/S _5756_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4707_ _5420_/A3 _5269_/A2 _4708_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_147_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5687_ hold375/Z _5852_/I0 _5691_/S _5687_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4638_ _4436_/B _4638_/A2 _5356_/C _5356_/A1 _4638_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold630 _4349_/Z _6850_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold641 _6695_/Q hold641/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4569_ _5364_/B _5438_/A1 _5356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_150_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold652 _5775_/Z _7117_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold663 _7215_/Q hold663/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6308_ _6554_/A1 _6307_/Z _6271_/Z _6308_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_150_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold674 _5717_/Z _7066_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold685 _7197_/Q hold685/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7288_ _7288_/D _6642_/Z _7304_/CLK hold38/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold696 _5603_/Z _6964_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_134_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6239_ _6300_/A4 _6285_/A2 _7237_/Q _3329_/I _6239_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7238__751 _7238_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_72_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__18 _4073__42/I _7207_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_150_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__29 _4073__4/I _7196_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3940_ _3940_/I _3941_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_189_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3871_ _6697_/Q _4146_/A1 _3936_/B1 _6691_/Q _3873_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_189_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5610_ _5784_/I0 hold769/Z _5610_/S _5610_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6590_ _6590_/I0 _7273_/Q _6602_/S _7273_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5541_ hold54/Z hold74/Z _5547_/S hold75/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_16__1359_ net1152_430/I _4073__7/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_118_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5472_ _5472_/A1 _5472_/A2 _4841_/B _5472_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_145_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7211_ _7211_/D _7211_/RN _7211_/CLK _7211_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xclkbuf_leaf_79__1359_ clkbuf_4_7_0__1359_/Z net802_62/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4423_ _4373_/Z _4385_/Z _4922_/A3 _4423_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_160_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7142_ _7142_/D fanout658/Z _7142_/CLK _7142_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_113_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4354_ _4103_/I hold883/Z _4355_/S _4354_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout406 _5248_/A3 _5442_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout417 _3478_/Z _5620_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3305_ _3305_/I _3500_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout428 _6452_/A3 _6484_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout439 _5848_/A3 _5875_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7073_ hold47/Z _7075_/RN _7073_/CLK hold46/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4285_ _6568_/I0 _6795_/Q _4288_/S _6795_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6024_ _6981_/Q _5988_/Z _6015_/Z _7005_/Q _6024_/C _6026_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_100_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6926_ _6926_/D _7211_/RN _6926_/CLK _6926_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6857_ _6857_/D _7154_/RN _6857_/CLK _6857_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_50_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5808_ _5808_/I0 hold729/Z _5811_/S _5808_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6788_ _6788_/D _6886_/RN _6788_/CLK _6788_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_10_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5739_ _5811_/I0 hold865/Z _5739_/S _5739_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold460 _6951_/Q hold460/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold471 _7015_/Q hold471/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold482 _7025_/Q hold482/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_2_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold493 _6762_/Q hold493/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_132_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_2__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _7304_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4070_ _7240_/Q _6896_/Q _6900_/Q _4070_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_3__1359_ net1152_451/I net1202_474/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4972_ _4496_/Z _5262_/A2 _5248_/A3 _4982_/A2 _4972_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6711_ _6711_/D _6894_/RN _6711_/CLK _6711_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3923_ _6972_/Q _3923_/A2 _3923_/B1 _6837_/Q _3923_/C1 _7078_/Q _3926_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_60_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6642_ _6644_/A1 _6650_/A2 _6642_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_60_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3854_ _7191_/Q _3909_/A2 _4210_/S input44/Z _3854_/C _3855_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_32_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet952_205 net952_248/I _7020_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet952_216 net952_216/I _7009_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet952_227 net952_227/I _6998_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet952_238 net952_238/I _6987_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6573_ _6575_/A2 _6573_/A2 _6607_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xnet952_249 net952_250/I _6976_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3785_ _6934_/Q _3910_/A2 _3959_/C1 _7184_/Q _3785_/C _3786_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_30_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5524_ _5524_/I0 _5797_/I0 _5527_/S _5524_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5455_ _5455_/I _5485_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_59_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4406_ _4428_/A2 _4395_/B _4719_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_160_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5386_ _5386_/A1 _5432_/A1 _5386_/A3 _5434_/A1 _5386_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_114_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7125_ _7125_/D _7125_/RN _7125_/CLK _7125_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4337_ _4361_/I1 hold590/Z _4337_/S _4337_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7056_ _7056_/D _7163_/RN _7056_/CLK _7056_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4268_ hold367/Z _5881_/I0 _4270_/S _4268_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6007_ _7036_/Q _6005_/Z _6006_/Z _7166_/Q _6008_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4199_ _4198_/Z hold295/Z _4211_/S _4199_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6909_ hold75/Z _7193_/RN _6909_/CLK hold74/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_126_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_62__1359_ clkbuf_4_15_0__1359_/Z net1152_419/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_152_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_142__1359_ net1152_451/I net1202_453/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_6_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold290 _5765_/Z _7108_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3570_ _5776_/A1 _5794_/A2 _3956_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_128_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet902_157 net902_157/I _7068_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet902_168 net902_168/I _7057_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5240_ _5368_/A1 _5389_/A2 _5240_/B _5451_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xnet902_179 net902_179/I _7046_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5171_ _5169_/Z _5170_/Z _5175_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4122_ _5842_/I0 hold162/Z _4127_/S _4122_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4053_ _6763_/Q input80/Z _4055_/S _4053_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput3 debug_out input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet1052_307 net1152_416/I _6918_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_318 net1202_487/I _6907_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_329 net952_251/I _6896_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4955_ _4419_/Z _4951_/Z _4955_/B _5068_/B _4959_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3906_ _5884_/A1 _3578_/Z _3920_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_20_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4886_ _4880_/Z _4886_/A2 _4884_/Z _4885_/Z _4886_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_32_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6625_ _6771_/RN _6648_/A2 _6625_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3837_ input47/Z _4227_/S _3855_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_165_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6556_ _6529_/S _7259_/Q _6556_/B _6557_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3768_ _5510_/A2 _3540_/Z _5532_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5507_ hold287/Z _5834_/I0 _5509_/S _5507_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_4_5_0__1359_ clkbuf_0__1359_/Z clkbuf_4_5_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_3_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6487_ _7101_/Q _6250_/Z _6299_/Z _7059_/Q _6995_/Q _6237_/Z _6492_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3699_ _6887_/Q _3912_/B1 _3916_/B1 _6882_/Q _3701_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_134_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5438_ _5438_/A1 _5475_/A4 _5438_/B _5438_/C _5439_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
Xoutput340 _6818_/Q wb_dat_o[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_126_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5369_ _5369_/A1 _5369_/A2 _5369_/B _5369_/C _5421_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_59_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7108_ _7108_/D _7220_/RN _7108_/CLK _7108_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_19_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7039_ _7039_/D _7185_/RN _7039_/CLK _7039_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_142_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4740_ _5478_/A3 _4695_/Z _5226_/A1 _5226_/C _4740_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_1591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4671_ _4530_/I _3404_/I _5137_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xnet1002_259 net952_228/I _6966_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6410_ _7146_/Q _6292_/Z _6300_/Z _7106_/Q _7082_/Q _6290_/Z _6411_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3622_ _7180_/Q _3945_/A2 _3913_/A2 input18/Z _3941_/B1 _7172_/Q _3647_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_128_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6341_ _6934_/Q _6263_/Z _6266_/Z _7014_/Q _6355_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3553_ _3525_/Z _3732_/A4 _3945_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_155_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6272_ _6300_/A2 _6285_/A2 _7237_/Q _6282_/A4 _6272_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_131_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3484_ _4317_/A1 _3483_/Z _3484_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_5223_ _5094_/B _5223_/A2 _5223_/B _5223_/C _5400_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_116_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5154_ _4568_/Z _4624_/Z _5376_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_96_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4105_ hold52/Z _7271_/Q _4117_/S hold53/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5085_ _4987_/Z _5085_/A2 _5260_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4036_ _4036_/I _4045_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5987_ _6068_/A2 _7230_/Q _3389_/I _6210_/B _5987_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XPHY_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4938_ _4998_/A2 _5389_/A2 _5442_/A1 _5323_/B _4938_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_36_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4869_ _4869_/A1 _4866_/Z _4867_/Z _4868_/Z _4872_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_123_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6608_ _6608_/I0 _6608_/I1 _6832_/Q _6608_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6539_ _6729_/Q _6247_/Z _6297_/Z _7077_/Q _6547_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_137_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput170 _4089_/Z irq[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput181 _3360_/ZN mgmt_gpio_oeb[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput192 _3350_/ZN mgmt_gpio_oeb[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_130_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet802_101 net802_81/I _7124_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5910_ _5951_/B _4006_/Z _5910_/B _5910_/C _5911_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_6890_ _6890_/D _6892_/RN _6890_/CLK _6890_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_34_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5841_ _5886_/I0 _5841_/I1 _5847_/S _5841_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5772_ _5889_/I0 hold130/Z _5775_/S _5772_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4723_ _4982_/A2 _3408_/I _5248_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_187_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4654_ _4944_/A1 _5315_/A2 _4589_/Z _5458_/A4 _4654_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3605_ _7085_/Q _3923_/C1 _3956_/A2 _7125_/Q _3606_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xinput50 mgmt_gpio_in[22] input50/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput61 mgmt_gpio_in[32] input61/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold801 _7083_/Q hold801/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xinput72 mgmt_gpio_in[9] input72/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4585_ _4887_/A1 _5399_/A2 _5276_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold812 _5662_/Z _7017_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold823 _6800_/Q hold823/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xinput83 spimemio_flash_clk input83/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput94 uart_enabled _4059_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6324_ _7143_/Q _6292_/Z _6300_/Z _7103_/Q _6325_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_116_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold834 _5792_/Z _7132_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3536_ _5517_/A2 _4350_/A2 _3927_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold845 _6723_/Q hold845/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold856 _5641_/Z _6998_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold867 _7155_/Q hold867/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold878 _4303_/Z _6810_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6255_ _7134_/Q _6253_/Z _6254_/Z _7174_/Q _6259_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold889 _6963_/Q hold889/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_115_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3467_ _3467_/I _7282_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5206_ _5189_/Z _5203_/Z _5357_/A2 _5440_/A1 _5206_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6186_ _6845_/Q _6211_/A2 _6211_/B1 _6837_/Q _6187_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_112_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3398_ _3398_/I _6595_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_29_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5137_ _5276_/C _5137_/A2 _5137_/B1 _5279_/A2 _5370_/B _5138_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_84_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5068_ _5260_/A1 _4761_/I _5068_/B _5334_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_83_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4019_ _4006_/Z _4019_/A2 _4014_/Z _4019_/B _6745_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_25_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold108 _7098_/Q hold108/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_176_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold119 _4254_/Z _6769_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_99_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4370_ _4836_/A3 _4456_/B _4456_/C _4884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_99_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3321_ _7226_/Q _5911_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ _6040_/I _6041_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6942_ _6942_/D _7238_/RN _6942_/CLK _6942_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xclkbuf_leaf_119__1359_ net952_221/I _4073__23/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_81_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6873_ _6873_/D _6631_/Z _4075_/I1 _6873_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_50_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5824_ _5869_/I0 _5824_/I1 _5829_/S _5824_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5755_ _5881_/I0 hold771/Z _5757_/S _5755_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4706_ _4765_/A1 _4782_/A1 _5302_/B _5218_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_5686_ hold957/Z _5869_/I0 _5691_/S _5686_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4637_ _4565_/Z _5293_/B _5039_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold620 _4190_/Z _6727_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold631 _6933_/Q hold631/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4568_ _5129_/A3 _4835_/A2 _5129_/A4 _3402_/I _4568_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold642 _4145_/Z _6695_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_2_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold653 _6995_/Q hold653/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6307_ _6307_/A1 _6307_/A2 _6307_/A3 _6306_/Z _6307_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold664 _5886_/Z _7215_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3519_ _3653_/A1 _3500_/Z _3904_/A3 _3680_/A3 _3519_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold675 _7221_/Q hold675/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7287_ _7287_/D _6641_/Z _7304_/CLK hold18/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_103_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold686 _5865_/Z _7197_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4499_ _4759_/A2 _4759_/A3 _4718_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold697 _6790_/Q hold697/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6238_ _7020_/Q _6549_/A2 _6237_/Z _6988_/Q _6260_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_89_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6169_ _6169_/A1 _6169_/A2 _6169_/A3 _6169_/A4 _6169_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__19 net802_82/I _7206_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3870_ _7103_/Q _5758_/A1 _3947_/A2 _7095_/Q _3873_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_182_1065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5540_ hold64/Z hold82/Z _5547_/S hold83/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5471_ _5471_/A1 _5276_/B _4555_/C _5471_/B2 _5472_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_69_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7210_ _7210_/D _7211_/RN _7210_/CLK _7210_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_145_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4422_ _4402_/B _4026_/B _4026_/C _4422_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_172_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7141_ hold13/Z _7141_/RN _7141_/CLK _7141_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_132_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4353_ _4353_/A1 _5520_/C _5517_/A3 _5517_/A1 _4355_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xfanout407 _4721_/ZN _5248_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout418 _6268_/Z _6550_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_3304_ _3304_/I _4041_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
X_7072_ _7072_/D _7163_/RN _7072_/CLK _7072_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4284_ _6567_/I0 _6794_/Q _4288_/S _6794_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout429 _5947_/ZN _6452_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6023_ _6941_/Q _5972_/Z _6021_/Z _6997_/Q _6026_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_140_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6925_ _6925_/D _7098_/RN _6925_/CLK _6925_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6856_ _6856_/D _6856_/RN _6856_/CLK _6856_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5807_ _5852_/I0 hold815/Z _5811_/S _5807_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6787_ _6787_/D _6886_/RN _6787_/CLK _6787_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3999_ _3999_/I _6835_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5738_ _5837_/I0 hold835/Z _5739_/S _5738_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5669_ hold252/Z _5879_/I0 _5673_/S _5669_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold450 _7183_/Q hold450/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold461 _7028_/Q hold461/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold472 _5660_/Z _7015_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_1_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold483 _5671_/Z _7025_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold494 _4245_/Z _6762_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_38_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_102__1359_ clkbuf_4_5_0__1359_/Z net802_89/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_54_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_22__1359_ _4073__49/I net802_98/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_85__1359_ clkbuf_4_13_0__1359_/Z net902_199/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4971_ _5201_/A1 _4905_/Z _4975_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_51_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6710_ _6710_/D _6854_/RN _6710_/CLK _6710_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_32_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3922_ _6855_/Q _3922_/A2 _3922_/B1 _6692_/Q _3922_/C _3963_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_189_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3853_ _3853_/I _3854_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6641_ _6644_/A1 _6650_/A2 _6641_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_177_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet952_206 net952_206/I _7019_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet952_217 net952_225/I _7008_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet952_228 net952_228/I _6997_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3784_ _3784_/I _3785_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet952_239 net952_239/I _6986_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ _6575_/A2 _6572_/A2 _6608_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5523_ hold357/Z _5798_/I0 _5527_/S _5523_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5454_ _5454_/A1 _5454_/A2 _5454_/A3 _5453_/Z _5455_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_161_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4405_ _4489_/B _4395_/B _4722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5385_ _5385_/A1 _5389_/C _5439_/B1 _5393_/A1 _5385_/C _5434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_132_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4336_ _4360_/I1 hold535/Z _4337_/S _4336_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7124_ _7124_/D _7124_/RN _7124_/CLK _7124_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_59_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7055_ _7055_/D _7075_/RN _7055_/CLK _7055_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4267_ hold187/Z _5781_/I0 _4270_/S _4267_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6006_ _3385_/I _3386_/I _6021_/A4 _6164_/A2 _6006_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_189_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4198_ hold94/Z hold54/Z _4202_/S _4198_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6908_ hold83/Z _7193_/RN _6908_/CLK hold82/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6839_ _6839_/D _6839_/RN _6839_/CLK _6839_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_50_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold280 _5690_/Z _7042_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold291 _7043_/Q hold291/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_172_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet902_158 net802_94/I _7067_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet902_169 net902_184/I _7056_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5170_ _5172_/B _5170_/A2 _5170_/A3 _5172_/C _5170_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_170_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4121_ _4343_/I0 hold633/Z _4127_/S _4121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4052_ _4052_/I _4052_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput4 mask_rev_in[0] input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1052_308 net902_194/I _6917_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1052_319 net1202_452/I _6906_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4954_ _5464_/A1 _5324_/A1 _4759_/Z _5263_/A4 _5068_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_178_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3905_ _6894_/Q _3904_/Z _3944_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4885_ _4887_/A1 _5315_/A2 _4990_/A1 _5380_/B2 _4885_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_178_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6624_ _7225_/RN _6656_/A2 _6624_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3836_ _5884_/A2 _3932_/A2 _3914_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_119_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6555_ _6548_/Z _6554_/Z _6555_/B1 _6286_/Z _6555_/C _6556_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3767_ _6700_/Q _3927_/A2 _3786_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_118_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5506_ hold102/Z _5842_/I0 _5509_/S _5506_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3698_ _7056_/Q _5701_/A1 _5674_/A1 _7032_/Q _3952_/A2 _7048_/Q _3701_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6486_ _6486_/A1 _6486_/A2 _6486_/A3 _6486_/A4 _6486_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_69_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput330 _7265_/Q wb_dat_o[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_105_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5437_ _5437_/A1 _5437_/A2 _5436_/Z _5437_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xoutput341 _6801_/Q wb_dat_o[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5368_ _5368_/A1 _5276_/C _5368_/B _5368_/C _5369_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_7107_ _7107_/D _7211_/RN _7107_/CLK _7107_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_113_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4319_ _4318_/Z _6833_/Q _6832_/Q _6601_/A2 _6819_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5299_ _5210_/Z _5396_/A1 _5267_/Z _5298_/Z _5299_/C _5300_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_101_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7038_ _7038_/D _7211_/RN _7038_/CLK _7038_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_75_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout590 _6500_/C _3324_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_65_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4670_ _4670_/A1 _4667_/Z _4669_/Z _4670_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_174_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3621_ _6946_/Q _5575_/A1 _3642_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_116_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6340_ _7176_/Q _6254_/Z _6355_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3552_ hold256/Z _3552_/A2 _3484_/Z hold137/Z _3552_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_51_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6271_ _6260_/Z _6271_/A2 _6271_/A3 _6271_/A4 _6271_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3483_ _3483_/I0 _3470_/B _3978_/S _3483_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5222_ _5222_/A1 _5310_/A2 _5223_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_130_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5153_ _5150_/Z _5487_/A2 _5153_/A3 _5289_/A3 _5153_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_111_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4104_ _5795_/I0 hold797/Z _4118_/S _4104_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5084_ _5359_/A1 _4982_/Z _5085_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4035_ _4034_/Z _4035_/A2 _4035_/A3 _4035_/A4 _4036_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_38_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ _7110_/Q _5984_/Z _5985_/Z _7060_/Q _6009_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XPHY_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4937_ _4998_/A2 _5328_/A1 _5442_/A1 _5323_/B _4937_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4868_ _4868_/A1 _5399_/A1 _4873_/A3 _5478_/A2 _4868_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_177_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6607_ _4900_/B _6607_/A2 _6610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3819_ _5821_/A2 _3560_/Z _4182_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_165_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4799_ _5173_/A2 _4534_/Z _5438_/A1 _5312_/A1 _4799_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_119_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6538_ _6723_/Q _6292_/Z _6299_/Z _6858_/Q _6548_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_107_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6469_ _7010_/Q _6549_/B1 _6552_/A2 _7034_/Q _6469_/C _6472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput171 _4065_/Z mgmt_gpio_oeb[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_82_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput182 _4064_/Z mgmt_gpio_oeb[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput193 _3377_/ZN mgmt_gpio_oeb[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_43_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5840_ _5867_/I0 _5840_/I1 _5847_/S _5840_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5771_ _5852_/I0 hold821/Z _5775_/S _5771_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4722_ _5083_/C _4722_/A2 _4923_/A2 _5080_/B _4976_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_175_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4653_ _4653_/A1 _5040_/C _4653_/A3 _5041_/B _4657_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_147_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput40 mgmt_gpio_in[13] input40/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3604_ _7149_/Q _3951_/C1 _5638_/A1 _7003_/Q _3606_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xinput51 mgmt_gpio_in[23] input51/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold802 _5737_/Z _7083_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xinput62 mgmt_gpio_in[33] input62/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4584_ _4584_/A1 _4584_/A2 _5349_/B _4591_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xinput73 pad_flash_io0_di input73/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput84 spimemio_flash_csb input84/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold813 _7003_/Q hold813/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_115_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold824 _4291_/Z _6800_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6323_ _7095_/Q _6250_/Z _6257_/Z _7061_/Q _6536_/B1 _7037_/Q _6328_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_116_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput95 wb_adr_i[0] input95/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3535_ _3904_/A3 hold144/I _3500_/Z hold221/I _3535_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold835 _7084_/Q hold835/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold846 _4184_/Z _6723_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold857 _7149_/Q hold857/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold868 _5818_/Z _7155_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_88_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6254_ _7237_/Q _6533_/A3 _6452_/A4 _6285_/A2 _6254_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_131_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold879 _7164_/Q hold879/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3466_ _3465_/Z _3466_/A2 _4056_/I1 _3430_/S _3467_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5205_ _5205_/A1 _5468_/A1 _5205_/B1 _5356_/C _5205_/C _5440_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_69_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6185_ _7248_/Q _6185_/I1 _6558_/S _7248_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3397_ _3397_/I _6592_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_57_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5136_ _5287_/C _4570_/Z _4598_/Z _5164_/A4 _5374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_96_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5067_ _4951_/Z _5078_/A2 _5070_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4018_ _6743_/Q _6901_/Q _4019_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_26_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5969_ _6117_/A2 _6211_/B1 _6021_/A2 _6021_/A4 _5969_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_32_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold109 _5754_/Z _7098_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_137_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3320_ _7224_/Q _5954_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6941_ _6941_/D fanout659/Z _6941_/CLK _6941_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_6872_ _6872_/D _6630_/Z _4075_/I1 _6872_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_179_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5823_ _5832_/I0 hold995/Z _5829_/S _5823_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5754_ hold20/Z hold108/Z _5757_/S _5754_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4705_ _5220_/B2 _4536_/Z _4491_/B _4705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_147_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5685_ hold422/Z _5886_/I0 _5691_/S _5685_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4636_ _4636_/A1 _5034_/B _4635_/Z _4639_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_135_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold610 _5890_/Z _7219_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_118_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold621 _6706_/Q hold621/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_2_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4567_ _5270_/A1 _5270_/A2 _5389_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold632 _5568_/Z _6933_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold643 _6694_/Q hold643/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6306_ _6306_/A1 _6306_/A2 _6306_/A3 _6306_/A4 _6306_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold654 _5637_/Z _6995_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_162_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold665 _7211_/Q hold665/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3518_ hold144/Z hold211/I hold145/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_89_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold676 _5892_/Z _7221_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7286_ _7286_/D _6640_/Z _7304_/CLK hold58/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_104_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4498_ _4494_/Z _4496_/Z _4998_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold687 _7204_/Q hold687/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold698 _4279_/Z _6790_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6237_ _7235_/Q _6275_/A4 _6533_/A3 _5942_/S _6237_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3449_ _7292_/Q _3449_/A2 _3450_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_76_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6168_ _7059_/Q _5924_/Z _6015_/Z _7011_/Q _6168_/C _6169_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5119_ _4773_/Z _4874_/C _5238_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6099_ _7138_/Q _5994_/I _6015_/Z _7008_/Q _6944_/Q _5972_/Z _6101_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_27_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_125__1359_ net952_221/I net1102_379/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_45__1359_ clkbuf_4_14_0__1359_/Z _4073__17/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_68_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5470_ _5470_/A1 _5372_/Z _5470_/A3 _5489_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_172_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4421_ _4960_/A1 _5055_/A2 _4589_/A4 _4456_/C _4421_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_99_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7140_ hold17/Z _7140_/RN _7140_/CLK _7140_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4352_ _6613_/I1 hold596/Z _4352_/S _4352_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout408 _5056_/C _5442_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_3303_ _4113_/S _4317_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4283_ _6566_/I0 _6793_/Q _4288_/S _6793_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout419 _6263_/Z _6545_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_7071_ _7071_/D _7071_/RN _7071_/CLK _7071_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_113_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6022_ _7079_/Q _5996_/Z _6005_/Z _7037_/Q _6965_/Q _5979_/Z _6031_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_66_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6924_ _6924_/D _7179_/RN _6924_/CLK _6924_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_81_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6855_ _6855_/D _6856_/RN _6855_/CLK _6855_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5806_ _5806_/I0 hold955/Z _5811_/S _5806_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6786_ _6786_/D _6786_/RN _6786_/CLK _6786_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_167_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3998_ _6600_/B2 _4097_/A1 _6829_/Q _3999_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_183_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5737_ _5881_/I0 hold801/Z _5739_/S _5737_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5668_ hold396/Z _5797_/I0 _5673_/S _5668_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4619_ _4565_/Z _5290_/A3 _5029_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5599_ _5782_/I0 hold515/Z _5601_/S _5599_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold440 _7153_/Q hold440/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_150_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold451 _5850_/Z _7183_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold462 _5675_/Z _7028_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold473 _6943_/Q hold473/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold484 _6866_/Q hold484/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold495 _6923_/Q hold495/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7269_ _7269_/D _7269_/CLK _7269_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4970_ _4970_/A1 _4967_/Z _4968_/Z _4969_/Z _4975_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_63_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3921_ _3921_/I _3922_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_189_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6640_ _6650_/A1 _6650_/A2 _6640_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3852_ _7215_/Q _3912_/A2 _3922_/A2 _6856_/Q _3853_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_32_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet952_207 net802_95/I _7018_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet952_218 net952_218/I _7007_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6571_ _6571_/I0 _7269_/Q _6571_/S _7269_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet952_229 net952_229/I _6996_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3783_ _7022_/Q _5665_/A1 _3959_/B1 _6668_/Q _3923_/C1 hold84/I _3784_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5522_ hold430/Z _5724_/I0 _5527_/S _5522_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5453_ _5126_/I _5452_/Z _5129_/Z _5453_/A4 _5453_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_132_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4404_ _4424_/B _4428_/A2 _4922_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5384_ _6577_/C _5267_/Z _5382_/Z _5384_/B _6862_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_5_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7123_ _7123_/D _7260_/RN _7123_/CLK _7123_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4335_ _4350_/A3 _4353_/A1 hold146/Z _5857_/A2 _4337_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_101_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7054_ _7054_/D _7211_/RN _7054_/CLK _7054_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_140_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4266_ hold195/Z _5798_/I0 _4270_/S _4266_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_91__1359_ clkbuf_4_5_0__1359_/Z net952_248/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_189_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6005_ _7230_/Q _3389_/I _6117_/A4 _6139_/A2 _6005_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_189_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4197_ _4196_/Z hold335/Z _4211_/S _4197_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6907_ _6907_/D _6907_/RN _6907_/CLK _6907_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6838_ _6838_/D _6892_/RN _6838_/CLK _6838_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_126_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6769_ _6769_/D _6771_/RN _6769_/CLK _6769_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_137_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold270 _5501_/Z _6881_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_123_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold281 _7193_/Q hold281/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_78_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold292 _5691_/Z _7043_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_77_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout750 _4547_/A4 _4836_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_93_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_opt_5_0__1359_ _4073__24/I clkbuf_opt_5_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet902_159 net802_94/I _7066_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_151_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4120_ _5537_/I1 hold805/Z _4127_/S _4120_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4051_ _7201_/Q input82/Z _4055_/S _4052_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput5 mask_rev_in[10] input5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1052_309 net1152_419/I _6916_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4953_ _4953_/A1 _5065_/B _4953_/A3 _4955_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_51_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3904_ hold221/Z _3904_/A2 _3904_/A3 _3904_/A4 _3904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_60_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4884_ _4884_/A1 _4659_/Z _4675_/Z _5426_/A1 _4884_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6623_ _7224_/RN _6648_/A2 _6623_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_20_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3835_ _5884_/A1 _3560_/Z _3922_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_178_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6554_ _6554_/A1 _6554_/A2 _6554_/A3 _6553_/Z _6554_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3766_ input26/Z _3927_/C2 _3794_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5505_ hold424/Z _5538_/I1 _5509_/S _5505_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6485_ _7117_/Q _6240_/Z _6297_/Z _6705_/Q _6485_/C _6486_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3697_ _6944_/Q _5575_/A1 _3707_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_161_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5436_ _4576_/C _5472_/A2 _5009_/Z _5435_/Z _5436_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xoutput320 _6793_/Q wb_dat_o[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_10_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput331 _7266_/Q wb_dat_o[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput342 _6802_/Q wb_dat_o[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_126_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5367_ _5438_/A1 _5367_/A2 _5368_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_160_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7106_ _7106_/D _7202_/RN _7106_/CLK _7106_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4318_ _4316_/Z _4318_/A2 _6833_/D _6828_/Q _4318_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5298_ _5296_/Z _5382_/A3 _5173_/Z _5464_/B _5298_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_87_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7037_ _7037_/D _7098_/RN _7037_/CLK _7037_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_87_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4249_ _5860_/I0 hold90/Z _4252_/S hold91/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout580 _6834_/Q _3315_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout591 _6744_/Q _6500_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_18_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3620_ _6954_/Q _5584_/A1 _3630_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3551_ _3525_/Z _5767_/A3 _3917_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_115_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6270_ _6948_/Q _6550_/C1 _6552_/A2 _7028_/Q _6271_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3482_ _4041_/B1 _6662_/Q _3975_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_170_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5221_ _5221_/I _5401_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_102_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5152_ _5287_/B _5290_/A3 _5164_/A4 _4624_/Z _4570_/Z _5153_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_155_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4103_ _4103_/I _5520_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_29_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5083_ _4977_/Z _4981_/Z _5083_/B _5083_/C _5337_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_4034_ _4033_/Z _4034_/A2 _4388_/A2 _4388_/A1 _4034_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_64_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5985_ _7231_/Q _6210_/C _6002_/A3 _5914_/S _5985_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XPHY_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4936_ _4936_/I _5410_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_162_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_10 hold77/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4867_ _5269_/A2 _4530_/I _4873_/A3 _5293_/B _4867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_36_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6606_ _4686_/B _6606_/A2 _6610_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3818_ _4350_/A2 _5794_/A2 _3960_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_123_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4798_ _5438_/A1 _4793_/Z _5452_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_165_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6537_ _6717_/Q _6250_/Z _6290_/Z _6709_/Q _6302_/Z _6713_/Q _6548_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_146_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3749_ _7129_/Q _3930_/A2 _5758_/A1 _7105_/Q _3941_/B1 _7169_/Q _3751_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_174_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6468_ _6468_/I _6469_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5419_ _5419_/A1 _5419_/A2 _5418_/Z _5431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6399_ hold86/I _6543_/A2 _6285_/Z hold80/I _7178_/Q _6254_/Z _6401_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_82_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput172 _3369_/ZN mgmt_gpio_oeb[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_121_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput183 _3359_/ZN mgmt_gpio_oeb[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput194 _3349_/ZN mgmt_gpio_oeb[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_56_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet1102_390 net902_199/I _6784_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ _5833_/I0 hold897/Z _5775_/S _5770_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ _4721_/A1 _4721_/A2 _4721_/B _4721_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_148_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4652_ _4652_/A1 _5139_/A2 _5471_/B2 _4652_/A4 _5041_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xinput30 mask_rev_in[4] input30/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3603_ _7117_/Q _3917_/A2 _5758_/A1 _7109_/Q _5674_/A1 _7035_/Q _3606_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xinput41 mgmt_gpio_in[14] input41/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput52 mgmt_gpio_in[24] input52/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4583_ _4570_/Z _5016_/B2 _5349_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput63 mgmt_gpio_in[34] input63/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold803 _7035_/Q hold803/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xinput74 pad_flash_io1_di _3337_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6322_ _6322_/A1 _6322_/A2 _6322_/A3 _6322_/A4 _6322_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold814 _5646_/Z _7003_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold825 _7296_/Q hold825/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3534_ _3680_/A3 hold211/Z hold212/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xinput85 spimemio_flash_io0_do input85/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput96 wb_adr_i[10] input96/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold836 _5738_/Z _7084_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_171_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold847 _6939_/Q hold847/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_171_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold858 _5811_/Z _7149_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold869 _7019_/Q hold869/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6253_ _7236_/Q _6300_/A2 _6533_/A4 _6253_/A4 _6253_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_89_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3465_ _3464_/Z _3442_/B _3465_/A3 _3465_/A4 _3465_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xclkbuf_leaf_9__1359_ net1152_430/I net802_66/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_130_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5204_ _5346_/A2 _5387_/A1 _5403_/B2 _5205_/A1 _5204_/C _5357_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6184_ _6364_/C _6181_/Z _6184_/A3 _6184_/B _6185_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_112_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3396_ _3396_/I _6589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_130_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5135_ _4589_/Z _5142_/A3 _5287_/C _5487_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_85_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5066_ _4944_/Z _5078_/A2 _5066_/B _5481_/C _5070_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_4017_ _4006_/Z _4019_/A2 _4020_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5968_ _6014_/A2 _3389_/I _5968_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_40_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4919_ _5343_/A1 _4496_/Z _5442_/A1 _5323_/B _4927_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5899_ _5910_/B _5899_/I1 _7223_/Q _7223_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_68__1359_ clkbuf_4_13_0__1359_/Z net952_239/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_148__1359_ net1152_451/I net1152_410/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6940_ _6940_/D fanout659/Z _6940_/CLK _6940_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_47_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6871_ _6871_/D _6629_/Z _4075_/I1 _6871_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_34_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5822_ _5822_/I0 _5822_/I1 _5829_/S _5822_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5753_ _5834_/I0 hold240/Z _5757_/S _5753_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4704_ _4687_/Z _4704_/A2 _5255_/A2 _5092_/A1 _5098_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_31_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5684_ hold339/Z _5822_/I0 _5691_/S _5684_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4635_ _4868_/A1 _5399_/A1 _5146_/A1 _4635_/A4 _4635_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_162_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold600 hold600/I hold600/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _5290_/A1 _5278_/C _5290_/A2 _4877_/A2 _4576_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold611 _6701_/Q hold611/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold622 _4159_/Z _6706_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold633 _6675_/Q hold633/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold644 _4144_/Z _6694_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6305_ _7198_/Q _6540_/A2 _6536_/B1 _7036_/Q _6306_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_162_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3517_ _3489_/I _3492_/Z _3517_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold655 _7075_/Q hold655/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7285_ _7285_/D _6639_/Z _7302_/CLK hold1/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold666 _5881_/Z _7211_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4497_ _3408_/I _4497_/A2 _4497_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
Xhold677 _6693_/Q hold677/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_103_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold688 _5873_/Z _7204_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold699 _7196_/Q hold699/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6236_ _5943_/S _3329_/I _6484_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3448_ _3448_/I _7293_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6167_ _6947_/Q _5972_/Z _6021_/Z _7003_/Q _6169_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3379_ _6929_/Q _6447_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ _5115_/Z _5117_/Z _5118_/A3 _5215_/C _5118_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6098_ _7090_/Q _6002_/Z _6019_/Z _7048_/Q _6098_/C _6101_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_27_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5049_ _5049_/A1 _5210_/A4 _5180_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_2805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4420_ _5170_/A2 _4836_/A4 _5258_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4351_ _6612_/I1 hold588/Z _4352_/S _4351_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3302_ hold31/I _6608_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout409 _5731_/A2 _4185_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7070_ _7070_/D _7220_/RN _7070_/CLK _7070_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_141_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4282_ _6565_/I0 _6792_/Q _4288_/S _6792_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6021_ _6164_/B1 _6021_/A2 _6210_/A2 _6021_/A4 _6021_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_86_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6923_ _6923_/D _7221_/RN _6923_/CLK _6923_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6854_ _6854_/D _6854_/RN _6854_/CLK _6854_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_62_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5805_ _5877_/I0 _5805_/I1 _5811_/S _5805_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6785_ _6785_/D _6786_/RN _6785_/CLK _6785_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3997_ _3997_/I _6834_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_51__1359_ clkbuf_4_14_0__1359_/Z net852_150/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5736_ _5808_/I0 hold725/Z _5739_/S _5736_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_131__1359_ net1152_446/I net852_106/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5667_ hold603/Z _5877_/I0 _5673_/S _5667_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4618_ _4618_/A1 _5151_/B _4616_/Z _4617_/Z _4622_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_164_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5598_ _5871_/I0 hold404/Z _5601_/S _5598_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold430 _6895_/Q hold430/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold441 _5816_/Z _7153_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4549_ _5288_/B _4944_/A1 _3407_/I _4549_/A4 _4549_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_2_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold452 _6973_/Q hold452/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold463 _6975_/Q hold463/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold474 _5579_/Z _6943_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold485 _5492_/Z _6866_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7268_ _7268_/D _7269_/CLK _7268_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold496 _5556_/Z _6923_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6219_ _6844_/Q _5971_/Z _5981_/Z _6788_/Q _6005_/Z _6850_/Q _6220_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_7199_ _7199_/D _7207_/RN _7199_/CLK _7199_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_58_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3920_ input71/Z _4244_/S _3920_/B1 _6866_/Q _6902_/Q _3920_/C2 _3921_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_44_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3851_ _7159_/Q _3941_/A2 _3912_/C1 _6707_/Q _4170_/A1 _6715_/Q _3855_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_177_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet952_208 net952_208/I _7017_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6570_ _6570_/I0 _7268_/Q _6571_/S _7268_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet952_219 net952_227/I _7006_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3782_ _7014_/Q _5656_/A1 _5638_/A1 _6998_/Q _3951_/C1 _7144_/Q _3786_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5521_ hold28/Z _5521_/A2 _5647_/A2 _5620_/A4 _5521_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_158_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5452_ _4791_/Z _5452_/A2 _5452_/A3 _4801_/Z _5452_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_8_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4403_ _4424_/B _4428_/A2 _4923_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_126_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5383_ _6862_/Q _6577_/C _5212_/Z _5320_/Z _5383_/C _5384_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_7122_ _7122_/D _7122_/RN _7122_/CLK _7122_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4334_ _5778_/I0 hold767/Z _4334_/S _4334_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7053_ _7053_/D _6821_/RN _7053_/CLK _7053_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_114_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4265_ hold189/Z _5797_/I0 _4270_/S _4265_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6004_ _7086_/Q _6002_/Z _6003_/Z _7158_/Q _6008_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4196_ hold118/Z hold64/I _4202_/S _4196_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6906_ _6906_/D _6907_/RN _6906_/CLK _6906_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_165_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6837_ _6837_/D _6892_/RN _6837_/CLK _6837_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_7_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6768_ _6768_/D _7193_/RN _6768_/CLK _6768_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_148_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5719_ _5857_/A2 _5785_/A3 _5731_/A2 _5866_/A3 _5727_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6699_ _6699_/D _6892_/RN _6699_/CLK _6699_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_109_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold260 _5516_/Z _6892_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_105_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold271 _7123_/Q hold271/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold282 _5861_/Z _7193_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_160_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold293 _6784_/Q hold293/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_132_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout740 _5051_/S _3404_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_49_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_10_0__1359_ clkbuf_0__1359_/Z _4073__24/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_2432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4050_ _4050_/I0 input90/Z _4050_/S _4050_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 mask_rev_in[11] input6/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4952_ _5020_/A2 _4951_/Z _4953_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3903_ _3903_/A1 _5517_/A1 hold146/I _5517_/A2 _3903_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4883_ _4881_/Z _4882_/Z _4886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_32_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3834_ hold258/I _4350_/A2 _3956_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6622_ _7224_/RN _6648_/A2 _6622_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_6553_ _6553_/A1 _6553_/A2 _6553_/A3 _6553_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_177_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3765_ _7046_/Q _3952_/A2 _3916_/B1 hold76/I _3790_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_158_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5504_ hold337/Z _5537_/I1 _5509_/S _5504_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6484_ _7133_/Q _6484_/A2 _6484_/A3 _6484_/A4 _6485_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3696_ _7008_/Q _3934_/A2 _3701_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_173_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5435_ _5438_/C _5435_/A2 _5475_/A3 _5475_/A4 _5435_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xoutput310 _7261_/Q wb_ack_o VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_145_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput321 _6794_/Q wb_dat_o[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput332 _7267_/Q wb_dat_o[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_156_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5366_ _5366_/A1 _5366_/A2 _5365_/Z _5469_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_142_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7105_ _7105_/D _7177_/RN _7105_/CLK _7105_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4317_ _4317_/A1 _6826_/Q _4318_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_59_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5297_ _4882_/Z _5170_/Z _5382_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7036_ _7036_/D _6786_/RN _7036_/CLK _7036_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_75_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4248_ _5538_/I1 hold501/Z _4252_/S _4248_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4179_ _5517_/A1 _5517_/A3 _4185_/A2 _5520_/C _4181_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_56_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout570 _5991_/A2 _3386_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_93_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout581 _4113_/S _3500_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_47_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout592 _3304_/I _3984_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_20_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3550_ _5875_/A1 _3507_/Z _3955_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_127_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3481_ _3481_/I _3552_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_127_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5220_ _4694_/Z _5310_/A2 _5220_/B1 _5220_/B2 _5221_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
Xnet1152_450 net802_67/I _6715_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5151_ _5287_/C _5287_/B _5164_/A4 _5151_/B _5487_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_130_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4102_ input58/Z hold62/Z _4117_/S hold63/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5082_ _4980_/Z _5081_/Z _5412_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_110_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4033_ _4028_/Z _4030_/Z _4026_/B _4026_/C _4033_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_84_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ _5984_/A1 _6210_/B _6068_/A2 _7230_/Q _5984_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_52_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4935_ _5442_/A2 _4497_/Z _4982_/A2 _5056_/C _4936_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_20_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_11 _3477_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4866_ _4868_/A1 _5399_/A1 _5364_/A1 _4873_/A3 _4866_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_178_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6605_ _4415_/B _6605_/A2 _6610_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3817_ _5510_/A2 _5830_/A1 _5536_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4797_ _4791_/Z _5452_/A2 _5453_/A4 _4797_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_6536_ _6691_/Q _6257_/Z _6536_/B1 _6850_/Q _6300_/Z _6721_/Q _6548_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3748_ _6677_/Q _3546_/Z _3947_/A2 _7097_/Q _6896_/Q _5528_/S _3758_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_180_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3679_ hold152/Z _4347_/A3 _5503_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6467_ _7026_/Q _6549_/A2 _6531_/A2 _6970_/Q _6549_/C1 _7002_/Q _6468_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_161_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5418_ _5418_/A1 _5418_/A2 _5417_/Z _5418_/A4 _5418_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6398_ _7098_/Q _6250_/Z _6302_/Z _7090_/Q _6401_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_115_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput173 _3368_/ZN mgmt_gpio_oeb[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput184 _3358_/ZN mgmt_gpio_oeb[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5349_ _5349_/A1 _5387_/A2 _5349_/B _5350_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_87_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput195 _3348_/ZN mgmt_gpio_oeb[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7019_ _7019_/D _7019_/RN _7019_/CLK _7019_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_46_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_28__1359_ clkbuf_opt_2_0__1359_/Z net1152_409/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_108__1359_ clkbuf_4_4_0__1359_/Z net1202_494/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_78_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1102_380 net1202_481/I _6810_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1102_391 net1152_410/I _6783_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4720_ _5083_/C _5080_/B _5259_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_1391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4651_ _4903_/A1 _5458_/A4 _5295_/A2 _5295_/A3 _4651_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_159_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput20 mask_rev_in[24] input20/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3602_ _7213_/Q _3960_/A2 _3955_/A2 _7205_/Q _6955_/Q _5584_/A1 _3607_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xinput31 mask_rev_in[5] input31/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4582_ _4638_/A2 _5345_/A2 _4438_/B _4944_/A1 _5016_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xinput42 mgmt_gpio_in[15] input42/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput53 mgmt_gpio_in[25] input53/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput64 mgmt_gpio_in[35] input64/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput75 porb input75/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6321_ _7069_/Q _6248_/Z _6297_/Z _6699_/Q _6321_/C _6322_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3533_ hold27/Z hold137/Z _3481_/I _3484_/Z _3533_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold804 _5682_/Z _7035_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xinput86 spimemio_flash_io0_oeb input86/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold815 _7145_/Q hold815/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold826 _6612_/Z _7296_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold837 _7172_/Q hold837/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xinput97 wb_adr_i[11] input97/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold848 _5574_/Z _6939_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6252_ _7094_/Q _6250_/Z _6550_/B1 _6980_/Q _6259_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_66_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold859 _6714_/Q hold859/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_131_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3464_ _7283_/Q _3441_/C _6664_/Q _6663_/Q _3464_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_103_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5203_ _5199_/Z _5354_/A2 _5202_/Z _5203_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6183_ _6364_/C _7247_/Q _6184_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3395_ _3395_/I _6586_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_97_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5134_ _5293_/A1 _4624_/Z _5275_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_69_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ _5403_/A1 _5252_/B _5065_/B _5481_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4016_ _3324_/I _5896_/I0 _4019_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_65_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5967_ _3385_/I _5991_/A2 _5914_/S _6002_/A2 _5967_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4918_ _4927_/A1 _4927_/A2 _5444_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_166_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5898_ _5901_/B _5899_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_179_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4849_ _4598_/Z _4681_/Z _4849_/B _5373_/B _4852_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_138_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6519_ _6716_/Q _6250_/Z _6293_/Z _6718_/Q _6521_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_10_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6870_ _6870_/D _6628_/Z _4075_/I1 _6870_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_62_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5821_ _5821_/A1 _5821_/A2 _5821_/A3 _5857_/A3 _5829_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_50_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5752_ _5869_/I0 hold943/Z _5757_/S _5752_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4703_ _5420_/A2 _4930_/A1 _4835_/A2 _5129_/A4 _4703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_33_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5683_ _5683_/A1 hold33/Z _5691_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_148_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4634_ _4868_/A1 _5399_/A1 _5373_/A2 _5287_/B _5034_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_163_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold601 _7101_/Q hold601/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4565_ _4635_/A4 _4456_/C _4456_/B _5269_/A1 _4565_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_162_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold612 _4153_/Z _6701_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_128_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold623 _6705_/Q hold623/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold634 _4121_/Z _6675_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6304_ _7166_/Q _6544_/A2 _6273_/Z _6972_/Q _6306_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3516_ _5857_/A1 _5884_/A2 _3912_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_89_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold645 _6931_/Q hold645/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold656 _5727_/Z _7075_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4496_ _4944_/A1 _4497_/A2 _4496_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_7284_ _7284_/D _6638_/Z _7304_/CLK hold52/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold667 _6838_/Q hold667/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold678 _4142_/Z _6693_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_103_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold689 _7168_/Q hold689/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6235_ _3328_/I _6300_/A1 _6275_/A4 _6533_/A3 _6235_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3447_ _3447_/A1 _3449_/A2 _3447_/B1 _7292_/Q _3448_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_98_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3378_ _6928_/Q _6418_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6166_ _6987_/Q _5988_/Z _6019_/Z _7051_/Q _6169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xclkbuf_leaf_11__1359_ net1152_430/I net802_63/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5117_ _5117_/A1 _5117_/A2 _5117_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
X_6097_ _6097_/I _6098_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5048_ _5395_/A1 _4991_/C _5210_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_66_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6999_ _6999_/D _7027_/RN _6999_/CLK _6999_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_43_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4350_ hold258/Z _4350_/A2 _4350_/A3 _4352_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_181_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3301_ _6663_/Q _3971_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_4_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4281_ _6564_/I0 _6791_/Q _4288_/S _6791_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6020_ _6933_/Q _5981_/Z _6019_/Z _7045_/Q _6037_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_79_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6922_ _6922_/D _7255_/RN _6922_/CLK _6922_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6853_ _6853_/D _6854_/RN _6853_/CLK _6853_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_168_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5804_ _5804_/I0 hold893/Z _5811_/S _5804_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6784_ _6784_/D _6967_/RN _6784_/CLK _6784_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3996_ _3315_/I _4097_/A1 _6828_/Q _3997_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_22_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5735_ _5888_/I0 hold438/Z _5739_/S _5735_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5666_ hold277/Z _5876_/I0 _5673_/S _5666_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4617_ _5290_/A1 _5146_/A1 _5478_/A1 _4483_/B _4617_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5597_ hold60/Z hold88/Z _5601_/S hold89/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold420 _6758_/Q hold420/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold431 _5522_/Z _6895_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4548_ _5365_/A3 _5281_/C _4652_/A1 _4449_/B _4555_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold442 _6849_/Q hold442/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold453 _5613_/Z _6973_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xclkbuf_4_8_0__1359_ clkbuf_0__1359_/Z _4073__6/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xhold464 _5615_/Z _6975_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_8_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold475 _6928_/Q hold475/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold486 _6969_/Q hold486/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7267_ _7267_/D _7269_/CLK _7267_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4479_ _4786_/A1 _4786_/A2 _4786_/A3 _5094_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xhold497 _6763_/Q hold497/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_77_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6218_ _6790_/Q _5972_/Z _6021_/Z _6840_/Q _6220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_131_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7198_ _7198_/D fanout656/Z _7198_/CLK _7198_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XTAP_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6149_ _6986_/Q _5988_/Z _5996_/Z _7084_/Q _6152_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3850_ _7069_/Q _3943_/A2 _4244_/S input72/Z _4161_/A1 _6709_/Q _3855_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_149_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet952_209 net952_209/I _7016_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3781_ _6974_/Q _3923_/A2 _3957_/A2 _6958_/Q _3956_/A2 _7120_/Q _3786_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5520_ hold222/Z _5520_/A2 _5520_/B _5520_/C hold223/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_118_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5451_ _4492_/Z _4536_/Z _5451_/B _5451_/C _5454_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_172_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4402_ _4580_/C _4489_/A1 _4402_/B _4412_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_99_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5382_ _5379_/Z _5464_/B _5382_/A3 _5382_/A4 _5382_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_7121_ _7121_/D _7179_/RN _7121_/CLK _7121_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4333_ _6612_/I1 hold647/Z _4334_/S _4333_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7052_ _7052_/D _6821_/RN _7052_/CLK _7052_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4264_ hold297/Z _5877_/I0 _4270_/S _4264_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6003_ _6015_/A3 _6164_/A2 _3385_/I _3386_/I _6003_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4195_ _4210_/S _4194_/Z _6652_/A2 _3540_/Z hold33/Z _4211_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_95_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6905_ _6905_/D _7179_/RN _6905_/CLK _6905_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_24_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6836_ _6836_/D _7279_/RN _7279_/CLK _6836_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_126_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6767_ _6767_/D _7193_/RN _6767_/CLK _6767_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3979_ _3978_/Z _3979_/I1 _3988_/S _6661_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5718_ _5775_/I0 hold627/Z _5718_/S _5718_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6698_ _6698_/D _7090_/RN _6698_/CLK _6698_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5649_ hold361/Z _5859_/I0 _5655_/S _5649_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold250 _7059_/Q hold250/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold261 _7063_/Q hold261/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_85_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold272 _5782_/Z _7123_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold283 _6911_/Q hold283/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold294 _4270_/Z _6784_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_120_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout730 _4752_/A2 _3408_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout741 _5051_/S _4456_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_93_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 mask_rev_in[12] input7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4951_ _4407_/Z _5259_/A1 _4759_/Z _5263_/A4 _4951_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3902_ _6889_/Q _3902_/A2 _3960_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_51_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4882_ _4367_/Z _4555_/B _5172_/B _5172_/C _4882_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_178_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6621_ _6644_/A1 _6650_/A2 _6621_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3833_ _3844_/A1 _3578_/Z _3936_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6552_ _6848_/Q _6552_/A2 _6273_/Z _6823_/Q _6553_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_119_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3764_ _6676_/Q _3546_/Z _3776_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_9_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5503_ hold28/Z _5503_/A2 _5647_/A2 _5620_/A4 _5509_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_146_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6483_ _7205_/Q _6540_/A2 _6296_/Z _7165_/Q _7067_/Q _6257_/Z _6486_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3695_ _7106_/Q _5758_/A1 _3719_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xoutput300 _3990_/I serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5434_ _5434_/A1 _5434_/A2 _5432_/Z _5433_/Z _5441_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_10_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput311 _6811_/Q wb_dat_o[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput322 _6812_/Q wb_dat_o[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_105_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput333 _6813_/Q wb_dat_o[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5365_ _5468_/B1 _5288_/B _5365_/A3 _4363_/Z _5365_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_0_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7104_ _7104_/D _7202_/RN _7104_/CLK _7104_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4316_ _6830_/Q _6829_/Q _6831_/Q _4316_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_101_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5296_ _5271_/Z _5296_/A2 _5295_/Z _5467_/B _5296_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_7035_ _7035_/D _7125_/RN _7035_/CLK _7035_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4247_ _4103_/I hold497/Z _4252_/S _4247_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4178_ _6613_/I1 hold951/Z _4178_/S _4178_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6819_ _6819_/D _7278_/RN _7279_/CLK _6819_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout560 _5943_/S _6300_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout571 _7228_/Q _5991_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout582 _4113_/S _4117_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_59_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout593 _3304_/I _3978_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_18_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3480_ _3479_/Z hold387/Z _3500_/S _3480_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_142_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1152_440 net1202_487/I _6725_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_451 net1152_451/I _6714_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5150_ _5374_/A2 _5148_/Z _5374_/A1 _5487_/A1 _5150_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_151_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4101_ _5517_/A2 _5794_/A3 _5517_/A3 _5629_/A3 _4118_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_116_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5081_ _5340_/A1 _5262_/A2 _5343_/A2 _5442_/A4 _5081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_57_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4032_ _4032_/A1 _4032_/A2 _4031_/Z _4035_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_110_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5983_ _3385_/I _5983_/A2 _5983_/B _5983_/C _6010_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_52_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4934_ _5464_/A1 _5325_/B _5061_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_61_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4865_ _4865_/A1 _4865_/A2 _5156_/B _4869_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA_12 hold19/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6604_ _4316_/Z _6604_/A2 _6833_/D _6828_/Q _7278_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3816_ _5776_/A1 _5510_/A2 _3902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_20_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4796_ _4793_/Z _5394_/A2 _5453_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6535_ _6856_/Q _6535_/A2 _6546_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3747_ _3747_/A1 _3747_/A2 _3747_/A3 _3747_/A4 _3747_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6466_ _6466_/A1 _6466_/A2 _6466_/A3 _6465_/Z _6466_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3678_ input31/Z _3927_/C2 _3951_/A2 _7139_/Q _3686_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_12_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5417_ _5417_/A1 _5417_/A2 _5263_/Z _5417_/A4 _5417_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_161_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6397_ _7186_/Q _6532_/A2 _6299_/Z _7056_/Q _6992_/Q _6237_/Z _6401_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xoutput174 _3367_/ZN mgmt_gpio_oeb[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5348_ _5348_/I _5437_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput185 _3357_/ZN mgmt_gpio_oeb[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_130_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput196 _3732_/A1 mgmt_gpio_oeb[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5279_ _5288_/A1 _5279_/A2 _4555_/C _5439_/A1 _5279_/C _5284_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_7018_ _7018_/D _7207_/RN _7018_/CLK _7018_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_101_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet1102_370 net1202_489/I _6840_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1102_381 net1202_481/I _6809_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout390 hold258/I _5875_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet1102_392 net902_179/I _6782_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4650_ _5365_/A3 _5288_/B _4652_/A4 _4652_/A1 _4650_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_159_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput10 mask_rev_in[15] input10/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3601_ _3601_/A1 _3601_/A2 _3601_/A3 _3601_/A4 _3601_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xinput21 mask_rev_in[25] input21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput32 mask_rev_in[6] input32/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4581_ _4557_/Z _5435_/A2 _5349_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xinput43 mgmt_gpio_in[16] input43/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput54 mgmt_gpio_in[26] input54/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6320_ _6320_/A1 _6239_/Z _6321_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_116_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold805 _6674_/Q hold805/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3532_ _3508_/Z hold137/Z _3904_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xinput65 mgmt_gpio_in[36] _7308_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput76 qspi_enabled _4050_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold816 _5807_/Z _7145_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xinput87 spimemio_flash_io1_do _7307_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold827 _6722_/Q hold827/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput98 wb_adr_i[12] input98/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold838 _5837_/Z _7172_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_6_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold849 _6709_/Q hold849/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6251_ _6300_/A2 _6300_/A4 _6300_/A1 _6533_/A2 _6251_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_143_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3463_ _7283_/Q _3462_/Z _3463_/S _7283_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5202_ _4626_/Z _5201_/Z _5202_/A3 _5202_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6182_ _6201_/A3 _6931_/Q _6184_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3394_ _3394_/I _6583_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_5133_ _5165_/A2 _5278_/B _5288_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5064_ _5064_/A1 _5410_/B _5063_/I _5064_/A4 _5066_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4015_ _5957_/S _3990_/I _5953_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_53_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5966_ _6972_/Q _5964_/Z _5965_/Z _6698_/Q _5974_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_12_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4917_ _5328_/A1 _5442_/A1 _5323_/B _5442_/A4 _4927_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_33_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5897_ _3324_/I _3990_/I _5901_/A1 _5950_/A1 _5901_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_178_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4848_ _4853_/A1 _5364_/A1 _5287_/B _3406_/I _5373_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xclkbuf_leaf_114__1359_ clkbuf_4_4_0__1359_/Z net802_83/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_34__1359_ clkbuf_4_11_0__1359_/Z _4073__48/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_148_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_97__1359_ clkbuf_4_5_0__1359_/Z net1052_328/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_148_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4779_ _5478_/B1 _4778_/Z _5456_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_180_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6518_ _6824_/Q _6550_/B1 _6535_/A2 _6855_/Q _6521_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_146_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6449_ _6449_/I _6450_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5820_ _5892_/I0 hold989/Z _5820_/S _5820_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5751_ _5751_/I0 hold979/Z _5757_/S _5751_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4702_ _4884_/A1 _3401_/I _5255_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5682_ hold803/Z _5811_/I0 _5682_/S _5682_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4633_ _4633_/A1 _5035_/A4 _5387_/B _4636_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_147_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4564_ _5290_/A2 _4643_/A4 _5439_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_156_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold602 _5757_/Z _7101_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold613 _6991_/Q hold613/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6303_ _7214_/Q _6543_/A2 _6302_/Z _7086_/Q _6306_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold624 _4157_/Z _6705_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold635 _6712_/Q hold635/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3515_ _3653_/A1 _3492_/Z _3680_/A3 hold211/Z _3515_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7283_ _7283_/D _6637_/Z _7302_/CLK _7283_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold646 _5565_/Z _6931_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4495_ _5458_/A4 _4884_/A1 _4495_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
Xhold657 _6692_/Q hold657/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold668 _4331_/Z _6838_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold679 _7212_/Q hold679/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_131_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6234_ _7233_/Q _7232_/Q _6299_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3446_ _3449_/A2 _3450_/A1 _3447_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_98_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6165_ _7019_/Q _5971_/Z _6005_/Z _7043_/Q _6169_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3377_ _6943_/Q _3377_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5116_ _5117_/A1 _5117_/A2 _5316_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6096_ _7146_/Q _5987_/Z _6003_/Z hold78/I _6097_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5047_ _5047_/A1 _5360_/B _5049_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6998_ _6998_/D _7247_/RN _6998_/CLK _6998_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_41_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5949_ _6282_/A1 _6544_/A2 _5950_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_40_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_80__1359_ clkbuf_4_7_0__1359_/Z net902_184/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_172_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3300_ _6664_/Q _3465_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_4280_ _6831_/Q _6563_/A2 _4288_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_98_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6921_ _6921_/D _7179_/RN _6921_/CLK _6921_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6852_ _6852_/D _6907_/RN _6852_/CLK _6852_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5803_ _3523_/Z _5839_/A2 _5866_/A3 _5811_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_90_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6783_ _6783_/D _6854_/RN _6783_/CLK _6783_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_167_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3995_ _3994_/Z _3995_/A2 _4097_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_22_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5734_ _5842_/I0 hold84/Z _5739_/S hold85/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5665_ _5665_/A1 _5674_/A2 _5673_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_4616_ _5290_/A1 _5373_/A2 _5478_/A1 _4483_/B _4616_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_163_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5596_ _5833_/I0 hold705/Z _5601_/S _5596_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold410 _6738_/Q hold410/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold421 _4237_/Z _6758_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4547_ _5278_/C _4878_/A2 _5426_/A1 _4547_/A4 _4547_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold432 _7104_/Q hold432/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold443 _4348_/Z _6849_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_150_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold454 _7182_/Q hold454/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold465 _6690_/Q hold465/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7266_ _7266_/D _7269_/CLK _7266_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold476 _5562_/Z _6928_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4478_ _4786_/A2 _4786_/A3 _4782_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold487 _5608_/Z _6969_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold498 _4247_/Z _6763_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6217_ _6217_/A1 _6217_/A2 _6217_/A3 _6217_/A4 _6217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_132_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3429_ _3971_/A1 _6730_/Q _3441_/C _6664_/Q _3430_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_58_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7197_ _7197_/D _7221_/RN _7197_/CLK _7197_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6148_ _6970_/Q _5979_/Z _5999_/Z _7034_/Q _6152_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6079_ _7129_/Q _6000_/Z _6019_/Z _7047_/Q _6967_/Q _5979_/Z _6085_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_2604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3780_ _7208_/Q _3960_/A2 _3955_/A2 _7200_/Q _3796_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_13_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5450_ _5450_/I _5463_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4401_ _4412_/A1 _4399_/Z _5083_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
X_5381_ _5381_/I _5382_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_160_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7120_ _7120_/D _6967_/RN _7120_/CLK _7120_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_125_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4332_ _4332_/A1 _5629_/A3 _5517_/A3 _5794_/A3 _4334_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_141_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7051_ _7051_/D _7125_/RN _7051_/CLK _7051_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_99_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4263_ hold173/Z _4103_/I _4270_/S _4263_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6002_ _7231_/Q _6002_/A2 _6002_/A3 _5914_/S _6002_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_140_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4194_ _4194_/A1 _3994_/Z _4194_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_39_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6904_ _6904_/D _7179_/RN _6904_/CLK _6904_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6835_ _6835_/D _7279_/RN _7279_/CLK _6835_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_165_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6766_ _6766_/D _6894_/RN _6766_/CLK _6766_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3978_ _3977_/Z _6660_/Q _3978_/S _3978_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5717_ _5855_/I0 hold673/Z _5718_/S _5717_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6697_ _6697_/D _6850_/RN _6697_/CLK _6697_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xclkbuf_2_1__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _4072_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5648_ hold575/Z _5804_/I0 _5648_/S _5648_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5579_ hold473/Z _5798_/I0 _5583_/S _5579_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold240 _7097_/Q hold240/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_105_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold251 _5709_/Z _7059_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold262 _5714_/Z _7063_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold273 _6996_/Q hold273/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_46_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold284 _5543_/Z _6911_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_172_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7249_ _7249_/D _7259_/RN _7260_/CLK _7249_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_131_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold295 _6736_/Q hold295/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xfanout720 input160/Z _6563_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_120_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout731 _5322_/A1 _4752_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout742 input117/Z _5051_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_131_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput8 mask_rev_in[13] input8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_188_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4950_ _5248_/A3 _4982_/A2 _4496_/Z _4958_/A4 _5252_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_91_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3901_ _6980_/Q _3901_/A2 _3926_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_33_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4881_ _5104_/A1 _4555_/B _4650_/Z _5172_/C _4881_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_2990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6620_ _6644_/A1 _6648_/A2 _6620_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3832_ _3519_/Z _3844_/A1 _4359_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6551_ _6790_/Q _6551_/A2 _6288_/Z _7297_/Q _6553_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_158_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3763_ input54/Z _4194_/A1 _3795_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5502_ _5502_/I0 hold20/Z hold29/Z hold30/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6482_ _7075_/Q _6248_/Z _6253_/Z _7141_/Q _7157_/Q _6293_/Z _6486_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3694_ _7064_/Q _3927_/B1 _3715_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5433_ _5433_/A1 _5433_/A2 _5433_/A3 _4662_/B _5433_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xoutput301 _3683_/Z serial_data_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput312 _6803_/Q wb_dat_o[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput323 _6795_/Q wb_dat_o[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput334 _7268_/Q wb_dat_o[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5364_ _5364_/A1 _5373_/A2 _5364_/B _5468_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_160_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7103_ _7103_/D _6856_/RN _7103_/CLK _7103_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_99_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4315_ _3315_/I _6600_/B2 _6597_/C1 _6832_/Q _5299_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_113_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5295_ _5295_/A1 _5295_/A2 _5295_/A3 _5315_/A1 _5295_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_87_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7034_ _7034_/D _7034_/RN _7034_/CLK _7034_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_141_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4246_ hold258/Z _5517_/A1 hold146/Z _5520_/C _4252_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4177_ _6612_/I1 hold911/Z _4178_/S _4177_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6818_ _6818_/D _7262_/CLK _6818_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6749_ _6749_/D _7122_/RN _6749_/CLK _6749_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_177_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout550 hold64/Z _5876_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout561 _7236_/Q _5946_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout572 _5914_/S _3387_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout583 hold1076/Z _4113_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_58_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout594 _6733_/Q _3304_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_101_892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1152_430 net1152_430/I _6740_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_441 net1152_441/I _6724_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4100_ hold8/Z hold31/Z _4117_/S hold32/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5080_ _4977_/Z _4981_/Z _5080_/B _5080_/C _5412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_1_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4031_ _4031_/A1 _4031_/A2 _4031_/A3 _4031_/A4 _4031_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_96_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5982_ _6964_/Q _5979_/Z _5981_/Z _6932_/Q _5980_/Z _7068_/Q _5983_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_18_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4933_ _4933_/A1 _4930_/Z _4933_/A3 _4933_/A4 _4939_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_52_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4864_ _4624_/Z _4844_/Z _5156_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_13 _7283_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3815_ _5821_/A2 _3617_/Z _4188_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6603_ _5299_/C _6833_/Q _6826_/Q _6603_/A4 _6604_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_119_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4795_ _5328_/A1 _5403_/A1 _5394_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6534_ _6727_/Q _6253_/Z _6296_/Z _6715_/Q _6542_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_158_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3746_ _7185_/Q _3959_/C1 _3901_/A2 _6983_/Q _3747_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_146_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6465_ _6465_/A1 _6465_/A2 _6465_/A3 _6464_/Z _6465_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3677_ input49/Z _4210_/S _5521_/A2 _3904_/A2 _3947_/A2 _7099_/Q _3687_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5416_ _5416_/I _5417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6396_ _7064_/Q _6257_/Z _6408_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_161_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5347_ _5347_/A1 _5347_/A2 _5347_/A3 _5347_/A4 _5348_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_99_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput175 _3366_/ZN mgmt_gpio_oeb[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput186 _3356_/ZN mgmt_gpio_oeb[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_130_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput197 _3346_/ZN mgmt_gpio_oeb[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5278_ _5290_/A2 _5287_/A2 _5278_/B _5278_/C _5279_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_101_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7017_ _7017_/D _7258_/RN _7017_/CLK _7017_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_130_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4229_ _4244_/S _4194_/Z _4060_/S _5830_/A1 hold33/Z _4245_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_75_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_137__1359_ net1152_446/I net852_149/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_68_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_57__1359_ clkbuf_4_15_0__1359_/Z net1152_434/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_55_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1102_360 net802_63/I _6850_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout380 _5821_/A3 _5517_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xnet1102_371 net1202_485/I _6839_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet1102_382 net1102_382/I _6800_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout391 hold257/Z hold258/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_19_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1102_393 net952_225/I _6781_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_188_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3600_ _7181_/Q _3945_/A2 _3945_/B1 _7093_/Q _3601_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xinput11 mask_rev_in[16] input11/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput22 mask_rev_in[26] input22/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4580_ _4604_/A2 _4604_/A3 _4580_/B _4580_/C _5435_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xinput33 mask_rev_in[7] input33/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput44 mgmt_gpio_in[17] input44/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3531_ _3505_/Z _5692_/A1 _3934_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_122_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput55 mgmt_gpio_in[27] input55/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput66 mgmt_gpio_in[37] _7309_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput77 ser_tx input77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold806 _4120_/Z _6674_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold817 _7129_/Q hold817/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold828 _4183_/Z _6722_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xinput88 spimemio_flash_io1_oeb input88/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold839 _6848_/Q hold839/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6250_ _5946_/S _6484_/A2 _6311_/A3 _6302_/A4 _6250_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_155_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput99 wb_adr_i[13] input99/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3462_ _3465_/A3 _3441_/C _4056_/I1 _3462_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_171_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5201_ _5201_/A1 _5438_/C _4557_/Z _4604_/Z _5201_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_170_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6181_ _6169_/Z _6181_/A2 _6181_/A3 _6180_/Z _6181_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_171_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3393_ _3393_/I _6580_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_130_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5132_ _5205_/A1 _5132_/A2 _5293_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_97_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5063_ _5063_/I _5330_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4014_ _7237_/Q _6484_/A2 _6311_/A3 _6285_/A2 _4014_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_26_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5965_ _6068_/A2 _5991_/A2 _5914_/S _6210_/C _5965_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_40_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4916_ _5324_/A1 _5263_/A4 _5056_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5896_ _5896_/I0 _5951_/B _5957_/S _5910_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4847_ _4530_/I _5399_/A2 _5104_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4778_ _4468_/Z _4782_/A1 _5307_/A3 _4778_/A4 _4778_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_120_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6517_ _6706_/Q _6254_/Z _6273_/Z _6822_/Q _6521_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3729_ _7201_/Q _3955_/A2 _3747_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_119_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6448_ _3324_/I _7255_/Q _6448_/B _6449_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_106_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6379_ _7137_/Q _6253_/Z _6297_/Z _6701_/Q _6380_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_88_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_40__1359_ _4073__46/I net802_53/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_120__1359_ net952_221/I net902_197/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_19_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5750_ _5822_/I0 hold971/Z _5757_/S _5750_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4701_ _4687_/Z _5097_/A1 _5403_/A1 _5092_/A1 _5459_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_176_924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5681_ hold763/Z _5681_/I1 _5682_/S _5681_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4632_ _5365_/A3 _4449_/B _3407_/I _4652_/A1 _5293_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_116_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4563_ _4402_/B _4395_/B _4026_/B _4026_/C _4563_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold603 _7021_/Q hold603/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_128_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3514_ _6979_/Q _3923_/A2 _3592_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_116_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6302_ _5946_/S _6311_/A3 _6302_/A3 _6302_/A4 _6302_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold614 _5633_/Z _6991_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold625 _7048_/Q hold625/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7282_ _7282_/D _6636_/Z _7304_/CLK _7282_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold636 _4168_/Z _6712_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4494_ _4652_/A4 _4884_/A1 _4494_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
Xhold647 _6839_/Q hold647/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_6_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold658 _4141_/Z _6692_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6233_ _5946_/S _7237_/Q _6233_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold669 _6837_/Q hold669/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3445_ _3452_/S _7291_/Q _3450_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6164_ _7027_/Q _6164_/A2 _6164_/B1 _6995_/Q _6176_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3376_ _6951_/Q _3376_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ _5113_/Z _5403_/C _5233_/A1 _5156_/B _5115_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6095_ _6968_/Q _5979_/Z _5996_/Z _7082_/Q _6095_/C _6101_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_97_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5046_ _5044_/Z _5433_/A1 _5047_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_85_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6997_ _6997_/D _7141_/RN _6997_/CLK _6997_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_53_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5948_ _7235_/Q _3329_/I _6300_/A2 _6484_/A3 _5948_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_159_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5879_ _5879_/I0 hold444/Z _5883_/S _5879_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6920_ _6920_/D _7255_/RN _6920_/CLK _6920_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6851_ _6851_/D _7297_/RN _6851_/CLK _6851_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_90_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5802_ hold6/Z _7141_/Q hold12/Z hold13/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6782_ _6782_/D _7247_/RN _6782_/CLK _6782_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3994_ _3994_/A1 _6902_/Q input67/Z _3994_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_50_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5733_ _5859_/I0 _5733_/I1 _5739_/S _5733_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5664_ hold869/Z _5784_/I0 _5664_/S _5664_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4615_ _5290_/A1 _5438_/A1 _5290_/A3 _4483_/B _5151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5595_ _5859_/I0 hold985/Z _5601_/S _5595_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold400 _6702_/Q hold400/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_117_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4546_ _4835_/A2 _3403_/I _3402_/I _5129_/A4 _4546_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold411 _4203_/Z _6738_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold422 _7037_/Q hold422/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_172_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold433 _5761_/Z _7104_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold444 _7209_/Q hold444/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold455 _5849_/Z _7182_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold466 _4138_/Z _6690_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7265_ _7265_/D _7269_/CLK _7265_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4477_ _4692_/B _4692_/C _4786_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold477 _6691_/Q hold477/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold488 _6740_/Q hold488/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6216_ _6723_/Q _5987_/Z _6015_/Z _6842_/Q _6217_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold499 _6760_/Q hold499/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_132_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3428_ _3427_/Z _6734_/Q _3428_/A3 _3428_/B _7301_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_7196_ _7196_/D _7221_/RN _7196_/CLK _7196_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_48_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6147_ _6147_/A1 _6147_/A2 _6147_/A3 _6147_/A4 _6147_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3359_ _7081_/Q _3359_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6078_ _6078_/A1 _6078_/A2 _6078_/A3 _6078_/A4 _6078_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_73_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5029_ _5353_/A1 _5439_/B2 _5029_/B _5354_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_2605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4400_ _4412_/A1 _4399_/Z _4491_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5380_ _4568_/Z _4892_/B _4821_/Z _5380_/B2 _5380_/C _5381_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_154_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4331_ _5796_/I0 hold667/Z _4331_/S _4331_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7050_ _7050_/D _7125_/RN _7050_/CLK _7050_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4262_ _4225_/S _3994_/Z hold33/Z _4270_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_141_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6001_ _7028_/Q _5999_/Z _6000_/Z _7126_/Q _6008_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_68_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4193_ hold639/Z _4361_/I1 _4193_/S _4193_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6903_ _6903_/D _7179_/RN _6903_/CLK _6903_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_39_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6834_ _6834_/D _7261_/RN _7279_/CLK _6834_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_39_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6765_ hold91/Z _7193_/RN _6765_/CLK hold90/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3977_ _6661_/Q _3973_/Z _3977_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5716_ _5782_/I0 hold923/Z _5718_/S _5716_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6696_ _6696_/D _6850_/RN _6696_/CLK _6696_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5647_ hold153/Z _5647_/A2 hold28/Z hold137/Z _5648_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_136_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5578_ hold398/Z _5797_/I0 _5583_/S _5578_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold230 _7195_/Q hold230/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold241 _5753_/Z _7097_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_117_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold252 _7023_/Q hold252/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4529_ _5420_/A2 _5097_/B2 _4672_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_160_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold263 _7122_/Q hold263/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold274 _5639_/Z _6996_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold285 _7109_/Q hold285/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7248_ _7248_/D _7259_/RN _7260_/CLK _7248_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_132_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold296 _4199_/Z _6736_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_132_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout710 _7224_/RN _6771_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout721 input124/Z _3406_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_59_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout732 _5458_/A4 _4460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_172_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout743 input108/Z _4402_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7179_ _7179_/D _7179_/RN _7179_/CLK _7179_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_59_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput9 mask_rev_in[14] input9/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3900_ _6728_/Q _4191_/A1 _3919_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_91_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4880_ _4880_/A1 _4877_/Z _4879_/Z _5167_/B _4880_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_2980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3831_ _4185_/A2 _3578_/Z _6611_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_189_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3762_ _3761_/Z _3762_/I1 _3899_/S _6871_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6550_ _6854_/Q _6550_/A2 _6550_/B1 _6825_/Q _6550_/C1 _6800_/Q _6553_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_118_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5501_ hold269/Z _5834_/I0 hold29/Z _5501_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3693_ _7000_/Q _5638_/A1 _3724_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6481_ _7213_/Q _6535_/A2 _6545_/A2 _6939_/Q _6493_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_145_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5432_ _5432_/A1 _5189_/Z _5209_/Z _4985_/Z _5432_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xoutput302 _3619_/Z serial_data_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput313 _6804_/Q wb_dat_o[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_127_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput324 _6796_/Q wb_dat_o[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5363_ _5363_/A1 _5342_/I _5363_/B1 _5396_/A1 _5383_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
Xoutput335 _7269_/Q wb_dat_o[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7102_ _7102_/D _6786_/RN _7102_/CLK _7102_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_141_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4314_ _6601_/A2 _6832_/Q _6577_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5294_ _5294_/A1 _5366_/A2 _5296_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_114_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7033_ _7033_/D _7259_/RN _7033_/CLK _7033_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4245_ _4244_/Z hold493/Z _4245_/S _4245_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4176_ _4350_/A2 _5821_/A2 _4350_/A3 _4178_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_82_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6817_ _6817_/D _7262_/CLK _6817_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6748_ _6748_/D _6967_/RN _6748_/CLK _6748_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_52_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_17__1359_ net1152_430/I _4073__35/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_137_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6679_ hold67/Z _6839_/RN _6679_/CLK hold66/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_176_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout540 _4360_/I1 _5537_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout551 hold63/Z hold64/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout562 _7235_/Q _3328_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout573 _5914_/S _6021_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_101_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout584 _6746_/Q _5951_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_47_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout595 _6665_/Q _3441_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_18_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1152_420 net902_199/I _6754_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet1152_431 net1152_431/I _6739_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_442 net852_149/I _6723_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_155_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4030_ _4386_/A3 _4386_/A4 _4391_/A1 _4391_/A2 _4030_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_49_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5981_ _6210_/C _6021_/A2 _6210_/A2 _3387_/I _5981_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_92_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4932_ _5258_/B2 _5442_/A1 _5323_/B _5248_/A2 _4933_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_33_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4863_ _4624_/Z _4833_/Z _4865_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_60_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_14 input75/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_6602_ _6602_/I0 _7277_/Q _6602_/S _7277_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3814_ _6729_/Q _4191_/A1 _3876_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4794_ _4673_/Z _4793_/Z _5452_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6533_ _6838_/Q _6533_/A2 _6533_/A3 _6533_/A4 _6540_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3745_ _7209_/Q _3960_/A2 _5665_/A1 _7023_/Q _3747_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_158_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6464_ _6464_/A1 _6464_/A2 _6464_/A3 _6464_/A4 _6464_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3676_ hold44/I _3917_/A2 _5683_/A1 _7041_/Q _3687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5415_ _5415_/A1 _4982_/Z _5415_/B1 _5083_/C _5416_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_6395_ _7254_/Q _6395_/I1 _6450_/S _7254_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5346_ _5393_/A2 _5346_/A2 _5346_/B _5347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_115_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput176 _3365_/ZN mgmt_gpio_oeb[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_87_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput187 _3355_/ZN mgmt_gpio_oeb[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput198 _3345_/ZN mgmt_gpio_oeb[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5277_ _5277_/I _5421_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7016_ _7016_/D _7140_/RN _7016_/CLK _7016_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4228_ _4227_/Z hold311/Z _4228_/S _4228_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4159_ _5822_/I0 hold621/Z _4160_/S _4159_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_4__1359_ net1152_451/I net802_55/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout370 _3535_/Z _4350_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet1102_361 net1202_468/I _6849_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1102_372 net802_90/I _6838_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout381 _3511_/ZN _5821_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xnet1102_383 net852_106/I _6799_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout392 _6282_/Z _6532_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xnet1102_394 net1102_394/I _6780_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 mask_rev_in[17] input12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput23 mask_rev_in[27] input23/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput34 mask_rev_in[8] input34/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput45 mgmt_gpio_in[18] input45/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3530_ _3507_/Z _3844_/A1 _5656_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xinput56 mgmt_gpio_in[28] input56/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput67 mgmt_gpio_in[3] input67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xhold807 _7033_/Q hold807/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xinput78 spi_csb input78/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput89 spimemio_flash_io2_do input89/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold818 _5789_/Z _7129_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_183_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold829 _7163_/Q hold829/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xclkbuf_leaf_63__1359_ clkbuf_4_13_0__1359_/Z net902_194/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_116_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3461_ _3441_/C _6663_/Q _6730_/Q _3463_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xclkbuf_leaf_143__1359_ net1152_451/I net1202_490/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_170_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5200_ _5205_/A1 _5291_/B _5200_/B1 _5346_/A2 _5200_/C _5354_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3392_ _6891_/Q _3903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6180_ _6180_/A1 _6180_/A2 _6180_/A3 _6180_/A4 _6180_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_130_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5131_ _5172_/A1 _5291_/A2 _5165_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_69_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5062_ _5403_/A1 _5330_/B2 _5062_/B _5063_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_42_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4013_ _5942_/S _3328_/I _6311_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_38_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5964_ _6117_/A4 _6014_/A2 _6139_/A2 _3389_/I _5964_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_52_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4915_ _4496_/Z _4982_/A2 _5263_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5895_ _5951_/B _3324_/I _5901_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_166_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4846_ _4846_/A1 _4846_/A2 _5090_/A2 _4849_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_178_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ _4782_/A1 _5099_/A1 _5456_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6516_ _6512_/Z _6516_/A2 _6516_/A3 _6516_/A4 _6516_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3728_ input46/Z _4210_/S _3739_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_146_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6447_ _6440_/Z _6446_/Z _6447_/B1 _6286_/Z _6529_/S _6448_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3659_ _7091_/Q _3945_/B1 _3927_/B1 _7065_/Q _3663_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_161_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6378_ _7071_/Q _6248_/Z _6293_/Z _7153_/Q _6380_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_103_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5329_ _5359_/A1 _5329_/A2 _5445_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_185_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4700_ _5420_/A2 _5129_/A3 _3404_/I _5129_/A4 _4700_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_1191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5680_ hold807/Z _5881_/I0 _5682_/S _5680_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4631_ _4868_/A1 _5399_/A1 _5403_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_8_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4562_ _5290_/A1 _4483_/B _5291_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_129_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold604 _5667_/Z _7021_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6301_ _7052_/Q _6299_/Z _6300_/Z _7102_/Q _6306_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold615 _6844_/Q hold615/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3513_ _5611_/A1 _3512_/Z _3923_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold626 _5697_/Z _7048_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7281_ _7281_/D _6635_/Z _7302_/CLK _7281_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
XFILLER_183_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4493_ _4808_/A2 _4492_/Z _5240_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_171_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold637 _6967_/Q hold637/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold648 _4333_/Z _6839_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6232_ _7250_/Q _6232_/I1 _6558_/S _7250_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold659 _6976_/Q hold659/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_170_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3444_ _3442_/B _3452_/S _3449_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_98_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3375_ hold88/I _3375_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6163_ _7125_/Q _5969_/Z _6176_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _4762_/Z _4867_/Z _5403_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6094_ _6094_/I _6095_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5045_ _5214_/A2 _5389_/A1 _5172_/B _5045_/C _5433_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_84_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6996_ _6996_/D _7155_/RN _6996_/CLK _6996_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_5947_ _6285_/A2 _7237_/Q _5947_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_22_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5878_ hold2/Z _7208_/Q _5883_/S _5878_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4829_ _4673_/Z _5287_/A2 _5276_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_166_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_13_0__1359_ clkbuf_0__1359_/Z clkbuf_4_13_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_71_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold1 hold1/I hold1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_66_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6850_ _6850_/D _6850_/RN _6850_/CLK _6850_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5801_ hold16/Z _7140_/Q hold12/Z hold17/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6781_ _6781_/D _7260_/RN _6781_/CLK _6781_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3993_ _3994_/A1 hold469/Z input67/Z _4064_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5732_ _5732_/I0 hold919/Z _5739_/S _5732_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5663_ hold891/Z _5837_/I0 _5664_/S _5663_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4614_ _5365_/A3 _4944_/A1 _4460_/B _3406_/I _4614_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_163_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5594_ _5804_/I0 hold963/Z _5601_/S _5594_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold401 _4154_/Z _6702_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4545_ _5269_/A1 _4878_/A2 _5172_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold412 _7016_/Q hold412/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold423 _5685_/Z _7037_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold434 _6668_/Q hold434/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold445 _5879_/Z _7209_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_172_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7264_ _7264_/D _7269_/CLK _7264_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold456 _7206_/Q hold456/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4476_ _4853_/A1 _4481_/A2 _5288_/B _4692_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xhold467 _6926_/Q hold467/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold478 _4139_/Z _6691_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6215_ _6713_/Q _6002_/Z _6003_/Z _6715_/Q _6217_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold489 _4207_/Z _6740_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3427_ _3304_/I _6732_/Q _6730_/Q _3427_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_7195_ _7195_/D _7219_/RN _7195_/CLK _7195_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_131_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6146_ _7124_/Q _5969_/Z _6146_/B _6147_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3358_ _7089_/Q _3358_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6077_ _7055_/Q _5924_/Z _5988_/Z _6983_/Q _6118_/B _6078_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_72_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5028_ _5023_/Z _5476_/A1 _5027_/I _5028_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_85_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6979_ _6979_/D _7124_/RN _6979_/CLK _6979_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_110_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold990 _5820_/Z _7157_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_0_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4330_ _5795_/I0 hold669/Z _4331_/S _4330_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4261_ _5547_/I0 hold265/Z _4261_/S _4261_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6000_ _6015_/A3 _6164_/B1 _3385_/I _3386_/I _6000_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_119_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4192_ hold546/Z _4360_/I1 _4193_/S _4192_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6902_ _6902_/D _7194_/RN _6902_/CLK _6902_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_36_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6833_ _6833_/D _7261_/RN _7279_/CLK _6833_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6764_ _6764_/D _6854_/RN _6764_/CLK _6764_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3976_ _3975_/Z _6662_/Q _3988_/S _6662_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5715_ _5871_/I0 hold406/Z _5718_/S _5715_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6695_ _6695_/D _6886_/RN _6695_/CLK _6695_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5646_ hold813/Z _5784_/I0 _5646_/S _5646_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5577_ hold931/Z _5796_/I0 _5583_/S _5577_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold220 _3488_/Z _3489_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold231 _5863_/Z _7195_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4528_ _5020_/A2 _4524_/Z _4549_/A4 _4501_/B _4528_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold242 _7161_/Q hold242/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold253 _5669_/Z _7023_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold264 _5781_/Z _7122_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_6_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7247_ _7247_/D _7247_/RN _7258_/CLK _7247_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold275 _6915_/Q hold275/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_49_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4459_ _4555_/B _5270_/A1 _4652_/A4 _4459_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
Xfanout700 _7253_/RN _7257_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xhold286 _5766_/Z _7109_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold297 _6778_/Q hold297/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xfanout711 _6650_/A1 _7224_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout722 input124/Z _5295_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout733 _5458_/A4 _3407_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7178_ _7178_/D _7215_/RN _7178_/CLK _7178_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout744 input108/Z _4428_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6129_ _6977_/Q _5964_/Z _6014_/Z _6961_/Q _6000_/Z _7131_/Q _6134_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3830_ _4353_/A1 _3540_/Z _3942_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_38_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3761_ _6567_/I0 _6870_/Q _3898_/S _3761_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5500_ hold76/Z _5842_/I0 hold29/Z hold77/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6480_ _7221_/Q _6543_/A2 _6285_/Z _7197_/Q _7181_/Q _6254_/Z _6493_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3692_ _3505_/Z _3527_/Z _3916_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_146_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5431_ _5431_/A1 _5299_/C _5431_/B _5431_/C _6863_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_127_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput303 _4070_/Z serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput314 _6805_/Q wb_dat_o[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5362_ _5362_/A1 _5362_/A2 _5362_/A3 _5363_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xoutput325 _6797_/Q wb_dat_o[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput336 _6814_/Q wb_dat_o[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_154_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7101_ _7101_/D _7220_/RN _7101_/CLK _7101_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4313_ _6600_/A1 _3316_/I _3317_/I _4313_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_142_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5293_ _5293_/A1 _5295_/A1 _5293_/B _5366_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_7032_ _7032_/D _7259_/RN _7032_/CLK _7032_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4244_ _6923_/Q _5547_/I0 _4244_/S _4244_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4175_ _4361_/I1 hold492/Z _4175_/S _6717_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6816_ _6816_/D _7262_/CLK _6816_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6747_ _6747_/D _6854_/RN _6747_/CLK _6747_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3959_ _7012_/Q _5656_/A1 _3959_/B1 _6666_/Q _3959_/C1 _7182_/Q _3961_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_149_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6678_ hold21/Z _6894_/RN _6678_/CLK _6678_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_109_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5629_ _5629_/A1 _5794_/A3 _5629_/A3 _5785_/A3 _5637_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_136_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout530 _5850_/I0 _5778_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout541 _4180_/I0 _4360_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_120_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout552 _5647_/A2 _6611_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout563 _3329_/I _6300_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_59_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout574 _7227_/Q _5914_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout585 _6745_/Q _5957_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout596 _4873_/A3 _5287_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_47_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_1_0__1359_ clkbuf_0__1359_/Z net1152_446/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_1521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1152_410 net1152_410/I _6764_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_157_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1152_421 net1152_421/I _6753_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet1152_432 net1152_434/I _6738_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_443 net852_149/I _6722_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5980_ _6015_/A3 _6210_/C _3385_/I _3386_/I _5980_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xclkbuf_leaf_103__1359_ clkbuf_4_5_0__1359_/Z net952_229/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_24_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_23__1359_ _4073__49/I _4073__51/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4931_ _5389_/A2 _5442_/A1 _5323_/B _5248_/A2 _4933_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xclkbuf_leaf_86__1359_ clkbuf_4_13_0__1359_/Z net952_251/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4862_ _4862_/A1 _4859_/Z _4861_/Z _4819_/Z _4865_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_36_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6601_ _6601_/A1 _6601_/A2 _6601_/B _6602_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_3813_ _5821_/A2 _3680_/Z _4191_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_177_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_15 hold541/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4793_ _4534_/Z _5312_/A1 _4491_/B _4402_/B _4793_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6532_ _6697_/Q _6532_/A2 _6542_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3744_ hold88/I _3957_/A2 _3927_/A2 _6701_/Q _3747_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6463_ _6938_/Q _6545_/A2 _6545_/B1 _7018_/Q _6464_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3675_ _7179_/Q _3945_/A2 _5758_/A1 _7107_/Q _3687_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_137_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5414_ _4997_/B _5414_/A2 _4659_/Z _5414_/B _5418_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_174_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6394_ _6394_/I _6395_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5345_ _5389_/C _5345_/A2 _5356_/B _5389_/A2 _5346_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_99_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput177 _3364_/ZN mgmt_gpio_oeb[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput188 _3354_/ZN mgmt_gpio_oeb[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_142_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5276_ _5276_/A1 _5276_/A2 _5276_/B _5276_/C _5277_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xoutput199 _4052_/ZN mgmt_gpio_oeb[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7015_ _7015_/D _7024_/RN _7015_/CLK _7015_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4227_ hold293/Z _5811_/I0 _4227_/S _4227_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4158_ _5821_/A1 _5839_/A2 _4347_/A3 _5629_/A3 _4160_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4089_ _6907_/Q input39/Z _4089_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_37_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout360 _5315_/A4 _4774_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xnet1102_362 net1102_382/I _6848_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout371 _3533_/Z _5517_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_87_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout382 _5629_/A1 _4332_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet1102_373 net802_90/I _6837_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout393 _6275_/Z _6536_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_19_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1102_384 net852_106/I _6790_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1102_395 net1152_425/I _6779_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput13 mask_rev_in[18] input13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput24 mask_rev_in[28] input24/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput35 mask_rev_in[9] input35/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput46 mgmt_gpio_in[19] input46/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput57 mgmt_gpio_in[29] input57/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput68 mgmt_gpio_in[5] input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_156_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold808 _5680_/Z _7033_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xinput79 spi_enabled _4055_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_6_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold819 _7071_/Q hold819/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_171_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3460_ hold52/Z _4056_/I1 _3460_/S _7284_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3391_ _7222_/Q _5894_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5130_ _5240_/B _5328_/A2 _5130_/B1 _5130_/B2 _5321_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_97_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5061_ _5403_/A1 _4936_/I _5061_/B _5410_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_96_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4012_ _6302_/A4 _5946_/S _6282_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_111_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5963_ _6021_/A2 _3387_/I _6117_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_80_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4914_ _4497_/Z _4494_/Z _5442_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5894_ _5894_/A1 _5894_/A2 _5894_/A3 _4019_/B _5951_/B _7222_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_4845_ _4596_/Z _5142_/A3 _5090_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_179_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4776_ _5401_/A2 _5236_/B _5121_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_148_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6515_ _6845_/Q _6549_/A2 _6237_/Z _6837_/Q _6516_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3727_ _3726_/Z _6872_/Q _3899_/S _6872_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6446_ _6554_/A1 _6446_/A2 _6446_/A3 _6446_/A4 _6446_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_161_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3658_ _7147_/Q _3951_/C1 _3924_/A2 _6969_/Q input25/Z _3954_/B1 _3688_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_106_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6377_ _7201_/Q _6272_/Z _6282_/Z _7185_/Q _6296_/Z _7161_/Q _6384_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_162_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3589_ _3589_/A1 _3589_/A2 _3589_/A3 _3589_/A4 _3589_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5328_ _5328_/A1 _5328_/A2 _5481_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_76_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5259_ _5259_/A1 _5259_/A2 _5337_/A2 _5449_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_29_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4630_ _4367_/Z _4555_/B _5291_/C _5387_/A1 _5387_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_175_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4561_ _4556_/Z _4561_/A2 _5003_/A2 _4561_/B _4584_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_156_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6300_ _6300_/A1 _6300_/A2 _6484_/A3 _6300_/A4 _6300_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_144_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3512_ _3653_/A1 hold144/I hold211/I _3492_/Z _3512_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_155_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold605 _7093_/Q hold605/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7280_ _7280_/D _6634_/Z _7302_/CLK hold8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
Xhold616 _4340_/Z _6844_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4492_ _4402_/B _4026_/B _4026_/C _5312_/A1 _4492_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_171_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold627 _7067_/Q hold627/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold638 _5606_/Z _6967_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6231_ _6231_/I _6232_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold649 _6713_/Q hold649/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3443_ _3438_/S _3440_/S _3443_/A3 _3443_/A4 _3452_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_144_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6162_ _7247_/Q _6162_/I1 _6450_/S _7247_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3374_ _6967_/Q _3374_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5113_ _5113_/A1 _5113_/A2 _5313_/A1 _5313_/A3 _5113_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ _7000_/Q _6021_/Z _6090_/Z _5924_/Z _6094_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5044_ _5044_/A1 _5386_/A1 _5044_/A3 _5432_/A1 _5044_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_66_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6995_ _6995_/D _7253_/RN _6995_/CLK _6995_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_53_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5946_ _5950_/B1 _5945_/B _5946_/S _7236_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5877_ _5877_/I0 hold721/Z _5883_/S _5877_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4828_ _5287_/B _5367_/A2 _5164_/A4 _4598_/Z _5364_/A1 _5421_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_138_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4759_ _4501_/B _4759_/A2 _4759_/A3 _4759_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_181_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6429_ _7139_/Q _6253_/Z _6296_/Z _7163_/Q _6434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_108_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold2 hold2/I hold2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_181_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5800_ _5818_/I0 hold600/Z hold12/Z _7139_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6780_ _6780_/D _7002_/RN _6780_/CLK _6780_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_90_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3992_ _7298_/Q hold8/I _3995_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5731_ _3523_/Z _5731_/A2 _5866_/A3 _5739_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_95_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5662_ hold811/Z _5827_/I0 _5664_/S _5662_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4613_ _5288_/B _5281_/C _4652_/A1 _5295_/A3 _5291_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_30_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5593_ _5875_/A3 _3523_/Z hold389/Z _5620_/A4 _5601_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_157_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4544_ _5270_/A2 _5420_/A4 _5276_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_128_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold402 _6936_/Q hold402/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold413 _5661_/Z _7016_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold424 _6884_/Q hold424/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold435 _4108_/Z _6668_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7263_ _7263_/D _7269_/CLK _7263_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold446 _7121_/Q hold446/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_132_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4475_ _5288_/C _4454_/Z _4367_/Z _4449_/B _4692_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold457 _5876_/Z _7206_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold468 _5560_/Z _6926_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6214_ _6825_/Q _5988_/Z _6019_/Z _6854_/Q _6217_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_89_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold479 hold479/I hold479/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3426_ _3304_/I _6732_/Q _6730_/Q _3434_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_7194_ hold81/Z _7194_/RN _7194_/CLK hold80/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6145_ _6954_/Q _5958_/Z _5994_/I _7140_/Q _6147_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3357_ _7097_/Q _3357_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6076_ _7089_/Q _6002_/Z _6015_/Z _7007_/Q _6076_/C _6078_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_39_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5027_ _5027_/I _5200_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6978_ _6978_/D _7124_/RN _6978_/CLK _6978_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_94_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5929_ _5925_/Z _6117_/A2 _6168_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_167_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold980 _5751_/Z _7095_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold991 _7150_/Q hold991/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_88_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4260_ _5645_/I1 hold246/Z _4261_/S _4260_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4191_ _4191_/A1 _6611_/A2 _4193_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_79_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6901_ _6901_/D _7225_/RN _6901_/CLK _6901_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6832_ _6832_/D _7261_/RN _7279_/CLK _6832_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_91_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6763_ _6763_/D _6854_/RN _6763_/CLK _6763_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3975_ _3483_/Z _3975_/I1 _3975_/S _3975_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5714_ _5879_/I0 hold261/Z _5718_/S _5714_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6694_ _6694_/D _6886_/RN _6694_/CLK _6694_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_50_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5645_ hold166/Z _5645_/I1 _5646_/S _5645_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5576_ hold983/Z _5795_/I0 _5583_/S _5576_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold210 _3501_/Z hold210/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold221 hold221/I hold221/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4527_ _5020_/A2 _4889_/A1 _5243_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold232 hold232/I hold232/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold243 _5825_/Z _7161_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold254 _6661_/Q _3470_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold265 _6776_/Q hold265/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7246_ _7246_/D _7258_/RN _7260_/CLK _7246_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4458_ _4467_/A1 _4555_/B _4736_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold276 _5547_/Z _6915_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_160_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold287 _6886_/Q hold287/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_172_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout701 fanout714/Z _7253_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold298 _4264_/Z _6778_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_120_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout712 _7071_/RN _6650_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_131_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3409_ _3441_/C _6664_/Q _6663_/Q _3409_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xfanout723 input124/Z _4449_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7177_ _7177_/D _7177_/RN _7177_/CLK _7177_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout734 input121/Z _5458_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4389_ _4427_/A2 _4427_/A3 _4485_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xfanout745 _4877_/A2 _4483_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6128_ _7065_/Q _5985_/Z _5997_/Z _7099_/Q _6128_/C _6134_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_100_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6059_ _7030_/Q _5999_/Z _6014_/Z _6958_/Q _6000_/Z _7128_/Q _6061_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_3116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3760_ _3760_/A1 _3739_/Z _3759_/Z _6567_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_13_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3691_ _3690_/Z _3691_/I1 _3899_/S _6873_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5430_ _5268_/Z _5430_/A2 _5428_/Z _5429_/Z _5431_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_69_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput304 _4069_/Z serial_resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5361_ _5361_/A1 _5209_/Z _5362_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xoutput315 _6806_/Q wb_dat_o[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_58_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput326 _6798_/Q wb_dat_o[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput337 _6815_/Q wb_dat_o[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4312_ _6571_/I0 _6818_/Q _4312_/S _6818_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_126__1359_ _4073__49/I net852_138/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7100_ _7100_/D _7179_/RN _7100_/CLK _7100_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xclkbuf_leaf_46__1359_ clkbuf_4_14_0__1359_/Z net802_68/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_141_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5292_ _5423_/A2 _5292_/A2 _5292_/A3 _5292_/A4 _5294_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_142_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7031_ _7031_/D _7034_/RN _7031_/CLK _7031_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4243_ _4242_/Z hold408/Z _4245_/S _4243_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4174_ _4180_/I0 _4174_/I1 _4175_/S _4174_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6815_ _6815_/D _7258_/CLK _6815_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6746_ _6746_/D _7225_/RN _4067_/I1 _6746_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3958_ _3958_/A1 _3958_/A2 _3958_/A3 _3958_/A4 _3958_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_177_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3889_ _3889_/A1 _3889_/A2 _3889_/A3 _3889_/A4 _3889_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6677_ _6677_/D _6839_/RN _6677_/CLK _6677_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_109_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5628_ _5784_/I0 hold779/Z _5628_/S _5628_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5559_ _5859_/I0 hold799/Z _5565_/S _5559_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7229_ _7229_/D _7255_/RN _7257_/CLK _7229_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout520 _5842_/I0 _5797_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout531 _5751_/I0 _5832_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout542 _5732_/I0 _6612_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout553 _5674_/A2 _5647_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_116_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout564 _3329_/I _6296_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout575 _6597_/C1 _3317_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xfanout586 _6745_/Q _4009_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout597 _5369_/A1 _4873_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_74_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet1152_411 net1152_427/I _6763_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet1152_422 net902_179/I _6752_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1152_433 net1152_434/I _6737_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_444 net1202_474/I _6721_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4930_ _4930_/A1 _5325_/B _3404_/I _5170_/A2 _4930_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_75_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4861_ _4887_/A1 _4868_/A1 _5364_/A1 _4873_/A3 _4861_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_2790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6600_ _6600_/A1 _6600_/A2 _6600_/B1 _6600_/B2 _3317_/I _6600_/C2 _6601_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3812_ _5821_/A2 _3578_/Z _4146_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4792_ _4492_/Z _4534_/Z _5129_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6531_ _6821_/Q _6531_/A2 _6554_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_20_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3743_ _7063_/Q _3927_/B1 _3924_/A2 _6967_/Q _3743_/C _3759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_119_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3674_ _3674_/A1 _3674_/A2 _3674_/A3 _3673_/Z _3674_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6462_ _7172_/Q _6544_/A2 _6544_/B1 _6962_/Q _6464_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_118_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5413_ _5448_/A1 _5483_/A1 _5412_/Z _5414_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6393_ _3324_/I _7253_/Q _6393_/B _6394_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5344_ _5438_/C _5475_/A4 _5387_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_114_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput167 _4087_/Z debug_in VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_115_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput178 _3363_/ZN mgmt_gpio_oeb[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput189 _3353_/ZN mgmt_gpio_oeb[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5275_ _5376_/B2 _5468_/A2 _5275_/B _5423_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_130_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4226_ _4225_/Z hold183/Z _4228_/S _4226_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7014_ _7014_/D _7124_/RN _7014_/CLK _7014_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_101_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4157_ _5775_/I0 hold623/Z _4157_/S _4157_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4088_ _6906_/Q input70/Z _4088_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_83_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6729_ _6729_/D _7170_/RN _6729_/CLK _6729_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_20_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_92__1359_ clkbuf_4_7_0__1359_/Z net952_216/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_28_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout350 _6657_/A2 _6656_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout361 _4689_/ZN _5315_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xnet1102_352 net1152_437/I _6858_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1102_363 net1102_382/I _6847_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout372 _3533_/Z _3932_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout383 _5611_/A1 _5629_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xnet1102_374 net1202_486/I _6825_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1102_385 net1202_486/I _6789_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout394 _6274_/Z _6543_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_115_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1102_396 net902_199/I _6778_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput14 mask_rev_in[19] input14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput25 mask_rev_in[29] input25/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput36 mgmt_gpio_in[0] input36/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput47 mgmt_gpio_in[1] input47/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput58 mgmt_gpio_in[2] input58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_10_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput69 mgmt_gpio_in[6] input69/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold809 _6682_/Q hold809/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3390_ _7241_/Q _6011_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ _5058_/Z _5060_/A2 _4928_/Z _5060_/A4 _5064_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_84_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4011_ _6282_/A2 _7232_/Q _6402_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_111_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5962_ _5984_/A1 _7230_/Q _6002_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_80_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4913_ _4376_/Z _5323_/B _4909_/Z _4927_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_5893_ _5945_/A1 _5951_/B _5894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4844_ _4873_/A3 _5420_/A4 _4530_/I _4873_/A2 _4844_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_33_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4775_ _4775_/A1 _4772_/Z _4773_/Z _4774_/Z _4781_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6514_ _6787_/Q _6545_/A2 _6545_/B1 _6843_/Q _6516_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_147_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3726_ _4297_/I0 _6871_/Q _3898_/S _3726_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6445_ _7049_/Q _6550_/A2 _6550_/C1 _6953_/Q _6535_/A2 _7211_/Q _6446_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3657_ _3657_/A1 _3657_/A2 _3657_/A3 _3657_/A4 _3657_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_134_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3588_ _7133_/Q _3930_/A2 _3941_/B1 _7173_/Q _3588_/C _3589_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6376_ _7113_/Q _6240_/Z _6376_/B _6384_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_103_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5327_ _4928_/Z _5326_/Z _5327_/A3 _5327_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_102_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5258_ _4890_/I _5258_/A2 _4972_/Z _5258_/B2 _5258_/C _5412_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_87_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4209_ _4208_/Z hold319/Z _4211_/S _4209_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5189_ _5386_/A1 _5386_/A3 _5189_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_68_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4560_ _5002_/A3 _5002_/A4 _5080_/B _5393_/B1 _4561_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_184_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3511_ _3904_/A3 hold221/I _3511_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_128_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold606 _5748_/Z _7093_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4491_ _4491_/A1 _4491_/A2 _4491_/B _5312_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_6_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold617 _6707_/Q hold617/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold628 _5718_/Z _7067_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6230_ _6529_/S _7249_/Q _6230_/B _6231_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold639 _6729_/Q hold639/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3442_ _3991_/A1 _4042_/A3 _3304_/I _3442_/B _3443_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_40_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6161_ _6161_/I _6162_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3373_ _6975_/Q _3373_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5112_ _5478_/A1 _5478_/A3 _5228_/A3 _5230_/B _5226_/A1 _5113_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XTAP_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6092_ _6092_/A1 _5991_/Z _6102_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5043_ _5385_/A1 _5043_/A2 _5043_/B _5432_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_0_wbbd_sck _7278_/Q clkbuf_0_wbbd_sck/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_25_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6994_ _6994_/D _7188_/RN _6994_/CLK _6994_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5945_ _5945_/A1 _4009_/B _5945_/B _5950_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_179_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5876_ _5876_/I0 hold456/Z _5883_/S _5876_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4827_ _5367_/A2 _5228_/A3 _5223_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_178_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4758_ _4973_/A4 _4500_/Z _4958_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_105_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3709_ _7210_/Q _3960_/A2 _3955_/A2 _7202_/Q _7186_/Q _3959_/C1 _3724_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_162_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4689_ _4687_/Z _5092_/A1 _4689_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_135_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6428_ _7009_/Q _6549_/B1 _6552_/A2 _7033_/Q _6440_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_134_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6359_ _6359_/I _6360_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_173_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold3 hold3/I hold3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_94_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3991_ _3991_/A1 _3412_/Z _3442_/B _3409_/Z _6730_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_5730_ hold735/Z _5778_/I0 _5730_/S _5730_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5661_ hold412/Z _5871_/I0 _5664_/S _5661_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4612_ _4612_/A1 _4612_/A2 _5025_/B _4618_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5592_ _5592_/I0 hold6/Z hold34/Z hold35/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4543_ _5129_/A3 _4873_/A2 _4878_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_117_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold403 _5571_/Z _6936_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold414 _7052_/Q hold414/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold425 _5505_/Z _6884_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_7_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold436 _6990_/Q hold436/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7262_ _7262_/D _7262_/CLK _7262_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4474_ _5288_/C _5269_/A1 _4367_/Z _4501_/B _4474_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold447 _5780_/Z _7121_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold458 _7061_/Q hold458/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6213_ _6821_/Q _5979_/Z _5996_/Z _6709_/Q _6217_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold469 _6902_/Q hold469/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3425_ _4041_/A3 _7302_/Q _3425_/S _7302_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7193_ _7193_/D _7193_/RN _7193_/CLK _7193_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_171_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6144_ _7066_/Q _5985_/Z _6000_/Z _7132_/Q _6144_/C _6147_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3356_ _7105_/Q _3356_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6075_ _7015_/Q _5971_/Z _6003_/Z _7161_/Q _6078_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5026_ _5471_/B2 _5291_/B _5002_/Z _5200_/B1 _5027_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_2608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6977_ _6977_/D _7083_/RN _6977_/CLK _6977_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_55_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5928_ _6068_/A2 _5941_/A1 _5931_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_110_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5859_ _5859_/I0 _5859_/I1 _5865_/S _5859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold970 _5814_/Z _7151_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold981 _7111_/Q hold981/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold992 _5813_/Z _7150_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_77_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4190_ hold619/Z _4361_/I1 _4190_/S _4190_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6900_ _6900_/D _7238_/RN _6900_/CLK _6900_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_78_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6831_ _6831_/D _7261_/RN _7279_/CLK _6831_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6762_ _6762_/D _7177_/RN _6762_/CLK _6762_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_126_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3974_ _6661_/Q _6660_/Q _6659_/Q _3972_/Z _3975_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_165_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5713_ _5860_/I0 hold179/Z _5718_/S _5713_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6693_ _6693_/D _6786_/RN _6693_/CLK _6693_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_188_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5644_ hold554/Z _5818_/I0 _5646_/S _5644_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5575_ _5575_/A1 _5674_/A2 _5583_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_145_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold200 _4220_/Z _6750_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold211 hold211/I hold211/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4526_ _4440_/B _4501_/B _5458_/A4 _3408_/I _4526_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold222 _3904_/Z hold222/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold233 hold233/I hold233/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold244 _7047_/Q hold244/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_132_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold255 hold255/I _3471_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7245_ _7245_/D _7258_/RN _7260_/CLK _7245_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold266 _4261_/Z _6776_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4457_ _5420_/A4 _4873_/A2 _4460_/B _4467_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xhold277 _7020_/Q hold277/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold288 _5507_/Z _6886_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold299 _6680_/Q hold299/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xfanout702 _7185_/RN _7188_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout713 fanout714/Z _7071_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3408_ _3408_/I _4903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_7176_ _7176_/D fanout655/Z _7176_/CLK _7176_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xfanout724 input124/Z _4501_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_59_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout735 _4589_/A4 _3403_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4388_ _4388_/A1 _4388_/A2 input97/Z input96/Z _4427_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xfanout746 _4877_/A2 _4395_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6127_ _6127_/A1 _6124_/Z _6127_/A3 _6127_/A4 _6127_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3339_ _3339_/I _3932_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6058_ _7062_/Q _5985_/Z _5997_/Z _7096_/Q _6061_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_22_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5009_ _4517_/Z _5020_/A2 _5435_/A2 _5475_/A3 _5009_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_38_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3690_ _6569_/I0 _6872_/Q _3898_/S _3690_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_187_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput305 _4086_/Z spi_sdi VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5360_ _5045_/C _5393_/B1 _5360_/B _5360_/C _5361_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_160_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput316 _6807_/Q wb_dat_o[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput327 _7262_/Q wb_dat_o[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput338 _6816_/Q wb_dat_o[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4311_ _6570_/I0 _6817_/Q _4312_/S _6817_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5291_ _4542_/Z _5291_/A2 _5291_/B _5291_/C _5377_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_142_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7030_ _7030_/D _6967_/RN _7030_/CLK _7030_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_142_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4242_ hold331/Z _5555_/I0 _4242_/S _4242_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_opt_1_0__1359_ _4073__6/I clkbuf_opt_1_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4173_ _5517_/A1 hold146/Z _4185_/A2 _5821_/A1 _4173_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_132_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6814_ _6814_/D _7262_/CLK _6814_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6745_ _6745_/D _7225_/RN _4067_/I1 _6745_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3957_ _6956_/Q _3957_/A2 _4289_/A1 _6799_/Q _3958_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_50_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6676_ _6676_/D _6839_/RN _6676_/CLK _6676_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_164_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3888_ _6989_/Q _3954_/A2 _3956_/A2 _7119_/Q _3889_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5627_ _5681_/I1 hold759/Z _5628_/S _5627_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5558_ hold64/Z hold226/Z _5565_/S _5558_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4509_ _5087_/A1 _5051_/S _5343_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5489_ _5489_/A1 _5489_/A2 _5472_/Z _5489_/A4 _5489_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_120_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7228_ _7228_/D _7255_/RN _7257_/CLK _7228_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
Xfanout510 _5808_/I0 _5781_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout521 _5833_/I0 _5869_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout532 _5751_/I0 _5859_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout543 _4180_/I0 _5732_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7159_ _7159_/D _6786_/RN _7159_/CLK _7159_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_76_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout554 hold33/I _5674_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout565 _7234_/Q _3329_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout576 _6836_/Q _6597_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout587 _6364_/C _6529_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xfanout598 _4563_/Z _5369_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_86_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_52__1359_ clkbuf_4_14_0__1359_/Z net802_94/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_187_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_132__1359_ net1152_446/I net1202_481/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_23_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1152_412 net852_120/I _6762_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_157_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1152_423 net952_225/I _6751_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_434 net1152_434/I _6736_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_155_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet1152_445 net1202_474/I _6720_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4860_ _5104_/A1 _4860_/A2 _5276_/B _5291_/B _5376_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_2780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3811_ _5629_/A1 _3578_/Z _3925_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_60_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4791_ _5312_/A2 _5214_/A2 _5456_/A1 _5220_/B2 _4791_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6530_ _7259_/Q _6529_/Z _6558_/S _7259_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3742_ _3742_/I _3743_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_186_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6461_ _7220_/Q _6274_/Z _6285_/Z _7196_/Q _7180_/Q _6254_/Z _6464_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3673_ _3673_/A1 _3673_/A2 _3673_/A3 _3673_/A4 _3673_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5412_ _5412_/A1 _5412_/A2 _5412_/A3 _4984_/B _5412_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_173_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6392_ _6385_/Z _6391_/Z _6392_/B1 _6286_/Z _6500_/C _6393_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_161_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5343_ _5343_/A1 _5343_/A2 _5343_/B _5418_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xoutput168 _6894_/Q irq[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput179 _3362_/ZN mgmt_gpio_oeb[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_82_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5274_ _5370_/A1 _5312_/A4 _5276_/B _5295_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_87_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7013_ _7013_/D fanout658/Z _7013_/CLK _7013_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4225_ hold158/Z _5645_/I1 _4225_/S _4225_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4156_ _5855_/I0 hold709/Z _4157_/S _4156_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4087_ input1/Z input36/Z _4087_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_56_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4989_ _5340_/A1 _5262_/A2 _5328_/A2 _5248_/A2 _4991_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6728_ _6728_/D _7170_/RN _6728_/CLK _6728_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_108_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6659_ _6659_/D _6614_/Z _4072_/B2 _6659_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_164_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout351 _4064_/S _6657_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xnet1102_353 net1152_437/I _6857_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout362 _5302_/B _5307_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout373 _3844_/A1 _4353_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet1102_364 net802_55/I _6846_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout384 _3509_/Z _5611_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet1102_375 net1202_486/I _6824_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1102_386 net1202_471/I _6788_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout395 _6272_/Z _6540_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xnet1102_397 net1152_427/I _6777_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_46_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput15 mask_rev_in[1] input15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 mask_rev_in[2] input26/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput37 mgmt_gpio_in[10] input37/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput48 mgmt_gpio_in[20] input48/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput59 mgmt_gpio_in[30] input59/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4010_ _4010_/I _6744_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5961_ _6948_/Q _5958_/Z _5960_/Z _7150_/Q _5974_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4912_ _5464_/A1 _5443_/A1 _5193_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5892_ _5892_/I0 hold675/Z _5892_/S _5892_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4843_ _4873_/A3 _5228_/A3 _5231_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_178_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4774_ _4782_/A1 _5236_/A1 _4774_/A3 _4695_/Z _4774_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_187_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6513_ _6809_/Q _6544_/B1 _6550_/C1 _6799_/Q _6549_/C1 _6839_/Q _6516_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_20_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3725_ _3708_/Z _3724_/Z _3725_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_146_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6444_ _7219_/Q _6543_/A2 _6285_/Z _7195_/Q _7179_/Q _6254_/Z _6446_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3656_ hold66/I _3546_/Z _3945_/C2 hold50/I _3657_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_146_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6375_ _7129_/Q _6452_/A2 _6452_/A3 _6484_/A4 _6376_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3587_ _3587_/I _3588_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5326_ _5246_/Z _5442_/A4 _5442_/A2 _5442_/A1 _5326_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_103_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5257_ _5257_/A1 _5246_/Z _5257_/B _5257_/C _5264_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_57_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4208_ hold246/Z _5645_/I1 _4210_/S _4208_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5188_ _5243_/A1 _5043_/B _5205_/A1 _4650_/Z _5386_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4139_ _4361_/I1 hold477/Z _4139_/S _4139_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3510_ _3507_/Z _5611_/A1 _5584_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4490_ _4491_/A1 _4491_/A2 _5092_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold607 _7173_/Q hold607/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_128_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold618 _4160_/Z _6707_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold629 _6850_/Q hold629/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_7_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3441_ _6664_/Q _6663_/Q _6730_/Q _3441_/C _3443_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_143_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6160_ _6364_/C _7246_/Q _6160_/B _6161_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3372_ _6983_/Q _3372_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5111_ _5478_/A1 _5142_/A3 _5111_/B _5111_/C _5113_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ _7024_/Q _6211_/A2 _6211_/B1 _6992_/Q _6092_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5042_ _5385_/A1 _5389_/C _5439_/B1 _5393_/A1 _5044_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6993_ _6993_/D _7155_/RN _6993_/CLK _6993_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_41_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5944_ _4009_/B _7235_/Q _3329_/I _6300_/A2 _5945_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5875_ _5875_/A1 _3523_/Z _5875_/A3 _5883_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_4826_ _4826_/A1 _5370_/B _4826_/A3 _4826_/B _4834_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_179_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4757_ _4757_/I _4766_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3708_ _3701_/Z _3708_/A2 _3708_/A3 _3707_/Z _3708_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_146_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4688_ _5080_/B _5092_/A1 _5312_/A1 _5094_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_119_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6427_ _6945_/Q _6551_/A2 _6288_/Z _7123_/Q _6440_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_146_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3639_ _7140_/Q _3951_/A2 _5665_/A1 _7026_/Q _7018_/Q _5656_/A1 _3642_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_108_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6358_ _7022_/Q _6549_/A2 _6549_/B1 _7006_/Q _6549_/C1 _6998_/Q _6359_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_88_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5309_ _5403_/A1 _5309_/A2 _5456_/A2 _5309_/B2 _5309_/C _5310_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6289_ _7182_/Q _6532_/A2 _6288_/Z _7118_/Q _6307_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_57_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold4 hold4/I hold4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_63_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3990_ _3990_/I _5896_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_15_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5660_ hold471/Z _5798_/I0 _5664_/S _5660_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4611_ _4446_/Z _4565_/Z _5025_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_175_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5591_ hold170/Z _5645_/I1 hold34/Z _6954_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4542_ _5055_/A2 _5129_/A3 _4873_/A2 _4542_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_156_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold404 _6960_/Q hold404/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_172_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold415 _5702_/Z _7052_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7261_ _7261_/D _7261_/RN _7279_/CLK _7261_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold426 _6927_/Q hold426/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4473_ _4472_/B _4473_/A2 _4481_/A2 _4853_/A1 _4786_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
Xhold437 _5632_/Z _6990_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold448 _7089_/Q hold448/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold459 _5712_/Z _7061_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6212_ _6212_/A1 _5991_/Z _6226_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_89_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3424_ _3465_/A4 _3465_/A3 _3971_/A1 _3442_/B _3425_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7192_ _7192_/D _7221_/RN _7192_/CLK _7192_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xclkbuf_leaf_29__1359_ clkbuf_opt_3_0__1359_/Z _4073__32/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_131_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_109__1359_ clkbuf_4_4_0__1359_/Z net1202_463/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6143_ _6143_/I _6144_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3355_ _7113_/Q _3355_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6074_ _7081_/Q _5996_/Z _6005_/Z _7039_/Q _6078_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5025_ _5439_/B2 _5200_/B1 _5025_/B _5476_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_54_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6976_ _6976_/D _7260_/RN _6976_/CLK _6976_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_54_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5927_ _5919_/Z _6014_/A2 _5941_/A1 _5925_/Z _5950_/A1 _7230_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_179_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5858_ _5885_/I0 _5858_/I1 _5865_/S _5858_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4809_ _4809_/A1 _4805_/Z _4807_/Z _4808_/Z _4812_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5789_ _5852_/I0 hold817/Z _5793_/S _5789_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold960 _5630_/Z _6988_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold971 _7094_/Q hold971/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_1_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold982 _5769_/Z _7111_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_150_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold993 _7110_/Q hold993/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_1_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6830_ _6833_/Q _7261_/RN _7279_/CLK _6830_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_36_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6761_ _6761_/D _7240_/RN _6761_/CLK _6761_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3973_ _6660_/Q _6659_/Q _3972_/Z _3973_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_189_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5712_ _5850_/I0 hold458/Z _5718_/S _5712_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6692_ _6692_/D _6786_/RN _6692_/CLK _6692_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5643_ hold550/Z _5781_/I0 _5646_/S _5643_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5574_ _5811_/I0 hold847/Z _5574_/S _5574_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold201 _6749_/Q hold201/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4525_ _5315_/A2 _4524_/Z _5130_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold212 hold212/I hold212/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold223 hold223/I _6894_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold234 _7011_/Q hold234/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7244_ _7244_/D _7258_/RN _7260_/CLK _7244_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold245 _5696_/Z _7047_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold256 _3473_/Z hold256/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4456_ _3401_/I _4547_/A4 _4456_/B _4456_/C _4481_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xhold267 _6999_/Q hold267/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold278 _5666_/Z _7020_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold289 _7108_/Q hold289/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xfanout703 _7185_/RN _6656_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3407_ _3407_/I _3407_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7175_ _7175_/D _7215_/RN _7175_/CLK _7175_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xfanout714 input75/Z fanout714/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_113_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4387_ _4388_/A1 _4388_/A2 input97/Z input96/Z _4387_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xfanout725 _4440_/B _4472_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout736 _4589_/A4 _5420_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6126_ _7083_/Q _5996_/Z _5999_/Z _7033_/Q _6969_/Q _5979_/Z _6127_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout747 input107/Z _4877_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3338_ _6927_/Q _6392_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XTAP_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6057_ _6057_/A1 _6057_/A2 _6057_/A3 _6057_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XTAP_3107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5008_ _5438_/C _5020_/A2 _5439_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_39_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6959_ hold89/Z _7247_/RN _6959_/CLK hold88/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_179_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold790 _5673_/Z _7027_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xclkbuf_leaf_12__1359_ net1152_430/I _4073__31/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_75__1359_ net902_187/I net802_95/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_39_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_0__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _4075_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_164_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput306 _4081_/Z spimemio_flash_io0_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput317 _6808_/Q wb_dat_o[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_126_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4310_ _6569_/I0 _6816_/Q _4312_/S _6816_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput328 _7263_/Q wb_dat_o[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput339 _6817_/Q wb_dat_o[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5290_ _5290_/A1 _5290_/A2 _5290_/A3 _4483_/B _5290_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4241_ _4240_/Z hold499/Z _4245_/S _4241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4172_ hold863/Z _5832_/I0 _4172_/S _4172_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6813_ _6813_/D _7262_/CLK _6813_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3956_ _7118_/Q _3956_/A2 _3956_/B1 _6712_/Q _3956_/C1 _6851_/Q _3958_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6744_ _6744_/D _7240_/RN _4067_/I1 _6744_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_52_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6675_ _6675_/D _6882_/RN _6675_/CLK _6675_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3887_ _6840_/Q _3925_/C2 _3956_/C1 _6852_/Q _3889_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_177_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5626_ _5818_/I0 hold490/Z _5628_/S _5626_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5557_ _5866_/A3 _3527_/Z _5839_/A3 _5857_/A3 _5565_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_105_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4508_ _4698_/B _5087_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_104_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _5374_/Z _5487_/Z _5489_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_104_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7227_ _7227_/D _7255_/RN _7257_/CLK _7227_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4439_ _4363_/Z _4369_/Z _4440_/B _4759_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xfanout500 _5782_/I0 _5818_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout511 _5724_/I0 _5808_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_59_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout522 _5833_/I0 _5806_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout533 _5751_/I0 _5886_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_104_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7158_ _7158_/D _6786_/RN _7158_/CLK _7158_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xfanout544 _5885_/I0 _5822_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_76_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout555 hold32/Z hold33/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout566 _6068_/A2 _3385_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6109_ _6101_/Z _6106_/Z _6109_/A3 _6109_/A4 _6109_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout577 _6600_/B2 _3316_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xfanout588 _6555_/C _6364_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7089_ _7089_/D _7219_/RN _7089_/CLK _7089_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
Xfanout599 _4643_/A4 _5364_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_18_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1152_402 net1152_434/I _6772_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1152_413 net1152_415/I _6761_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_424 net1152_425/I _6750_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_435 net1152_435/I _6735_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_446 net1152_446/I _6719_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3810_ _4332_/A1 _3560_/Z _4301_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_60_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4790_ _4790_/A1 _5213_/C _4787_/Z _4789_/Z _4803_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_162_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3741_ _7081_/Q _3923_/C1 _5575_/A1 _6943_/Q _3925_/A2 input6/Z _3742_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6460_ _6994_/Q _6237_/Z _6247_/Z _7132_/Q _6460_/C _6465_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_146_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3672_ hold46/I _3943_/A2 _3941_/A2 _7163_/Q _3673_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_173_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5411_ _5248_/Z _5327_/Z _5411_/A3 _5483_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_63_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6391_ _6554_/A1 _6391_/A2 _6391_/A3 _6390_/Z _6391_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_174_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5342_ _5342_/I _5418_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput169 _4088_/Z irq[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_88_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5273_ _5290_/A2 _5287_/A2 _5364_/B _5468_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_7012_ _7012_/D _7140_/RN _7012_/CLK _7012_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_101_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4224_ _4223_/Z hold383/Z _4228_/S _4224_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4155_ hold40/Z hold42/Z _4157_/S hold43/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4086_ _4055_/S input63/Z _4086_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_83_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4988_ _5083_/C _4568_/Z _4659_/Z _5173_/A2 _4988_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6727_ _6727_/D _7170_/RN _6727_/CLK _6727_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3939_ _6696_/Q _4146_/A1 _4359_/A1 _6857_/Q _3939_/C1 _6710_/Q _3940_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6658_ _6658_/D _4098_/Z _4072_/B2 _6658_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_125_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ _5837_/I0 hold567/Z _5610_/S _5609_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6589_ _6589_/A1 _6601_/A2 _6589_/B _6590_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_180_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout352 _3543_/ZN _4244_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_87_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet1102_354 _4073__35/I _6856_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout363 _4689_/ZN _5302_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_115_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout374 _5692_/A1 _3844_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet1102_365 net802_55/I _6845_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1102_376 net1202_481/I _6823_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout385 _5785_/A3 _5857_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_143_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet1102_387 net802_71/I _6787_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout396 _6269_/Z _6552_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_19_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet1102_398 net1152_431/I _6776_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput16 mask_rev_in[20] input16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput27 mask_rev_in[30] input27/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput38 mgmt_gpio_in[11] input38/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput49 mgmt_gpio_in[21] input49/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5960_ _3385_/I _6164_/A2 _6021_/A2 _3387_/I _5960_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4911_ _5464_/A1 _4903_/Z _5205_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5891_ _5891_/I0 hold711/Z _5892_/S _5891_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4842_ _5104_/A1 _4860_/A2 _4555_/C _5276_/B _4842_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4773_ _4782_/A1 _4774_/A3 _4695_/Z _5226_/A1 _4773_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_159_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6512_ _6512_/A1 _6512_/A2 _6512_/A3 _6511_/Z _6512_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3724_ _3715_/Z _3724_/A2 _3724_/A3 _3723_/Z _3724_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_147_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6443_ _7025_/Q _6549_/A2 _6544_/B1 _6961_/Q _6443_/C _6446_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3655_ _7219_/Q _3912_/A2 _3948_/C1 _7309_/I _3657_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_162_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6374_ _7209_/Q _6535_/A2 _6545_/A2 _6935_/Q _6385_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_173_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3586_ _6931_/Q _3935_/A2 _3943_/A2 _7075_/Q _7157_/Q _3916_/A2 _3587_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5325_ _5329_/A2 _5394_/A2 _5325_/B _5327_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_130_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5256_ _5262_/A2 _4902_/Z _5246_/Z _5257_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_69_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4207_ _4206_/Z hold488/Z _4211_/S _4207_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5187_ _5392_/B _5339_/A4 _5417_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4138_ _4360_/I1 hold465/Z _4139_/S _4138_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4069_ _7238_/Q _6897_/Q _6900_/Q _4069_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold608 _5838_/Z _7173_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold619 _6727_/Q hold619/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3440_ _4056_/I1 _3440_/I1 _3440_/S _7294_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3371_ _6991_/Q _3371_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5110_ _5478_/A1 _5142_/A3 _5111_/C _5479_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6090_ _6210_/A2 _7056_/Q _6090_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_88_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5041_ _5439_/B1 _5002_/Z _5041_/B _5386_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_0_wb_clk_i wb_clk_i clkbuf_0_wb_clk_i/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_38_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6992_ _6992_/D _7141_/RN _6992_/CLK _6992_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_92_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5943_ _5943_/I0 _5940_/Z _5943_/S _7235_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5874_ _5892_/I0 hold719/Z _5874_/S _5874_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4825_ _4539_/I _5287_/A2 _4826_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_138_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4756_ _5236_/A1 _4752_/Z _4757_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_105_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3707_ _3707_/A1 _3707_/A2 _3707_/A3 _3707_/A4 _3707_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4687_ _5080_/B _4687_/A2 _4687_/A3 _4687_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_147_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6426_ _6969_/Q _6531_/A2 _6545_/B1 _7017_/Q _6426_/C _6440_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_108_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3638_ _3638_/A1 _3638_/A2 _3638_/A3 _3638_/A4 _3638_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_161_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6357_ _6357_/A1 _6357_/A2 _6356_/Z _6357_/A4 _6357_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3569_ _5884_/A2 _5692_/A1 _5674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_103_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5308_ _5303_/Z _5308_/A2 _5221_/I _5480_/A1 _5308_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6288_ _5946_/S _6302_/A3 _6533_/A4 _6302_/A4 _6288_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_130_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _5238_/Z _4801_/Z _5453_/A4 _5452_/A2 _5241_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_124_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_140_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold5 hold5/I hold5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_181_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4610_ _5287_/C _4589_/Z _4612_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5590_ hold541/Z _5818_/I0 hold34/Z _6953_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4541_ _5278_/C _5279_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_156_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold405 _5598_/Z _6960_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7260_ _7260_/D _7260_/RN _7260_/CLK _7260_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold416 _7053_/Q hold416/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4472_ _4464_/Z _5270_/A2 _4472_/B _4764_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold427 _5561_/Z _6927_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold438 _7081_/Q hold438/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6211_ _6846_/Q _6211_/A2 _6211_/B1 _6838_/Q _6212_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold449 _5744_/Z _7089_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_132_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3423_ _3422_/Z _7303_/Q _3988_/S _7303_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7191_ _7191_/D _7215_/RN _7191_/CLK _7191_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XTAP_710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6142_ _6978_/Q _5964_/Z _5981_/Z _6938_/Q _6014_/Z _6962_/Q _6143_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_48_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3354_ _7121_/Q _3354_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6073_ _6073_/A1 _6073_/A2 _6073_/A3 _6073_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XTAP_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _4604_/Z _5475_/A3 _5200_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_39_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet852_150 net852_150/I _7075_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6975_ _6975_/D _7024_/RN _6975_/CLK _6975_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_5926_ _5950_/A1 _5925_/Z _5931_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_22_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5857_ _5857_/A1 _5857_/A2 _5857_/A3 _5857_/A4 _5865_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_181_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4808_ _5173_/A2 _4808_/A2 _5312_/A1 _5475_/A4 _4808_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_21_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5788_ _5869_/I0 hold913/Z _5793_/S _5788_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4739_ _4739_/A1 _5106_/A1 _4738_/Z _4743_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_175_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6409_ hold22/I _6544_/A2 _6544_/B1 _6960_/Q _6545_/B1 _7016_/Q _6411_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold950 _5614_/Z _6974_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold961 _7126_/Q hold961/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold972 _5750_/Z _7094_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold983 _6940_/Q hold983/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold994 _5768_/Z _7110_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_131_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_4_0__1359_ clkbuf_0__1359_/Z clkbuf_4_4_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_9_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_115__1359_ clkbuf_4_4_0__1359_/Z net952_245/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_35__1359_ _4073__46/I _4073__8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_8_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_98__1359_ clkbuf_4_5_0__1359_/Z net952_228/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_9_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6760_ _6760_/D _7179_/RN _6760_/CLK _6760_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_90_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3972_ _7305_/Q _7304_/Q _7303_/Q _6658_/Q _3972_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5711_ _5804_/I0 hold905/Z _5718_/S _5711_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6691_ _6691_/D _7170_/RN _6691_/CLK _6691_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_176_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5642_ hold267/Z _5879_/I0 _5646_/S _5642_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5573_ _5837_/I0 hold582/Z _5574_/S _5573_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold202 _4218_/Z _6749_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4524_ _4460_/B _4752_/A2 _4524_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_117_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold213 _5521_/Z _5527_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold224 _6913_/Q hold224/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold235 _5655_/Z _7011_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7243_ _7243_/D _7258_/RN _7260_/CLK _7243_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold246 _6775_/Q hold246/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4455_ _4555_/B _4455_/A2 _5170_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold257 _3485_/Z hold257/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold268 _5642_/Z _6999_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_160_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold279 _7042_/Q hold279/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3406_ _3406_/I _4522_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_7174_ _7174_/D _7215_/RN _7174_/CLK _7174_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xfanout704 _7071_/RN _7185_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4386_ input99/Z input98/Z _4386_/A3 _4386_/A4 _4427_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xfanout715 input58/Z _4056_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_59_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout726 _4440_/B _5295_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout737 _4589_/A4 _4456_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6125_ _6945_/Q _5972_/Z _6021_/Z _7001_/Q _6127_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3337_ _3337_/I _4082_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout748 _4878_/A4 _3402_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6056_ _7070_/Q _5980_/Z _6005_/Z _7038_/Q _6057_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_105_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5007_ _5435_/A2 _5475_/A3 _5194_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_67_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6958_ _6958_/D _7019_/RN _6958_/CLK _6958_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_157_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5909_ _7226_/Q _5908_/Z _5910_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6889_ _6889_/D _6892_/RN _6889_/CLK _6889_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_139_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold780 _5628_/Z _6987_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_1_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold791 _6667_/Q hold791/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_110_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput307 _4082_/ZN spimemio_flash_io1_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput318 _6791_/Q wb_dat_o[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput329 _7264_/Q wb_dat_o[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ hold377/Z _5890_/I0 _4244_/S _4240_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4171_ hold859/Z _5822_/I0 _4172_/S _4171_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6812_ _6812_/D _7262_/CLK _6812_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6743_ _6743_/D _7225_/RN _4067_/I1 _6743_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3955_ _7198_/Q _3955_/A2 _3955_/B1 _6847_/Q _3958_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_91_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6674_ _6674_/D _6894_/RN _6674_/CLK _6674_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3886_ _6790_/Q _3928_/B1 _4289_/A1 _6800_/Q _6810_/Q _4301_/A1 _3889_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5625_ _5781_/I0 hold519/Z _5628_/S _5625_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5556_ _5892_/I0 hold495/Z _5556_/S _5556_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4507_ _5420_/A3 _5129_/A3 _3402_/I _4698_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_144_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5487_ _5487_/A1 _5487_/A2 _5487_/A3 _5487_/A4 _5487_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_104_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7226_ _7226_/D _7240_/RN _4067_/I1 _7226_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4438_ _4648_/A1 _4648_/A2 _4438_/B _4438_/C _5190_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xfanout501 _5836_/I0 _5782_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout512 _5880_/I0 _5724_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout523 _5842_/I0 _5833_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_160_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout534 _5850_/I0 _5751_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7157_ _7157_/D _7205_/RN _7157_/CLK _7157_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout545 _5867_/I0 _5885_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4369_ _4836_/A3 _4456_/B _4456_/C _4369_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xfanout556 _6002_/A3 _6021_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_101_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6108_ hold24/I _5960_/Z _5964_/Z _6976_/Q _5981_/Z _6936_/Q _6109_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xfanout567 _6068_/A2 _6117_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout578 _6835_/Q _6600_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout589 _6744_/Q _6555_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7088_ _7088_/D _7202_/RN _7088_/CLK _7088_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_6039_ _6364_/C _7241_/Q _6039_/B _6040_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_73_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1152_403 net1152_434/I _6771_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_414 net1152_414/I _6760_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_182_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1152_425 net1152_425/I _6749_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_163_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1152_436 net802_55/I _6729_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1152_447 _4073__3/I _6718_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3740_ _6935_/Q _3910_/A2 _3927_/C2 input29/Z _3954_/A2 _6991_/Q _3759_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_159_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3671_ _6977_/Q _3923_/A2 _5665_/A1 _7025_/Q _3673_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_185_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5410_ _5410_/A1 _5481_/B1 _5410_/B _5411_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6390_ _6390_/A1 _6390_/A2 _6390_/A3 _6390_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_133_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5341_ _4997_/B _4878_/Z _5341_/B _5341_/C _5342_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_142_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5272_ _5165_/Z _5270_/Z _4877_/Z _5425_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7011_ _7011_/D _7125_/RN _7011_/CLK _7011_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4223_ hold367/Z _5881_/I0 _4227_/S _4223_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4154_ _5871_/I0 hold400/Z _4157_/S _4154_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4085_ _4059_/S input68/Z _4085_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_55_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4987_ _4367_/Z _5340_/A1 _4555_/B _5172_/B _4987_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6726_ _6726_/D _7170_/RN _6726_/CLK _6726_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3938_ _3929_/Z _3938_/A2 _3938_/A3 _3937_/Z _3938_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_20_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6657_ _7185_/RN _6657_/A2 _6657_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3869_ _3869_/A1 _3869_/A2 _3869_/A3 _3868_/Z _3869_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_165_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5608_ _5782_/I0 hold486/Z _5610_/S _5608_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6588_ _6600_/A1 _6588_/A2 _6588_/B1 _3316_/I _3317_/I _6588_/C2 _6589_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5539_ _5857_/A1 _5857_/A3 _5821_/A3 _5857_/A4 _5547_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_145_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7209_ _7209_/D _7221_/RN _7209_/CLK _7209_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xfanout353 _3543_/ZN _4242_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_120_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1102_355 net802_66/I _6855_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout364 _4517_/Z _5438_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout375 _3529_/Z _5692_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet1102_366 net1152_441/I _6844_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1102_377 net852_106/I _6822_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout386 _3503_/ZN _5785_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_115_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1102_388 net902_185/I _6786_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout397 _6266_/Z _6545_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xnet1102_399 net1102_400/I _6775_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput17 mask_rev_in[21] input17/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 mask_rev_in[31] input28/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput39 mgmt_gpio_in[12] input39/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_122_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4910_ _5442_/A2 _4909_/Z _5443_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_33_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5890_ _5890_/I0 hold609/Z _5892_/S _5890_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4841_ _5369_/A1 _4836_/Z _4841_/B _4841_/C _4846_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_2590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4772_ _4782_/A1 _5315_/A4 _4695_/Z _5478_/B1 _4772_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6511_ _6511_/A1 _6511_/A2 _6511_/A3 _6511_/A4 _6511_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3723_ _3719_/Z _3723_/A2 _3723_/A3 _3723_/A4 _3723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_187_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6442_ _6442_/I _6443_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3654_ _5857_/A1 _3653_/Z _3948_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_174_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6373_ _7217_/Q _6543_/A2 _6285_/Z _7193_/Q _7177_/Q _6254_/Z _6385_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3585_ _7221_/Q _3912_/A2 _3959_/C1 _7189_/Q _3589_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_138_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5324_ _5324_/A1 _5324_/A2 _5324_/B _5324_/C _5444_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_177_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5255_ _5258_/B2 _5255_/A2 _5051_/Z _5255_/B _5446_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_4206_ hold205/Z _5890_/I0 _4210_/S _4206_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5186_ _4506_/Z _5260_/A1 _5339_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_111_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4137_ _4353_/A1 _5821_/A1 _5517_/A3 _5629_/A3 _4139_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_28_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4068_ _6760_/Q _3339_/I _6905_/Q _4068_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6709_ _6709_/D _6856_/RN _6709_/CLK _6709_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_184_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold609 _7219_/Q hold609/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_128_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3370_ _6999_/Q _3370_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5040_ _5439_/B1 _5439_/B2 _5040_/B _5040_/C _5044_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6991_ _6991_/D _7075_/RN _6991_/CLK _6991_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_81_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5942_ _5943_/I0 _5936_/Z _5942_/S _7234_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_92_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5873_ _5891_/I0 hold687/Z _5874_/S _5873_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4824_ _4997_/C _5415_/A1 _5370_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_119_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4755_ _4755_/A1 _5313_/A2 _5233_/A1 _4766_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_147_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3706_ _6952_/Q _5584_/A1 _3951_/C1 _7146_/Q _3707_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_88_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4686_ _5240_/B _5214_/A2 _4686_/B _4812_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_162_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6425_ _6425_/I _6426_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3637_ input59/Z _4194_/A1 _3917_/A2 _7116_/Q _5528_/S _3619_/Z _3638_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_134_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6356_ _6356_/A1 _6356_/A2 _6356_/A3 _6355_/Z _6356_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_143_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3568_ _3512_/Z _3732_/A4 _3941_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_89_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5307_ _5367_/A2 _5478_/A2 _5307_/A3 _5307_/B _5480_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_142_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6287_ _6287_/A1 _6287_/A2 _6287_/A3 _6499_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_3499_ _3499_/I _3500_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5238_ _5238_/A1 _5454_/A1 _5238_/A3 _5238_/A4 _5238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_103_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5169_ _5169_/A1 _5425_/A1 _5425_/A3 _5169_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_72_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_138__1359_ net1152_451/I net802_71/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold6 hold6/I hold6/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xclkbuf_leaf_58__1359_ clkbuf_4_15_0__1359_/Z net1152_435/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_48_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4540_ _5365_/A3 _4449_/B _3407_/I _4652_/A1 _5278_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_144_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold406 _7064_/Q hold406/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_7_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4471_ _4853_/A1 _4481_/A2 _4735_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold417 _5703_/Z _7053_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold428 _7136_/Q hold428/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6210_ _6858_/Q _6210_/A2 _6210_/B _6210_/C _6220_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xhold439 _5735_/Z _7081_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3422_ _3422_/I0 _4056_/I1 _3978_/S _3422_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7190_ _7190_/D _6856_/RN _7190_/CLK _7190_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_125_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6141_ _6141_/A1 _5991_/Z _6146_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3353_ _7129_/Q _3353_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_152_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6072_ _7121_/Q _5969_/Z _6072_/B _6073_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5023_ _5019_/Z _5020_/Z _5023_/A3 _5285_/B _5023_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet852_140 net802_76/I _7085_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_151 _4073__37/I _7074_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6974_ _6974_/D _6967_/RN _6974_/CLK _6974_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_53_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5925_ _5991_/A2 _5914_/S _7230_/Q _3389_/I _5925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_80_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5856_ _5892_/I0 hold701/Z _5856_/S _5856_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4807_ _5173_/A2 _4534_/Z _5312_/A1 _5414_/A2 _4807_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_166_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5787_ _5886_/I0 _5787_/I1 _5793_/S _5787_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4738_ _5403_/A1 _5309_/A2 _4738_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_108_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4669_ _4397_/Z _5209_/A3 _4889_/A1 _5464_/A1 _4669_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6408_ _6408_/A1 _6408_/A2 _6408_/A3 _6408_/A4 _6408_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold940 _5694_/Z _7045_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_150_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold951 _6719_/Q hold951/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_122_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold962 _5786_/Z _7126_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold973 _6979_/Q hold973/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold984 _5576_/Z _6940_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6339_ _7252_/Q _6339_/I1 _6450_/S _7252_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold995 _7159_/Q hold995/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_131_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3971_ _3971_/A1 _3434_/B _6663_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_62_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5710_ _5776_/A1 _5767_/A3 _5866_/A3 _5718_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_189_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6690_ _6690_/D _7170_/RN _6690_/CLK _6690_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_149_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5641_ hold855/Z _5806_/I0 _5646_/S _5641_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5572_ _5818_/I0 hold542/Z _5574_/S _5572_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4523_ _5458_/A4 _4752_/A2 _5139_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold203 _7131_/Q hold203/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_156_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold214 _5524_/Z _6897_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7242_ _7242_/D _7247_/RN _7258_/CLK _7242_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold225 _5545_/Z _6913_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold236 _7192_/Q hold236/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4454_ _5426_/A1 _4836_/A3 _4454_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_132_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold247 _4260_/Z _6775_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold258 hold258/I hold258/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold269 _6881_/Q hold269/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3405_ _4472_/B _4441_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_7173_ _7173_/D _7173_/RN _7173_/CLK _7173_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout705 _7237_/RN _7075_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_4385_ input99/Z input98/Z _4386_/A3 _4386_/A4 _4385_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xfanout716 _7279_/RN _7278_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6124_ _6124_/A1 _6124_/A2 _6124_/A3 _6124_/A4 _6124_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout727 _4549_/A4 _4440_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3336_ _7209_/Q _4050_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout738 input120/Z _4589_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout749 _4836_/A3 _4878_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6055_ _7014_/Q _5971_/Z _5979_/Z _6966_/Q _5996_/Z hold84/I _6057_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5006_ _5389_/C _5170_/A2 _5170_/A3 _5130_/B2 _5347_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xclkbuf_leaf_121__1359_ net952_221/I net802_82/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_41__1359_ clkbuf_4_11_0__1359_/Z _4073__28/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6957_ _6957_/D fanout655/Z _6957_/CLK _6957_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_121_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5908_ _7223_/Q _7224_/Q _7225_/Q _5908_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6888_ hold41/Z _7296_/RN _6888_/CLK _6888_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_14_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5839_ _5884_/A3 _5839_/A2 _5839_/A3 _5857_/A3 _5847_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_139_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold770 _5610_/Z _6971_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold781 _7091_/Q hold781/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold792 _4106_/Z _6667_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_150_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput308 _7308_/Z spimemio_flash_io2_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_154_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput319 _6792_/Q wb_dat_o[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4170_ _4170_/A1 _5647_/A2 _4172_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_110_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6811_ _6811_/D _7262_/CLK _6811_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6742_ _6742_/D _7194_/RN _6742_/CLK _6742_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_189_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3954_ _6988_/Q _3954_/A2 _3954_/B1 input20/Z _4301_/A1 _6809_/Q _3958_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_50_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6673_ hold69/Z fanout659/Z _6673_/CLK hold68/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_176_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3885_ _3876_/Z _3885_/A2 _3885_/A3 _3884_/Z _3885_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5624_ hold60/Z _5624_/I1 _5628_/S hold61/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5555_ _5555_/I0 hold331/Z _5556_/S _5555_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4506_ _4997_/B _4494_/Z _4496_/Z _5263_/A2 _4506_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5486_ _4616_/Z _4855_/C _5487_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_133_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7225_ _7225_/D _7225_/RN _4067_/I1 _7225_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_132_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4437_ _4438_/B _4438_/C _4648_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xfanout502 _5836_/I0 _5881_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout513 hold19/Z _5880_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout524 hold2/Z _5842_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7156_ _7156_/D _7221_/RN _7156_/CLK _7156_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4368_ _4456_/B _4456_/C _4455_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xfanout535 _5877_/I0 _5796_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout546 _4180_/I0 _5867_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_141_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6107_ _7064_/Q _5985_/Z _5997_/Z _7098_/Q hold22/I _6006_/Z _6109_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xfanout557 _3385_/ZN _6210_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_100_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout568 _7231_/Q _6068_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3319_ _7223_/Q _5900_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7087_ _7087_/D fanout656/Z _7087_/CLK _7087_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xfanout579 _3315_/I _6600_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4299_ _6570_/I0 _6807_/Q _4300_/S _6807_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6038_ _6031_/Z _6037_/Z _6336_/B1 _6118_/B _6555_/C _6039_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_55_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1152_404 net1152_434/I _6770_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_415 net1152_415/I _6759_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_426 net952_251/I _6748_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_437 net1152_437/I _6728_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_151_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1152_448 net1202_474/I _6717_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3670_ hold42/I _3927_/A2 _3952_/A2 _7049_/Q _3673_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_173_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5340_ _5340_/A1 _5370_/B _5340_/B _5340_/C _5363_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_115_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5271_ _5165_/Z _5270_/Z _4877_/Z _5271_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_130_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7010_ _7010_/D _7125_/RN _7010_/CLK _7010_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4222_ _4221_/Z hold197/Z _4228_/S _4222_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4153_ _5852_/I0 hold611/Z _4157_/S _4153_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4084_ _4084_/I0 _4084_/I1 _6732_/Q _7281_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4986_ _4986_/A1 _4980_/Z _4986_/A3 _4993_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3937_ _3937_/A1 _3937_/A2 _3937_/A3 _3903_/Z _3937_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6725_ _6725_/D _6854_/RN _6725_/CLK _6725_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_51_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6656_ _6656_/A1 _6656_/A2 _6656_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3868_ _3868_/A1 _3868_/A2 _3868_/A3 _3868_/A4 _3868_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_20_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5607_ _5781_/I0 hold503/Z _5610_/S _5607_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6587_ _6587_/I0 _7272_/Q _6602_/S _7272_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3799_ _3798_/Z _3799_/I1 _3899_/S _6870_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5538_ hold777/Z _5538_/I1 _5538_/S _5538_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5469_ _5469_/A1 _5423_/Z _5469_/A3 _5469_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_121_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7208_ hold3/Z _7220_/RN _7208_/CLK _7208_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout343 _6499_/A1 _6554_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7139_ _7139_/D _7141_/RN _7139_/CLK _7139_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout354 _3541_/ZN _4210_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_101_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet1102_356 net1152_410/I _6854_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout365 _5794_/A2 _5821_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet1102_367 net1152_441/I _6843_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout376 _3527_/Z _5510_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet1102_378 net1102_379/I _6821_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout387 hold152/Z _5857_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_19_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout398 _6265_/Z _6549_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xnet1102_389 net1152_430/I _6785_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput18 mask_rev_in[22] input18/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput29 mask_rev_in[3] input29/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4840_ _5281_/B _5132_/A2 _4840_/B1 _5214_/A2 _4841_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_2580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4771_ _4944_/A1 _4463_/Z _4782_/A1 _5307_/A3 _5236_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_1890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6510_ _6841_/Q _6549_/B1 _6288_/Z _7296_/Q _6511_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_159_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3722_ hold80/I _3909_/A2 _3948_/C1 _7308_/I _4225_/S _4075_/I1 _3723_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_119_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6441_ _6985_/Q _6550_/B1 _6273_/Z _6977_/Q _6549_/C1 _7001_/Q _6442_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3653_ _3653_/A1 _3492_/Z _3680_/A3 _3500_/Z _3653_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6372_ _7169_/Q _5948_/Z _6544_/B1 hold88/I _6545_/B1 _7015_/Q _6385_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3584_ _7197_/Q _3909_/A2 _4225_/S input70/Z _4194_/A1 input60/Z _3589_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_173_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5323_ _5323_/A1 _4920_/Z _5322_/Z _5323_/B _5324_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_5254_ _4761_/I _5245_/Z _5254_/B _5254_/C _5257_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_130_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4205_ _4204_/Z hold305/Z _4211_/S _4205_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5185_ _5185_/A1 _5185_/A2 _6577_/C _5185_/B2 _6860_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_68_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4136_ hold6/Z hold70/Z _4136_/S hold71/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4067_ _6761_/Q _4067_/I1 _6903_/Q _4067_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4969_ _4718_/B _4903_/Z _4973_/A4 _5010_/A1 _4969_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6708_ _6708_/D _6856_/RN _6708_/CLK _6708_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_132_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ _6650_/A1 _6650_/A2 _6639_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_137_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_18__1359_ net1152_430/I net902_189/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_10_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6990_ _6990_/D _7141_/RN _6990_/CLK _6990_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_66_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5941_ _5941_/A1 _5940_/Z _5943_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5872_ _5890_/I0 hold584/Z _5874_/S _5872_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4823_ _5270_/A1 _5269_/A1 _4889_/A1 _4554_/Z _4659_/Z _4826_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_21_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1002_300 net902_157/I _6925_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4754_ _5226_/A1 _4752_/Z _5233_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_144_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3705_ _6960_/Q _3957_/A2 _3959_/B1 _6670_/Q _3707_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_119_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4685_ _4685_/A1 _4685_/A2 _5180_/A3 _5211_/C _5001_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_146_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6424_ _7171_/Q _6544_/A2 _6545_/A2 _6937_/Q _6425_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3636_ _7196_/Q _3909_/A2 _4227_/S input69/Z _3945_/B1 _7092_/Q _3638_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_162_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6355_ _6355_/A1 _6355_/A2 _6355_/A3 _6355_/A4 _6355_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3567_ _3512_/Z _5692_/A1 _5683_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_115_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5306_ _5306_/I _5307_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6286_ _6287_/A1 _6287_/A2 _6287_/A3 _6286_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_102_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3498_ _3498_/I0 _4056_/I1 _3984_/S _3499_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5237_ _5238_/A1 _5238_/A4 _5457_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_111_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5168_ _5270_/A2 _4997_/C _4820_/Z _5420_/A4 _5425_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_111_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4119_ _5520_/C _5517_/A2 _5629_/A3 _5785_/A3 _4127_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_17_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5099_ _5099_/A1 _5099_/A2 _5226_/A1 _5228_/A3 _4549_/Z _5100_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_95_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_1_1__f__1062_ clkbuf_0__1062_/Z _6568_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_116_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold7 hold7/I hold7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_59_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_5__1359_ net1152_451/I net1152_437/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_48_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4470_ _4463_/Z _4468_/Z _4765_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold407 _5715_/Z _7064_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold418 _7125_/Q hold418/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_7_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold429 _5797_/Z _7136_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_99_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3421_ _3421_/A1 _3421_/A2 _7304_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_171_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6140_ _7026_/Q _6164_/A2 _6164_/B1 _6994_/Q _6141_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3352_ _7137_/Q _3352_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_171_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6071_ _7153_/Q _5960_/Z _5965_/Z _6701_/Q _5981_/Z _6935_/Q _6073_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_opt_4_0__1359_ _4073__24/I clkbuf_opt_4_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_135_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5022_ _5198_/C _5023_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet852_130 _4073__35/I _7095_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_141 _4073__9/I _7084_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6973_ _6973_/D _7207_/RN _6973_/CLK _6973_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_53_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5924_ _6021_/A2 _6015_/A3 _6014_/A2 _5984_/A1 _5924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_181_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5855_ _5855_/I0 hold717/Z _5856_/S _5855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4806_ _4492_/Z _4536_/Z _5319_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_142_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5786_ _5867_/I0 hold961/Z _5793_/S _5786_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4737_ _5226_/C _5226_/B _5309_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_175_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_64__1359_ clkbuf_4_13_0__1359_/Z net952_218/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_135_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4668_ _4411_/Z _5343_/A1 _5393_/A2 _5165_/A4 _5360_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xclkbuf_leaf_144__1359_ net1152_451/I net1202_452/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_119_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6407_ _7072_/Q _6248_/Z _6293_/Z hold24/I _6407_/C _6408_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3619_ _7260_/Q _6899_/Q _6900_/Q _3619_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold930 _5585_/Z _6948_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold941 _6809_/Q hold941/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4599_ _5129_/A3 _4598_/Z _4873_/A2 _5269_/A1 _4599_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold952 _4178_/Z _6719_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold963 _6956_/Q hold963/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold974 _5619_/Z _6979_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6338_ _6338_/I _6339_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold985 _6957_/Q hold985/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold996 _5823_/Z _7159_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_135_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6269_ _3328_/I _6300_/A1 _6302_/A3 _6275_/A4 _6269_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_48_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3970_ _3967_/Z _3970_/A2 _6664_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_189_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5640_ hold598/Z _5877_/I0 _5646_/S _5640_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5571_ _5871_/I0 hold402/Z _5574_/S _5571_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4522_ _5365_/A3 _4522_/A2 _5164_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_157_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold204 _5791_/Z _7131_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_172_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold215 _6900_/Q hold215/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_102_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7241_ _7241_/D _7258_/RN _7258_/CLK _7241_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold226 _6924_/Q hold226/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4453_ _5129_/A4 _3402_/I _4555_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold237 _5860_/Z _7192_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold248 _7031_/Q hold248/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_172_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold259 _5515_/Z _5516_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3404_ _3404_/I _3404_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7172_ _7172_/D _7173_/RN _7172_/CLK _7172_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_125_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4384_ _4376_/Z _4381_/Z _4580_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_98_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout706 _7071_/RN _7237_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6123_ _7147_/Q _5987_/Z _6015_/Z _7009_/Q _6124_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout717 _7279_/RN _7261_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_3335_ _7217_/Q _4049_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout728 _3408_/I _4652_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout739 _3404_/I _4873_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6054_ _6934_/Q _5981_/Z _5988_/Z _6982_/Q _7046_/Q _6019_/Z _6057_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_61_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ _5043_/A2 _5389_/C _5393_/B1 _5043_/B _5347_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_22_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3340__1 _3340__1/I _6603_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6956_ _6956_/D _7140_/RN _6956_/CLK _6956_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_41_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5907_ _5906_/Z _5904_/B _7225_/Q _7225_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6887_ _6887_/D _6886_/RN _6887_/CLK _6887_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_139_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5838_ _5865_/I0 hold607/Z _5838_/S _5838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5769_ _5886_/I0 hold981/Z _5775_/S _5769_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold760 _5627_/Z _6986_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold771 _7099_/Q hold771/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_150_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold782 _5746_/Z _7091_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold793 _6683_/Q hold793/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet802_90 net802_90/I _7135_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput309 _7309_/Z spimemio_flash_io3_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_5_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6810_ _6810_/D _6847_/RN _6810_/CLK _6810_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6741_ _6741_/D _7194_/RN _6741_/CLK _6741_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3953_ _3953_/A1 _3953_/A2 _3953_/A3 _3953_/A4 _3953_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_177_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6672_ hold49/Z fanout659/Z _6672_/CLK hold48/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3884_ _3884_/A1 _3884_/A2 _3884_/A3 _3884_/A4 _3884_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_137_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5623_ _5806_/I0 hold937/Z _5628_/S _5623_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5554_ _5890_/I0 hold377/Z _5556_/S _5554_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4505_ _5340_/A1 _4982_/A2 _4497_/Z _5262_/A2 _5343_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5485_ _5480_/Z _5485_/A2 _5485_/B _5490_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_117_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7224_ _7224_/D _7224_/RN _4067_/I1 _7224_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4436_ _4652_/A4 _5201_/A1 _4436_/B _4438_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_99_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout503 _5836_/I0 _5827_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7155_ _7155_/D _7155_/RN _7155_/CLK _7155_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout514 _5834_/I0 _5798_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_4367_ _4456_/B _4456_/C _4367_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
Xfanout525 hold2/Z _5860_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_59_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout536 _5850_/I0 _5877_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_86_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout547 hold64/Z _4180_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6106_ _6106_/A1 _6106_/A2 _6106_/A3 _6106_/A4 _6106_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3318_ _6743_/Q _5945_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_7086_ _7086_/D _7098_/RN _7086_/CLK _7086_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_86_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout558 _3385_/ZN _6139_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4298_ _6569_/I0 _6806_/Q _4300_/S _6806_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout569 _7229_/Q _3389_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6037_ _6037_/A1 _6037_/A2 _6037_/A3 _6037_/A4 _6037_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_132_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6939_ _6939_/D _7149_/RN _6939_/CLK _6939_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XPHY_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1152_405 net1152_435/I _6769_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1152_416 net1152_416/I _6758_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_151_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1152_427 net1152_427/I _6747_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_438 net802_71/I _6727_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_449 net1202_468/I _6716_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold590 _6842_/Q hold590/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_110_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5270_ _5270_/A1 _5270_/A2 _4997_/C _4820_/Z _5270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4221_ hold187/Z _5781_/I0 _4227_/S _4221_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4152_ _5869_/I0 hold925/Z _4157_/S _4152_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4083_ _6734_/Q _6731_/Q _4084_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_64_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4985_ _4397_/Z _5209_/A3 _4659_/Z _5415_/A1 _4985_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_168_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6724_ _6724_/D _6854_/RN _6724_/CLK _6724_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_189_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3936_ _7028_/Q _5674_/A1 _3936_/B1 _6690_/Q _3937_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_177_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6655_ _6656_/A1 _6657_/A2 _6655_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3867_ _7079_/Q _3923_/C1 _3956_/B1 _6713_/Q _3867_/C _3868_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_20_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5606_ _5798_/I0 hold637/Z _5610_/S _5606_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6586_ _6586_/A1 _6601_/A2 _6586_/B _6587_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_3798_ _6566_/I0 _6869_/Q _3898_/S _3798_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5537_ hold795/Z _5537_/I1 _5538_/S _5537_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5468_ _5468_/A1 _5468_/A2 _5468_/B1 _4650_/Z _5468_/C _5469_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_133_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7207_ _7207_/D _7207_/RN _7207_/CLK _7207_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4419_ _4960_/A1 _5055_/A2 _4589_/A4 _4419_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_5399_ _5399_/A1 _5399_/A2 _5478_/A2 _5302_/B _5399_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_99_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7138_ _7138_/D _7140_/RN _7138_/CLK _7138_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout344 _6450_/S _6558_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_87_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout355 _3541_/ZN _4202_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout366 _5794_/A2 _5839_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet1102_357 net1152_410/I _6853_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1102_368 net1152_421/I _6842_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout377 hold145/Z hold146/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xnet1102_379 net1102_379/I _6820_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout388 _5875_/A1 _5857_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_28_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7069_ _7069_/D _7098_/RN _7069_/CLK _7069_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xfanout399 _6262_/Z _6531_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_98_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput19 mask_rev_in[23] input19/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ _4770_/A1 _5118_/A3 _4770_/A3 _5117_/A1 _4775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_1880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3721_ _6678_/Q _3546_/Z _3916_/A2 hold24/I hold22/I _3941_/B1 _3723_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_158_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6440_ _6440_/A1 _6440_/A2 _6440_/A3 _6439_/Z _6440_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3652_ input68/Z _4227_/S _4244_/S input40/Z _3657_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_61_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3583_ _6971_/Q _3924_/A2 _3607_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6371_ _7063_/Q _6257_/Z _6299_/Z _7055_/Q _6383_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_155_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5322_ _5322_/A1 _4494_/Z _5328_/A2 _5442_/A1 _5322_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_142_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5253_ _5254_/C _5334_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4204_ hold98/Z _5889_/I0 _4210_/S _4204_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5184_ _3315_/I _5182_/Z _5184_/B _5184_/C _5185_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_69_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4135_ _5645_/I1 hold313/Z _4136_/S _4135_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4066_ _6762_/Q user_clock _6904_/Q _4066_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4968_ _4903_/Z _4973_/A4 _4718_/B _4666_/Z _4968_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6707_ _6707_/D _6786_/RN _6707_/CLK _6707_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_149_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3919_ _3919_/A1 _3919_/A2 _3919_/A3 _3919_/A4 _3919_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_138_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4899_ _6577_/C _4899_/A2 _5000_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_137_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6638_ _6644_/A1 _6650_/A2 _6638_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_118_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6569_ _6569_/I0 _7267_/Q _6571_/S _7267_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4073__2 _4073__3/I _7297_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5940_ _4009_/B _7233_/Q _7232_/Q _3329_/I _5940_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_81_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5871_ _5871_/I0 hold507/Z _5874_/S _5871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4822_ _4554_/Z _4659_/Z _4820_/Z _5278_/B _4826_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_33_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1002_301 net1152_414/I _6924_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_178_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4753_ _5478_/B1 _4752_/Z _5313_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_30_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3704_ _7138_/Q _3951_/A2 _3901_/A2 _6984_/Q input30/Z _3927_/C2 _3707_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_174_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4684_ _4414_/Z _4452_/Z _4666_/Z _4892_/B _5287_/A2 _4685_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_175_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6423_ _7099_/Q _6250_/Z _6439_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_88_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3635_ input50/Z _4202_/S _3947_/A2 _7100_/Q _3638_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_128_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6354_ _7168_/Q _6544_/A2 _6261_/Z _6958_/Q _6355_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3566_ _3507_/Z _5517_/A2 _3954_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5305_ _5367_/A2 _4673_/Z _5307_/A3 _5305_/B _5306_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_88_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3497_ _3497_/I hold144/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
X_6285_ _6452_/A2 _6285_/A2 _7237_/Q _6452_/A4 _6285_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_130_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5236_ _5236_/A1 _5414_/A2 _5236_/B _5238_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_102_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5167_ _4546_/Z _4651_/Z _5380_/B2 _5167_/B _5425_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_84_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4118_ hold6/Z hold68/Z _4118_/S hold69/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5098_ _5098_/A1 _5302_/B _5098_/B _5098_/C _5101_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_84_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_104__1359_ clkbuf_4_7_0__1359_/Z net802_54/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4049_ _4049_/I0 input92/Z _4050_/S _4049_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_87__1359_ clkbuf_4_7_0__1359_/Z net902_179/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold8 hold8/I hold8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_74_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold408 _6761_/Q hold408/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold419 _5784_/Z _7125_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3420_ _3988_/S _3422_/I0 _3421_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_125_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3351_ _7145_/Q _3351_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6070_ _6951_/Q _5958_/Z _5967_/Z _7105_/Q _7137_/Q _5994_/I _6073_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5021_ _4604_/Z _4606_/Z _5003_/Z _5021_/B _5198_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_79_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet852_120 net852_120/I _7105_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet852_131 net852_131/I _7094_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_142 net902_168/I _7083_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6972_ _6972_/D _7098_/RN _6972_/CLK _6972_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_80_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5923_ _7230_/Q _3389_/I _6210_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_62_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5854_ _5881_/I0 hold683/Z _5856_/S _5854_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4805_ _4835_/A2 _4492_/Z _4534_/Z _4681_/Z _4805_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_179_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5785_ _5866_/A3 _5839_/A2 _5785_/A3 _5857_/A2 _5793_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4736_ _4736_/A1 _5307_/A3 _4736_/A3 _4467_/B _5226_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_119_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4667_ _4414_/Z _5038_/A1 _4557_/Z _5475_/A4 _4667_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_162_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6406_ _6406_/I _6407_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold920 _5732_/Z _7078_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3618_ _5510_/A2 _3617_/Z _5528_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold931 _6941_/Q hold931/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4598_ _5287_/B _4460_/B _5399_/A2 _4752_/A2 _4598_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold942 _4302_/Z _6809_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold953 _6699_/Q hold953/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold964 _5594_/Z _6956_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6337_ _6500_/C _7251_/Q _6337_/B _6338_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold975 _6972_/Q hold975/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3549_ hold258/I _3512_/Z _4194_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold986 _5595_/Z _6957_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold997 _6854_/Q hold997/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_131_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6268_ _7233_/Q _7232_/Q _6533_/A2 _6452_/A4 _6268_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_103_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5219_ _5303_/A1 _5303_/A3 _5224_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_29_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6199_ _6789_/Q _5972_/Z _6021_/Z _6839_/Q _6201_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_28_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_70__1359_ clkbuf_4_15_0__1359_/Z net802_76/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_44_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5570_ _5888_/I0 hold533/Z _5574_/S _5570_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4521_ _4440_/B _4449_/B _5139_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_156_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold205 _6774_/Q hold205/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7240_ _7240_/D _7240_/RN _4067_/I1 _7240_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold216 _5527_/Z _6900_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_171_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4452_ _5038_/A1 _4648_/B _4638_/A2 _4452_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
Xhold227 _5558_/Z _6924_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold238 _7169_/Q hold238/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold249 _5678_/Z _7031_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3403_ _3403_/I _3403_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7171_ _7171_/D _7171_/RN _7171_/CLK _7171_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_171_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4383_ _5201_/A1 _4383_/A2 _5385_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6122_ _7091_/Q _6002_/Z _6003_/Z _7163_/Q _6124_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout707 _7240_/RN _7225_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout718 _6865_/RN _7279_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3334_ _3334_/I _4029_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout729 _3408_/I _4436_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ _6053_/A1 _6053_/A2 _6053_/A3 _6053_/A4 _6053_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_85_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5004_ _5368_/A1 _5420_/A1 _5002_/Z _5389_/B _5191_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_85_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6955_ hold35/Z _7002_/RN _6955_/CLK _6955_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5906_ _7223_/Q _7224_/Q _5910_/B _5906_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6886_ _6886_/D _6886_/RN _6886_/CLK _6886_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_34_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5837_ _5837_/I0 hold837/Z _5838_/S _5837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5768_ _5867_/I0 hold993/Z _5775_/S _5768_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4719_ _5083_/B _4719_/A2 _4721_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_107_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5699_ _5837_/I0 hold592/Z _5700_/S _5699_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold750 _5852_/Z _7185_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold761 _6962_/Q hold761/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_1_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold772 _5755_/Z _7099_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold783 _7076_/Q hold783/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold794 _4130_/Z _6683_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_118_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet802_80 _4073__4/I _7145_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet802_91 net802_91/I _7134_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6740_ _6740_/D _7194_/RN _6740_/CLK _6740_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3952_ _7044_/Q _3952_/A2 _5638_/A1 _6996_/Q _6948_/Q _5584_/A1 _3953_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_51_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6671_ _6671_/D fanout659/Z _6671_/CLK _6671_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_149_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3883_ input53/Z _4194_/A1 _3948_/C1 input62/Z _3941_/B1 _7167_/Q _3884_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_91_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5622_ _5796_/I0 hold739/Z _5628_/S _5622_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5553_ _5880_/I0 hold160/Z _5556_/S _5553_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ _4759_/A2 _4759_/A3 _4504_/B _4504_/C _5263_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_144_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5484_ _5483_/Z _5450_/I _5477_/Z _5441_/B _5485_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_6_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7223_ _7223_/D _7225_/RN _4067_/I1 _7223_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4435_ _4652_/A4 _4455_/A2 _5170_/A2 _4436_/B _4438_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_132_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7154_ hold25/Z _7154_/RN _7154_/CLK hold24/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout504 hold40/Z _5836_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout515 hold60/Z _5834_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_98_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4366_ _4440_/B _3407_/I _4652_/A1 _4501_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xfanout526 _4343_/I0 _5538_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6105_ _7114_/Q _5984_/Z _6000_/Z _7130_/Q _6106_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xfanout537 hold54/Z _5850_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_98_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout548 _5876_/I0 _5795_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_141_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3317_ _3317_/I _4686_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_7085_ _7085_/D _7149_/RN _7085_/CLK _7085_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_112_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout559 _6253_/A4 _6302_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_140_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4297_ _4297_/I0 _6805_/Q _4300_/S _6805_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _6973_/Q _5964_/Z _5984_/Z _7111_/Q _6036_/C _6037_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_55_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6938_ _6938_/D _7173_/RN _6938_/CLK _6938_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XPHY_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6869_ _6869_/D _6627_/Z _4075_/I1 _6869_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_22_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1152_406 net1152_409/I _6768_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_157_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet1152_417 net1152_419/I _6757_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_428 net1152_431/I _6742_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_439 net802_71/I _6726_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold580 _5779_/Z _7120_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold591 _4337_/Z _6842_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4220_ _4219_/Z hold199/Z _4228_/S _4220_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4151_ _5796_/I0 hold953/Z _4157_/S _4151_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4082_ _4082_/A1 _7299_/Q _4082_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_110_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4984_ _5260_/A1 _4982_/Z _4984_/B _4986_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6723_ _6723_/D _7170_/RN _6723_/CLK _6723_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3935_ _6924_/Q _3935_/A2 _3935_/B1 _6849_/Q _3937_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_189_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6654_ _7225_/RN _6656_/A2 _6654_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3866_ _3866_/A1 _5731_/A2 _3617_/Z _3866_/B _3867_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_137_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5605_ _5797_/I0 _5605_/I1 _5610_/S _5605_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6585_ _6600_/A1 _6585_/A2 _6585_/B1 _3316_/I _3317_/I _6585_/C2 _6586_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3797_ _3776_/Z _3797_/A2 _3797_/A3 _3796_/Z _6566_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_118_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5536_ _5536_/A1 _6611_/A2 _5538_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_127_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5467_ _4570_/Z _4651_/Z _5467_/B _5467_/C _5468_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_117_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7206_ _7206_/D _6821_/RN _7206_/CLK _7206_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_133_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4418_ _5170_/A2 _4456_/B _5343_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_114_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5398_ _5391_/Z _5398_/A2 _5419_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7137_ _7137_/D _7146_/RN _7137_/CLK _7137_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4349_ _5832_/I0 hold629/Z _4349_/S _4349_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout345 _6476_/S _6450_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout356 _4225_/S _4227_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xnet1102_358 net802_75/I _6852_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout367 _5794_/A2 _3732_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xnet1102_369 net1152_421/I _6841_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout378 hold145/Z _4347_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7068_ _7068_/D _7098_/RN _7068_/CLK _7068_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xfanout389 _5875_/A1 _5884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_115_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6019_ _3386_/I _3387_/I _6164_/A2 _6210_/A2 _6019_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_100_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3720_ _7114_/Q _3917_/A2 _3947_/A2 _7098_/Q _3945_/A2 _7178_/Q _3723_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_187_963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3651_ _7187_/Q _3959_/C1 _3960_/A2 _7211_/Q _3657_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6370_ _6991_/Q _6237_/Z _6380_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xnet902_200 net952_250/I _7025_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3582_ _5611_/A1 _5884_/A2 _3924_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_54_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5321_ _5321_/A1 _5212_/Z _5454_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_154_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5252_ _5343_/A1 _5343_/A2 _5255_/A2 _5252_/B _5254_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_170_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4203_ _4202_/Z hold410/Z _4211_/S _4203_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5183_ _5181_/Z _4686_/B _5299_/C _5184_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_111_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4134_ hold40/Z hold50/Z _4136_/S hold51/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4065_ _6392_/B1 input2/Z input1/Z _4065_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4967_ _4903_/Z _4973_/A4 _4718_/B _5359_/A1 _4967_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3918_ input36/Z _4225_/S _4143_/A1 _6694_/Q _3919_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6706_ _6706_/D _7162_/RN _6706_/CLK _6706_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_149_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4898_ _5097_/B2 _4893_/Z _4898_/B _4898_/C _4899_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_164_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6637_ _6771_/RN _6648_/A2 _6637_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3849_ _7175_/Q _3945_/A2 _3939_/C1 _6711_/Q _3897_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_165_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6568_ _6568_/I0 _7266_/Q _6571_/S _7266_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_47__1359_ clkbuf_4_14_0__1359_/Z _4073__37/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_127__1359_ clkbuf_4_4_0__1359_/Z net852_147/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5519_ _6894_/Q hold222/Z _5520_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_146_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6499_ _6499_/A1 _6499_/A2 _6499_/A3 _6498_/Z _6499_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_87_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4073__3 _4073__3/I _7296_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_7_0__1359_ clkbuf_0__1359_/Z clkbuf_4_7_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_11_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5870_ hold60/Z hold301/Z _5874_/S _5870_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4821_ _5290_/A2 _5295_/A3 _4887_/A1 _5295_/A2 _4821_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_61_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4752_ _5315_/A4 _4752_/A2 _4463_/Z _5226_/C _4752_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_187_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3703_ input48/Z _4210_/S _4244_/S input39/Z _3708_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_147_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4683_ _5420_/A3 _4715_/A1 _3403_/I _4878_/A4 _4683_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6422_ _7065_/Q _6257_/Z _6434_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_174_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3634_ _7220_/Q _3912_/A2 _4242_/S input41/Z _3930_/A2 _7132_/Q _3638_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_162_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6353_ _7208_/Q _6535_/A2 _6285_/Z _7192_/Q _6543_/A2 hold36/I _6355_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_162_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3565_ _5611_/A1 _5830_/A1 _3901_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_108_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5304_ _5478_/A2 _5478_/A3 _5456_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_89_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6284_ _6281_/Z _6283_/Z _6550_/B1 _6273_/Z _6287_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3496_ _3495_/Z hold142/Z _3500_/S _3496_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5235_ _5316_/A2 _5234_/Z _5238_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_25_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5166_ _5166_/A1 _5467_/B _5166_/A3 _5165_/Z _5169_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_25_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4117_ hold4/Z _7277_/Q _4117_/S hold5/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5097_ _5097_/A1 _5328_/A2 _5368_/B _5097_/B2 _5098_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4048_ _6767_/Q input89/Z _4050_/S _4048_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5999_ _6211_/A2 _6021_/A2 _6210_/A2 _3387_/I _5999_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XPHY_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput290 _6685_/Q pll_trim[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_58_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold9 hold9/I hold9/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_101_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold409 _4243_/Z _6761_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_87_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_110__1359_ clkbuf_4_4_0__1359_/Z net802_91/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_30__1359_ clkbuf_opt_4_0__1359_/Z net1052_315/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3350_ _7153_/Q _3350_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_93__1359_ clkbuf_4_5_0__1359_/Z net952_225/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5020_ _5438_/C _5020_/A2 _4604_/Z _4606_/Z _5020_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet852_110 net952_234/I _7115_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet852_121 net802_62/I _7104_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet852_132 net802_52/I _7093_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_143 net802_89/I _7082_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6971_ _6971_/D _7124_/RN _6971_/CLK _6971_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_93_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5922_ _5922_/I _7229_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5853_ _5880_/I0 hold122/Z _5856_/S _5853_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4804_ _4681_/Z _4793_/Z _5319_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5784_ _5784_/I0 hold418/Z _5784_/S _5784_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4735_ _3406_/I _4735_/A2 _4764_/A3 _5226_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_119_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4666_ _4960_/A1 _5420_/A2 _4835_/A2 _3403_/I _4666_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_163_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6405_ _7138_/Q _6253_/Z _6297_/Z _6702_/Q _6406_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_135_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3617_ hold144/I _3500_/Z hold221/I _3492_/Z _3617_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold910 _5569_/Z _6934_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold921 _7134_/Q hold921/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4597_ _5369_/A1 _4596_/Z _5420_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold932 _5577_/Z _6941_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold943 _7096_/Q hold943/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold954 _4151_/Z _6699_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6336_ _6329_/Z _6335_/Z _6336_/B1 _6286_/Z _6555_/C _6337_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3548_ _3519_/Z _3932_/A2 _3945_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold965 _6710_/Q hold965/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_1_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold976 _5612_/Z _6972_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold987 _7184_/Q hold987/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold998 _4355_/Z _6854_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_88_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6267_ _6996_/Q _6549_/C1 _6545_/B1 _7012_/Q _6271_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_130_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3479_ _6659_/Q _6658_/Q _3984_/S _3479_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5218_ _4673_/Z _5478_/B1 _5218_/B _5303_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6198_ _6198_/A1 _6198_/A2 _6198_/A3 _6198_/A4 _6198_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_97_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5149_ _5165_/A2 _4598_/Z _5374_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_28_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4520_ _4835_/A2 _3403_/I _3402_/I _5097_/B2 _5093_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_129_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold206 _4259_/Z _6774_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_172_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4451_ _4604_/A2 _4604_/A3 _4451_/B _4451_/C _5038_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xhold217 _6898_/Q hold217/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_7_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold228 _6768_/Q hold228/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold239 _5834_/Z _7169_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3402_ _3402_/I _3402_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7170_ hold23/Z _7170_/RN _7170_/CLK hold22/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_144_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4382_ _4440_/B _4501_/B _5458_/A4 _4436_/B _4383_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6121_ _6985_/Q _5988_/Z _6019_/Z _7049_/Q _6124_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_4_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout708 _7071_/RN _7240_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_3333_ _4395_/B _4424_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
Xfanout719 _6563_/A2 _6865_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6052_ _6950_/Q _5958_/Z _5967_/Z _7104_/Q _6052_/C _6053_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _5165_/A4 _5003_/A2 _5010_/A1 _4491_/B _5003_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_0__1062_ _3725_/ZN clkbuf_0__1062_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_61_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6954_ _6954_/D _7141_/RN _6954_/CLK _6954_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_53_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5905_ _5905_/I _7224_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6885_ _6885_/D _7296_/RN _6885_/CLK _6885_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_179_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5836_ _5836_/I0 hold317/Z _5838_/S _5836_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5767_ _5785_/A3 _5839_/A3 _5767_/A3 _5866_/A3 _5775_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_108_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4718_ _4504_/B _4504_/C _4718_/B _5056_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5698_ _5782_/I0 hold513/Z _5700_/S _5698_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4649_ _4570_/Z _5438_/B _4653_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_162_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold740 _5622_/Z _6981_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold751 _6788_/Q hold751/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold762 _5600_/Z _6962_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold773 _7133_/Q hold773/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold784 _5729_/Z _7076_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6319_ _7127_/Q _6402_/A2 _6533_/A3 _7111_/Q _6320_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold795 _6906_/Q hold795/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_131_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7299_ _7299_/D _6651_/Z _7302_/CLK _7299_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_103_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet802_70 net802_87/I _7155_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet802_81 net802_81/I _7144_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet802_92 net802_94/I _7133_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3951_ _7134_/Q _3951_/A2 _5665_/A1 _7020_/Q _3951_/C1 _7142_/Q _3953_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_50_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6670_ _6670_/D fanout659/Z _6670_/CLK _6670_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3882_ _6925_/Q _3935_/A2 _3933_/B1 _6786_/Q _3942_/C1 _6854_/Q _3884_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_32_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ _5804_/I0 hold723/Z _5628_/S _5621_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5552_ _5879_/I0 hold359/Z _5556_/S _5552_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4503_ _4718_/B _4973_/A4 _5262_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5483_ _5483_/A1 _5483_/A2 _5483_/A3 _5483_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_4434_ _4467_/B _4460_/B _4887_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7222_ _7222_/D _7240_/RN _4067_/I1 _7222_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_160_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7153_ _7153_/D _7219_/RN _7153_/CLK _7153_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4365_ _4440_/B _3407_/I _4652_/A1 _5288_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_113_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout505 hold40/Z _5890_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout516 hold60/Z _5888_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6104_ _7106_/Q _5967_/Z _5980_/Z _7072_/Q _5969_/Z _7122_/Q _6106_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xfanout527 _4343_/I0 _4361_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_112_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout538 hold53/Z hold54/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3316_ _3316_/I _4415_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_7084_ _7084_/D _7173_/RN _7084_/CLK _7084_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout549 _5876_/I0 _5804_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4296_ _6567_/I0 _6804_/Q _4300_/S _6804_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6035_ _6035_/I _6036_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6937_ _6937_/D _7141_/RN _6937_/CLK _6937_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XPHY_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_179_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6868_ _6868_/D _6626_/Z _4075_/I1 _6868_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_50_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5819_ _5891_/I0 hold917/Z _5820_/S _5819_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6799_ _6799_/D _6847_/RN _6799_/CLK _6799_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_109_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1152_407 net1152_409/I _6767_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_418 net902_194/I _6756_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_429 net1152_431/I _6741_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold570 _4322_/Z _6821_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold581 _7137_/Q hold581/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold592 _7050_/Q hold592/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_77_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150_ _5804_/I0 hold903/Z _4157_/S _4150_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4081_ _4081_/A1 input73/Z _4081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_96_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4983_ _5083_/C _4659_/Z _5415_/A1 _5173_/A2 _4984_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6722_ _6722_/D _7170_/RN _6722_/CLK _6722_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3934_ _7004_/Q _3934_/A2 _3934_/B1 _6845_/Q _5532_/A1 _6905_/Q _3937_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_149_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3865_ _6900_/Q _5528_/S _6611_/A1 _7297_/Q _3868_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6653_ _6771_/RN _6656_/A2 _6653_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_149_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5604_ _5859_/I0 hold901/Z _5610_/S _5604_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3796_ _3796_/A1 _3796_/A2 _3786_/Z _3795_/Z _3796_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6584_ _6584_/I0 _7271_/Q _6602_/S _7271_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5535_ hold177/Z hold64/Z _5535_/S _5535_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5466_ _5425_/Z _5428_/Z _5429_/Z _5465_/Z _5466_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_160_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7205_ _7205_/D _7205_/RN _7205_/CLK _7205_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4417_ _4930_/A1 _4715_/A1 _4836_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_121_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5397_ _5433_/A2 _5433_/A3 _5434_/A2 _5209_/Z _5398_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_160_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4348_ _5822_/I0 hold442/Z _4349_/S _4348_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7136_ _7136_/D _7141_/RN _7136_/CLK _7136_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_101_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout346 _4060_/S _6652_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xfanout357 _3520_/ZN _4225_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_143_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet1102_359 _4073__3/I _6851_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout368 _3552_/Z _5794_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_7067_ _7067_/D _7237_/RN _7067_/CLK _7067_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4279_ _6613_/I1 hold697/Z _4279_/S _4279_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout379 _3515_/Z _5884_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_98_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6018_ _7143_/Q _3385_/I _6210_/B _6211_/A2 _6024_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_74_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3650_ _7195_/Q _3909_/A2 _4194_/A1 input57/Z _3955_/A2 _7203_/Q _3689_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_174_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3581_ _3523_/Z _3932_/A2 _3925_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_127_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet902_201 net952_250/I _7024_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5320_ _5320_/A1 _5319_/Z _5452_/A2 _5453_/A4 _5320_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_177_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5251_ _5330_/B2 _5246_/Z _5251_/B _5254_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_47_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4202_ hold96/Z _5852_/I0 _4202_/S _4202_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5182_ _5182_/A1 _5340_/C _5265_/A4 _4511_/Z _5182_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4133_ hold20/Z hold114/Z _4136_/S _4133_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4064_ _6392_/B1 _7281_/Q _4064_/S _4064_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4966_ _4966_/A1 _4966_/A2 _5073_/B _4970_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6705_ _6705_/D _7237_/RN _6705_/CLK _6705_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3917_ _7110_/Q _3917_/A2 _6611_/A1 _7296_/Q _3919_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_20_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4897_ _3315_/I _6600_/B2 _6597_/C1 _4897_/A4 _4898_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_22_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6636_ _7075_/RN _6656_/A2 _6636_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_177_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3848_ _7127_/Q _3930_/A2 _3920_/B1 _6867_/Q _3922_/B1 _6693_/Q _3897_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_34_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6567_ _6567_/I0 _7265_/Q _6571_/S _7265_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3779_ _6982_/Q _3901_/A2 _3927_/B1 _7062_/Q _3796_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_180_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5518_ _4103_/I hold559/Z _5518_/S _5518_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6498_ _6498_/A1 _6498_/A2 _6498_/A3 _6498_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_106_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5449_ _5449_/A1 _5342_/I _5416_/I _5449_/A4 _5450_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_78_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7119_ _7119_/D _6933_/RN _7119_/CLK _7119_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_74_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/Z _4072_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_31_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__4 _4073__4/I _7221_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4820_ _4489_/B _4395_/B _4026_/B _4026_/C _4820_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_179_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_133__1359_ net1152_446/I net1202_483/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_61_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_53__1359_ clkbuf_4_14_0__1359_/Z net802_60/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_21_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4751_ _4751_/A1 _4748_/Z _4750_/Z _4755_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XTAP_1690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3702_ hold86/I _3912_/A2 _4194_/A1 input56/Z _3941_/A2 hold78/I _3708_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_4682_ _4530_/I _4878_/A2 _5312_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_147_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3633_ _6978_/Q _3923_/A2 _3960_/A2 _7212_/Q _3633_/C _3646_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6421_ _7255_/Q _6421_/I1 _6450_/S _7255_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6352_ _6990_/Q _6237_/Z _6240_/Z _7112_/Q _6352_/C _6356_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3564_ _5884_/A2 _5767_/A3 _3945_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_143_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5303_ _5303_/A1 _5303_/A2 _5303_/A3 _5303_/A4 _5303_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6283_ _6550_/A2 _6536_/B1 _6532_/A2 _6283_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_3495_ _7304_/Q _7303_/Q _3984_/S _3495_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5234_ _5234_/A1 _5314_/A1 _5404_/A1 _5234_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_130_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5165_ _5209_/A3 _5165_/A2 _4651_/Z _5165_/A4 _5165_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_151_1032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4116_ hold16/Z hold48/Z _4118_/S hold49/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5096_ _4539_/I _5369_/A1 _4673_/Z _5458_/A4 _5098_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_110_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4047_ _6768_/Q input91/Z _4050_/S _4047_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5998_ _7078_/Q _5996_/Z _5997_/Z _7094_/Q _6008_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XPHY_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4949_ _5464_/A1 _4944_/Z _5065_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_32_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6619_ _6644_/A1 _6648_/A2 _6619_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_137_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput280 _6668_/Q pll_trim[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput291 _6686_/Q pll_trim[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet852_111 _4073__51/I _7114_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_122 _4073__35/I _7103_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_133 _4073__9/I _7092_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_144 _4073__8/I _7081_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6970_ _6970_/D _7124_/RN _6970_/CLK _6970_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_81_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ _5920_/Z _5957_/I1 _7229_/Q _5913_/I _5922_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5852_ _5852_/I0 hold749/Z _5856_/S _5852_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4803_ _4803_/A1 _4797_/Z _4803_/B _4809_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_5783_ _5837_/I0 hold563/Z _5784_/S _5783_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4734_ _5401_/A2 _4728_/Z _5106_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_175_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4665_ _5170_/A2 _4878_/A2 _5389_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_119_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6404_ _7202_/Q _6540_/A2 _6536_/B1 _7040_/Q _6296_/Z hold78/I _6408_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_147_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold900 _4166_/Z _6711_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3616_ _5857_/A2 hold212/I _5521_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold911 _6718_/Q hold911/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold922 _5795_/Z _7134_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4596_ _5288_/B _4460_/B _4752_/A2 _4472_/B _4596_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold933 _7012_/Q hold933/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_127_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6335_ _6554_/A1 _6335_/A2 _6335_/A3 _6335_/A4 _6335_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold944 _5752_/Z _7096_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold955 _7144_/Q hold955/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3547_ _5875_/A1 _3523_/Z _3960_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold966 _4165_/Z _6710_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold977 _7013_/Q hold977/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold988 _5851_/Z _7184_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold999 _7069_/Q hold999/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6266_ _6300_/A2 _6533_/A4 _6285_/A2 _6302_/A4 _6266_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3478_ _3478_/I0 _5474_/A1 _3500_/S _3478_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5217_ _5460_/A1 _5460_/A4 _5224_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_130_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6197_ _6722_/Q _5987_/Z _6015_/Z _6841_/Q _6198_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5148_ _5147_/Z _5139_/Z _5148_/A3 _5470_/A3 _5148_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_85_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5079_ _5079_/A1 _5258_/C _5086_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_44_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4450_ _4607_/A1 _4451_/B _4451_/C _5356_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xhold207 _6756_/Q hold207/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold218 _5525_/Z _6898_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold229 _4252_/Z _6768_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3401_ _3401_/I _3401_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4381_ _4440_/B _4501_/B _3407_/I _4436_/B _4381_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_153_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6120_ _7017_/Q _5971_/Z _6005_/Z _7041_/Q _6124_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3332_ _4402_/B _4489_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XTAP_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout709 _6650_/A1 _6644_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ _6051_/A1 _6051_/A2 _6051_/B1 _5991_/Z _6052_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XTAP_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _4411_/Z _5258_/B2 _5002_/A3 _5002_/A4 _5002_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_94_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6953_ _6953_/D _7141_/RN _6953_/CLK _6953_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5904_ _7224_/Q _5903_/Z _5904_/B _5905_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6884_ _6884_/D _6886_/RN _6884_/CLK _6884_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_5835_ hold20/Z hold22/Z _5838_/S hold23/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5766_ hold285/Z _5865_/I0 _5766_/S _5766_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4717_ _5222_/A1 _5095_/B1 _5223_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5697_ _5808_/I0 hold625/Z _5700_/S _5697_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4648_ _4648_/A1 _4648_/A2 _4648_/B _5356_/C _5438_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_146_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold730 _5808_/Z _7146_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold741 _6787_/Q hold741/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_122_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4579_ _4380_/Z _4579_/A2 _4451_/B _4451_/C _5345_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold752 _4276_/Z _6788_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_150_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold763 _7034_/Q hold763/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6318_ _7199_/Q _6540_/A2 _6293_/Z _7151_/Q _6318_/C _6322_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold774 _5793_/Z _7133_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold785 _6825_/Q hold785/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold796 _5537_/Z _6906_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_118_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7298_ _7298_/D _6650_/Z _7302_/CLK _7298_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_89_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6249_ _7126_/Q _6247_/Z _6248_/Z _7068_/Q _6259_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_104_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet802_60 net802_60/I _7165_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet802_71 net802_71/I _7154_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet802_82 net802_82/I _7143_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet802_93 net802_93/I _7132_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold90 hold90/I hold90/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_75_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3950_ _6726_/Q _4188_/A1 _3950_/B1 _6724_/Q _3950_/C1 _6843_/Q _3953_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_189_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3881_ _7037_/Q _5683_/A1 _5674_/A1 _7029_/Q _3881_/C _3884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_91_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5620_ _5875_/A3 _5830_/A1 hold389/Z _5620_/A4 _5628_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_176_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5551_ _5860_/I0 hold132/Z _5556_/S _5551_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4502_ _4504_/B _4504_/C _5072_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5482_ _5482_/A1 _5482_/A2 _5483_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_172_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7221_ _7221_/D _7221_/RN _7221_/CLK _7221_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_160_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4433_ _4648_/A1 _4648_/A2 _4638_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_104_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7152_ _7152_/D _7207_/RN _7152_/CLK _7152_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_99_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4364_ _4460_/B _4752_/A2 _5315_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_141_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout506 hold39/Z hold40/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6103_ _6702_/Q _5965_/Z _6014_/Z _6960_/Q _6106_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xfanout517 _5879_/I0 _5852_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout528 _5850_/I0 _4343_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3315_ _3315_/I _4900_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_7083_ _7083_/D _7083_/RN _7083_/CLK _7083_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout539 _4360_/I1 _4103_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4295_ _6566_/I0 _6803_/Q _4300_/S _6803_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6034_ _7029_/Q _5999_/Z _6014_/Z _6957_/Q _6000_/Z _7127_/Q _6035_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6936_ _6936_/D _7140_/RN _6936_/CLK _6936_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XPHY_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6867_ _6867_/D _7162_/RN _6867_/CLK _6867_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5818_ _5818_/I0 hold867/Z _5820_/S _5818_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6798_ _6798_/D _7269_/CLK _6798_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5749_ _5857_/A3 _5821_/A3 _5767_/A3 _5857_/A4 _5757_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xnet1152_408 net1152_427/I _6766_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1152_419 net1152_419/I _6755_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold560 _5518_/Z _6893_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_2_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold571 _6820_/Q hold571/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold582 _6938_/Q hold582/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold593 _5699_/Z _7050_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_103_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4080_ input85/Z input58/Z _7300_/Q _4080_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4982_ _4997_/B _4982_/A2 _5263_/A2 _5322_/A1 _4982_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_63_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6721_ _6721_/D _6844_/RN _6721_/CLK _6721_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_189_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3933_ _7222_/Q _5528_/S _3933_/B1 _6785_/Q _3933_/C _3938_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_60_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6652_ _6850_/RN _6652_/A2 _6652_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3864_ _6723_/Q _4182_/A1 _3946_/A2 _6721_/Q input12/Z _3913_/A2 _3868_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5603_ _5804_/I0 hold695/Z _5610_/S _5603_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6583_ _6583_/A1 _6601_/A2 _6583_/B _6584_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_3795_ _3795_/A1 _3790_/Z _3794_/Z _3795_/A4 _3795_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5534_ hold171/Z hold54/Z _5535_/S _5534_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5465_ _5465_/A1 _5170_/Z _4882_/Z _4881_/Z _5465_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_105_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7204_ _7204_/D _7205_/RN _7204_/CLK _7204_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_160_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4416_ _5420_/A4 _4873_/A2 _5104_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_28_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5396_ _5396_/A1 _5395_/Z _5434_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_28_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7135_ _7135_/D _6892_/RN _7135_/CLK _7135_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4347_ _5821_/A1 _4353_/A1 _4347_/A3 _5821_/A3 _4349_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_59_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout347 _4064_/S _4060_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout358 _4976_/A3 _5324_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xfanout369 _3542_/Z _5830_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7066_ _7066_/D _7188_/RN _7066_/CLK _7066_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4278_ _5732_/I0 hold691/Z _4279_/S _4278_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6017_ _7167_/Q _6006_/Z _6030_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_67_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/Z _3340__1/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6919_ _6919_/D _7255_/RN _6919_/CLK _6919_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_74_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold390 _5602_/Z _5610_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_78_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3580_ _3505_/Z _5611_/A1 _5575_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_155_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5250_ _5250_/A1 _5247_/Z _5248_/Z _5250_/A4 _5251_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_170_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_13__1359_ net1152_430/I net1102_400/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4201_ _4200_/Z hold353/Z _4211_/S _4201_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5181_ _5127_/Z _5181_/A2 _5321_/A1 _5242_/A3 _5181_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xclkbuf_leaf_76__1359_ net902_187/I net802_73/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4132_ _5834_/I0 hold327/Z _4136_/S _4132_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4063_ _6747_/Q input3/Z input1/Z _4063_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4965_ _5076_/A1 _4908_/Z _5073_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6704_ _6704_/D _7188_/RN _6704_/CLK _6704_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_33_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3916_ _7150_/Q _3916_/A2 _3916_/B1 _6878_/Q _4274_/A1 _6787_/Q _3919_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_178_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4896_ _5290_/A2 _4892_/B _4897_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_177_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6635_ _7225_/RN _6656_/A2 _6635_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3847_ _5821_/A2 _3653_/Z _4170_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6566_ _6566_/I0 _7264_/Q _6571_/S _7264_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3778_ input37/Z _4244_/S _3948_/C1 input63/Z _3797_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5517_ _5517_/A1 _5517_/A2 _5517_/A3 _5520_/C _5518_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_133_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6497_ _7035_/Q _6269_/Z _6273_/Z _6979_/Q _6498_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5448_ _5448_/A1 _5483_/A2 _5448_/A3 _5463_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_161_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5379_ _5469_/A1 _5379_/A2 _5377_/Z _5379_/A4 _5379_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_160_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7118_ _7118_/D _6933_/RN _7118_/CLK _7118_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_75_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7049_ _7049_/D _7083_/RN _7049_/CLK _7049_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_41_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__5 _4073__5/I _7220_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4750_ _5478_/A3 _5099_/A1 _5401_/A2 _5226_/C _4750_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_1680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_0__1359_ net1152_451/I net1152_441/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3701_ _3701_/A1 _3701_/A2 _3701_/A3 _3701_/A4 _3701_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_30_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4681_ _5420_/A3 _4878_/A4 _3403_/I _4681_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_187_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6420_ _6420_/I _6421_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3632_ _3632_/I _3633_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_175_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6351_ _6351_/I _6352_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3563_ _5767_/A3 _3542_/Z _5758_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5302_ _4536_/Z _5283_/B _5302_/B _5303_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_143_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6282_ _6282_/A1 _6282_/A2 _7232_/Q _6282_/A4 _6282_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3494_ _3653_/A1 hold151/Z hold152/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_115_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5233_ _5233_/A1 _4757_/I _5156_/B _5233_/A4 _5404_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_170_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5164_ _5315_/A1 _5164_/A2 _5278_/B _5164_/A4 _5467_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_29_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4115_ hold14/Z _7276_/Q _4117_/S hold15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5095_ _5278_/C _5307_/A3 _5228_/A3 _5095_/B1 _4697_/Z _5460_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_112_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4046_ _4046_/I _6832_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ _6068_/A2 _6117_/A4 _6014_/A2 _3389_/I _5997_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XPHY_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4948_ _4948_/A1 _4945_/Z _4946_/Z _4947_/Z _4953_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_178_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4879_ _5315_/A2 _4524_/Z _5146_/A1 _4820_/Z _4879_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_177_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6618_ _6644_/A1 _6650_/A2 _6618_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_119_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6549_ _6846_/Q _6549_/A2 _6549_/B1 _6842_/Q _6549_/C1 _6840_/Q _6554_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_180_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput270 _6885_/Q pll_sel[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput281 _6669_/Q pll_trim[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput292 hold50/I pll_trim[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_58_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet852_112 net802_93/I _7113_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_123 net802_66/I _7102_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_134 _4073__39/I _7091_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_145 net802_89/I _7080_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5920_ _7229_/Q _6210_/B _5920_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_81_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5851_ _5869_/I0 hold987/Z _5856_/S _5851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4802_ _5453_/A4 _5420_/A3 _5456_/A1 _5130_/B1 _5129_/A2 _5389_/A1 _4803_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_21_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5782_ _5782_/I0 hold271/Z _5784_/S _5782_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4733_ _4733_/A1 _4729_/Z _4731_/Z _4732_/Z _4739_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_187_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4664_ _4664_/A1 _4664_/A2 _4663_/Z _4670_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_175_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6403_ _7114_/Q _6240_/Z _6403_/B _6408_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3615_ _5857_/A2 _5857_/A3 _3508_/Z _3477_/Z _3866_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_128_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold901 _6965_/Q hold901/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4595_ _5190_/A2 _4635_/A4 _5438_/A1 _5435_/A2 _4595_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold912 _4177_/Z _6718_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold923 _7065_/Q hold923/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold934 _5657_/Z _7012_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6334_ _7045_/Q _6550_/A2 _6550_/C1 _6949_/Q _6543_/A2 _7215_/Q _6335_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3546_ hold221/I _3492_/Z _3904_/A4 _3904_/A2 _3546_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold945 _7030_/Q hold945/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold956 _5806_/Z _7144_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold967 _7014_/Q hold967/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold978 _5658_/Z _7013_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_171_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6265_ _6302_/A3 _6533_/A4 _6285_/A2 _6302_/A4 _6265_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold989 _7157_/Q hold989/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_88_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3477_ _3475_/Z _3309_/I _3500_/S _3477_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_88_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5216_ _4697_/Z _5310_/A2 _5460_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_131_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6196_ _6712_/Q _6002_/Z _6003_/Z _6714_/Q _6198_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_9_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5147_ _4842_/Z _5147_/A2 _5147_/A3 _5147_/A4 _5147_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_28_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5078_ _5324_/A1 _5078_/A2 _5263_/A4 _5263_/A2 _5337_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_38_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4029_ _4029_/A1 _4029_/A2 _4391_/A3 _4391_/A4 _4031_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_44_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold208 _4233_/Z _6756_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold219 _6862_/Q hold219/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3400_ _3400_/I _6601_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_4380_ _4501_/A1 _4455_/A2 _5170_/A2 _4380_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_3331_ _7237_/Q _6253_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _7152_/Q _5960_/Z _5965_/Z _6700_/Q _5969_/Z _7120_/Q _6053_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5001_ _5000_/Z _5001_/A2 _5001_/B _6859_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6952_ _6952_/D _7002_/RN _6952_/CLK _6952_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_81_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5903_ _5901_/B _5902_/Z _7223_/Q _5903_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6883_ _6883_/D _6886_/RN _6883_/CLK _6883_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_62_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5834_ _5834_/I0 hold238/Z _5838_/S _5834_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5765_ hold289/Z _5891_/I0 _5766_/S _5765_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4716_ _5420_/A2 _4835_/A2 _5420_/A4 _5129_/A4 _4716_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5696_ _5879_/I0 hold244/Z _5700_/S _5696_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4647_ _5038_/A1 _5475_/A3 _5439_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold720 _5874_/Z _7205_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold731 _6858_/Q hold731/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4578_ _5201_/A1 _5438_/C _5346_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold742 _4275_/Z _6787_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold753 _6824_/Q hold753/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6317_ _7135_/Q _6253_/Z _6296_/Z _7159_/Q _6322_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold764 _5681_/Z _7034_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3529_ _3478_/Z _3552_/A2 _3484_/Z hold27/Z _3529_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_131_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7297_ _7297_/D _7297_/RN _7297_/CLK _7297_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold775 _6669_/Q hold775/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_1_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold786 _4328_/Z _6825_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold797 _6666_/Q hold797/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_115_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6248_ _5946_/S _6452_/A2 _6452_/A4 _6253_/A4 _6248_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_162_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6179_ _7117_/Q _5984_/Z _5997_/Z _7101_/Q _7075_/Q _5980_/Z _6180_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_45_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet802_61 net802_93/I _7164_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet802_72 _4073__8/I _7153_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet802_83 net802_83/I _7142_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet802_94 net802_94/I _7131_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold80 hold80/I hold80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_91_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold91 hold91/I hold91/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_17_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3880_ _3880_/I _3881_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_189_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5550_ hold54/Z _5550_/I1 _5556_/S hold55/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4501_ _4501_/A1 _4884_/A1 _4501_/B _4504_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_144_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5481_ _4944_/Z _5245_/Z _5481_/B1 _4951_/Z _5481_/C _5482_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_184_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7220_ _7220_/D _7220_/RN _7220_/CLK _7220_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4432_ _3407_/I _4376_/Z _4648_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_126_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7151_ _7151_/D _7218_/RN _7151_/CLK _7151_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_126_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4363_ _3407_/I _4652_/A1 _4363_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_98_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6102_ _6952_/Q _5958_/Z _5999_/Z _7032_/Q _6102_/C _6106_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xfanout507 hold19/Z hold20/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_141_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3314_ _6950_/Q _3994_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
Xfanout518 hold60/Z _5879_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_7082_ _7082_/D _7155_/RN _7082_/CLK _7082_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout529 _5778_/I0 _6613_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4294_ _6565_/I0 _6802_/Q _4300_/S _6802_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6033_ _7061_/Q _5985_/Z _5997_/Z _7095_/Q _6037_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6935_ _6935_/D _7177_/RN _6935_/CLK _6935_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XPHY_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6866_ _6866_/D _7162_/RN _6866_/CLK _6866_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5817_ hold20/Z hold24/Z _5820_/S hold25/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6797_ _6797_/D _7269_/CLK _6797_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5748_ _5865_/I0 hold605/Z _5748_/S _5748_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5679_ hold552/Z _5808_/I0 _5682_/S _5679_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1152_409 net1152_409/I _6765_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold550 _7000_/Q hold550/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold561 _6890_/Q hold561/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold572 _4321_/Z _6820_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_132_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold583 _5573_/Z _6938_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_173_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold594 _6930_/Q hold594/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_173_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4981_ _5262_/A2 _5255_/A2 _4982_/A2 _4497_/Z _4981_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6720_ _6720_/D _6844_/RN _6720_/CLK _6720_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3932_ _3932_/A1 _3932_/A2 _5830_/A1 _3932_/B _3933_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_108_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_36__1359_ _4073__6/I net1152_414/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_116__1359_ net952_221/I net902_181/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6651_ _7225_/RN _6656_/A2 _6651_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_20_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3863_ _6973_/Q _3923_/A2 _3959_/C1 _7183_/Q _3869_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_177_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_99__1359_ clkbuf_4_5_0__1359_/Z net952_241/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_176_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5602_ _5866_/A3 _3515_/Z hold389/Z _5620_/A4 _5602_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6582_ _6600_/A1 _6582_/A2 _6582_/B1 _3316_/I _3317_/I _6582_/C2 _6583_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3794_ _3794_/A1 _3794_/A2 _3794_/A3 _3794_/A4 _3794_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_164_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5533_ hold191/Z _5860_/I0 _5535_/S _5533_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5464_ _5464_/A1 _4659_/Z _4675_/Z _5464_/B _5465_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_145_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7203_ _7203_/D _7219_/RN _7203_/CLK _7203_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4415_ _5385_/A1 _5045_/C _4415_/B _5211_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_132_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5395_ _5395_/A1 _4991_/C _5428_/A2 _5395_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_67_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7134_ _7134_/D _6892_/RN _7134_/CLK _7134_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_87_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4346_ _6613_/I1 hold839/Z _4346_/S _4346_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout348 _6657_/A2 _6650_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7065_ _7065_/D _7083_/RN _7065_/CLK _7065_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_101_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4277_ _4332_/A1 _5794_/A3 hold146/Z _5857_/A2 _4279_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xfanout359 _5315_/A4 _5478_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_101_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6016_ _7013_/Q _5971_/Z _6031_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_55_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6918_ _6918_/D _7257_/RN _6918_/CLK _6918_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6849_ _6849_/D _6850_/RN _6849_/CLK _6849_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_50_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold380 _5777_/Z _7118_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold391 _5605_/Z _6966_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_117_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold1080 _7282_/Q _4041_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4200_ hold128/Z _5860_/I0 _4202_/S _4200_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5180_ _5180_/A1 _5180_/A2 _5180_/A3 _5211_/C _5185_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_111_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4131_ _5842_/I0 hold140/Z _4136_/S _4131_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_4_12_0__1359_ clkbuf_0__1359_/Z net902_187/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4062_ _4061_/Z _3337_/I _7299_/Q _4062_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4964_ _5010_/A1 _4908_/Z _4966_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6703_ hold43/Z _7075_/RN _6703_/CLK hold42/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3915_ _3915_/A1 _3915_/A2 _3915_/A3 _3915_/A4 _3915_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4895_ _4886_/Z _4887_/Z _4891_/Z _4895_/A4 _4898_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_32_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3846_ _3540_/Z _5821_/A2 _3939_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6634_ _6644_/A1 _6650_/A2 _6634_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_20_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet1202_490 net1202_490/I _6675_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6565_ _6565_/I0 _7263_/Q _6571_/S _7263_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3777_ _7176_/Q _3945_/A2 _5532_/A1 _6903_/Q _3797_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5516_ _5795_/I0 _5516_/I1 _5516_/S _5516_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6496_ _6947_/Q _6551_/A2 _6288_/Z _7125_/Q _6498_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_146_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5447_ _5447_/A1 _5447_/A2 _5448_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_133_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5378_ _5425_/A2 _5425_/A3 _5379_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4329_ _4332_/A1 _5629_/A3 hold146/Z _5794_/A3 _4331_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7117_ _7117_/D _7237_/RN _7117_/CLK _7117_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_102_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7048_ _7048_/D _7260_/RN _7048_/CLK _7048_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_101_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4073__6 _4073__6/I _7219_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_156_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_82__1359_ net902_187/I net952_206/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_7_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout690 fanout714/Z _6915_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_65_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3700_ _6686_/Q _3945_/C2 _5683_/A1 _7040_/Q _3701_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4680_ _4414_/Z _4452_/Z _4666_/Z _5395_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_175_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3631_ _6938_/Q _3910_/A2 _3954_/A2 _6994_/Q _7204_/Q _3955_/A2 _3632_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6350_ _7128_/Q _6247_/Z _6297_/Z _6700_/Q _6351_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3562_ _3507_/Z _5731_/A2 _3927_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_128_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5301_ _5301_/I _6861_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6281_ _6484_/A3 _6535_/A2 _6540_/A2 _6543_/A2 _6281_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_142_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3493_ _3493_/I0 hold150/Z _3500_/S _3493_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5232_ _5364_/A1 _4752_/Z _5233_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_64_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5163_ _5356_/A1 _4650_/Z _5231_/A2 _5468_/A1 _5166_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_97_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4114_ _5836_/I0 hold303/Z _4118_/S _4114_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5094_ _5328_/A1 _5389_/A1 _5094_/B _5094_/C _5347_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_151_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4045_ _6832_/Q _4097_/A1 _4045_/B1 _6826_/Q _4046_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_37_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5996_ _6068_/A2 _6210_/B _6014_/A2 _3389_/I _5996_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XPHY_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4947_ _5072_/A4 _4903_/Z _5010_/A1 _4500_/Z _4947_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_138_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4878_ _4889_/A1 _4878_/A2 _5426_/A1 _4878_/A4 _4878_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_166_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6617_ _7071_/RN _6657_/A2 _6617_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3829_ _5767_/A3 _3560_/Z _4161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6548_ _6548_/A1 _6548_/A2 _6548_/A3 _6547_/Z _6548_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_116_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6479_ _7189_/Q _6532_/A2 _6492_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_161_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput260 _6891_/Q pll_bypass VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput271 _6682_/Q pll_trim[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput282 _6683_/Q pll_trim[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput293 _6688_/Q pll_trim[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet852_102 net952_229/I _7123_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_113 net902_187/I _7112_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_124 _4073__12/I _7101_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet852_135 _4073__39/I _7090_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet852_146 net852_146/I _7079_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5850_ _5850_/I0 hold450/Z _5856_/S _5850_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4801_ _5312_/A2 _5312_/A4 _5456_/A1 _5220_/B2 _4801_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_2190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5781_ _5781_/I0 hold263/Z _5784_/S _5781_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4732_ _4765_/A1 _5236_/A1 _4774_/A3 _5099_/A2 _4732_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_187_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4663_ _4411_/Z _5214_/A2 _5172_/B _5165_/A4 _4663_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6402_ _7130_/Q _6402_/A2 _6452_/A3 _6533_/A4 _6403_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3614_ _3505_/Z _3932_/A2 _3770_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4594_ _5190_/A2 _5435_/A2 _5389_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold902 _5604_/Z _6965_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold913 _7128_/Q hold913/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold924 _5716_/Z _7065_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6333_ _7207_/Q _6535_/A2 _6544_/B1 _6957_/Q _6285_/Z _7191_/Q _6335_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3545_ _5875_/A1 _5776_/A1 _3959_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold935 _7135_/Q hold935/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold946 _5677_/Z _7030_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold957 _7038_/Q hold957/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold968 _5659_/Z _7014_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_115_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6264_ _6956_/Q _6544_/B1 _6545_/A2 _6932_/Q _6531_/A2 _6964_/Q _6271_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_115_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold979 _7095_/Q hold979/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_88_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3476_ _3476_/I _3478_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5215_ _4698_/B _5403_/A2 _5215_/B _5215_/C _5316_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_6195_ _6824_/Q _5988_/Z _6019_/Z _6853_/Q _6198_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_9_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5146_ _5146_/A1 _5364_/B _4586_/Z _4598_/Z _5438_/A1 _5147_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_97_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5077_ _4973_/Z _5078_/A2 _5258_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_56_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4028_ input97/Z input96/Z input99/Z input98/Z _4028_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_44_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5979_ _6002_/A2 _6021_/A2 _6210_/A2 _6021_/A4 _5979_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_139_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold209 _6859_/Q _3305_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_172_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3330_ _5946_/S _6285_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_152_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_0_0__1359_ clkbuf_0__1359_/Z net1152_451/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5000_ _5000_/A1 _5000_/A2 _5000_/A3 _5000_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XTAP_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6951_ _6951_/D _7002_/RN _6951_/CLK _6951_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_53_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5902_ _5911_/A1 _5951_/B _7225_/Q _5902_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_81_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6882_ hold30/Z _6882_/RN _6882_/CLK _6882_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_179_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5833_ _5833_/I0 hold689/Z _5838_/S _5833_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5764_ hold345/Z _5881_/I0 _5766_/S _5764_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4715_ _4715_/A1 _5087_/A1 _5328_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5695_ _5806_/I0 _5695_/I1 _5700_/S _5695_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4646_ _4648_/A1 _4648_/A2 _4648_/B _5475_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_30_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold710 _4156_/Z _6704_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_162_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold721 _7207_/Q hold721/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4577_ _5002_/A3 _5002_/A4 _5080_/B _5003_/A2 _5043_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold732 _4361_/Z _6858_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold743 _6785_/Q hold743/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_1_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold754 _4327_/Z _6824_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6316_ _7167_/Q _6544_/A2 _6551_/A2 _6941_/Q _6545_/A2 _6933_/Q _6329_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold765 _6993_/Q hold765/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3528_ _3525_/Z _5510_/A2 _3935_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_103_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7296_ _7296_/D _7296_/RN _7296_/CLK _7296_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold776 _4110_/Z _6669_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold787 _6822_/Q hold787/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_130_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold798 _4104_/Z _6666_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_130_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6247_ _5946_/S _6452_/A2 _6533_/A4 _6253_/A4 _6247_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3459_ hold1/Z hold52/Z _3460_/S _7285_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6178_ _7157_/Q _5960_/Z _5965_/Z _6705_/Q _6006_/Z _7173_/Q _6180_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_69_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5129_ _5420_/A2 _5129_/A2 _5129_/A3 _5129_/A4 _5129_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_2904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet802_62 net802_62/I _7163_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet802_73 net802_73/I _7152_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet802_84 net802_84/I _7141_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet802_95 net802_95/I _7130_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold70 hold70/I hold70/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold81 hold81/I hold81/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_91_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold92 hold92/I hold92/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_63_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4500_ _4759_/A2 _4759_/A3 _4500_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
X_5480_ _5480_/A1 _5480_/A2 _5480_/A3 _5479_/Z _5480_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_172_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_1 _5498_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4431_ _4414_/Z _5010_/A1 _5393_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_144_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7150_ _7150_/D _6907_/RN _7150_/CLK _7150_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4362_ _5299_/C _6859_/Q _5001_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_113_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6101_ _6101_/A1 _6101_/A2 _6101_/A3 _6101_/A4 _6101_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3313_ _6830_/Q _4038_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7081_ _7081_/D _7179_/RN _7081_/CLK _7081_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xfanout508 hold19/Z _5889_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4293_ _6564_/I0 _6801_/Q _4300_/S _6801_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout519 hold59/Z hold60/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_140_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6032_ _7069_/Q _5980_/Z _6003_/Z _7159_/Q _6037_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xclkbuf_leaf_59__1359_ clkbuf_4_15_0__1359_/Z net1152_415/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_139__1359_ net1152_451/I net1202_471/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_112_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6934_ _6934_/D _7019_/RN _6934_/CLK _6934_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XPHY_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6865_ _6865_/D _6865_/RN _6865_/CLK hold26/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5816_ _5888_/I0 hold440/Z _5820_/S _5816_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6796_ _6796_/D _7269_/CLK _6796_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5747_ _5837_/I0 hold831/Z _5748_/S _5747_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5678_ hold248/Z _5879_/I0 _5682_/S _5678_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4629_ _5190_/A2 _4604_/Z _5387_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_151_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold540 _5617_/Z _6977_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold551 _5643_/Z _7000_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_1_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold562 _5512_/Z _6890_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold573 _6891_/Q hold573/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold584 _7203_/Q hold584/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold595 _5564_/Z _6930_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7279_ _7279_/D _7279_/RN _7279_/CLK hold31/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_131_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput160 wb_rstn_i input160/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4980_ _4998_/A2 _5262_/A2 _5255_/A2 _5323_/B _4980_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_91_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3931_ _7052_/Q _5701_/A1 _5536_/A1 _6906_/Q _3932_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_60_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6650_ _6650_/A1 _6650_/A2 _6650_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_31_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3862_ _6957_/Q _3957_/A2 _3928_/C1 _6823_/Q _3925_/B1 _6825_/Q _3869_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_31_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5601_ _5784_/I0 hold889/Z _5601_/S _5601_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6581_ _6581_/I0 hold62/I _6602_/S _7270_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3793_ _7136_/Q _3951_/A2 _3924_/A2 _6966_/Q _3794_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_176_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5532_ _5532_/A1 hold33/I _5535_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_173_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5463_ _5463_/A1 _5463_/A2 _5485_/A2 _5463_/B2 _5463_/C _5474_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_7202_ _7202_/D _7202_/RN _7202_/CLK _7202_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4414_ _4397_/Z _4491_/B _5003_/A2 _4414_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_5394_ _4892_/B _5394_/A2 _5428_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_113_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7133_ _7133_/D _7188_/RN _7133_/CLK _7133_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4345_ _6612_/I1 hold851/Z _4346_/S _4345_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7064_ _7064_/D _7090_/RN _7064_/CLK _7064_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4276_ hold751/Z _5538_/I1 _4276_/S _4276_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout349 _6656_/A2 _6648_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_113_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6015_ _7228_/Q _6164_/B1 _6015_/A3 _6139_/A2 _6015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_55_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6917_ hold55/Z _7034_/RN _6917_/CLK _6917_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6848_ _6848_/D _7297_/RN _6848_/CLK _6848_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_52_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6779_ _6779_/D _7002_/RN _6779_/CLK _6779_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold370 _4235_/Z _6757_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold381 _6670_/Q hold381/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_77_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold392 _6950_/Q hold392/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_122__1359_ net952_221/I _4073__42/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_42__1359_ clkbuf_4_11_0__1359_/Z _4073__4/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_58_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold1070 _7294_/Q _3433_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1081 _7294_/Q _3440_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4130_ _6613_/I1 hold793/Z _4136_/S _4130_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4061_ _4060_/Z input38/Z _7301_/Q _4061_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4963_ _4963_/A1 _4960_/Z _4961_/Z _4962_/Z _4966_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6702_ _6702_/D _7140_/RN _6702_/CLK _6702_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3914_ _7102_/Q _5758_/A1 _3914_/B1 _6876_/Q _3915_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4894_ _4894_/A1 _4893_/Z _4895_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_189_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6633_ _7162_/RN _6652_/A2 _6633_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3845_ _7061_/Q _3927_/B1 _3955_/B1 _6848_/Q _3895_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xnet1202_480 net1202_481/I _6685_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1202_491 net1202_491/I _6674_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6564_ _6564_/I0 _7262_/Q _6571_/S _7262_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3776_ _3773_/Z _3776_/A2 _3776_/A3 _3776_/A4 _3776_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5515_ hold258/Z _5785_/A3 _5629_/A3 hold11/Z _5515_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_145_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6495_ _7051_/Q _6241_/Z _6550_/B1 _6987_/Q _6550_/C1 _6955_/Q _6498_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_121_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5446_ _5446_/A1 _5446_/A2 _5447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_173_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5377_ _5377_/A1 _5290_/Z _5377_/A3 _5377_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_7116_ _7116_/D _7185_/RN _7116_/CLK _7116_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4328_ _6613_/I1 hold785/Z _4328_/S _4328_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7047_ _7047_/D _7125_/RN _7047_/CLK _7047_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4259_ _5890_/I0 hold205/Z _4261_/S _4259_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__7 _4073__7/I _7218_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_169_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_170_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout680 fanout685/Z _7163_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_19_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout691 _7205_/RN _7221_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_93_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3630_ _3630_/A1 _3630_/A2 _3630_/A3 _3630_/A4 _3630_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_159_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3561_ _3932_/A2 _3560_/Z _3913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_115_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5300_ _5242_/Z _5266_/Z _5300_/A3 _5299_/C _6861_/Q _5301_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_128_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3492_ _3491_/I _3307_/I _3500_/S _3492_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_6280_ _6551_/A2 _6531_/A2 _6545_/A2 _6279_/Z _6287_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_154_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5231_ _5291_/B _5231_/A2 _5231_/B _5231_/C _5314_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_103_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5162_ _5165_/A2 _5278_/B _5164_/A2 _5315_/A1 _5467_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4113_ hold38/Z _7275_/Q _4113_/S hold39/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5093_ _5093_/A1 _5438_/A1 _5218_/B _5303_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_96_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4044_ _4044_/I _6732_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5995_ _7052_/Q _5924_/Z _5994_/I _7134_/Q _5995_/C _6009_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XPHY_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4946_ _4500_/Z _4903_/Z _5072_/A4 _5475_/A4 _4946_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_21_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4877_ _4651_/Z _4877_/A2 _5173_/A2 _5287_/A2 _4877_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_20_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6616_ _6656_/A1 _6657_/A2 _6616_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3828_ _4350_/A2 _5731_/A2 _3956_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_165_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6547_ _6547_/A1 _6547_/A2 _6542_/Z _6546_/Z _6547_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3759_ _3759_/A1 _3759_/A2 _3747_/Z _3758_/Z _3759_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_152_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6478_ _7043_/Q _6536_/B1 _6486_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_173_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5429_ _4898_/C _4991_/C _5392_/B _4893_/Z _5429_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_134_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput250 _4092_/ZN pad_flash_csb_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput261 _6877_/Q pll_dco_ena VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput272 _6676_/Q pll_trim[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput283 _6670_/Q pll_trim[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput294 hold70/I pll_trim[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_88_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet852_103 net952_241/I _7122_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_114 net802_98/I _7111_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet852_125 _4073__48/I _7100_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_136 net852_136/I _7089_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_147 net852_147/I _7078_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_171_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4800_ _5380_/B2 _5287_/A2 _5130_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_21_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5780_ _5888_/I0 hold446/Z _5784_/S _5780_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _4765_/A1 _4774_/A3 _5099_/A2 _5226_/A1 _4731_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_187_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4662_ _5464_/A1 _4414_/Z _4659_/Z _4662_/B _4664_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_30_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6401_ _6401_/A1 _6401_/A2 _6401_/A3 _6401_/A4 _6401_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_70_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3613_ _7074_/Q _3943_/A2 _3647_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_174_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4593_ _4593_/A1 _5018_/B _4601_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_31_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold903 _6698_/Q hold903/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6332_ _6981_/Q _6550_/B1 _6254_/Z _7175_/Q _6332_/C _6335_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold914 _5788_/Z _7128_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold925 _6700_/Q hold925/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3544_ input51/Z _4202_/S _4244_/S input42/Z _3589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold936 _5796_/Z _7135_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold947 _7051_/Q hold947/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold958 _5686_/Z _7038_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold969 _7151_/Q hold969/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6263_ _7232_/Q _6275_/A4 _6452_/A4 _6282_/A2 _6263_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_142_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3475_ _6660_/Q _3475_/I1 _3984_/S _3475_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5214_ _5343_/A2 _5214_/A2 _5310_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6194_ _6820_/Q _5979_/Z _5996_/Z _6708_/Q _6198_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_96_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5145_ _4570_/Z _5145_/A2 _4878_/Z _5278_/B _4820_/Z _4821_/Z _5147_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai222_4
XFILLER_56_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5076_ _5076_/A1 _4905_/Z _4973_/Z _5260_/A1 _5076_/C _5079_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_4027_ _4027_/A1 _4027_/A2 _4031_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_53_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5978_ _5924_/Z _5975_/Z _5976_/Z _5977_/Z _5983_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_139_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4929_ _4929_/A1 _4928_/Z _4929_/A3 _4933_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_138_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6950_ _6950_/D _7002_/RN _6950_/CLK _6950_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_53_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5901_ _5901_/A1 _5951_/A3 _5901_/B _5904_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_35_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6881_ _6881_/D _6882_/RN _6881_/CLK _6881_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_90_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5832_ _5832_/I0 _5832_/I1 _5838_/S _5832_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5763_ hold347/Z _5871_/I0 _5766_/S _5763_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_19__1359_ _4073__49/I net902_185/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4714_ _4709_/Z _4711_/Z _5305_/B _4714_/A4 _4727_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5694_ _5859_/I0 hold939/Z _5700_/S _5694_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4645_ _4565_/Z _4641_/Z _5040_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_147_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold700 _5864_/Z _7196_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold711 _7220_/Q hold711/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_162_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4576_ _4549_/Z _4570_/Z _5192_/B _4576_/C _4584_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xhold722 _5877_/Z _7207_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold733 _7180_/Q hold733/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold744 _4272_/Z _6785_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6315_ _7183_/Q _6532_/A2 _6322_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold755 _6929_/Q hold755/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3527_ _3552_/A2 _3484_/Z hold27/Z hold137/Z _3527_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_104_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7295_ _7295_/D _6649_/Z _7302_/CLK _7295_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold766 _5635_/Z _6993_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold777 _6907_/Q hold777/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold788 _4324_/Z _6822_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6246_ _7004_/Q _6549_/B1 _6551_/A2 _6940_/Q _6260_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold799 _6925_/Q hold799/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_103_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3458_ hold58/Z hold1/Z _3460_/S _7286_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6177_ _7109_/Q _5967_/Z _6177_/B _6180_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3389_ _3389_/I _5984_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_58_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5128_ _5453_/A4 _5319_/A3 _5181_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_73_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5059_ _5260_/A1 _5325_/B _5060_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet802_52 net802_52/I _7173_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet802_63 net802_63/I _7162_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet802_74 _4073__7/I _7151_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet802_85 net802_87/I _7140_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet802_96 net802_96/I _7129_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold60 hold60/I hold60/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold71 hold71/I hold71/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold82 hold82/I hold82/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold93 hold93/I hold93/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_75_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4430_ _4402_/B _4026_/B _4026_/C _5083_/C _4997_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_172_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_2 _5518_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4361_ hold731/Z _4361_/I1 _4361_/S _4361_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6100_ _7016_/Q _5971_/Z _5988_/Z _6984_/Q _6005_/Z _7040_/Q _6101_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_113_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3312_ _3312_/I _3428_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7080_ hold85/Z _7155_/RN _7080_/CLK hold84/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xfanout509 _5880_/I0 _5871_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4292_ _6828_/Q _6563_/A2 _4300_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_141_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6031_ _6031_/A1 _6026_/Z _6030_/Z _6031_/A4 _6031_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_98_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6933_ _6933_/D _6933_/RN _6933_/CLK _6933_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_70_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6864_ _6864_/D _6865_/RN _6865_/CLK _6864_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_168_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5815_ _5869_/I0 hold885/Z _5820_/S _5815_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6795_ _6795_/D _7258_/CLK _6795_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ _5881_/I0 hold781/Z _5748_/S _5746_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5677_ hold945/Z _5806_/I0 _5682_/S _5677_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4628_ _4565_/Z _4624_/Z _5035_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_163_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold530 _5493_/Z _6867_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold541 hold541/I hold541/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_144_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4559_ _5464_/A1 _4889_/A1 _5393_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold552 _7032_/Q hold552/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_2_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold563 _7124_/Q hold563/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold574 _5514_/Z _6891_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_131_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold585 _5872_/Z _7203_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7278_ _7278_/D _7278_/RN _7279_/CLK _7278_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold596 _6852_/Q hold596/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_103_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6229_ _6220_/Z _6228_/Z _6555_/B1 _6118_/B _6555_/C _6230_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_145__1359_ net1152_451/I net1202_487/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_65__1359_ clkbuf_4_13_0__1359_/Z net952_226/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_154_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput150 wb_dat_i[2] _3395_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput161 wb_sel_i[0] _6572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3930_ _7126_/Q _3930_/A2 _3930_/B1 _6841_/Q _4170_/A1 _6714_/Q _3938_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_147_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3861_ _7207_/Q _3960_/A2 _3955_/A2 _7199_/Q _3924_/A2 _6965_/Q _3869_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_32_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5600_ _5681_/I1 hold761/Z _5601_/S _5600_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6580_ _6580_/A1 _6601_/A2 _6580_/B _6581_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_3792_ _6990_/Q _3954_/A2 _3954_/B1 input22/Z _3794_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5531_ _5885_/I0 hold469/Z _5531_/S _5531_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5462_ _5404_/Z _5457_/Z _5461_/I _5463_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_145_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7201_ _7201_/D _7201_/RN _7201_/CLK _7201_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4413_ _5209_/A3 _4397_/Z _5045_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5393_ _5393_/A1 _5393_/A2 _5393_/B1 _5045_/C _5433_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_132_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7132_ _7132_/D _7188_/RN _7132_/CLK _7132_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_154_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4344_ _4353_/A1 _4350_/A2 _4350_/A3 _4346_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_114_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7063_ _7063_/D _7075_/RN _7063_/CLK _7063_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4275_ hold741/Z _5537_/I1 _4276_/S _4275_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6014_ _6210_/B _6014_/A2 _6139_/A2 _3389_/I _6014_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_39_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6916_ _6916_/D _7257_/RN _6916_/CLK _6916_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6847_ _6847_/D _6847_/RN _6847_/CLK _6847_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_11_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6778_ _6778_/D _6967_/RN _6778_/CLK _6778_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5729_ hold783/Z _5732_/I0 _5730_/S _5729_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold360 _5552_/Z _6919_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold371 _7006_/Q hold371/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold382 _4112_/Z _6670_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold393 _5587_/Z _6950_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_105_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1060 _6661_/Q _3979_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold1071 _7008_/Q _5652_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4060_ _6748_/Q _6875_/Q _4060_/S _4060_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4962_ _4500_/Z _4906_/Z _5072_/A4 _4666_/Z _4962_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3913_ input11/Z _3913_/A2 _3913_/B1 _6892_/Q _3915_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_51_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6701_ _6701_/D _7075_/RN _6701_/CLK _6701_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_189_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4893_ _5139_/A2 _5139_/A3 _4542_/Z _5172_/C _4893_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_149_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6632_ _7162_/RN _6652_/A2 _6632_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3844_ _3844_/A1 _4350_/A2 _3955_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_20_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet1202_470 net1202_471/I _6695_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1202_481 net1202_481/I _6684_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6563_ _6833_/D _6563_/A2 _6571_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_158_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet1202_492 net1202_494/I _6673_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3775_ _7112_/Q _3917_/A2 _3913_/A2 input13/Z _3916_/A2 _7152_/Q _3776_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_158_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5514_ _4103_/I hold573/Z _5514_/S _5514_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6494_ _7027_/Q _6235_/Z _6243_/Z _7011_/Q _6549_/C1 _7003_/Q _6499_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_145_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5445_ _4376_/Z _5255_/B _4972_/Z _5445_/B2 _5056_/B _5445_/C2 _5446_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_145_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5376_ _5276_/B _5376_/A2 _5468_/B1 _5376_/B2 _5376_/C _5377_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_87_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7115_ hold45/Z _7237_/RN _7115_/CLK hold44/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4327_ _5732_/I0 hold753/Z _4328_/S _4327_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7046_ _7046_/D _7247_/RN _7046_/CLK _7046_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4258_ _5889_/I0 hold98/Z _4261_/S hold99/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4189_ hold523/Z _4360_/I1 _4190_/S _4189_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073__8 _4073__8/I _7217_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_169_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold190 _4265_/Z _6779_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout670 _7083_/RN _7259_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_77_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout681 _7027_/RN _7124_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout692 _7205_/RN _7201_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_93_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3560_ _3904_/A3 _3680_/A3 _3500_/Z hold221/I _3560_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_115_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3491_ _3491_/I _3493_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5230_ _5236_/A1 _5364_/A1 _5230_/B _5231_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_154_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_170_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5161_ _5161_/A1 _5161_/A2 _5366_/A1 _5166_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_142_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4112_ _5871_/I0 hold381/Z _4118_/S _4112_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5092_ _5092_/A1 _4705_/Z _5218_/B _5228_/A3 _5303_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_56_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4043_ _4043_/A1 _6732_/Q _3304_/I _3409_/Z _4044_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_83_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5994_ _5994_/I _6051_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_178_710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4945_ _4500_/Z _4903_/Z _4973_/A4 _5020_/A2 _4945_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_33_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4876_ _4650_/Z _4876_/A2 _4876_/B _4876_/C _4880_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_166_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3827_ _4185_/A2 _3540_/Z _3946_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6615_ _6656_/A1 _6657_/A2 _6615_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_177_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6546_ _6546_/A1 _6546_/A2 _6546_/A3 _6546_/A4 _6546_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_119_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3758_ _3758_/A1 _3751_/Z _3757_/Z _3758_/A4 _3758_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_174_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6477_ _6971_/Q _6262_/Z _6499_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_118_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3689_ _3689_/A1 _3657_/Z _3688_/Z _6569_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_5428_ _5381_/I _5428_/A2 _6577_/C _5428_/A4 _5428_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_160_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput240 _6750_/Q mgmt_gpio_out[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput251 _4080_/Z pad_flash_io0_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput262 _6878_/Q pll_div[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput273 _6677_/Q pll_trim[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput284 _6671_/Q pll_trim[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_87_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5359_ _5359_/A1 _4892_/B _5360_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xoutput295 _6674_/Q pll_trim[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_58_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7029_ _7029_/D _6821_/RN _7029_/CLK _7029_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_75_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet852_104 net852_136/I _7121_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_115 _4073__51/I _7110_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet852_126 _4073__23/I _7099_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_137 _4073__41/I _7088_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_148 net852_149/I _7077_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4730_ _5226_/A1 _4728_/Z _5105_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_1480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4661_ _4414_/Z _5038_/A1 _5020_/A2 _4557_/Z _4662_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_159_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6400_ _7210_/Q _6535_/A2 _6545_/A2 _6936_/Q _6401_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3612_ _6680_/Q _3546_/Z _3625_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_156_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4592_ _4565_/Z _4586_/Z _5018_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold904 _4150_/Z _6698_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6331_ _6331_/I _6332_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3543_ _5857_/A1 _5830_/A1 _3543_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold915 _7029_/Q hold915/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold926 _4152_/Z _6700_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold937 _6982_/Q hold937/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold948 _5700_/Z _7051_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold959 _6988_/Q hold959/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6262_ _6302_/A3 _6300_/A4 _6300_/A1 _6275_/A4 _6262_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3474_ _4041_/B1 _6660_/Q _3981_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_131_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5213_ _4673_/Z _5124_/B _5213_/B _5213_/C _5454_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_131_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6193_ _6193_/A1 _6193_/A2 _6193_/A3 _6193_/A4 _6193_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_142_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5144_ _4555_/C _5276_/C _5145_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_85_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5075_ _5255_/B _5051_/Z _5075_/B _5076_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4026_ _4402_/B _4395_/B _4026_/B _4026_/C _4412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_52_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5977_ _6996_/Q _6211_/B1 _6021_/A2 _3387_/I _5977_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_80_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4928_ _4376_/Z _5442_/A1 _5323_/B _5442_/A4 _4928_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_60_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4859_ _5478_/A1 _4873_/A2 _4873_/A3 _4681_/Z _4859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_165_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6529_ _6529_/I0 _7258_/Q _6529_/S _6529_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5900_ _5900_/A1 _5954_/A3 _5951_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_34_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6880_ hold77/Z _6882_/RN _6880_/CLK hold76/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_5831_ _5885_/I0 hold873/Z _5838_/S _5831_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5762_ hold479/Z _5888_/I0 _5766_/S _7105_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4713_ _4713_/A1 _5094_/B _4691_/Z _5403_/A1 _5305_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_147_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5693_ _5804_/I0 _5693_/I1 _5700_/S _5693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4644_ _4644_/A1 _5038_/B _4643_/Z _4653_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_129_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold701 _7189_/Q hold701/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4575_ _4652_/A4 _4539_/I _5373_/A2 _4643_/A4 _5192_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold712 _5891_/Z _7220_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold723 _6980_/Q hold723/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6314_ _7053_/Q _6299_/Z _6328_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3526_ _3552_/A2 _3484_/Z hold27/Z hold28/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xhold734 _5846_/Z _7180_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold745 _6932_/Q hold745/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7294_ _7294_/D _6648_/Z _7304_/CLK _7294_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_1_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold756 _5563_/Z _6929_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold767 _6840_/Q hold767/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_118_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold778 _5538_/Z _6907_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_157_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6245_ _7233_/Q _6275_/A4 _6452_/A4 _6279_/A3 _6245_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_157_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold789 _7027_/Q hold789/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3457_ hold18/Z hold58/Z _3460_/S _7287_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6176_ _5991_/Z _6176_/A2 _6176_/B _6176_/C _6177_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3388_ _7230_/Q _6014_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_57_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5127_ _5127_/A1 _5457_/A1 _5213_/B _5127_/A4 _5127_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5058_ _5058_/A1 _5055_/Z _5193_/A2 _5058_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XTAP_2906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4009_ _4009_/A1 _3324_/I _4009_/B _4010_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_2928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet802_53 net802_53/I _7172_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet802_64 net802_64/I _7161_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet802_75 net802_75/I _7150_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet802_86 net802_87/I _7139_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet802_97 net802_97/I _7128_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold50 hold50/I hold50/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_76_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold61 hold61/I hold61/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xclkbuf_leaf_25__1359_ _4073__6/I net852_136/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold72 hold72/I hold72/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xclkbuf_leaf_105__1359_ clkbuf_4_4_0__1359_/Z net952_209/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold83 hold83/I hold83/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_48_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold94 hold94/I hold94/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xclkbuf_leaf_88__1359_ clkbuf_4_7_0__1359_/Z net952_227/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_91_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_3 _5645_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4360_ hold544/Z _4360_/I1 _4361_/S _4360_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3311_ _6730_/Q _3442_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_4291_ hold823/Z _6613_/I1 _4291_/S _4291_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6030_ _6030_/A1 _6030_/A2 _6030_/A3 _6030_/A4 _6030_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_39_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6932_ _6932_/D _7140_/RN _6932_/CLK _6932_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_35_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6863_ _6863_/D _6865_/RN _6865_/CLK _6863_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5814_ _5832_/I0 hold969/Z _5820_/S _5814_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6794_ _6794_/D _7258_/CLK _6794_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5745_ _5871_/I0 hold511/Z _5748_/S _5745_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5676_ hold915/Z _5877_/I0 _5682_/S _5676_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4627_ _4627_/A1 _4625_/Z _4626_/Z _4633_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xhold520 _5625_/Z _6984_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold531 _6843_/Q hold531/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4558_ _5038_/A1 _4557_/Z _5393_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold542 _6937_/Q hold542/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold553 _5679_/Z _7032_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_1_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold564 _5783_/Z _7124_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_132_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold575 _7004_/Q hold575/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3509_ _5620_/A4 _3481_/I _3484_/Z hold27/Z _3509_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_143_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold586 _7179_/Q hold586/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4489_ _4489_/A1 _4692_/B _4489_/B _4491_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7277_ _7277_/D _7278_/RN _7279_/CLK _7277_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold597 _4352_/Z _6852_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ _6228_/A1 _6228_/A2 _6228_/A3 _6227_/Z _6228_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_106_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6159_ _6147_/Z _6158_/Z _6473_/B1 _6118_/B _6500_/C _6160_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_66_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput140 wb_dat_i[20] _6591_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput151 wb_dat_i[30] _6597_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput162 wb_sel_i[1] _6574_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3860_ _3860_/A1 _3860_/A2 _3860_/A3 _3860_/A4 _3860_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_147_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3791_ _6950_/Q _5584_/A1 _5575_/A1 _6942_/Q _3925_/A2 input5/Z _3794_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XPHY_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5530_ _5857_/A1 _5839_/A3 hold212/Z _5857_/A4 _5531_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_185_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5461_ _5461_/I _5480_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7200_ _7200_/D fanout677/Z _7200_/CLK _7200_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_173_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4412_ _4412_/A1 _4399_/Z _4412_/B _4412_/C _5209_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_5392_ _5051_/S _5360_/B _5392_/B _5433_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_132_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4343_ _4343_/I0 hold557/Z _4343_/S _4343_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7131_ _7131_/D _7188_/RN _7131_/CLK _7131_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_67_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7062_ _7062_/D _7075_/RN _7062_/CLK _7062_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4274_ _4274_/A1 _6611_/A2 _4276_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_59_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6013_ _6013_/A1 _5991_/Z _6027_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_98_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_71__1359_ clkbuf_4_14_0__1359_/Z _4073__12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6915_ _6915_/D _6915_/RN _6915_/CLK _6915_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6846_ _6846_/D _6886_/RN _6846_/CLK _6846_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_50_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6777_ _6777_/D _6894_/RN _6777_/CLK _6777_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3989_ _7239_/Q _6895_/Q _6900_/Q _3990_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_5728_ _5728_/A1 _6611_/A2 _5730_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_148_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5659_ hold967/Z _5806_/I0 _5664_/S _5659_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold350 _4123_/Z _6677_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold361 _7005_/Q hold361/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold372 _5650_/Z _7006_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold383 _6752_/Q hold383/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold394 _7119_/Q hold394/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_104_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1050 _6966_/Q _5605_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1061 _6917_/Q _4232_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold1072 _7293_/Q _3447_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XTAP_3234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4961_ _4500_/Z _4906_/Z _4973_/A4 _5020_/A2 _4961_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_45_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6700_ _6700_/D _7207_/RN _6700_/CLK _6700_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_3912_ _7214_/Q _3912_/A2 _3912_/B1 _6883_/Q _3912_/C1 _6706_/Q _3915_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_4892_ _4990_/A1 _5329_/A2 _4892_/B _4894_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_32_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6631_ _7162_/RN _6652_/A2 _6631_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3843_ _4353_/A1 _3617_/Z _3950_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xnet1202_460 net802_94/I _6705_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1202_471 net1202_471/I _6694_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1202_482 net1202_483/I _6683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3774_ _6926_/Q _3935_/A2 _3945_/C2 _6684_/Q _5701_/A1 _7054_/Q _3776_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6562_ _6562_/I _7261_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet1202_493 net802_84/I _6672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5513_ _5520_/C _5517_/A2 hold146/Z _5517_/A1 _5514_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_146_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6493_ _6493_/A1 _6493_/A2 _6486_/Z _6492_/Z _6493_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_173_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5444_ _5444_/A1 _5444_/A2 _5442_/Z _5444_/A4 _5483_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_172_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5375_ _5421_/A2 _5470_/A1 _5372_/Z _5374_/Z _5379_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_160_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7114_ _7114_/D _7215_/RN _7114_/CLK _7114_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4326_ _4332_/A1 _5517_/A1 _5517_/A3 _5794_/A3 _4328_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7045_ _7045_/D _7098_/RN _7045_/CLK _7045_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4257_ hold60/Z hold96/Z _4261_/S hold97/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4188_ _4188_/A1 _6611_/A2 _4190_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_41_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4073__9 _4073__9/I _7216_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6829_ _6829_/D _7261_/RN _7279_/CLK _6829_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold180 _5713_/Z _7062_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold191 _6903_/Q hold191/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_2_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout660 _7146_/RN _7140_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout671 _7171_/RN _7083_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xfanout682 _7019_/RN _6967_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_59_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout693 _7205_/RN _7220_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_92_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3490_ _7305_/Q _3490_/I1 _3984_/S _3491_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5160_ _5287_/B _5293_/B _5164_/A4 _5160_/B _5366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_170_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4111_ hold18/Z _7274_/Q _4113_/S hold19/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5091_ _5367_/A2 _5307_/A3 _5228_/A3 _5095_/B1 _5222_/A1 _5103_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_68_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4042_ _7291_/Q _3409_/Z _4042_/A3 _4043_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_68_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5993_ _3385_/I _3386_/I _3387_/I _6164_/B1 _5994_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_64_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4944_ _4944_/A1 _4495_/Z _4976_/A3 _4759_/Z _4944_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_80_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4875_ _4651_/Z _5142_/A3 _4876_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_32_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6614_ _7188_/RN _6657_/A2 _6614_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3826_ _3844_/A1 _3560_/Z _3934_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_178_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6545_ _6788_/Q _6545_/A2 _6545_/B1 _6844_/Q _6546_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3757_ _3757_/A1 _3757_/A2 _3757_/A3 _3757_/A4 _3757_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_118_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6476_ _7257_/Q _6476_/I1 _6476_/S _7257_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3688_ _3688_/A1 _3663_/Z _3674_/Z _3687_/Z _3688_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_161_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5427_ _5427_/A1 _5425_/Z _5426_/Z _4881_/Z _5430_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xoutput230 _6913_/Q mgmt_gpio_out[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput241 _6751_/Q mgmt_gpio_out[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_88_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput252 _4079_/ZN pad_flash_io0_ie VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput263 _6879_/Q pll_div[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput274 _6678_/Q pll_trim[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput285 hold48/I pll_trim[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5358_ _5432_/A1 _5189_/Z _5355_/Z _5357_/Z _5362_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput296 _6675_/Q pll_trim[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4309_ _6568_/I0 _6815_/Q _4312_/S _6815_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5289_ _5029_/B _5289_/A2 _5289_/A3 _5292_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_102_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7028_ _7028_/D _7090_/RN _7028_/CLK _7028_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_101_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet852_105 net802_81/I _7120_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet852_116 _4073__12/I _7109_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_127 net902_157/I _7098_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout490 _5547_/I0 _5775_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xnet852_138 net852_138/I _7087_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet852_149 net852_149/I _7076_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4660_ _4376_/Z _4411_/Z _5172_/B _5165_/A4 _5385_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_159_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3611_ _3610_/Z _3611_/I1 _3899_/S _6875_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4591_ _4591_/A1 _4587_/Z _4590_/Z _4593_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_162_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6330_ _7005_/Q _6549_/B1 _6552_/A2 _7029_/Q _7119_/Q _6288_/Z _6331_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_155_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold905 _7060_/Q hold905/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3542_ _3653_/A1 _3904_/A3 _3680_/A3 hold211/I _3542_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold916 _5676_/Z _7029_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_183_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold927 _7088_/Q hold927/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_143_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold938 _5623_/Z _6982_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold949 _6974_/Q hold949/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_89_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6261_ _6300_/A1 _6275_/A4 _6533_/A3 _6300_/A4 _6261_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3473_ _3471_/I _5490_/A1 _3500_/S _3473_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5212_ _5242_/A3 _4810_/B _4812_/B _5212_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_142_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ _6718_/Q _5960_/Z _6192_/B _6193_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_9_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5143_ _4820_/Z _4821_/Z _4878_/Z _5278_/B _5372_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_9_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5074_ _5074_/A1 _5408_/C _5072_/Z _5335_/C _5075_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_69_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4025_ _4489_/B _4424_/B _4034_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_37_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5976_ _6015_/A3 _6211_/B1 _7004_/Q _3386_/I _5976_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_40_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4927_ _4927_/A1 _4927_/A2 _4927_/A3 _4929_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_100_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4858_ _4858_/A1 _4858_/A2 _5289_/A2 _4862_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_166_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3809_ _4332_/A1 _3617_/Z _4289_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_121_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4789_ _5270_/A1 _4808_/A2 _4530_/I _5302_/B _4789_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_119_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6528_ _6516_/Z _6527_/Z _6528_/B1 _6286_/Z _6529_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_181_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6459_ _6459_/I _6460_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_48__1359_ clkbuf_4_11_0__1359_/Z net802_93/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_128__1359_ clkbuf_4_4_0__1359_/Z net1202_485/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_109_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5830_ _5830_/A1 _5839_/A2 _5857_/A4 _5838_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_61_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5761_ hold432/Z _5806_/I0 _5766_/S _5761_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4712_ _4687_/Z _5092_/A1 _4713_/A1 _4691_/Z _5222_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5692_ _5692_/A1 _5830_/A1 _5866_/A3 _5700_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_175_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4643_ _5315_/A1 _5164_/A2 _5146_/A1 _4643_/A4 _4643_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_163_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4574_ _5278_/C _4990_/A1 _5370_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold702 _5856_/Z _7189_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold713 _7074_/Q hold713/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold724 _5621_/Z _6980_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6313_ _6997_/Q _6549_/C1 _6545_/B1 _7013_/Q _6329_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_144_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold735 _7077_/Q hold735/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3525_ _3653_/A1 _3904_/A3 hold144/I hold211/I _3525_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold746 _5567_/Z _6932_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_7293_ _7293_/D _6647_/Z _7302_/CLK _7293_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold757 _6786_/Q hold757/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_131_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold768 _4334_/Z _6840_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_131_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold779 _6987_/Q hold779/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6244_ _3328_/I _6296_/A2 _6282_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3456_ hold38/Z hold18/Z _3460_/S _7288_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3387_ _3387_/I _6015_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_6175_ _6955_/Q _5958_/Z _5994_/I _7141_/Q _6176_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_85_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5126_ _5126_/I _5127_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5057_ _5078_/A2 _5443_/A1 _5057_/B _5324_/C _5058_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_44_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4008_ _4008_/I _4009_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_2918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet802_54 net802_54/I _7171_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet802_65 net802_97/I _7160_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet802_76 net802_76/I _7149_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet802_87 net802_87/I _7138_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet802_98 net802_98/I _7127_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5959_ _6014_/A2 _5984_/A1 _5959_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_138_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold40 hold40/I hold40/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_29_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold51 hold51/I hold51/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold62 hold62/I hold62/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold73 hold73/I hold73/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold84 hold84/I hold84/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_60_1070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold95 hold95/I hold95/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_63_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_4 _3477_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3310_ hold26/Z _5490_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_140_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4290_ hold853/Z _6612_/I1 _4291_/S _4290_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_15_0__1359_ clkbuf_0__1359_/Z clkbuf_4_15_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_13_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6931_ _6931_/D _7034_/RN _6931_/CLK _6931_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6862_ _6862_/D _6865_/RN _6865_/CLK _6862_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_179_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5813_ _4103_/I hold991/Z _5820_/S _5813_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6793_ _6793_/D _7258_/CLK _6793_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5744_ _5888_/I0 hold448/Z _5748_/S _5744_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5675_ hold461/Z _5876_/I0 _5682_/S _5675_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4626_ _4887_/A1 _4868_/A1 _5146_/A1 _4635_/A4 _4626_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold510 _4187_/Z _6725_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold521 _6945_/Q hold521/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xclkbuf_leaf_111__1359_ clkbuf_4_4_0__1359_/Z net1202_499/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_31__1359_ clkbuf_opt_5_0__1359_/Z net1052_312/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4557_ _4436_/B _4648_/A1 _4648_/A2 _4557_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
Xhold532 _4339_/Z _6843_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold543 _5572_/Z _6937_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
XFILLER_116_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_94__1359_ clkbuf_4_5_0__1359_/Z net952_250/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold554 _7001_/Q hold554/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold565 _6889_/Q hold565/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_3508_ hold27/Z _3481_/I _3484_/Z _3508_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_7276_ _7276_/D _7278_/RN _7279_/CLK _7276_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold576 _5648_/Z _7004_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_4488_ _4392_/Z _4474_/Z _4722_/A2 _4923_/A2 _4491_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold587 _5845_/Z _7179_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
Xhold598 _6997_/Q hold598/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_4
X_6227_ _6227_/A1 _6227_/A2 _6227_/A3 _6227_/A4 _6227_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3439_ _3971_/A1 _3442_/B _6665_/Q _6664_/Q _3440_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_44_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6158_ _6152_/Z _6155_/Z _6158_/A3 _6158_/A4 _6158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5109_ _5108_/Z _4853_/Z _4740_/Z _5111_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6089_ _7244_/Q _6089_/I1 _6558_/S _7244_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput130 wb_dat_i[11] _6588_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput141 wb_dat_i[21] _6594_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput152 wb_dat_i[31] _6600_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput163 wb_sel_i[2] _6573_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3790_ _3790_/A1 _3790_/A2 _3790_/A3 _3790_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XPHY_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5460_ _5460_/A1 _5303_/Z _5460_/A3 _5460_/A4 _5461_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_8_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _5083_/B _4412_/B _4412_/C _4411_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_5391_ _5388_/Z _4985_/Z _5386_/Z _5390_/Z _5391_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_172_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7130_ _7130_/D _7207_/RN _7130_/CLK _7130_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_113_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4342_ _4360_/I1 hold517/Z _4343_/S _4342_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7061_ _7061_/D _7090_/RN _7061_/CLK _7061_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_113_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4273_ _5859_/I0 hold757/Z _4273_/S _4273_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6012_ _7021_/Q _6211_/A2 _6164_/B1 _6989_/Q _6013_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_154_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

