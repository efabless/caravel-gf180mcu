VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gpio_defaults_block_087
  CLASS BLOCK ;
  FOREIGN gpio_defaults_block_087 ;
  ORIGIN 0.430 0.430 ;
  SIZE 19.900 BY 16.540 ;
  PIN gpio_defaults[0]
    PORT
      LAYER Metal1 ;
        RECT 2.340 2.210 2.700 3.390 ;
        RECT 2.340 1.850 3.365 2.210 ;
        RECT 2.990 0.580 3.365 1.850 ;
      LAYER Via1 ;
        RECT 3.025 1.245 3.325 1.545 ;
      LAYER Metal2 ;
        RECT 2.860 1.235 5.020 1.555 ;
        RECT 3.500 -0.420 3.780 1.235 ;
    END
  END gpio_defaults[0]
  PIN gpio_defaults[4]
    PORT
      LAYER Metal1 ;
        RECT 11.300 0.530 11.675 1.650 ;
      LAYER Via1 ;
        RECT 11.335 1.245 11.635 1.545 ;
      LAYER Metal2 ;
        RECT 9.575 1.235 11.740 1.555 ;
        RECT 10.220 -0.420 10.500 1.235 ;
    END
  END gpio_defaults[4]
  PIN gpio_defaults[8]
    PORT
      LAYER Metal1 ;
        RECT 16.900 0.530 17.275 1.650 ;
      LAYER Via1 ;
        RECT 16.935 1.245 17.235 1.545 ;
      LAYER Metal2 ;
        RECT 15.215 1.235 17.310 1.555 ;
        RECT 16.940 -0.420 17.220 1.235 ;
    END
  END gpio_defaults[8]
  PIN gpio_defaults[7]
    PORT
      LAYER Metal1 ;
        RECT 14.660 10.050 15.020 11.230 ;
        RECT 14.660 9.690 15.685 10.050 ;
        RECT 15.310 8.420 15.685 9.690 ;
      LAYER Via1 ;
        RECT 15.345 9.085 15.645 9.385 ;
      LAYER Metal2 ;
        RECT 14.605 9.385 17.340 9.395 ;
        RECT 14.605 9.085 16.935 9.385 ;
        RECT 17.235 9.085 17.340 9.385 ;
        RECT 14.605 9.075 17.340 9.085 ;
        RECT 14.605 0.885 14.885 9.075 ;
        RECT 14.605 0.605 15.540 0.885 ;
        RECT 15.260 -0.420 15.540 0.605 ;
    END
  END gpio_defaults[7]
  PIN gpio_defaults[1]
    PORT
      LAYER Metal1 ;
        RECT 2.990 5.990 3.365 7.260 ;
        RECT 2.340 5.630 3.365 5.990 ;
        RECT 2.340 4.450 2.700 5.630 ;
      LAYER Via1 ;
        RECT 3.025 6.295 3.325 6.595 ;
      LAYER Metal2 ;
        RECT 2.925 6.285 5.660 6.605 ;
        RECT 5.380 0.785 5.660 6.285 ;
        RECT 5.180 0.485 5.660 0.785 ;
        RECT 5.180 -0.420 5.460 0.485 ;
    END
  END gpio_defaults[1]
  PIN gpio_defaults[5]
    PORT
      LAYER Metal1 ;
        RECT 11.300 6.190 11.675 7.310 ;
      LAYER Via1 ;
        RECT 11.335 6.295 11.635 6.595 ;
      LAYER Metal2 ;
        RECT 9.645 6.285 12.480 6.605 ;
        RECT 12.200 0.870 12.480 6.285 ;
        RECT 11.900 0.590 12.480 0.870 ;
        RECT 11.900 -0.420 12.180 0.590 ;
    END
  END gpio_defaults[5]
  PIN gpio_defaults[9]
    PORT
      LAYER Metal1 ;
        RECT 16.900 6.190 17.275 7.310 ;
      LAYER Via1 ;
        RECT 16.935 6.295 17.235 6.595 ;
      LAYER Metal2 ;
        RECT 15.205 6.285 18.900 6.605 ;
        RECT 18.620 -0.420 18.900 6.285 ;
    END
  END gpio_defaults[9]
  PIN gpio_defaults[3]
    PORT
      LAYER Metal1 ;
        RECT 4.580 14.030 4.955 15.150 ;
      LAYER Via1 ;
        RECT 4.615 14.135 4.915 14.435 ;
      LAYER Metal2 ;
        RECT 2.880 14.125 8.495 14.445 ;
        RECT 8.215 2.480 8.495 14.125 ;
        RECT 8.215 2.200 8.820 2.480 ;
        RECT 8.540 -0.420 8.820 2.200 ;
    END
  END gpio_defaults[3]
  PIN gpio_defaults[2]
    PORT
      LAYER Metal1 ;
        RECT 2.340 10.050 2.700 11.230 ;
        RECT 2.340 9.690 3.365 10.050 ;
        RECT 2.990 8.420 3.365 9.690 ;
      LAYER Via1 ;
        RECT 3.025 9.085 3.325 9.385 ;
      LAYER Metal2 ;
        RECT 2.925 9.075 7.140 9.395 ;
        RECT 6.860 -0.420 7.140 9.075 ;
    END
  END gpio_defaults[2]
  PIN gpio_defaults[6]
    PORT
      LAYER Metal1 ;
        RECT 11.300 8.370 11.675 9.490 ;
      LAYER Via1 ;
        RECT 11.335 9.085 11.635 9.385 ;
      LAYER Metal2 ;
        RECT 9.645 9.075 13.860 9.395 ;
        RECT 13.580 -0.420 13.860 9.075 ;
    END
  END gpio_defaults[6]
  PIN VDD
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0.370 12.060 0.710 13.760 ;
        RECT 1.370 12.060 1.600 13.320 ;
        RECT 3.705 12.060 3.935 13.335 ;
        RECT 7.365 12.060 7.595 13.190 ;
        RECT 9.605 12.060 9.835 13.190 ;
        RECT 11.845 12.060 12.075 13.190 ;
        RECT 12.690 12.060 13.030 13.760 ;
        RECT 15.205 12.060 15.435 13.190 ;
        RECT 17.445 12.060 17.675 13.190 ;
        RECT 18.290 12.060 18.630 13.760 ;
        RECT 0.000 11.460 19.040 12.060 ;
        RECT 0.370 9.760 0.710 11.460 ;
        RECT 1.370 10.200 1.600 11.460 ;
        RECT 3.705 10.185 3.935 11.460 ;
        RECT 7.365 10.330 7.595 11.460 ;
        RECT 8.090 10.200 8.320 11.460 ;
        RECT 10.425 10.185 10.655 11.460 ;
        RECT 12.690 9.760 13.030 11.460 ;
        RECT 13.690 10.200 13.920 11.460 ;
        RECT 16.025 10.185 16.255 11.460 ;
        RECT 18.290 9.760 18.630 11.460 ;
        RECT 0.390 4.220 0.730 5.910 ;
        RECT 1.370 4.220 1.600 5.480 ;
        RECT 3.705 4.220 3.935 5.495 ;
        RECT 7.365 4.220 7.595 5.350 ;
        RECT 8.090 4.220 8.320 5.480 ;
        RECT 10.425 4.220 10.655 5.495 ;
        RECT 12.710 4.220 13.050 5.910 ;
        RECT 13.690 4.220 13.920 5.480 ;
        RECT 16.025 4.220 16.255 5.495 ;
        RECT 18.310 4.220 18.650 5.910 ;
        RECT 0.000 3.620 19.040 4.220 ;
        RECT 0.370 1.920 0.710 3.620 ;
        RECT 1.370 2.360 1.600 3.620 ;
        RECT 3.705 2.345 3.935 3.620 ;
        RECT 7.365 2.490 7.595 3.620 ;
        RECT 8.090 2.360 8.320 3.620 ;
        RECT 10.425 2.345 10.655 3.620 ;
        RECT 12.710 1.930 13.050 3.620 ;
        RECT 13.690 2.360 13.920 3.620 ;
        RECT 16.025 2.345 16.255 3.620 ;
        RECT 18.310 1.930 18.650 3.620 ;
      LAYER Via1 ;
        RECT 8.965 11.650 11.810 11.950 ;
        RECT 8.965 3.750 11.810 4.050 ;
      LAYER Metal2 ;
        RECT 8.900 11.590 11.880 12.005 ;
        RECT 8.900 3.690 11.880 4.105 ;
      LAYER Via2 ;
        RECT 8.965 11.650 11.810 11.950 ;
        RECT 8.965 3.750 11.810 4.050 ;
      LAYER Metal3 ;
        RECT 8.865 -0.265 11.895 15.960 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 15.380 19.040 15.980 ;
        RECT 0.370 14.490 0.710 15.380 ;
        RECT 1.370 14.520 1.600 15.380 ;
        RECT 3.605 14.520 3.835 15.380 ;
        RECT 5.845 14.585 6.075 15.380 ;
        RECT 8.085 14.585 8.315 15.380 ;
        RECT 10.325 14.585 10.555 15.380 ;
        RECT 12.690 14.490 13.030 15.380 ;
        RECT 13.685 14.585 13.915 15.380 ;
        RECT 15.925 14.585 16.155 15.380 ;
        RECT 18.290 14.490 18.630 15.380 ;
        RECT 0.370 8.140 0.710 9.030 ;
        RECT 1.370 8.140 1.600 9.000 ;
        RECT 3.605 8.140 3.835 9.000 ;
        RECT 5.845 8.140 6.075 8.935 ;
        RECT 8.090 8.140 8.320 9.000 ;
        RECT 10.325 8.140 10.555 9.000 ;
        RECT 12.690 8.140 13.030 9.030 ;
        RECT 13.690 8.140 13.920 9.000 ;
        RECT 15.925 8.140 16.155 9.000 ;
        RECT 18.290 8.140 18.630 9.030 ;
        RECT 0.000 7.540 19.040 8.140 ;
        RECT 0.390 6.655 0.730 7.540 ;
        RECT 1.370 6.680 1.600 7.540 ;
        RECT 3.605 6.680 3.835 7.540 ;
        RECT 5.845 6.745 6.075 7.540 ;
        RECT 8.090 6.680 8.320 7.540 ;
        RECT 10.325 6.680 10.555 7.540 ;
        RECT 12.710 6.655 13.050 7.540 ;
        RECT 13.690 6.680 13.920 7.540 ;
        RECT 15.925 6.680 16.155 7.540 ;
        RECT 18.310 6.655 18.650 7.540 ;
        RECT 0.370 0.300 0.710 1.190 ;
        RECT 1.370 0.300 1.600 1.160 ;
        RECT 3.605 0.300 3.835 1.160 ;
        RECT 5.845 0.300 6.075 1.095 ;
        RECT 8.090 0.300 8.320 1.160 ;
        RECT 10.325 0.300 10.555 1.160 ;
        RECT 12.710 0.300 13.050 1.185 ;
        RECT 13.690 0.300 13.920 1.160 ;
        RECT 15.925 0.300 16.155 1.160 ;
        RECT 18.310 0.300 18.650 1.185 ;
        RECT 0.000 -0.300 19.040 0.300 ;
      LAYER Via1 ;
        RECT 0.415 15.550 3.260 15.850 ;
        RECT 0.415 7.700 3.260 8.000 ;
        RECT 0.460 -0.145 3.105 0.155 ;
      LAYER Metal2 ;
        RECT 0.350 15.490 3.330 15.905 ;
        RECT 0.350 7.640 3.330 8.055 ;
        RECT 0.400 -0.200 3.165 0.215 ;
      LAYER Via2 ;
        RECT 0.415 15.550 3.260 15.850 ;
        RECT 0.415 7.700 3.260 8.000 ;
        RECT 0.460 -0.145 3.105 0.155 ;
      LAYER Metal3 ;
        RECT 0.330 -0.265 3.360 15.960 ;
    END
  END VSS
  OBS
      LAYER Pwell ;
        RECT -0.430 13.920 19.470 16.110 ;
      LAYER Nwell ;
        RECT -0.430 9.600 19.470 13.920 ;
      LAYER Pwell ;
        RECT -0.430 6.080 19.470 9.600 ;
      LAYER Nwell ;
        RECT -0.430 1.760 19.470 6.080 ;
      LAYER Pwell ;
        RECT -0.430 -0.430 19.470 1.760 ;
      LAYER Metal1 ;
        RECT 2.490 14.345 2.720 15.150 ;
        RECT 1.995 14.110 2.720 14.345 ;
      LAYER Metal1 ;
        RECT 2.990 13.830 3.365 15.100 ;
        RECT 2.340 13.470 3.365 13.830 ;
      LAYER Metal1 ;
        RECT 5.845 14.125 7.120 14.355 ;
        RECT 4.230 13.495 4.955 13.730 ;
      LAYER Metal1 ;
        RECT 2.340 12.290 2.700 13.470 ;
      LAYER Metal1 ;
        RECT 4.725 12.290 4.955 13.495 ;
        RECT 5.845 12.290 6.075 14.125 ;
        RECT 7.365 13.720 7.595 15.150 ;
        RECT 6.330 13.490 7.595 13.720 ;
        RECT 8.085 14.125 9.360 14.355 ;
        RECT 8.085 12.290 8.315 14.125 ;
        RECT 9.605 13.720 9.835 15.150 ;
        RECT 8.570 13.490 9.835 13.720 ;
        RECT 10.325 14.125 11.600 14.355 ;
        RECT 10.325 12.290 10.555 14.125 ;
        RECT 11.845 13.720 12.075 15.150 ;
        RECT 10.810 13.490 12.075 13.720 ;
        RECT 13.685 14.125 14.960 14.355 ;
        RECT 13.685 12.290 13.915 14.125 ;
        RECT 15.205 13.720 15.435 15.150 ;
        RECT 14.170 13.490 15.435 13.720 ;
        RECT 15.925 14.125 17.200 14.355 ;
        RECT 15.925 12.290 16.155 14.125 ;
        RECT 17.445 13.720 17.675 15.150 ;
        RECT 16.410 13.490 17.675 13.720 ;
        RECT 4.725 10.025 4.955 11.230 ;
        RECT 4.230 9.790 4.955 10.025 ;
        RECT 1.995 9.175 2.720 9.410 ;
        RECT 2.490 8.370 2.720 9.175 ;
      LAYER Metal1 ;
        RECT 4.580 8.370 4.955 9.490 ;
      LAYER Metal1 ;
        RECT 5.845 9.395 6.075 11.230 ;
      LAYER Metal1 ;
        RECT 9.060 10.050 9.420 11.230 ;
      LAYER Metal1 ;
        RECT 6.330 9.800 7.595 10.030 ;
        RECT 5.845 9.165 7.120 9.395 ;
        RECT 7.365 8.370 7.595 9.800 ;
      LAYER Metal1 ;
        RECT 9.060 9.690 10.085 10.050 ;
      LAYER Metal1 ;
        RECT 11.445 10.025 11.675 11.230 ;
        RECT 17.045 10.025 17.275 11.230 ;
        RECT 10.950 9.790 11.675 10.025 ;
        RECT 16.550 9.790 17.275 10.025 ;
        RECT 8.715 9.175 9.440 9.410 ;
        RECT 9.210 8.370 9.440 9.175 ;
      LAYER Metal1 ;
        RECT 9.710 8.420 10.085 9.690 ;
      LAYER Metal1 ;
        RECT 14.315 9.175 15.040 9.410 ;
        RECT 14.810 8.370 15.040 9.175 ;
      LAYER Metal1 ;
        RECT 16.900 8.370 17.275 9.490 ;
      LAYER Metal1 ;
        RECT 2.490 6.505 2.720 7.310 ;
        RECT 1.995 6.270 2.720 6.505 ;
      LAYER Metal1 ;
        RECT 4.580 6.190 4.955 7.310 ;
      LAYER Metal1 ;
        RECT 5.845 6.285 7.120 6.515 ;
        RECT 4.230 5.655 4.955 5.890 ;
        RECT 4.725 4.450 4.955 5.655 ;
        RECT 5.845 4.450 6.075 6.285 ;
        RECT 7.365 5.880 7.595 7.310 ;
        RECT 9.210 6.505 9.440 7.310 ;
        RECT 8.715 6.270 9.440 6.505 ;
      LAYER Metal1 ;
        RECT 9.710 5.990 10.085 7.260 ;
      LAYER Metal1 ;
        RECT 14.810 6.505 15.040 7.310 ;
        RECT 14.315 6.270 15.040 6.505 ;
      LAYER Metal1 ;
        RECT 15.310 5.990 15.685 7.260 ;
      LAYER Metal1 ;
        RECT 6.330 5.650 7.595 5.880 ;
      LAYER Metal1 ;
        RECT 9.060 5.630 10.085 5.990 ;
      LAYER Metal1 ;
        RECT 10.950 5.655 11.675 5.890 ;
      LAYER Metal1 ;
        RECT 9.060 4.450 9.420 5.630 ;
      LAYER Metal1 ;
        RECT 11.445 4.450 11.675 5.655 ;
      LAYER Metal1 ;
        RECT 14.660 5.630 15.685 5.990 ;
      LAYER Metal1 ;
        RECT 16.550 5.655 17.275 5.890 ;
      LAYER Metal1 ;
        RECT 14.660 4.450 15.020 5.630 ;
      LAYER Metal1 ;
        RECT 17.045 4.450 17.275 5.655 ;
        RECT 4.725 2.185 4.955 3.390 ;
        RECT 4.230 1.950 4.955 2.185 ;
        RECT 1.995 1.335 2.720 1.570 ;
        RECT 2.490 0.530 2.720 1.335 ;
      LAYER Metal1 ;
        RECT 4.580 0.530 4.955 1.650 ;
      LAYER Metal1 ;
        RECT 5.845 1.555 6.075 3.390 ;
      LAYER Metal1 ;
        RECT 9.060 2.210 9.420 3.390 ;
      LAYER Metal1 ;
        RECT 6.330 1.960 7.595 2.190 ;
        RECT 5.845 1.325 7.120 1.555 ;
        RECT 7.365 0.530 7.595 1.960 ;
      LAYER Metal1 ;
        RECT 9.060 1.850 10.085 2.210 ;
      LAYER Metal1 ;
        RECT 11.445 2.185 11.675 3.390 ;
        RECT 10.950 1.950 11.675 2.185 ;
      LAYER Metal1 ;
        RECT 14.660 2.210 15.020 3.390 ;
        RECT 14.660 1.850 15.685 2.210 ;
      LAYER Metal1 ;
        RECT 17.045 2.185 17.275 3.390 ;
        RECT 16.550 1.950 17.275 2.185 ;
        RECT 8.715 1.335 9.440 1.570 ;
        RECT 9.210 0.530 9.440 1.335 ;
      LAYER Metal1 ;
        RECT 9.710 0.580 10.085 1.850 ;
      LAYER Metal1 ;
        RECT 14.315 1.335 15.040 1.570 ;
        RECT 14.810 0.530 15.040 1.335 ;
      LAYER Metal1 ;
        RECT 15.310 0.580 15.685 1.850 ;
  END
END gpio_defaults_block_087
END LIBRARY

