* NGSPICE file created from housekeeping.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_4 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_4 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_4 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_4 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_20 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_12 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 D RN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 D SETN CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_8 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

.subckt housekeeping VDD VSS debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oe
+ pad_flash_csb pad_flash_csb_oe pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ie
+ pad_flash_io0_oe pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ie pad_flash_io1_oe
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out qspi_enabled reset
+ ser_rx ser_tx serial_clock serial_data_1 serial_data_2 serial_load serial_resetn
+ spi_csb spi_enabled spi_sck spi_sdi spi_sdo spi_sdoenb spimemio_flash_clk spimemio_flash_csb
+ spimemio_flash_io0_di spimemio_flash_io0_do spimemio_flash_io0_oeb spimemio_flash_io1_di
+ spimemio_flash_io1_do spimemio_flash_io1_oeb spimemio_flash_io2_di spimemio_flash_io2_do
+ spimemio_flash_io2_oeb spimemio_flash_io3_di spimemio_flash_io3_do spimemio_flash_io3_oeb
+ trap uart_enabled user_clock wb_ack_o wb_adr_i[0] wb_adr_i[10] wb_adr_i[11] wb_adr_i[12]
+ wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17] wb_adr_i[18] wb_adr_i[19]
+ wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23] wb_adr_i[24] wb_adr_i[25]
+ wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2] wb_adr_i[30] wb_adr_i[31]
+ wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7] wb_adr_i[8] wb_adr_i[9]
+ wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11] wb_dat_i[12] wb_dat_i[13]
+ wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18] wb_dat_i[19] wb_dat_i[1]
+ wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24] wb_dat_i[25] wb_dat_i[26]
+ wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30] wb_dat_i[31] wb_dat_i[3]
+ wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8] wb_dat_i[9] wb_dat_o[0]
+ wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14] wb_dat_o[15] wb_dat_o[16]
+ wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20] wb_dat_o[21] wb_dat_o[22]
+ wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27] wb_dat_o[28] wb_dat_o[29]
+ wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4] wb_dat_o[5] wb_dat_o[6]
+ wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0] wb_sel_i[1] wb_sel_i[2]
+ wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_79_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6914_ _6914_/D _7193_/RN _6914_/CLK _6914_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6845_ _6845_/D _7193_/RN _6845_/CLK _6845_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_167_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3988_ _3988_/I0 _6658_/Q _3988_/S _6658_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6776_ hold96/Z _7193_/RN _6776_/CLK hold95/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5727_ hold2/Z hold195/Z _5727_/S _5727_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5658_ hold626/Z hold271/Z _5664_/S _5658_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4609_ _4601_/Z _5285_/B _4607_/Z _5021_/B _4612_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_105_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5589_ hold79/Z hold62/Z _5592_/S hold80/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold362 _7063_/Q hold362/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_117_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold351 _6886_/Q hold351/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold340 hold340/I _6894_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold373 _5878_/Z _7208_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold395 _7085_/Q hold395/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold384 _4110_/Z _6669_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7259_ _7259_/D _7260_/RN _7260_/CLK _7259_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_104_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_461 _4073__20/I _6704_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_472 net813_472/I _6693_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_494 net413_86/I _6671_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_483 net813_483/I _6682_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_1_0__f__1062_ clkbuf_0__1062_/Z _4309_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_95_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4960_ _5420_/A3 _5420_/A2 _5270_/A1 _4761_/I _4960_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_51_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4891_ _5315_/A2 _4524_/Z _4675_/Z _4700_/Z _4891_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_60_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3911_ _3485_/Z _3525_/Z _3913_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_177_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6630_ _7193_/RN _6652_/A2 _6630_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_20_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3842_ _3519_/Z _3537_/Z _3950_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6561_ _6561_/A1 _7261_/Q _6833_/D _6561_/B2 _6562_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_80_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3773_ _3773_/A1 _3773_/A2 _3773_/A3 _3773_/A4 _3773_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5512_ hold271/Z hold930/Z _5512_/S _5512_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6492_ _6492_/A1 _6492_/A2 _6492_/A3 _6492_/A4 _6492_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_172_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5443_ _5443_/A1 _5245_/Z _5444_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_146_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5374_ _5374_/A1 _5374_/A2 _5374_/A3 _5374_/A4 _5374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7113_ _7113_/D _7221_/RN _7113_/CLK _7113_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4325_ hold271/Z hold872/Z _4325_/S _4325_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4256_ hold86/Z hold312/Z _4261_/S _4256_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7044_ _7044_/D _7297_/RN _7044_/CLK _7044_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_110_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4187_ hold271/Z hold743/Z _4187_/S _4187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6828_ _6828_/D _7279_/RN _7279_/CLK _6828_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_50_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6759_ _6759_/D _7258_/RN _6759_/CLK _6759_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_109_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold170 _5556_/Z _6923_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold192 _6929_/Q hold192/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold181 _5783_/Z _7124_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_59_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_170_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5090_ _5090_/A1 _5090_/A2 _5400_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4110_ hold52/Z hold383/Z _4118_/S _4110_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4041_ _3425_/S _7283_/Q _4041_/A3 _4041_/B1 _3409_/Z _6733_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
Xclkbuf_4_3_0__1359_ clkbuf_0__1359_/Z net613_253/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_49_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5992_ _5992_/A1 _5991_/Z _5995_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4943_ _4759_/Z _4903_/Z _5330_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_33_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4874_ _4641_/Z _4833_/Z _4874_/B _4874_/C _4876_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_71_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6613_ hold886/Z hold271/Z _6613_/S _6613_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3825_ _3519_/Z _3527_/Z _3933_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_174_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3756_ _6685_/Q _3945_/C2 _3941_/A2 _7161_/Q _3757_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6544_ _6711_/Q _5948_/Z _6261_/Z _6810_/Q _6546_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_173_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6475_ _6475_/I _6476_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5426_ _3401_/I _4369_/Z _5172_/B _5172_/C _5426_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3687_ _3687_/A1 _3687_/A2 _3687_/A3 _3686_/Z _3687_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xoutput253 _4079_/I pad_flash_io0_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput242 _6752_/Q mgmt_gpio_out[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput220 _4062_/Z mgmt_gpio_out[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput231 _6749_/Q mgmt_gpio_out[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5357_ _5357_/A1 _5357_/A2 _5357_/A3 _5357_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xoutput275 _6679_/Q pll_trim[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput286 hold93/I pll_trim[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput264 _6880_/Q pll_div[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5288_ _5288_/A1 _5468_/A2 _5288_/B _5288_/C _5292_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_99_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ _6567_/I0 _6814_/Q _4312_/S _6814_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput297 _6892_/Q pwr_ctrl_out VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4239_ _4238_/Z hold787/Z _4245_/S _4239_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7027_ _7027_/D _7258_/RN _7027_/CLK _7027_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_101_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4590_ _4454_/Z _4878_/A2 _5364_/B _4586_/Z _4590_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_147_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3610_ _6571_/I0 _6874_/Q _3898_/S _3610_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3541_ _3485_/Z _3540_/Z _4210_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_171_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold917 _4151_/Z _6699_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_6_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold906 _6713_/Q hold906/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold928 _4275_/Z _6787_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_31_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3472_ _3472_/I0 hold31/Z hold21/Z hold32/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
Xhold939 _5877_/Z _7207_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6260_ _6260_/A1 _6260_/A2 _6260_/A3 _6259_/Z _6260_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_170_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5211_ _4892_/B _4683_/Z _5211_/B _5211_/C _5396_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_6191_ _7076_/Q _5965_/Z _5980_/Z _6694_/Q _5967_/Z _6720_/Q _6193_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_43_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5142_ _5281_/C _4539_/I _4817_/Z _5364_/B _4547_/Z _5470_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_97_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ _4699_/Z _5255_/B _5073_/B _5335_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_38_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4024_ _4024_/I _6731_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5975_ _7044_/Q _7228_/Q _7227_/Q wire348/Z _5975_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_178_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4926_ _5324_/A1 _4926_/A2 _4926_/B _4929_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_139_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4857_ _4614_/Z _4833_/Z _5289_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3808_ _3537_/Z _3617_/Z _5728_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xnet563_219 net563_248/I _7006_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_208 net563_225/I _7017_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_181_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4788_ _5414_/A2 _5218_/B _5125_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6527_ _6554_/A1 _6521_/Z _6526_/Z _6527_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_118_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3739_ _3739_/A1 _3739_/A2 _3739_/A3 _3739_/A4 _3739_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6458_ _7116_/Q _6240_/Z _6297_/Z _6704_/Q _6459_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_109_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5409_ _5334_/Z _5409_/A2 _5448_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_133_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6389_ _7031_/Q _6269_/Z _6273_/Z _6975_/Q _6390_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_102_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5760_ hold932/Z hold271/Z _5766_/S _5760_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5691_ hold178/Z hold2/Z _5691_/S _5691_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4711_ _5302_/B _5099_/A1 _5099_/A2 _4703_/Z _4711_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_1290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4642_ _5315_/A1 _5315_/A2 _4551_/Z _5364_/B _5038_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_175_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4573_ _4551_/Z _5364_/B _5471_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_116_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold703 _6858_/Q hold703/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7292_ _7292_/D _6646_/Z _7303_/CLK _7292_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_171_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold725 _5774_/Z _7116_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3524_ _3509_/Z _3523_/Z _3957_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6312_ _6989_/Q _6533_/A2 _6533_/A3 _6533_/A4 _6318_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold714 _4145_/Z _6695_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold736 _4340_/Z _6844_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold747 _6735_/Q hold747/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3455_ hold14/Z hold28/Z _3460_/S _7289_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6243_ _6484_/A2 _6533_/A4 _6285_/A2 _6302_/A4 _6243_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold769 _6785_/Q hold769/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold758 _5516_/Z _6892_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_130_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6174_ _7067_/Q _5985_/Z _6000_/Z _7133_/Q _6174_/C _6180_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3386_ _7228_/Q _6021_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_5125_ _5317_/A1 _5123_/Z _5125_/A3 _5126_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_69_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5056_ _4699_/Z _5051_/Z _5056_/B _5056_/C _5057_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_84_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4007_ _3990_/I _4006_/Z _4008_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_66_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_54__1359_ net663_324/I _4073__20/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_134__1359_ net613_293/I net463_147/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_26_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5958_ _7228_/Q _7227_/Q _6210_/C _6210_/A2 _5958_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_187_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4909_ _4500_/Z _5072_/A4 _4436_/B _4494_/Z _4909_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_40_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5889_ hold62/Z hold320/Z _5892_/S _5889_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold41 hold41/I hold41/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold30 hold30/I hold30/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold52 hold52/I hold52/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold63 hold63/I hold63/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold74 hold74/I hold74/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold85 hold85/I hold85/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_152_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold96 hold96/I hold96/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_84_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_7__f_wb_clk_i clkbuf_0_wb_clk_i/Z _4067_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_5 _4187_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6930_ _6930_/D _7258_/RN _6930_/CLK _6930_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6861_ _6861_/D _7279_/RN _7230_/CLK _6861_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5812_ _3515_/Z _3552_/Z _5520_/C _5820_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_63_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6792_ _6792_/D _7265_/CLK _6792_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5743_ hold86/Z hold604/Z _5748_/S _5743_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5674_ _5674_/A1 hold18/Z _5682_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_163_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4625_ _4887_/A1 _4868_/A1 _4551_/Z _5364_/B _4625_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4556_ _4528_/Z _4536_/Z _4556_/A3 _4547_/Z _4556_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold500 _7104_/Q hold500/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold511 _5635_/Z _6993_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold544 _5843_/Z _7177_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3507_ hold338/Z _3497_/I _3501_/Z _3489_/I _3507_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold533 _6782_/Q hold533/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold522 _7009_/Q hold522/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7275_ _7275_/D _7279_/RN _7279_/CLK _7275_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_171_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4487_ _4687_/A2 _4687_/A3 _5220_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold577 _5849_/Z _7182_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold588 _6753_/Q hold588/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold555 _7017_/Q hold555/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold566 _6895_/Q hold566/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3438_ input58/Z hold997/Z _3438_/S _7295_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold599 _5570_/Z _6935_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6226_ _6727_/Q _5994_/I _6226_/B _6227_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_112_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3369_ _7007_/Q _3369_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6157_ _7116_/Q _5984_/Z _5997_/Z _7100_/Q _7074_/Q _5980_/Z _6158_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5108_ _5400_/A1 _5108_/A2 _5310_/C _5107_/I _5108_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_66_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6088_ _6088_/I _6089_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5039_ _5035_/Z _5036_/Z _5205_/C _5039_/A4 _5040_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_2727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput120 wb_adr_i[3] _4456_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xinput142 wb_dat_i[22] _6597_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput131 wb_dat_i[12] _6591_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput153 wb_dat_i[3] _3396_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_88_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput164 wb_sel_i[3] _6575_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4410_ _4412_/B _4412_/C _5003_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_172_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5390_ _5390_/A1 _5390_/A2 _5350_/Z _5390_/A4 _5390_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_172_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4341_ _3529_/Z hold630/Z _5520_/C _4341_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_114_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4272_ _4103_/I hold769/Z _4273_/S _4272_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7060_ _7060_/D _7297_/RN _7060_/CLK _7060_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_6011_ _6011_/A1 _6558_/S _6011_/B1 _6310_/A3 _7241_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_113_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6913_ _6913_/D _7193_/RN _6913_/CLK _6913_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_130_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6844_ _6844_/D _7193_/RN _6844_/CLK _6844_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_189_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3987_ _6733_/Q _3972_/Z _3987_/A3 _3987_/B _3988_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_6775_ _6775_/D _7193_/RN _6775_/CLK _6775_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5726_ hold15/Z hold298/Z _5727_/S _5726_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5657_ hold129/Z hold113/Z _5664_/S _5657_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4608_ _4551_/Z _4501_/B _4853_/A1 _5364_/B _5021_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_123_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5588_ hold77/Z hold52/Z _5592_/S hold78/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold330 _6920_/Q hold330/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4539_ _4539_/I _5281_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
Xhold341 _7108_/Q hold341/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold352 _5507_/Z _6886_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold363 _5714_/Z _7063_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7258_ _7258_/D _7258_/RN _7258_/CLK _7258_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold396 _5739_/Z _7085_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold374 _7093_/Q hold374/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold385 _6668_/Q hold385/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_120_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6209_ _7297_/Q _5969_/Z _6227_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7189_ _7189_/D _7221_/RN _7189_/CLK _7189_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_131_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_462 net413_94/I _6703_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_473 net813_473/I _6692_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_484 net813_485/I _6681_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_495 net813_495/I _6670_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_13_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4890_ _4890_/I _5259_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3910_ _6932_/Q _3910_/A2 _3953_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_33_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3841_ _6695_/Q _4143_/A1 _3868_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_20_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6560_ _6561_/B2 _6559_/Z _6561_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3772_ _7216_/Q _3912_/A2 _3930_/A2 _7128_/Q _3773_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_186_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5511_ _4103_/I hold874/Z _5512_/S _5511_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6491_ _7173_/Q _5948_/Z _6261_/Z _6963_/Q _6266_/Z _7019_/Q _6492_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_173_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5442_ _5056_/C _5442_/A2 _5442_/A3 _5442_/A4 _5442_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_146_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5373_ _5287_/C _4551_/Z _5364_/B _5373_/B _5374_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_7112_ _7112_/D _7258_/RN _7112_/CLK _7112_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4324_ _4103_/I hold805/Z _4325_/S _4324_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7043_ _7043_/D _7258_/RN _7043_/CLK _7043_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4255_ hold271/Z hold795/Z _4261_/S _4255_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4186_ _4103_/I hold670/Z _4187_/S _4186_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6827_ _6827_/D _7279_/RN _7279_/CLK _6833_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_24_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6758_ _6758_/D _7258_/RN _6758_/CLK _6758_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_6_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5709_ hold226/Z hold2/Z _5709_/S _5709_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6689_ _6689_/D _7297_/RN _6689_/CLK _6689_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_164_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold160 _7011_/Q hold160/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold171 _6994_/Q hold171/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold193 _5563_/Z _6929_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_78_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold182 _6978_/Q hold182/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_137_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4040_ _4040_/I _6734_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _7231_/Q _7228_/Q _7227_/Q _5991_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_24_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4942_ _4939_/Z _4942_/A2 _5062_/B _4948_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_177_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet413_90 net413_90/I _7135_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4873_ _4641_/Z _5051_/S _5287_/B _4681_/Z _4874_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_21_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6612_ hold819/Z _4103_/I _6613_/S _6612_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3824_ _3529_/Z _3653_/Z _3935_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3755_ hold77/I _5584_/A1 _3956_/A2 _7121_/Q _7145_/Q _3951_/C1 _3757_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6543_ _6852_/Q _6274_/Z _6285_/Z _6693_/Q _6707_/Q _6254_/Z _6546_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6474_ _6744_/Q _7256_/Q _6474_/B _6475_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_119_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3686_ _3686_/A1 _3686_/A2 _3686_/A3 _3686_/A4 _3686_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_161_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5425_ _5425_/A1 _5425_/A2 _5425_/A3 _5425_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
Xoutput210 _4056_/Z mgmt_gpio_out[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput232 _6914_/Q mgmt_gpio_out[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput221 _6739_/Q mgmt_gpio_out[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput243 _4059_/Z mgmt_gpio_out[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5356_ _5356_/A1 _5387_/A2 _5356_/B _5356_/C _5357_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xoutput254 _7307_/Z pad_flash_io1_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput276 _6680_/Q pll_trim[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput265 _6881_/Q pll_div[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5287_ _4554_/Z _4683_/Z _5287_/B _5287_/C _5487_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_101_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput287 _6889_/Q pll_trim[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4307_ _6566_/I0 _6813_/Q _4312_/S _6813_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput298 _3907_/Z reset VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4238_ hold330/Z hold62/Z _4244_/S _4238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7026_ _7026_/D _7260_/RN _7026_/CLK _7026_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_83_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4169_ hold271/Z hold906/Z _4169_/S _4169_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwire348 wire348/I wire348/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_7_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3540_ _3653_/A1 _3617_/A1 hold629/Z _3492_/Z _3540_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_155_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold918 _7014_/Q hold918/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold907 _4169_/Z _6713_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_31_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5210_ _5209_/Z _5208_/Z _5417_/A1 _5210_/A4 _5210_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_143_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3471_ _3471_/I _3472_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold929 _7135_/Q hold929/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6190_ _6716_/Q _5997_/Z _6014_/Z _6809_/Q _6193_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_130_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5141_ _5293_/A1 _4614_/Z _5289_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_111_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5072_ _4500_/Z _4906_/Z _5078_/A2 _5072_/A4 _5072_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_97_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4023_ hold995/Z _4022_/Z _4024_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_65_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5974_ _5974_/A1 _5974_/A2 _5974_/A3 _5974_/A4 _5983_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4925_ _5083_/B _5080_/C _5370_/B _4926_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_100_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4856_ _4614_/Z _4817_/Z _4858_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_178_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_209 net663_326/I _7016_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3807_ _3509_/Z _3519_/Z _3923_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_165_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4787_ _5220_/B2 _5092_/A1 _4787_/A3 _4491_/B _4787_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_20_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6526_ _6526_/A1 _6526_/A2 _6526_/A3 _6526_/A4 _6526_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_147_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3738_ input67/Z _4227_/S _4244_/S input38/Z _5701_/A1 _7055_/Q _3739_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_146_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6457_ _7188_/Q _6282_/Z _6293_/Z _7156_/Q _6296_/Z _7164_/Q _6465_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_107_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3669_ hold49/I _5584_/A1 _3959_/B1 _6671_/Q _3673_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5408_ _4761_/I _5245_/Z _5481_/B1 _4908_/Z _5408_/C _5409_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_6388_ hold65/I _6245_/Z _6288_/Z _7121_/Q _6390_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_86_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_14__1359_ net413_58/I net413_74/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5339_ _5261_/I _5338_/Z _5262_/Z _5339_/A4 _5340_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_87_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_77__1359_ net413_53/I net413_65/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7009_ _7009_/D _7260_/RN _7009_/CLK _7009_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xclkbuf_3_6__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7279_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5690_ hold278/Z hold15/Z _5691_/S _5690_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4710_ _4694_/Z _4703_/Z _5308_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_1291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4641_ _5281_/C _4467_/B _4472_/B _4501_/B _4641_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4572_ _4572_/I _5472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_129_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7291_ _7291_/D _6645_/Z _7303_/CLK _7291_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_128_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3523_ hold338/Z _3617_/A1 _3501_/Z _3489_/I _3523_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6311_ _6973_/Q _6484_/A2 _6311_/A3 _6533_/A2 _6327_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold737 _6729_/Q hold737/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold715 _6764_/Q hold715/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold726 _6846_/Q hold726/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold704 _4361_/Z _6858_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold748 _4197_/Z _6735_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3454_ hold1/Z hold14/Z _3460_/S _7290_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold759 _6674_/Q hold759/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6242_ _7110_/Q _6240_/Z _6241_/Z _7044_/Q _6260_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_170_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6173_ _6173_/I _6174_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3385_ _7231_/Q _6210_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_12
XFILLER_112_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5124_ _5414_/A2 _4784_/Z _5124_/B _5317_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_97_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5055_ _5130_/B2 _5420_/A2 _4367_/Z _5291_/C _5055_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_73_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4006_ _5900_/A1 _5911_/A1 _7225_/Q _7224_/Q _4006_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_37_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5957_ _3990_/I _6745_/Q _5957_/S _6558_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_111_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_1__1359_ net713_387/I net763_445/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4908_ _5324_/A1 _4759_/Z _4494_/Z _4496_/Z _4908_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_52_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5888_ hold52/Z hold644/Z _5892_/S _5888_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4839_ _4887_/A1 _5414_/A2 _5399_/A2 _5287_/B _5369_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_153_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6509_ _6692_/Q _6285_/Z _6299_/Z _6857_/Q _6511_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_162_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold31 hold31/I hold31/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_0_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold20 hold20/I hold20/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_48_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold64 hold64/I hold64/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold42 hold42/I hold42/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold53 hold53/I hold53/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_29_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold86 hold86/I hold86/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_63_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold97 hold97/I hold97/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_21_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold75 hold75/I hold75/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_90_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_6 _6803_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_60__1359_ clkbuf_4_15_0__1359_/Z net663_305/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_3_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_140__1359_ net563_220/I net763_447/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_66_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6860_ _6860_/D _7279_/RN _7230_/CLK _6860_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_47_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5811_ hold2/Z hold176/Z _5811_/S _5811_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6791_ _6791_/D _7243_/CLK _6791_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet613_290 _4073__45/I _6935_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5742_ hold271/Z hold986/Z _5748_/S _5742_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5673_ hold152/Z hold2/Z _5673_/S _5673_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ _4441_/B _5281_/C _4436_/B _4501_/B _4624_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_135_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4555_ _5129_/A3 _4835_/A2 _4555_/B _4555_/C _4556_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xhold501 _5761_/Z _7104_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold523 _7216_/Q hold523/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold512 _7089_/Q hold512/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold545 _7121_/Q hold545/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3506_ _3485_/Z _3505_/Z _3909_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold534 _4268_/Z _6782_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4486_ _4486_/A1 _4483_/B _4486_/B1 _4484_/Z _5312_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_7274_ _7274_/D _7279_/RN _7279_/CLK _7274_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_116_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold567 _7114_/Q hold567/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold578 _7198_/Q hold578/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold556 _5662_/Z _7017_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3437_ _3442_/B _6663_/Q _6664_/Q _6665_/Q _3438_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6225_ _6800_/Q _5958_/Z _5967_/Z _6721_/Q _6227_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold589 _4226_/Z _6753_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3368_ hold56/I _3368_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6156_ _7156_/Q _5960_/Z _5965_/Z _6704_/Q _6006_/Z _7172_/Q _6158_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ _5107_/I _5309_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3299_ _6665_/Q _3465_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6087_ _6555_/C _7243_/Q _6087_/B _6088_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5038_ _5038_/A1 _4606_/Z _5003_/Z _5038_/B _5205_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XTAP_2728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6989_ _6989_/D _7210_/RN _6989_/CLK _6989_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_167_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput110 wb_adr_i[23] _4026_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_150_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput143 wb_dat_i[23] _6600_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput132 wb_dat_i[13] _6594_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput154 wb_dat_i[4] _3397_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput121 wb_adr_i[4] _4460_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_163_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput165 wb_stb_i _4032_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_36_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4340_ hold271/Z hold735/Z _4340_/S _4340_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4271_ _5520_/C _3527_/Z _5513_/A3 _5839_/A3 _4273_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_140_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6010_ _6010_/A1 _6010_/A2 _6924_/Q _6201_/A3 _6011_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_100_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6912_ _6912_/D _7193_/RN _6912_/CLK _6912_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6843_ _6843_/D _7193_/RN _6843_/CLK _6843_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3986_ _7305_/Q _3415_/Z _6658_/Q _3987_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6774_ _6774_/D _7193_/RN _6774_/CLK _6774_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5725_ hold29/Z hold290/Z _5727_/S _5725_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5656_ _5656_/A1 hold18/Z _5664_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_4607_ _4607_/A1 _4570_/Z _4606_/Z _4501_/B _4607_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_175_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold320 _7218_/Q hold320/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5587_ hold108/Z hold86/Z _5592_/S _5587_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold331 _5553_/Z _6920_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold342 _5765_/Z _7108_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4538_ _5288_/B _4467_/B _4472_/B _4539_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_105_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold353 _7090_/Q hold353/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7257_ _7257_/D _7258_/RN _7258_/CLK _7257_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_117_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4469_ _4459_/Z _4469_/A2 _4690_/B _4690_/C _4786_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold375 _5748_/Z _7093_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold386 _4108_/Z _6668_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold364 _6820_/Q hold364/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold397 _6964_/Q hold397/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6208_ _7249_/Q _6208_/I1 _6558_/S _7249_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7188_ _7188_/D _7221_/RN _7188_/CLK _7188_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_131_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6139_ _7058_/Q _6210_/A2 _6210_/B _6210_/C _6155_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_485 net813_485/I _6680_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_452 _4073__2/I _6713_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_463 net413_89/I _6702_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet813_474 net813_475/I _6691_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_496 net413_88/I _6669_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3840_ _3537_/Z _3680_/Z _4143_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_186_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3771_ _7070_/Q _3943_/A2 _3945_/B1 _7088_/Q _3773_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_34_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5510_ _3521_/Z _3527_/Z _5520_/C _5512_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_173_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6490_ _7085_/Q _6290_/Z _6302_/Z _7093_/Q _6490_/C _6492_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_172_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5441_ _5437_/Z _5440_/Z _5441_/B _5463_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_145_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5372_ _5372_/A1 _5139_/Z _5055_/Z _5372_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_114_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7111_ _7111_/D _7219_/RN _7111_/CLK _7111_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4323_ _3509_/Z _5821_/A3 _5513_/A3 _5520_/C _4325_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7042_ _7042_/D _7258_/RN _7042_/CLK _7042_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_113_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4254_ hold113/Z hold238/Z _4261_/S _4254_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4185_ _5520_/C _3537_/Z _5513_/A3 _5839_/A3 _4187_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_94_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6826_ _6826_/D _7279_/RN _7279_/CLK _6826_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_149_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6757_ _6757_/D _7258_/RN _6757_/CLK _6757_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3969_ _3427_/Z _6663_/Q _6664_/Q _3970_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_176_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5708_ hold184/Z hold15/Z _5709_/S _5708_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6688_ _6688_/D _7297_/RN _6688_/CLK _6688_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_12_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_opt_3_0__1359_ net663_304/I clkbuf_opt_3_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_128_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5639_ hold120/Z hold113/Z hold19/Z _6996_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold161 _6915_/Q hold161/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7309_ _7309_/I _7309_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold150 _6979_/Q hold150/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_5_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold194 _7010_/Q hold194/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold183 _5618_/Z _6978_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold172 _5636_/Z _6994_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5990_ _7020_/Q wire348/Z _6002_/A2 _6956_/Q _6211_/B1 _6988_/Q _5992_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_4941_ _5464_/A1 _5410_/A1 _5062_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_52_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet413_80 net413_80/I _7145_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4872_ _4872_/A1 _5215_/C _5117_/A2 _5215_/B _4874_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4073__50 _4073__51/I _7175_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_91 net413_91/I _7134_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_178_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3823_ _6981_/Q _3901_/A2 _3889_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6611_ _6611_/A1 hold18/Z _6613_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_158_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3754_ _7137_/Q _3951_/A2 _3954_/B1 input23/Z _3754_/C _3757_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6542_ _6542_/A1 _6542_/A2 _6542_/A3 _6542_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6473_ _6466_/Z _6472_/Z _6473_/B1 _6286_/Z _6555_/C _6474_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3685_ hold58/I _3957_/A2 _3941_/B1 _7171_/Q _3686_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xoutput200 _4050_/Z mgmt_gpio_oeb[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_173_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5424_ _5489_/A1 _5423_/Z _5427_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_173_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput233 _6915_/Q mgmt_gpio_out[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput222 _6740_/Q mgmt_gpio_out[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput211 _6758_/Q mgmt_gpio_out[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput244 _6754_/Q mgmt_gpio_out[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5355_ _5437_/A2 _5350_/Z _5352_/Z _5354_/Z _5355_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_142_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput255 _4077_/ZN pad_flash_io1_ie VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput277 _6681_/Q pll_trim[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput266 _6882_/Q pll_div[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5286_ _5286_/A1 _5374_/A3 _5374_/A2 _5292_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_102_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput299 _4085_/Z ser_rx VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput288 _6890_/Q pll_trim[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4306_ _6565_/I0 _6812_/Q _4312_/S _6812_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4237_ _4236_/Z hold807/Z _4245_/S _4237_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7025_ hold44/Z _7260_/RN _7025_/CLK hold43/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_74_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_5__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7260_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4168_ _4103_/I hold817/Z _4169_/S _4168_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4099_ hold5/Z _6608_/I0 hold21/I hold6/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_83_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_37__1359_ net413_53/I _4073__22/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_51_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_117__1359_ net613_293/I net813_499/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_24_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6809_ _6809_/D _7210_/RN _6809_/CLK _6809_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold919 _6989_/Q hold919/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold908 _7079_/Q hold908/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3470_ _6660_/Q _6733_/Q _6661_/Q _3471_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_155_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5140_ _5293_/A1 _4549_/Z _5147_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5071_ _4376_/Z _5071_/A2 _5257_/A1 _4699_/Z _5408_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_29_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4022_ _7282_/Q _3409_/Z _4022_/A3 _6730_/Q _4022_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_56_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5973_ _7012_/Q _5971_/Z _5972_/Z _6940_/Q _5974_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4924_ _5259_/A1 _5337_/A2 _5258_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_21_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4855_ _5287_/C _4844_/Z _4855_/B _4855_/C _4858_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_20_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4786_ _4786_/A1 _4786_/A2 _4786_/A3 _5137_/B1 _4787_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3806_ _3509_/Z _3535_/Z _3924_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_181_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3737_ _6927_/Q _3935_/A2 _3916_/A2 _7153_/Q _3912_/B1 _6886_/Q _3739_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6525_ _6694_/Q _6248_/Z _6300_/Z _6720_/Q _6526_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_162_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6456_ hold25/I _6253_/Z _6272_/Z _7204_/Q _6456_/C _6465_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_118_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3668_ hold47/I _3923_/C1 _3956_/A2 hold59/I _3668_/C _3674_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_115_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5407_ _5406_/Z _5454_/A2 _5419_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6387_ _7047_/Q _6241_/Z _6251_/Z _6983_/Q _6268_/Z hold77/I _6390_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3599_ _7011_/Q _3934_/A2 _5683_/A1 _7043_/Q _7051_/Q _3952_/A2 _3601_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_173_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5338_ _5332_/Z _5334_/Z _5447_/A1 _5338_/A4 _5338_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_161_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5269_ _4454_/Z _5269_/A2 _4651_/Z _4675_/Z _5464_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_75_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7008_ _7008_/D _7297_/RN _7008_/CLK _7008_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_55_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_20__1359_ net613_253/I _4073__51/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_100__1359_ clkbuf_4_5_0__1359_/Z net563_212/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4640_ _5315_/A1 _5315_/A2 _5468_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4571_ _4549_/Z _4570_/Z _4572_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6310_ _6308_/Z _6310_/A2 _6310_/A3 _6558_/S _6310_/B2 _7251_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_128_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7290_ _7290_/D _6644_/Z _7303_/CLK hold1/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_155_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold705 _7192_/Q hold705/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3522_ _3509_/Z _3521_/Z _3910_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold716 _4248_/Z _6764_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold727 _6691_/Q hold727/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3453_ _4041_/B1 _3442_/B _6732_/Q _3460_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_144_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6241_ _7235_/Q _7234_/Q _6300_/A2 _6533_/A2 _6241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold749 _6721_/Q hold749/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold738 _4193_/Z _6729_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_157_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6172_ _6979_/Q _5964_/Z _6014_/Z _6963_/Q _5999_/Z _7035_/Q _6173_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5123_ _5456_/A1 _5220_/B2 _5312_/A2 _5137_/B1 _5123_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3384_ _6786_/Q _6555_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_5054_ _5370_/B _5258_/A2 _4977_/Z _5323_/B _5324_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_69_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4005_ _4005_/A1 _4003_/Z _5945_/A1 _6901_/Q _6743_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_84_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_350 net413_74/I _6867_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5956_ _5957_/S _6745_/Q _6310_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_187_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4907_ _4759_/Z _4906_/Z _5257_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_179_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5887_ hold86/Z hold523/Z _5892_/S _5887_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4838_ _4555_/C _4876_/A2 _4838_/B1 _5291_/C _4841_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_166_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4769_ _4703_/Z _4764_/Z _5117_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_5_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6508_ _6724_/Q _6240_/Z _6247_/Z _6728_/Q _6511_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_136_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6439_ _6434_/Z _6439_/A2 _6439_/A3 _6439_/A4 _6439_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_121_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold21 hold21/I hold21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold10 hold10/I hold10/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold32 hold32/I hold32/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_0_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold54 hold54/I hold54/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold43 hold43/I hold43/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold65 hold65/I hold65/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_91_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold76 hold76/I hold76/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold98 hold98/I hold98/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold87 hold87/I hold87/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_17_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_7 _5505_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5810_ hold15/Z hold426/Z _5811_/S _5810_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6790_ _6790_/D _7210_/RN _6790_/CLK _6790_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_96_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_291 net613_291/I _6934_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5741_ hold113/Z hold584/Z _5748_/S _5741_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet613_280 net663_326/I _6945_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5672_ hold186/Z hold15/Z _5673_/S _5672_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4623_ _4887_/A1 _4868_/A1 _5376_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold502 _6701_/Q hold502/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_129_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4554_ _3401_/I _3402_/I _4456_/B _5051_/S _4554_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7273_ _7273_/D _7279_/RN _7279_/CLK _7273_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_144_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold535 _7189_/Q hold535/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_128_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold524 _5887_/Z _7216_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_117_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold513 _5744_/Z _7089_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3505_ _3617_/A1 _3501_/Z _3489_/I _3492_/Z _3505_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4485_ _4381_/Z _4485_/A2 _4486_/B1 _4424_/B _4687_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_104_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold546 _5780_/Z _7121_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold568 _5772_/Z _7114_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold579 _5867_/Z _7198_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6224_ _6719_/Q _5960_/Z _5965_/Z _7077_/Q _6006_/Z _6711_/Q _6227_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold557 _6749_/Q hold557/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3436_ _6665_/Q _6664_/Q _6663_/Q _3898_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_131_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3367_ _7023_/Q _3367_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6155_ _6155_/A1 _6155_/A2 _6155_/A3 _6155_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_98_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ _6073_/Z _6085_/Z _6392_/B1 _6168_/C _6555_/C _6087_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_5106_ _5106_/A1 _5106_/A2 _5107_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5037_ _5039_/A4 _5036_/Z _5357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3298_ hold4/Z hold5/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6988_ _6988_/D _7297_/RN _6988_/CLK _6988_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5939_ _6745_/Q _5939_/A2 _5913_/I _6282_/A2 _7233_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_15_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput111 wb_adr_i[24] _4029_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput100 wb_adr_i[14] _4386_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_89_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput144 wb_dat_i[24] _6579_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput133 wb_dat_i[14] _6597_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput122 wb_adr_i[5] _4436_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_76_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput166 wb_we_i _6575_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xinput155 wb_dat_i[5] _3398_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_5_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4270_ hold440/Z hold2/Z _4270_/S _4270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6911_ _6911_/D _7193_/RN _6911_/CLK _6911_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_62_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6842_ _6842_/D input75/Z _6842_/CLK _6842_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_74_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3985_ _3984_/Z _6659_/Q _3988_/S _6659_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6773_ _6773_/D _7193_/RN _6773_/CLK _6773_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5724_ hold62/Z hold571/Z _5727_/S _5724_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5655_ hold160/Z hold2/Z _5655_/S _7011_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4606_ _4648_/A2 _4467_/B _4648_/A1 _4606_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_11_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold310 _6703_/Q hold310/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5586_ hold620/Z hold271/Z _5592_/S _5586_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold332 _6772_/Q hold332/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4537_ _4441_/B _4501_/B _5399_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_89_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold321 _5889_/Z _7218_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold343 _7186_/Q hold343/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7256_ _7256_/D _7258_/RN _7258_/CLK _7256_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4468_ _4467_/B _4736_/A1 _4468_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
Xhold354 _5745_/Z _7090_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold376 _6956_/Q hold376/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold387 _7118_/Q hold387/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold365 _4321_/Z _6820_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3419_ _4041_/B1 _6730_/Q _7304_/Q _3421_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7187_ _7187_/D _7258_/RN _7187_/CLK _7187_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold398 _7004_/Q hold398/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6207_ _6207_/I _6208_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4399_ _4402_/B _4483_/B _4026_/B _4026_/C _4399_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6138_ _7108_/Q _5967_/Z _6147_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_86_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ _7063_/Q _5985_/Z _6084_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_93_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_464 net413_96/I _6701_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_453 _4073__2/I _6712_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet813_475 net813_475/I _6690_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_187_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet813_497 net413_88/I _6668_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_486 net813_489/I _6679_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3770_ _7160_/Q _3941_/A2 _5503_/A2 _3904_/A2 _3770_/C _3773_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_160_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5440_ _5440_/A1 _5357_/Z _5388_/Z _5440_/A4 _5440_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_157_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5371_ _5371_/A1 _5287_/B _5470_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_59_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7110_ _7110_/D _7219_/RN _7110_/CLK _7110_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4322_ hold271/Z hold697/Z _4322_/S _4322_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4253_ _3485_/Z _3540_/Z _6652_/A2 hold6/Z _4261_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7041_ _7041_/D _7260_/RN _7041_/CLK _7041_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_101_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4184_ hold731/Z hold271/Z _4184_/S _4184_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_3_4__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7258_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_103_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6825_ _6825_/D _7210_/RN _6825_/CLK _6825_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3968_ _6665_/Q _3967_/Z _6665_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6756_ _6756_/D _7258_/RN _6756_/CLK _6756_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5707_ hold553/Z hold29/Z _5709_/S _5707_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3899_ _3898_/Z hold992/Z _3899_/S _6869_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6687_ _6687_/D _7297_/RN _6687_/CLK _6687_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_163_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5638_ _5638_/A1 hold18/Z hold19/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_152_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5569_ hold86/Z hold564/Z _5574_/S _5569_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold162 _5547_/Z _6915_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_151_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7308_ _7308_/I _7308_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold140 _6987_/Q hold140/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold151 _5619_/Z _6979_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold195 _7075_/Q hold195/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold184 _7058_/Q hold184/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_78_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold173 _6970_/Q hold173/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7239_ _7239_/D _7258_/RN _4067_/I1 _7239_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_104_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4940_ _4421_/Z _5410_/A1 _4942_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_64_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet413_70 net413_70/I _7155_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__40 net413_80/I _7185_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_92 net413_94/I _7133_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4871_ _4641_/Z _4817_/Z _5117_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4073__51 _4073__51/I _7174_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_81 net413_81/I _7144_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6610_ _6610_/A1 _6610_/A2 _6610_/A3 _6610_/A4 _7279_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_60_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3822_ _6788_/Q _4274_/A1 _3947_/B1 _6717_/Q _3873_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6541_ _6725_/Q _6240_/Z _6248_/Z _6695_/Q _6542_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_145_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3753_ _3753_/I _3754_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6472_ _6554_/A1 _6472_/A2 _6472_/A3 _6472_/A4 _6472_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3684_ _7155_/Q _3916_/A2 _5528_/S _3683_/Z _3686_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xoutput201 _4049_/Z mgmt_gpio_oeb[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_173_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5423_ _5423_/A1 _5423_/A2 _5377_/Z _5422_/Z _5423_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xoutput234 _4053_/Z mgmt_gpio_out[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5354_ _5354_/A1 _5354_/A2 _5354_/A3 _5354_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xoutput212 _6759_/Q mgmt_gpio_out[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput223 _6741_/Q mgmt_gpio_out[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput245 _4058_/Z mgmt_gpio_out[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_88_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput267 _6876_/Q pll_ena VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput256 _4077_/I pad_flash_io1_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4305_ _6564_/I0 _6811_/Q _4312_/S _6811_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5285_ _4598_/Z _4683_/Z _5285_/B _5374_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_99_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput278 _6666_/Q pll_trim[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput289 _6684_/Q pll_trim[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4236_ hold347/Z hold52/Z _4244_/S _4236_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7024_ hold90/Z _7260_/RN _7024_/CLK hold89/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_114_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4167_ _3535_/Z _3537_/Z _5520_/C _4169_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_67_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4098_ _7221_/RN _6656_/A2 _4098_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_24_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6808_ _6808_/D _7265_/CLK _6808_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6739_ _6739_/D _7193_/RN _6739_/CLK _6739_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_20_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold909 _5733_/Z _7079_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5070_ _5070_/A1 _5070_/A2 _5334_/A1 _5070_/A4 _5074_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xclkbuf_leaf_43__1359_ net613_299/I net463_133/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_96_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4021_ _4021_/I _6746_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_123__1359_ _4073__15/I net413_62/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5972_ _7228_/Q _6210_/C _6015_/A3 _6210_/A2 _5972_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4923_ _4423_/Z _4923_/A2 _4923_/B _5080_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_52_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4854_ _4422_/Z _5414_/A2 _4614_/Z _4483_/B _4855_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_60_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4785_ _4808_/A2 _5220_/B2 _5092_/A1 _4491_/B _5124_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3805_ _3519_/Z _3552_/Z _3912_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_21_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3736_ _7217_/Q _3912_/A2 _4194_/A1 input55/Z _3948_/C1 input64/Z _3739_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_118_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6524_ _6690_/Q _6257_/Z _6275_/Z _6849_/Q _6526_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_118_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6455_ _7084_/Q _6290_/Z _6299_/Z _7058_/Q _6466_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3667_ _3667_/I _3668_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5406_ _5406_/A1 _5404_/Z _5406_/A3 _4799_/Z _5406_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6386_ _7023_/Q _6235_/Z _6243_/Z _7007_/Q _6265_/Z _6999_/Q _6391_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3598_ _7165_/Q _3941_/A2 _3947_/A2 _7101_/Q _7059_/Q _5701_/A1 _3601_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5337_ _5337_/A1 _5337_/A2 _5337_/B _5337_/C _5449_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_87_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5268_ _5368_/A1 _4650_/Z _5172_/C _5268_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_141_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7007_ _7007_/D _7260_/RN _7007_/CLK _7007_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4219_ hold75/Z hold52/Z _4227_/S _4219_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5199_ _5191_/Z _5196_/Z _5390_/A2 _5476_/A2 _5199_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_69_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4570_ _5270_/A1 _4454_/Z _5364_/B _4570_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_128_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3521_ _3489_/I _3492_/Z _3497_/I _3501_/Z _3521_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_183_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold706 _5860_/Z _7192_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_7_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold717 _6717_/Q hold717/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold728 _4139_/Z _6691_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3452_ _3451_/Z _7291_/Q _3452_/S _7291_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6240_ _7236_/Q _6533_/A4 _6302_/A4 _6533_/A3 _6240_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold739 _6747_/Q hold739/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6171_ _7149_/Q _5987_/Z _6002_/Z _7093_/Q _6003_/Z _7165_/Q _6181_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_97_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3383_ _7077_/Q _3866_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5122_ _5456_/A1 _5231_/A2 _5122_/B _5213_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_69_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5053_ _5325_/B _5078_/A2 _5060_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4004_ _4005_/A1 _4003_/Z _5894_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_133_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_351 net413_74/I _6866_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_340 net663_341/I _6885_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_92_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5955_ _5954_/Z _7240_/Q _5955_/S _7240_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4906_ _4494_/Z _5259_/A1 _4496_/Z _4407_/Z _4906_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5886_ hold271/Z hold934/Z _5892_/S _5886_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4837_ _5278_/C _4784_/Z _4838_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4768_ _4510_/Z _4764_/Z _4770_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_135_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4699_ _5420_/A3 _4835_/A2 _4456_/B _3402_/I _4699_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3719_ _3719_/A1 _3719_/A2 _3719_/A3 _3719_/A4 _3719_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6507_ _6726_/Q _6253_/Z _6296_/Z _6714_/Q _6511_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_161_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6438_ hold47/I _6290_/Z _6302_/Z _7091_/Q _6438_/C _6439_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_161_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6369_ _6967_/Q _6262_/Z _6391_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_130_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold22 hold22/I hold22/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold11 hold11/I hold11/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_130_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold33 hold33/I hold33/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_75_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold55 hold55/I hold55/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold44 hold44/I hold44/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold66 hold66/I hold66/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold77 hold77/I hold77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold99 hold99/I hold99/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold88 hold88/I hold88/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_57_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_8 _5506_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5740_ _3515_/Z _3537_/Z hold6/Z _5748_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_62_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_281 net613_281/I _6944_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_292 net813_499/I _6933_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_270 net613_273/I _6955_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5671_ hold43/Z hold29/Z _5673_/S hold44/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4622_ _4622_/A1 _5029_/B _5353_/B _4627_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_156_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4553_ _4836_/A4 _4454_/Z _5370_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_128_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4484_ _4381_/Z _4385_/Z _4387_/Z _4424_/B _4484_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_7272_ _7272_/D _7279_/RN _7279_/CLK _7272_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold514 _7145_/Q hold514/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold525 _7039_/Q hold525/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold536 _5856_/Z _7189_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold503 _4153_/Z _6701_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3504_ _5857_/A2 _5857_/A3 _5647_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3435_ _3435_/A1 _3435_/A2 _7298_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_144_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold569 _7098_/Q hold569/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6223_ _6691_/Q _5985_/Z _6014_/Z _6810_/Q _6228_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold547 _6751_/Q hold547/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold558 _4218_/Z _6749_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_143_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3366_ _7031_/Q _3366_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6154_ _7018_/Q _5971_/Z _6005_/Z _7042_/Q _7050_/Q _6019_/Z _6155_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_58_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3297_ _7291_/Q _3451_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6085_ _6078_/Z _6085_/A2 _6085_/A3 _6084_/Z _6085_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_97_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5105_ _5105_/A1 _5104_/Z _5310_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_85_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5036_ _5356_/C _5389_/C _5328_/A1 _5356_/B _5036_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_73_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6987_ _6987_/D _7260_/RN _6987_/CLK _6987_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_81_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5938_ _6484_/A2 _6302_/A3 _5939_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_41_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5869_ hold86/Z hold646/Z _5874_/S _5869_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput101 wb_adr_i[15] _4386_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_122_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput145 wb_dat_i[25] _6582_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput134 wb_dat_i[15] _6600_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput123 wb_adr_i[6] _4472_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xinput112 wb_adr_i[25] _3334_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_131_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput156 wb_dat_i[6] _3399_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_91_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_3_3__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7230_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_39_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_6_0__1359_ clkbuf_0__1359_/Z _4073__15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6910_ _6910_/D _7193_/RN _6910_/CLK _6910_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_130_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6841_ _6841_/D input75/Z _6841_/CLK _6841_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3984_ _3983_/Z _6658_/Q _6733_/Q _3984_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6772_ _6772_/D _7258_/RN _6772_/CLK _6772_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5723_ hold52/Z hold358/Z _5727_/S _5723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5654_ hold194/Z hold15/Z _5655_/S _7010_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4605_ _4638_/A2 _4648_/B _5356_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_148_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold311 _4155_/Z _6703_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold300 _7097_/Q hold300/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5585_ hold122/Z hold113/Z _5592_/S _5585_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold333 _4257_/Z _6772_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4536_ _5414_/A2 _4501_/B _4472_/B _4524_/Z _4536_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold344 _5853_/Z _7186_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold322 _7211_/Q hold322/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7255_ _7255_/D _7258_/RN _7258_/CLK _7255_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold377 _7181_/Q hold377/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4467_ _4467_/A1 _4555_/B _4467_/B _4690_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xhold366 _6885_/Q hold366/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold355 _7008_/Q hold355/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4398_ _5002_/A3 _5002_/A4 _5165_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3418_ _3417_/Z _7305_/Q _3988_/S _7305_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7186_ _7186_/D _7210_/RN _7186_/CLK _7186_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold399 _6670_/Q hold399/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold388 _5777_/Z _7118_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6206_ _6555_/C _7248_/Q _6206_/B _6207_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold1000 _7294_/Q _3433_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3349_ _7161_/Q _3349_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6137_ _7246_/Q _6136_/Z _6558_/S _7246_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6068_ _7145_/Q _7231_/Q _6210_/B wire348/I _6076_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_85_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5019_ _5191_/A3 _5019_/A2 _5390_/A1 _5019_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XTAP_2527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_465 net813_465/I _6700_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_476 net813_483/I _6689_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_454 net813_470/I _6711_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_487 net813_491/I _6678_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_498 net813_499/I _6667_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5370_ _5370_/A1 _5172_/B _5370_/B _5370_/C _5371_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_160_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4321_ hold113/Z hold364/Z _4322_/S _4321_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4252_ hold29/Z hold452/Z _4252_/S _4252_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7040_ _7040_/D _7193_/RN _7040_/CLK _7040_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_68_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4183_ hold689/Z _4103_/I _4184_/S _4183_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6824_ _6824_/D _7210_/RN _6824_/CLK _6824_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3967_ _3427_/Z _6663_/Q _6664_/Q _3967_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6755_ _6755_/D _7258_/RN _6755_/CLK _6755_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5706_ hold356/Z hold62/Z _5709_/S _5706_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_177_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3898_ _6565_/I0 _6868_/Q _3898_/S _3898_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6686_ _6686_/D _7297_/RN _6686_/CLK _6686_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_31_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5637_ hold2/Z hold154/Z _5637_/S _5637_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5568_ hold271/Z hold835/Z _5574_/S _5568_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4519_ _5170_/A2 _5269_/A2 _5328_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_137_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold141 _5628_/Z _6987_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold152 _7027_/Q hold152/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7307_ _7307_/I _7307_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold130 _5657_/Z _7012_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold185 _5708_/Z _7058_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold163 _7125_/Q hold163/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold174 _6986_/Q hold174/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7238_ _7238_/D _7238_/RN _7260_/CLK _7238_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5499_ hold410/Z hold271/Z _5502_/S _5499_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold196 _5727_/Z _7075_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_137_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7169_ _7169_/D _7219_/RN _7169_/CLK _7169_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_58_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_7__1359_ net413_58/I net413_75/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet413_60 net413_77/I _7165_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_93 net413_96/I _7132_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4870_ _5293_/B _4844_/Z _5215_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4073__30 _4073__30/I _7195_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__41 _4073__41/I _7184_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet413_71 net413_71/I _7154_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_82 net413_83/I _7143_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3821_ _3537_/Z _3653_/Z _3947_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6540_ _6867_/Q _6272_/Z _6293_/Z _6719_/Q _6540_/C _6547_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_60_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_66__1359_ clkbuf_4_13_0__1359_/Z net613_297/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_146__1359_ net563_220/I net663_341/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3752_ _6975_/Q _3923_/A2 _3959_/B1 _6669_/Q _5656_/A1 hold56/I _3753_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_174_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6471_ _6946_/Q _6245_/Z _6273_/Z _6978_/Q _7124_/Q _6288_/Z _6472_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3683_ _7250_/Q _6898_/Q _6900_/Q _3683_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5422_ _5034_/B _4866_/Z _5422_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
Xoutput235 _4054_/Z mgmt_gpio_out[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_161_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5353_ _5353_/A1 _5387_/A2 _5353_/B _5354_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xoutput213 _4068_/Z mgmt_gpio_out[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput224 _6742_/Q mgmt_gpio_out[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput202 _3376_/ZN mgmt_gpio_oeb[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_126_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput246 _4057_/Z mgmt_gpio_out[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4304_ _6829_/Q _7279_/RN _4312_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xoutput257 _6886_/Q pll90_sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput268 _6883_/Q pll_sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5284_ _5284_/A1 _5369_/B _5284_/A3 _5277_/I _5286_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_101_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput279 _6667_/Q pll_trim[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4235_ _4234_/Z hold771/Z _4245_/S _4235_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7023_ _7023_/D _7260_/RN _7023_/CLK _7023_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_68_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4166_ hold271/Z hold745/Z _4166_/S _4166_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4097_ _4097_/A1 _4415_/B _6828_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6807_ _6807_/D _7243_/CLK _6807_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4999_ _4999_/A1 _4999_/A2 _4998_/Z _5341_/B _5000_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_23_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6738_ _6738_/D _7258_/RN _6738_/CLK _6738_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6669_ _6669_/D _7238_/RN _6669_/CLK _6669_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_152_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4020_ _4014_/Z _4020_/A2 _6746_/Q _4003_/Z _4021_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_38_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5971_ _7228_/Q _7227_/Q _6211_/B1 _6210_/A2 _5971_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4922_ _4373_/Z _4385_/Z _4922_/A3 _4922_/A4 _4923_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_64_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4853_ _4853_/A1 _5287_/B _4784_/Z _4501_/B _4853_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_60_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4784_ _5420_/A3 _3402_/I _4456_/B _5051_/S _4784_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3804_ _6842_/Q _3930_/B1 _3884_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_147_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3735_ _7113_/Q _3917_/A2 _5674_/A1 _7031_/Q _3735_/C _3760_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6523_ _6866_/Q _6272_/Z _6290_/Z _6708_/Q _6526_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_134_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6454_ _7100_/Q _6250_/Z _6302_/Z _7092_/Q _6292_/Z _7148_/Q _6466_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_106_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5405_ _5454_/A1 _4791_/Z _5126_/I _5406_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3666_ _6929_/Q _3935_/A2 _5656_/A1 _7017_/Q _3667_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_161_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6385_ _6385_/A1 _6385_/A2 _6385_/A3 _6384_/Z _6385_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3597_ _6681_/Q _3546_/Z _3945_/C2 _6689_/Q _3913_/A2 input19/Z _3601_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5336_ _5412_/A1 _5412_/A3 _5338_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5267_ _4898_/C _5428_/A4 _4893_/Z _5267_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_102_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4218_ _4217_/Z hold557/Z _4228_/S _4218_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7006_ _7006_/D _7260_/RN _7006_/CLK _7006_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5198_ _5309_/B2 _5205_/A1 _5351_/C _5205_/B1 _5198_/C _5476_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_96_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4149_ _3507_/Z _3537_/Z _5520_/C _4157_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_83_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3520_ _3485_/Z _3519_/Z _4225_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_155_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold707 _6907_/Q hold707/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_6_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold718 _4175_/Z _6717_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3451_ _3451_/I0 input58/Z _6730_/Q _3451_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold729 _7172_/Q hold729/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6170_ _6971_/Q _5979_/Z _5981_/Z _6939_/Q _5996_/Z _7085_/Q _6181_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3382_ _6785_/Q _6528_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_5121_ _5121_/A1 _4876_/C _5457_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_34_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5052_ _4936_/I _5051_/Z _5064_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_38_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4003_ _5954_/A3 _7225_/Q _7226_/Q _7223_/Q _4003_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_66_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_330 net763_422/I _6895_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_341 net663_341/I _6884_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5954_ _7223_/Q _5954_/A2 _5954_/A3 _6746_/Q _5954_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4905_ _4467_/B _4495_/Z _5263_/A2 _5324_/A1 _4905_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_178_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5885_ _4103_/I hold882/Z _5892_/S _5885_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4836_ _5420_/A3 _4549_/Z _3402_/I _4836_/A4 _4836_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_119_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4767_ _4716_/Z _4764_/Z _5118_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_14_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6506_ _6820_/Q _6262_/Z _6269_/Z _6847_/Q _6512_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_135_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4698_ _5097_/A1 _4704_/A2 _4698_/B _5094_/B _4714_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3718_ input16/Z _3913_/A2 _3945_/B1 _7090_/Q _3719_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3649_ _3648_/Z hold989/Z _3899_/S _6874_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6437_ _6437_/I _6438_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6368_ _7145_/Q _6292_/Z _6383_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_88_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5319_ _5392_/B _4801_/Z _5319_/A3 _5319_/A4 _5319_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_102_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6299_ _7236_/Q _6533_/A3 _6452_/A4 _6302_/A4 _6299_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold12 hold12/I hold12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold23 hold23/I hold23/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_69_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold34 hold34/I hold34/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold45 hold45/I hold45/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold56 hold56/I hold56/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_91_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold67 hold67/I hold67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold89 hold89/I hold89/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_29_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold78 hold78/I hold78/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_56_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_45_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_9 _5508_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_2__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7269_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_79_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet613_260 _4073__43/I _6965_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_271 net613_273/I _6954_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_282 net763_424/I _6943_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet613_293 net613_293/I _6932_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5670_ hold89/Z hold62/Z _5673_/S hold90/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4621_ _4367_/Z _4555_/B _5291_/C _5353_/A1 _5353_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_148_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4552_ _4549_/Z _4551_/Z _5011_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_117_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7271_ _7271_/D _7279_/RN _7279_/CLK _7271_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold515 _5807_/Z _7145_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold526 _5687_/Z _7039_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold504 _7129_/Q hold504/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4483_ _4489_/A1 _4692_/B _4483_/B _4687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_3503_ _3497_/I hold629/Z _5857_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_7_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3434_ _3442_/B _3409_/Z _3434_/B _3435_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold537 _6905_/Q hold537/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold548 _4222_/Z _6751_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold559 _6896_/Q hold559/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6222_ _6823_/Q _5964_/Z _5999_/Z _6848_/Q _6729_/Q _6000_/Z _6228_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3365_ _7039_/Q _3365_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6153_ _6946_/Q _5972_/Z _6021_/Z _7002_/Q _6155_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3296_ _7294_/Q _4084_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5104_ _5104_/A1 _5139_/A3 _5094_/B _5104_/A4 _5104_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6084_ _6084_/A1 _6084_/A2 _6084_/A3 _6084_/A4 _6084_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_98_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5035_ _5035_/A1 _5032_/Z _5204_/C _5035_/A4 _5035_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6986_ _6986_/D _7260_/RN _6986_/CLK _6986_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_179_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5937_ _6279_/A3 _7233_/Q _6302_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_53_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5868_ hold271/Z hold958/Z _5874_/S _5868_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4819_ _4422_/Z _4624_/Z _4673_/Z _4483_/B _4819_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5799_ hold62/Z hold223/Z hold7/Z _7138_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput102 wb_adr_i[16] _4391_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_103_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput135 wb_dat_i[16] _6579_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput113 wb_adr_i[26] _4031_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput124 wb_adr_i[7] _4501_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_163_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput146 wb_dat_i[26] _6585_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput157 wb_dat_i[7] _3400_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_172_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6840_ _6840_/D _7210_/RN _6840_/CLK _6840_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6771_ _6771_/D _7258_/RN _6771_/CLK _6771_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_90_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3983_ _6659_/Q _3972_/Z _3983_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5722_ hold86/Z hold508/Z _5727_/S _5722_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5653_ hold522/Z hold29/Z _5655_/S _7009_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4604_ _4501_/B _4604_/A2 _4604_/A3 _4604_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_175_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5584_ _5584_/A1 hold18/Z _5592_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_4535_ _5414_/A2 _4534_/Z _5323_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_144_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold301 _5753_/Z _7097_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_7_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold312 _6771_/Q hold312/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_117_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold334 _7194_/Q hold334/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold323 _5881_/Z _7211_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7254_ _7254_/D _7258_/RN _7258_/CLK _7254_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4466_ _4454_/Z _4367_/Z _4363_/Z _4690_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_117_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold378 _5847_/Z _7181_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold345 _7047_/Q hold345/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold356 _7056_/Q hold356/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold367 _5506_/Z _6885_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4397_ _5002_/A3 _5002_/A4 _4397_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3417_ _3416_/Z _7304_/Q _6733_/Q _3417_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7185_ _7185_/D _7221_/RN _7185_/CLK _7185_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold389 _7078_/Q hold389/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6205_ _6193_/Z _6204_/Z _6528_/B1 _6168_/C _6555_/C _6206_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3348_ _7169_/Q _3348_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6136_ _6136_/I0 _7245_/Q _6555_/C _6136_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xhold1001 _7282_/Q _4041_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XTAP_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6067_ _6067_/A1 _5991_/Z _6072_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_46_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5018_ _5389_/B _5439_/B2 _5018_/B _5390_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_2517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_455 net813_470/I _6710_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_466 net413_79/I _6699_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet813_477 net813_483/I _6688_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_488 net813_489/I _6677_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_499 net813_499/I _6666_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6969_ hold40/Z _7238_/RN _6969_/CLK _6969_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_146_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold890 _6840_/Q hold890/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_150_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4320_ hold6/Z _3535_/Z hold38/Z hold11/Z _4322_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_114_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4251_ hold62/Z hold560/Z _4252_/S _4251_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4182_ _4182_/A1 hold18/Z _4184_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_110_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_26__1359_ clkbuf_opt_1_0__1359_/Z net763_429/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_68_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_106__1359_ clkbuf_4_5_0__1359_/Z net613_273/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_89__1359_ clkbuf_4_13_0__1359_/Z net613_255/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_91_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6823_ _6823_/D _7210_/RN _6823_/CLK _6823_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6754_ _6754_/D _7260_/RN _6754_/CLK _6754_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3966_ _3966_/I _6868_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5705_ hold360/Z hold52/Z _5709_/S _5705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6685_ _6685_/D _7297_/RN _6685_/CLK _6685_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_176_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5636_ hold15/Z hold171/Z _5637_/S _5636_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3897_ _3897_/A1 _3897_/A2 _3855_/Z _3896_/Z _6565_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_148_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5567_ hold113/Z hold699/Z _5574_/S _5567_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4518_ _4835_/A2 _4456_/B _5269_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold142 _7051_/Q hold142/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold153 _5673_/Z _7027_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold131 _6678_/Q hold131/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5498_ hold424/Z _4103_/I _5502_/S _5498_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold120 _6996_/Q hold120/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4449_ _4853_/A1 _5464_/A1 _4501_/B _4451_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7237_ _7237_/D _7237_/RN _4067_/I1 _7237_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_105_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold164 _5784_/Z _7125_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold175 _5627_/Z _6986_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold186 _7026_/Q hold186/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold197 _6705_/Q hold197/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_137_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7168_ _7168_/D _7258_/RN _7168_/CLK _7168_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_59_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7099_ _7099_/D _7219_/RN _7099_/CLK _7099_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_85_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6119_ _7155_/Q _5960_/Z _6133_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_3037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet413_61 net413_61/I _7164_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_94 net413_94/I _7131_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__20 _4073__20/I _7205_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_72 net413_72/I _7153_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__42 net413_65/I _7183_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__31 net413_56/I _7194_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet413_83 net413_83/I _7142_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3820_ _3527_/Z _3578_/Z _4274_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3751_ _3751_/A1 _3751_/A2 _3732_/Z _3751_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_20_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6470_ _7050_/Q _6241_/Z _6251_/Z _6986_/Q _6268_/Z hold26/I _6472_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3682_ hold41/I _5638_/A1 _3912_/B1 _6888_/Q _3686_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_127_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5421_ _5420_/Z _5421_/A2 _5421_/A3 _5421_/A4 _5489_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_64_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5352_ _5191_/Z _5352_/A2 _5285_/B _5020_/Z _5352_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_160_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput214 _4067_/Z mgmt_gpio_out[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xoutput225 _6908_/Q mgmt_gpio_out[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput203 _3375_/ZN mgmt_gpio_oeb[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput236 _6765_/Q mgmt_gpio_out[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4303_ hold880/Z hold271/Z _4303_/S _4303_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput247 _4075_/Z pad_flash_clk VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xoutput258 _6887_/Q pll90_sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_142_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5283_ _5278_/C _4554_/Z _5283_/B _5471_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_87_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7022_ _7022_/D _7260_/RN _7022_/CLK _7022_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xoutput269 _6884_/Q pll_sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4234_ hold306/Z hold86/Z _4244_/S _4234_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4165_ _4103_/I hold672/Z _4166_/S _4165_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4096_ _4097_/A1 _4096_/A2 _6829_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_56_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6806_ _6806_/D _7265_/CLK _6806_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4998_ _5340_/A1 _4998_/A2 _5262_/A2 _5343_/A2 _4998_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_56_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6737_ _6737_/D _7258_/RN _6737_/CLK _6737_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3949_ _3949_/A1 _3949_/A2 _3949_/A3 _3949_/A4 _3949_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_136_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6668_ _6668_/D _7238_/RN _6668_/CLK _6668_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_20_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6599_ _6599_/I0 _7276_/Q _6602_/S _7276_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5619_ hold2/Z hold150/Z _5619_/S _5619_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_72__1359_ clkbuf_4_13_0__1359_/Z net513_191/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_74_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5970_ _7102_/Q _5967_/Z _5969_/Z _7118_/Q _5974_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4921_ _4920_/Z _4890_/I _4926_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4852_ _4852_/A1 _5106_/A2 _4852_/A3 _4855_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_178_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3803_ _3529_/Z _3680_/Z _3930_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_147_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4783_ _4836_/A4 _4530_/I _5137_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3734_ _3734_/I _3735_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6522_ _6696_/Q _6282_/Z _6302_/Z _6712_/Q _6526_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_158_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6453_ _7066_/Q _6257_/Z _6275_/Z _7042_/Q _6300_/Z _7108_/Q _6466_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3665_ _7009_/Q _3934_/A2 _3954_/A2 _6993_/Q _3674_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_146_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5404_ _5404_/A1 _5314_/Z _5404_/A3 _5404_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6384_ _6384_/A1 _6384_/A2 _6380_/Z _6383_/Z _6384_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3596_ _3592_/Z _3596_/A2 _3596_/A3 _3596_/A4 _3596_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5335_ _4908_/Z _5245_/Z _5481_/B1 _4905_/Z _5335_/C _5447_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_142_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5266_ _5265_/Z _5341_/B _4994_/Z _5266_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_141_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4217_ _6779_/Q hold86/Z _4227_/S _4217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7005_ _7005_/D _7210_/RN _7005_/CLK _7005_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5197_ _5346_/A2 _5349_/A1 _5276_/C _5205_/A1 _5197_/C _5390_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_84_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4148_ hold709/Z hold271/Z _4148_/S _4148_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4079_ _4079_/I _4079_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_1__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7265_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_78_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold708 _5538_/Z _6907_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold719 _6842_/Q hold719/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3450_ _3450_/A1 _3450_/A2 _7292_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_130_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3381_ _6931_/Q _6500_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5120_ _5118_/Z _5238_/A1 _5127_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5051_ _4698_/B _5343_/A1 _5051_/S _5051_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_97_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4002_ _7225_/Q _7226_/Q _5954_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_112_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_320 _4073__48/I _6905_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet663_342 net713_358/I _6883_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_331 net763_445/I _6894_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_92_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5953_ _5953_/I0 _7239_/Q _5955_/S _7239_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4904_ _5263_/A2 _4903_/Z _5255_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_178_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5884_ _3485_/Z _3515_/Z _5520_/C _5892_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_80_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4835_ _4555_/C _4835_/A2 _5129_/A3 _5420_/A2 _5368_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4766_ _4766_/A1 _4766_/A2 _4762_/Z _4765_/Z _4770_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_14_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3717_ _6928_/Q _3935_/A2 _3943_/A2 _7072_/Q _6895_/Q _5528_/S _3719_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6505_ _6853_/Q _6241_/Z _6297_/Z _7076_/Q _6512_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_107_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4697_ _4467_/B _4463_/Z _5302_/B _5099_/A2 _4697_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_134_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3648_ _6570_/I0 _6873_/Q _3898_/S _3648_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6436_ hold45/I _6292_/Z _6300_/Z _7107_/Q _6437_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_136_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6367_ _7253_/Q _6367_/I1 _6558_/S _7253_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3579_ _3533_/Z _3578_/Z _3959_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5318_ _5318_/A1 _5314_/Z _5316_/Z _5318_/A4 _5320_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_96_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6298_ _7158_/Q _6296_/Z _6297_/Z _6698_/Q _6298_/C _6307_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold13 hold13/I hold13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_29_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5249_ _5410_/A1 _5245_/Z _5250_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_103_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold24 hold24/I hold24/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold46 hold46/I hold46/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold35 hold35/I hold35/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_75_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold79 hold79/I hold79/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold68 hold68/I hold68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_28_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold57 hold57/I hold57/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_56_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet613_283 net713_394/I _6942_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_272 net613_276/I _6953_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet613_261 net413_83/I _6964_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet613_294 net613_295/I _6931_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4620_ _4557_/Z _4604_/Z _5353_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_163_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4551_ _5129_/A3 _5051_/S _3401_/I _3402_/I _4551_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_128_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4482_ _4381_/Z _4485_/A2 _4390_/Z _5170_/A3 _4486_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_7270_ _7270_/D _7279_/RN _7279_/CLK _7270_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold505 _5789_/Z _7129_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold527 _7105_/Q hold527/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3502_ _3617_/A1 _3501_/Z _3904_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold516 _6985_/Q hold516/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3433_ _3427_/Z _3433_/A2 _3433_/B _3435_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold549 _6903_/Q hold549/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold538 _5535_/Z _6905_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6221_ _6725_/Q _5984_/Z _5997_/Z _6717_/Q _6695_/Q _5980_/Z _6228_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_131_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6152_ _6152_/A1 _6152_/A2 _6152_/A3 _6152_/A4 _6152_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3364_ _7047_/Q _3364_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5103_ _5103_/A1 _5101_/Z _5103_/A3 _5308_/A2 _5108_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3295_ _7283_/Q _4022_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6083_ _6975_/Q _5964_/Z _5999_/Z _7031_/Q _6084_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ _5190_/A2 _4604_/Z _5003_/Z _5034_/B _5204_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_66_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6985_ _6985_/D _7260_/RN _6985_/CLK _6985_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5936_ _6745_/Q _7233_/Q _7232_/Q _5936_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_90_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5867_ hold113/Z hold578/Z _5874_/S _5867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4818_ _4624_/Z _4817_/Z _5313_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5798_ hold52/Z hold222/Z hold7/Z _7137_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4749_ _4703_/Z _5230_/B _5313_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_162_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6419_ _6744_/Q _7254_/Q _6419_/B _6420_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_89_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput136 wb_dat_i[17] _6582_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput103 wb_adr_i[17] _4391_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput114 wb_adr_i[27] _4027_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput125 wb_adr_i[8] _4388_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput147 wb_dat_i[27] _6588_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput158 wb_dat_i[8] _6579_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3982_ _3981_/Z _6660_/Q _3988_/S _6660_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6770_ _6770_/D _7237_/RN _6770_/CLK _6770_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_90_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_189_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5721_ hold271/Z hold964/Z _5727_/S _5721_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5652_ hold355/Z hold62/Z _5655_/S _7008_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4603_ _4580_/B _4604_/A3 _5351_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_175_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_49__1359_ net663_304/I _4073__36/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_129__1359_ net613_253/I _4073__43/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_50_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5583_ _6947_/Q hold2/Z hold23/I hold3/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4534_ _4782_/A1 _4736_/A3 _4736_/A1 _4436_/B _4534_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold302 _7155_/Q hold302/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold313 _4256_/Z _6771_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_117_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold335 _5862_/Z _7194_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold324 _7163_/Q hold324/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7253_ _7253_/D _7258_/RN _7258_/CLK _7253_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold346 _5696_/Z _7047_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4465_ _5315_/A1 _4481_/A2 _4473_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold368 _7106_/Q hold368/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold357 _5706_/Z _7056_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4396_ _5385_/A1 _4385_/Z _4922_/A3 _4424_/B _5002_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3416_ _7305_/Q _3415_/Z _3416_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xhold379 _7221_/Q hold379/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_98_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7184_ _7184_/D _7258_/RN _7184_/CLK _7184_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_6204_ _6198_/Z _6201_/Z _6204_/A3 _6204_/A4 _6204_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3347_ _7177_/Q _3732_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_98_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6135_ _6127_/Z _6134_/Z _6447_/B1 _6168_/C _6136_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold1002 _7294_/Q _3440_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6066_ _7023_/Q wire348/Z _6211_/B1 _6991_/Q _6067_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_58_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5017_ _5017_/A1 _5197_/C _5019_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_456 net413_58/I _6709_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_467 net813_467/I _6698_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_489 net813_489/I _6676_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_478 net813_483/I _6687_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6968_ _6968_/D _7238_/RN _6968_/CLK hold72/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_107_1032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5919_ _6021_/A2 _6015_/A3 _5984_/A1 _6745_/Q _5919_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_50_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6899_ hold16/Z _7238_/RN _6899_/CLK _6899_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_41_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold891 _4334_/Z _6840_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold880 _6810_/Q hold880/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4250_ hold52/Z hold118/Z _4252_/S _4250_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4181_ hold271/Z hold749/Z _4181_/S _4181_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6822_ _6822_/D _7210_/RN _6822_/CLK _6822_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_90_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3965_ _6564_/I0 _3965_/A2 hold993/Z _3899_/S _3966_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6753_ _6753_/D input75/Z _6753_/CLK _6753_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_32_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5704_ hold473/Z hold86/Z _5709_/S _5704_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6684_ _6684_/D _7297_/RN _6684_/CLK _6684_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3896_ _3860_/Z _3869_/Z _3885_/Z _3895_/Z _3896_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_109_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5635_ hold29/Z hold510/Z _5637_/S _5635_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5566_ hold6/Z _3521_/Z hold38/Z hold11/Z _5574_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold110 _6881_/Q hold110/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4517_ _5165_/A4 _5003_/A2 _4491_/B _5438_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_7305_ _7305_/D _6657_/Z _4072_/B2 _7305_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_117_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold143 _5700_/Z _7051_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5497_ _5647_/A1 hold33/Z hold18/Z hold11/Z _5502_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold132 _4124_/Z _6678_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold121 _6940_/Q hold121/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4448_ _3401_/I _5288_/C _4369_/Z _5288_/B _4451_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_160_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7236_ _7236_/D _7237_/RN _4067_/I1 _7236_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xhold176 _7149_/Q hold176/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold165 _6908_/Q hold165/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold154 _6995_/Q hold154/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold198 _4157_/Z _6705_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold187 _5672_/Z _7026_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4379_ _4853_/A1 _5464_/A1 _4604_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_99_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7167_ _7167_/D _7219_/RN _7167_/CLK _7167_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_86_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7098_ _7098_/D _7219_/RN _7098_/CLK _7098_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6118_ _7057_/Q _5924_/Z _6168_/C _6127_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_3027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6049_ _6942_/Q _5972_/Z _6021_/Z _6998_/Q _6049_/C _6053_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_58_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_112__1359_ clkbuf_4_5_0__1359_/Z net413_89/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_154_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_95 net413_96/I _7130_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__21 _4073__21/I _7204_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__32 net413_58/I _7193_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__10 _4073__47/I _7215_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet413_73 net413_73/I _7152_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_84 net413_86/I _7141_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet413_62 net413_62/I _7163_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__43 _4073__43/I _7182_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3750_ _7007_/Q _3934_/A2 _5638_/A1 _6999_/Q _3916_/B1 _6881_/Q _3751_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_186_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3681_ _3527_/Z _3680_/Z _3912_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_174_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5420_ _5420_/A1 _5420_/A2 _5420_/A3 _4456_/B _5420_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xnet713_400 net763_429/I _6774_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5351_ _5356_/A1 _5387_/A2 _5356_/B _5351_/C _5352_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xoutput215 _4066_/Z mgmt_gpio_out[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_142_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput226 _6909_/Q mgmt_gpio_out[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput204 _3374_/ZN mgmt_gpio_oeb[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_57_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput237 _4055_/Z mgmt_gpio_out[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5282_ _5281_/C _4467_/B _5399_/A2 _4683_/Z _5283_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_114_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput248 _4094_/ZN pad_flash_clk_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4302_ hold815/Z _4103_/I _4303_/S _4302_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput259 _6888_/Q pll90_sel[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4233_ _4232_/Z hold838/Z _4245_/S _4233_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7021_ _7021_/D _7260_/RN _7021_/CLK _7021_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_136_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4164_ _5520_/C _3552_/Z hold637/Z _5821_/A3 _4166_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4095_ _4097_/A1 _4900_/B _6831_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_96_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6805_ _6805_/D _7269_/CLK _6805_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6736_ _6736_/D _7258_/RN _6736_/CLK _6736_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4997_ _4546_/Z _4716_/Z _4997_/B _4997_/C _4999_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_183_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3948_ input43/Z _4210_/S _4194_/A1 input52/Z _3948_/C1 input61/Z _3949_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_20_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3879_ _7087_/Q _3945_/B1 _3952_/A2 _7045_/Q _3950_/C1 _6844_/Q _3880_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6667_ _6667_/D _7297_/RN _6667_/CLK _6667_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_6598_ _6598_/A1 _4313_/Z _6598_/B _6599_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_164_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5618_ hold15/Z hold182/Z _5619_/S _5618_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5549_ hold113/Z hold257/Z _5556_/S _5549_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_0__f_wb_clk_i clkbuf_0_wb_clk_i/Z _7243_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7219_ _7219_/D _7219_/RN _7219_/CLK _7219_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_48_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4920_ _5130_/B2 _5420_/A3 _4367_/Z _4920_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_61_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4851_ _5287_/C _4833_/Z _4852_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_127_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3802_ _3509_/Z _3540_/Z _3925_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_165_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4782_ _4782_/A1 _4510_/Z _5302_/B _5099_/A1 _5213_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_158_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3733_ _7193_/Q _3909_/A2 _5683_/A1 _7039_/Q _3952_/A2 _7047_/Q _3734_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6521_ _6521_/A1 _6521_/A2 _6521_/A3 _6521_/A4 _6521_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_174_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6452_ _7074_/Q _6484_/A2 _6484_/A3 _6452_/A4 _6456_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3664_ input17/Z _3913_/A2 _5674_/A1 _7033_/Q _3674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_162_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5403_ _4699_/Z _5403_/A2 _5456_/A2 _5403_/B2 _5403_/C _5404_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_173_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6383_ _6383_/A1 _6383_/A2 _6383_/A3 _6383_/A4 _6383_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3595_ _6995_/Q _3954_/A2 _3927_/A2 _6705_/Q _3596_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5334_ _5334_/A1 _5334_/A2 _5334_/A3 _5334_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_170_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5265_ _5265_/A1 _4991_/C _5392_/B _5265_/A4 _5265_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_141_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5196_ _5347_/A1 _5437_/A1 _5195_/Z _5347_/A3 _5196_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_134_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4216_ _4215_/Z hold827/Z _4228_/S _4216_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7004_ _7004_/D _7297_/RN _7004_/CLK _7004_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_69_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4147_ hold809/Z _4103_/I _4148_/S _4147_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4078_ _4081_/A1 input86/Z _4079_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_23_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6719_ _6719_/D _7210_/RN _6719_/CLK _6719_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_164_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold709 _6697_/Q hold709/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3380_ _6930_/Q _6473_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_124_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5050_ _5343_/A2 _5389_/A2 _5078_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_85_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4001_ _4001_/I _6836_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_310 net663_310/I _6915_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_321 _4073__48/I _6904_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_332 net713_387/I _6893_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_343 net813_471/I _6882_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5952_ _6746_/Q _6744_/Q _5952_/A3 _5952_/B _5955_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_81_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4903_ _4467_/B _4407_/Z _4495_/Z _5259_/A1 _4903_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_80_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5883_ hold2/Z hold242/Z _5883_/S _5883_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4834_ _4834_/A1 _4834_/A2 _4846_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_61_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4765_ _4765_/A1 _5302_/B _4700_/Z _5226_/C _4765_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_146_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3716_ _7130_/Q _3930_/A2 _3925_/A2 input7/Z _5647_/A1 _3904_/A2 _3719_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6504_ _6789_/Q _6245_/Z _6274_/Z _6851_/Q _6512_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4696_ _5099_/A2 _4695_/Z _4704_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_161_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3647_ _3647_/A1 _3625_/Z _3646_/Z _3647_/A4 _6570_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6435_ _7187_/Q _6282_/Z _6299_/Z _7057_/Q _6993_/Q _6237_/Z _6439_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_143_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6366_ _6366_/I _6367_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3578_ _3653_/A1 hold338/Z _3617_/A1 hold629/Z _3578_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_143_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5317_ _5317_/A1 _5454_/A1 _5318_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold14 hold14/I hold14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6297_ _6300_/A2 _6484_/A3 _5943_/S _5942_/S _6297_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5248_ _5246_/Z _5248_/A2 _5442_/A2 _5056_/C _5248_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_152_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold36 hold36/I hold36/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_130_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold25 hold25/I hold25/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold47 hold47/I hold47/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5179_ _5240_/B _5343_/A2 _5179_/B _5242_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_102_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold69 hold69/I hold69/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold58 hold58/I hold58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_72_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet613_262 net613_276/I _6963_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_273 net613_273/I _6952_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xnet613_295 net613_295/I _6930_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet613_284 net713_394/I _6941_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4550_ _4454_/Z _5269_/A2 _5368_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_4481_ _4481_/A1 _4481_/A2 _4486_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_143_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3501_ _3499_/I _3305_/I hold21/Z _3501_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_7_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold517 _5626_/Z _6985_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold506 _7049_/Q hold506/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3432_ _3432_/I _7299_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold528 _5762_/Z _7105_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold539 _7153_/Q hold539/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6220_ _6217_/Z _6220_/A2 _6220_/A3 _6220_/A4 _6220_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3363_ _7055_/Q _3363_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6151_ _7148_/Q _5987_/Z _6015_/Z _7010_/Q _6152_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5102_ _4586_/Z _4817_/Z _5103_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6082_ _7169_/Q _6006_/Z _6014_/Z _6959_/Q _6084_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3294_ _7300_/Q _4081_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5033_ _5035_/A4 _5032_/Z _5388_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6984_ _6984_/D _7297_/RN _6984_/CLK _6984_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5935_ _6282_/A2 _6279_/A3 _6300_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_80_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5866_ _3485_/Z _3507_/Z hold6/Z _5874_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_33_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4817_ _5420_/A3 _5287_/B _3402_/I _5269_/A2 _4817_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_21_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5797_ hold86/Z hold117/Z hold7/Z _7136_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_4_11_0__1359_ clkbuf_0__1359_/Z net463_109/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_119_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4748_ _4510_/Z _5302_/B _5099_/A1 _5226_/C _4748_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_174_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4679_ _4670_/Z _5451_/C _4685_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_134_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6418_ _6411_/Z _6417_/Z _6418_/B1 _6286_/Z _6555_/C _6419_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_162_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6349_ _7200_/Q _6272_/Z _6282_/Z _7184_/Q _6296_/Z _7160_/Q _6356_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_1_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput104 wb_adr_i[18] _4391_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput115 wb_adr_i[28] _4027_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput126 wb_adr_i[9] _4388_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_131_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_0__1359_ _4072_/ZN clkbuf_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput148 wb_dat_i[28] _6591_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput137 wb_dat_i[18] _6585_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput159 wb_dat_i[9] _6582_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_172_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3981_ _3981_/A1 _3981_/A2 _3981_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5720_ _4103_/I hold952/Z _5727_/S _5720_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5651_ hold251/Z hold52/Z _5655_/S _7007_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4602_ _4524_/Z _5399_/A2 _4554_/Z _5364_/B _5285_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5582_ _6946_/Q hold15/Z hold23/Z hold24/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4533_ _4736_/A3 _4690_/C _4713_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_156_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7252_ _7252_/D _7258_/RN _7258_/CLK _7252_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold303 _5818_/Z _7155_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold314 _7107_/Q hold314/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold325 _5827_/Z _7163_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold358 _7071_/Q hold358/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold347 _6919_/Q hold347/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold336 _6861_/Q _3307_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4464_ _4456_/B _5051_/S _4460_/B _4436_/B _4464_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold369 _5763_/Z _7106_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6203_ _6724_/Q _5984_/Z _6000_/Z _6728_/Q _6710_/Q _6006_/Z _6204_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_4395_ _4580_/C _4489_/A1 _4483_/B _5002_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_3415_ _7304_/Q _7303_/Q _3415_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_113_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7183_ _7183_/D _7210_/RN _7183_/CLK _7183_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3346_ _7185_/Q _3346_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6134_ _6134_/A1 _6134_/A2 _6134_/A3 _6133_/Z _6134_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_113_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6065_ _7243_/Q _6065_/I1 _6558_/S _7243_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5016_ _5438_/C _4551_/Z _4586_/Z _5003_/Z _5016_/B2 _5197_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_85_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_457 net813_472/I _6708_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _6967_/D _7260_/RN _6967_/CLK _6967_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xnet813_479 net813_482/I _6686_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet813_468 net413_71/I _6697_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5918_ _6745_/Q _5917_/Z _5913_/I _6021_/A2 _7228_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_167_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6898_ hold35/Z _7260_/RN _6898_/CLK _6898_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_167_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5849_ hold113/Z hold576/Z _5856_/S _5849_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold870 _6752_/Q hold870/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold881 _4303_/Z _6810_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_27_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold892 _7102_/Q hold892/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_55__1359_ net663_324/I net413_94/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_17_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_135__1359_ net613_293/I net813_485/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_45_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4180_ _4103_/I hold675/Z _4181_/S _4180_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6821_ _6821_/D _7210_/RN _6821_/CLK _6821_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_177_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3964_ _3898_/S _3899_/S _3965_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6752_ _6752_/D _7260_/RN _6752_/CLK _6752_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5703_ hold948/Z hold271/Z _5709_/S _5703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6683_ _6683_/D _7297_/RN _6683_/CLK _6683_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3895_ _3895_/A1 _3889_/Z _3895_/A3 _3894_/Z _3895_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_164_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5634_ hold62/Z hold83/Z _5637_/S hold84/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7304_ _7304_/D _6656_/Z _7304_/CLK _7304_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5565_ hold2/Z hold199/Z _5565_/S _5565_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold100 _4269_/Z _6783_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4516_ _5003_/A2 _4561_/A2 _5389_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_176_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold133 _6659_/Q hold133/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5496_ hold271/Z _6877_/Q _5496_/S _5496_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold111 _5501_/Z _6881_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold144 _7080_/Q hold144/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold122 _6948_/Q hold122/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4447_ _5420_/A2 _4853_/A1 _5270_/A1 _4501_/B _4504_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_176_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7235_ _7235_/D _7237_/RN _4067_/I1 _7235_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
Xhold177 _5811_/Z _7149_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold166 _5540_/Z _6908_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold155 _5637_/Z _6995_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_160_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold199 _6931_/Q hold199/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold188 _7018_/Q hold188/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7166_ _7166_/D _7219_/RN _7166_/CLK _7166_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4378_ _5281_/C _5464_/A1 _4648_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_101_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6117_ _7073_/Q _7231_/Q _6210_/C _6117_/A4 _6128_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3329_ _7234_/Q _5942_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_7097_ _7097_/D _7219_/RN _7097_/CLK _7097_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_59_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6048_ _5925_/Z _6048_/A2 _6048_/B _6048_/C _6049_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XTAP_3039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet413_52 net413_68/I _7173_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__22 _4073__22/I _7203_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__11 _4073__7/I _7214_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_74 net413_74/I _7151_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet413_63 net413_67/I _7162_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_85 net413_89/I _7140_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet413_96 net413_96/I _7129_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__33 _4073__36/I _7192_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__44 net413_61/I _7181_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3680_ _3489_/I _3492_/Z _3497_/I hold629/Z _3680_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xnet713_401 net763_431/I _6773_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5350_ _5350_/A1 _5350_/A2 _5350_/A3 _5350_/A4 _5350_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xoutput216 _6735_/Q mgmt_gpio_out[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_154_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput205 _3373_/ZN mgmt_gpio_oeb[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput238 _4048_/Z mgmt_gpio_out[36] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput227 _6910_/Q mgmt_gpio_out[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5281_ _5288_/A1 _5281_/A2 _5281_/B _5281_/C _5369_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xoutput249 _4074_/Z pad_flash_csb VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4301_ _4301_/A1 hold18/Z _4303_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_4232_ hold831/Z hold271/Z _4244_/S _4232_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7020_ _7020_/D _7260_/RN _7020_/CLK _7020_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_68_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4163_ hold974/Z hold271/Z _4163_/S _4163_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4094_ _4094_/I _4094_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4996_ _5083_/C _4997_/C _4716_/Z _4422_/Z _5341_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6804_ _6804_/D _7265_/CLK _6804_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6735_ _6735_/D _7258_/RN _6735_/CLK _6735_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3947_ _7094_/Q _3947_/A2 _3947_/B1 _6716_/Q _3949_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_104_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3878_ _6904_/Q _5532_/A1 _3935_/B1 _6850_/Q _3885_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6666_ _6666_/D _7297_/RN _6666_/CLK _6666_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_6597_ _6834_/Q _6597_/A2 _6597_/B1 _6835_/Q _6836_/Q _6597_/C2 _6598_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5617_ hold29/Z hold54/Z _5619_/S hold55/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5548_ _3485_/Z _3542_/Z _6652_/A2 hold6/Z _5556_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_173_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5479_ _5479_/A1 _5479_/A2 _5479_/A3 _5479_/A4 _5479_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7218_ _7218_/D _7219_/RN _7218_/CLK _7218_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_87_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7149_ _7149_/D _7237_/RN _7149_/CLK _7149_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_63_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4850_ _5287_/C _4817_/Z _5106_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_45_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3801_ _3509_/Z _3653_/Z _3928_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_1990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4781_ _4781_/A1 _5121_/A1 _5456_/B _5122_/B _4790_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_60_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6520_ _6710_/Q _5948_/Z _6292_/Z _6722_/Q _6521_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3732_ _3732_/A1 _5857_/A3 _5839_/A3 _3552_/Z _3732_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_174_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6451_ _7212_/Q _6256_/Z _6464_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_9_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3663_ _3663_/A1 _3663_/A2 _3663_/A3 _3663_/A4 _3663_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_173_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6382_ _7039_/Q _6275_/Z _6300_/Z _7105_/Q _6383_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5402_ _5480_/A1 _5480_/A2 _5406_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5333_ _4761_/I _5481_/B1 _5334_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_155_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3594_ _6963_/Q _3957_/A2 _3927_/C2 input33/Z _5575_/A1 _6947_/Q _3596_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_173_1034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5264_ _5264_/A1 _5412_/A3 _5264_/A3 _5263_/Z _5265_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5195_ _5350_/A1 _5350_/A3 _5195_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_130_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7003_ _7003_/D _7260_/RN _7003_/CLK _7003_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4215_ hold763/Z hold271/Z _4227_/S _4215_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4146_ _4146_/A1 hold18/Z _4148_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_56_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4077_ _4077_/I _4077_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4979_ _4419_/Z _4973_/Z _4979_/B _4979_/C _4986_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_137_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6718_ _6718_/D _7210_/RN _6718_/CLK _6718_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6649_ _7237_/RN _6657_/A2 _6649_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_165_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4000_ _6836_/Q _4097_/A1 _6831_/Q _4001_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xnet663_311 net663_313/I _6914_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet663_322 _4073__48/I _6903_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_344 net813_471/I _6881_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_333 net813_499/I _6892_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_9_0__1359_ clkbuf_0__1359_/Z net413_53/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_81_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5951_ _7225_/Q _7226_/Q _5951_/A3 _6746_/Q _5952_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_65_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4902_ _4436_/B _4494_/Z _5323_/B _4902_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_5882_ hold15/Z hold428/Z _5883_/S _5882_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4833_ _4422_/Z _4530_/I _4878_/A2 _4483_/B _4833_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4764_ _4765_/A1 _5302_/B _4764_/A3 _4692_/C _4764_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6503_ _7258_/Q _6503_/I1 _6558_/S _7258_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3715_ _3715_/A1 _3715_/A2 _3715_/A3 _3715_/A4 _3715_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_174_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4695_ _4736_/A3 _4467_/B _4736_/A1 _4695_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_6434_ _6434_/A1 _6434_/A2 _6434_/A3 _6434_/A4 _6434_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_162_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3646_ _3646_/A1 _3630_/Z _3646_/A3 _3645_/Z _3646_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_162_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6365_ _6744_/Q _7252_/Q _6365_/B _6366_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_115_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3577_ _3512_/Z _3537_/Z _3947_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_161_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6296_ _7235_/Q _7234_/Q _6484_/A2 _6484_/A3 _6296_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_130_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5316_ _5316_/A1 _5316_/A2 _5315_/Z _4772_/Z _5316_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5247_ _5246_/Z _5442_/A2 _5056_/C _4496_/Z _5247_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold37 hold37/I hold37/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold15 hold15/I hold15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_69_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold26 hold26/I hold26/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5178_ _5180_/A3 _5180_/A2 _5211_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_75_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold59 hold59/I hold59/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold48 hold48/I hold48/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_28_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4129_ _4103_/I hold912/Z _4136_/S _4129_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_263 net613_263/I _6962_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_252 _4073__18/I _6973_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet613_274 net613_285/I _6951_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_296 net613_297/I _6929_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_285 net613_285/I _6940_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3500_ _3500_/I0 _3500_/I1 hold21/Z _3500_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_128_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4480_ _4463_/Z _4468_/Z _4786_/A2 _4786_/A3 _4808_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold518 _7033_/Q hold518/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold507 _5698_/Z _7049_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3431_ _6734_/Q _3434_/B _7299_/Q _3432_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold529 _7202_/Q hold529/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3362_ _7063_/Q _3362_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6150_ _7092_/Q _6002_/Z _6003_/Z _7164_/Q _6152_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5101_ _5303_/A1 _5460_/A1 _5101_/A3 _5303_/A2 _5101_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_83_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3293_ _7301_/Q _3428_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6081_ _7113_/Q _5984_/Z _5997_/Z _7097_/Q _7071_/Q _5980_/Z _6084_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_98_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5032_ _4397_/Z _4411_/Z _5328_/A1 _5387_/A1 _5032_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6983_ _6983_/D _7260_/RN _6983_/CLK _6983_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5934_ _5934_/I _7232_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5865_ hold2/Z hold531/Z _5865_/S _5865_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4816_ _5287_/B _4673_/Z _5132_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_22_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5796_ hold271/Z hold929/Z hold7/Z _7135_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4747_ _4747_/A1 _4747_/A2 _5231_/C _4751_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_162_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4678_ _4997_/C _4673_/Z _4675_/Z _5451_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_150_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3629_ _7124_/Q _3956_/A2 _3927_/B1 _7066_/Q _3630_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6417_ _6554_/A1 _6417_/A2 _6417_/A3 _6417_/A4 _6417_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6348_ _7136_/Q _6253_/Z _6293_/Z _7152_/Q _6348_/C _6356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xinput127 wb_cyc_i _4032_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput116 wb_adr_i[29] _4031_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput105 wb_adr_i[19] _4391_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6279_ _6452_/A4 _6285_/A2 _6279_/A3 _7237_/Q _6279_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_130_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput149 wb_dat_i[29] _6594_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput138 wb_dat_i[19] _6588_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_15__1359_ net413_58/I _4073__7/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_107_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_78__1359_ net613_299/I net413_57/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3980_ _6733_/Q _3972_/Z _6659_/Q _3981_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_63_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_189_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5650_ _7006_/Q hold86/Z _5655_/S _5650_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4601_ _4601_/A1 _4595_/Z _4599_/Z _4600_/Z _4601_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5581_ _6945_/Q hold29/Z hold23/Z hold30/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_184_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4532_ _5420_/A2 _4456_/B _5051_/S _3401_/I _5414_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_7_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7251_ _7251_/D _7258_/RN _7258_/CLK _7251_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_117_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4463_ _4460_/B _4481_/A2 _4463_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
Xhold304 _7187_/Q hold304/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold326 _7171_/Q hold326/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold315 _5764_/Z _7107_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3414_ _6733_/Q _3413_/Z _3442_/B _3988_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_172_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold359 _5723_/Z _7071_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold348 _5552_/Z _6919_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold337 hold337/I hold337/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6202_ _6799_/Q _5958_/Z _5969_/Z _7296_/Q _6726_/Q _5994_/I _6204_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_4394_ _4427_/A3 _4481_/A1 _4922_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7182_ _7182_/D _7193_/RN _7182_/CLK _7182_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3345_ _7193_/Q _3345_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6133_ _6133_/A1 _6133_/A2 _6133_/A3 _6133_/A4 _6133_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_133_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6064_ _6064_/I _6065_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5015_ _5013_/Z _5350_/A2 _5017_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_100_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet813_458 net813_473/I _6707_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6966_ _6966_/D _7238_/RN _6966_/CLK _6966_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xnet813_469 net413_75/I _6696_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5917_ _7228_/Q _7227_/Q _5917_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_41_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6897_ _6897_/D _7238_/RN _6897_/CLK hold88/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_179_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5848_ _3485_/Z _3521_/Z hold6/Z _5856_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_10_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5779_ hold86/Z hold679/Z _5784_/S _5779_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold882 _7214_/Q hold882/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold871 _4224_/Z _6752_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold860 _6790_/Q hold860/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold893 _5759_/Z _7102_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_2__1359_ net713_387/I net763_437/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_160_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6820_ _6820_/D _7210_/RN _6820_/CLK _6820_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_17_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6751_ _6751_/D _7238_/RN _6751_/CLK _6751_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_32_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3963_ _3915_/Z _3919_/Z _3963_/A3 _3962_/Z _6564_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_176_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5702_ hold454/Z hold113/Z _5709_/S _5702_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6682_ _6682_/D _7297_/RN _6682_/CLK _6682_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3894_ _3894_/A1 _3894_/A2 _3894_/A3 _3894_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_5633_ hold52/Z hold252/Z _5637_/S _5633_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5564_ hold15/Z hold282/Z _5565_/S _5564_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4515_ _5002_/A3 _5002_/A4 _5083_/B _4561_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7303_ _7303_/D _6655_/Z _7303_/CLK _7303_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold101 _6671_/Q hold101/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold112 _7270_/Q hold112/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold134 _3476_/I hold134/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5495_ _4103_/I hold255/Z _5496_/S _5495_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold123 _5585_/Z _6948_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7234_ _7234_/D _7237_/RN _7258_/CLK _7234_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_144_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4446_ _4441_/B _5281_/C _4467_/B _4501_/B _5287_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold167 _6765_/Q hold167/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold156 _7019_/Q hold156/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold145 _5734_/Z _7080_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4377_ _3401_/I _3402_/I _4456_/B _5051_/S _5464_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_160_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_61__1359_ clkbuf_4_15_0__1359_/Z net763_416/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold178 _7043_/Q hold178/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7165_ _7165_/D _7221_/RN _7165_/CLK _7165_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold189 _5663_/Z _7018_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xclkbuf_leaf_141__1359_ net563_220/I net713_383/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3328_ _7235_/Q _5943_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_113_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6116_ _6116_/A1 _5991_/Z _6132_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_85_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7096_ _7096_/D _7258_/RN _7096_/CLK _7096_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_58_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6047_ _7144_/Q _5987_/Z _6015_/Z _7006_/Q _6047_/C _6048_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_27_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6949_ _6949_/D _7260_/RN _6949_/CLK _6949_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_168_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold690 _4183_/Z _6722_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__12 _4073__12/I _7213_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_53 net413_53/I _7172_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_64 _4073__7/I _7161_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__23 net413_57/I _7202_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_86 net413_86/I _7139_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet413_75 net413_75/I _7150_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet413_97 net413_97/I _7128_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__45 _4073__45/I _7180_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__34 _4073__47/I _7191_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput217 _6736_/Q mgmt_gpio_out[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput206 _3372_/ZN mgmt_gpio_oeb[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput239 _4047_/Z mgmt_gpio_out[37] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_182_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5280_ _5372_/A1 _5055_/Z _5284_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_142_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput228 _6911_/Q mgmt_gpio_out[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4300_ _6571_/I0 _6808_/Q _4300_/S _6808_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4231_ _4230_/Z hold755/Z _4245_/S _4231_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4162_ hold785/Z _4103_/I _4163_/S _4162_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4093_ _7299_/Q input75/Z _4094_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_82_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4995_ _4892_/B _4716_/Z _5428_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6803_ _6803_/D _7265_/CLK _6803_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6734_ _6734_/D _6625_/Z _7303_/CLK _6734_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_149_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3946_ _6720_/Q _3946_/A2 _4161_/A1 _6708_/Q _6674_/Q _3546_/Z _3949_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_182_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6665_ _6665_/D _6620_/Z _7303_/CLK _6665_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_143_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3877_ _7005_/Q _3934_/A2 _3916_/B1 _6879_/Q _3885_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_180_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6596_ _6596_/I0 _7275_/Q _6602_/S _7275_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5616_ hold62/Z hold73/Z _5619_/S hold74/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5547_ hold2/Z hold161/Z _5547_/S _5547_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5478_ _4614_/Z _4683_/Z _5302_/B _4700_/Z _5230_/B _5479_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_4429_ _5083_/C _4422_/Z _5340_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7217_ _7217_/D _7219_/RN _7217_/CLK _7217_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_7148_ _7148_/D _7221_/RN _7148_/CLK _7148_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_86_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7079_ _7079_/D _7210_/RN _7079_/CLK _7079_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_104_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet463_150 net513_159/I _7075_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4780_ _4716_/Z _4778_/Z _5122_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3800_ _3509_/Z _3680_/Z _3928_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_21_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3731_ input14/Z _3913_/A2 _3758_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_159_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6450_ _7256_/Q _6450_/I1 _6558_/S _7256_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3662_ _7131_/Q _3930_/A2 _3901_/A2 _6985_/Q _3663_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_162_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6381_ _7097_/Q _6250_/Z _6290_/Z _7081_/Q _6302_/Z _7089_/Q _6383_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3593_ _6939_/Q _3910_/A2 _3901_/A2 _6987_/Q _3596_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5401_ _4694_/Z _4703_/Z _5401_/B _5401_/C _5480_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_62_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5332_ _5444_/A2 _5327_/Z _5482_/A1 _5332_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_161_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5263_ _4997_/B _5263_/A2 _4716_/Z _5263_/A4 _5263_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_130_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5194_ _4555_/C _5205_/A1 _5194_/B1 _5346_/A2 _5350_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_7002_ hold20/Z _7238_/RN _7002_/CLK _7002_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4214_ _4213_/Z hold739/Z _4228_/S _4214_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4145_ hold713/Z hold271/Z _4145_/S _4145_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4076_ _7299_/Q input88/Z _4077_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_37_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4978_ _5258_/A2 _4977_/Z _4979_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_177_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3929_ _3926_/Z _3929_/A2 _3929_/A3 _3929_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6717_ _6717_/D input75/Z _6717_/CLK _6717_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6648_ _7237_/RN _6656_/A2 _6648_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_164_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6579_ _6834_/Q _6579_/A2 _6579_/B1 _6835_/Q _6836_/Q _6579_/C2 _6580_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_124_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_312 net663_313/I _6913_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_323 net413_74/I _6902_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_334 net813_491/I _6891_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_345 net713_358/I _6880_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5950_ _5950_/A1 _5950_/A2 _5950_/B1 _6302_/A4 _7237_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_34_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4901_ _4700_/Z _4716_/Z _5442_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_74_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5881_ hold29/Z hold322/Z _5883_/S _5881_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4832_ _5287_/B _4683_/Z _5281_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4763_ _4765_/A1 _5302_/B _5226_/C _5403_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_60_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6502_ _6502_/I _6503_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4694_ _5302_/B _4778_/A4 _4468_/Z _5099_/A2 _4694_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_53_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3714_ hold89/I _5665_/A1 _3923_/C1 hold68/I _3714_/C _3715_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_146_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6433_ _7073_/Q _6248_/Z _6297_/Z _6703_/Q _6433_/C _6434_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_146_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3645_ _3638_/Z _3642_/Z _3645_/A3 _3645_/A4 _3645_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6364_ _6357_/Z _6363_/Z _6364_/B1 _6286_/Z _6555_/C _6365_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3576_ _3521_/Z _3529_/Z _5638_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5315_ _5315_/A1 _5315_/A2 _4683_/Z _5302_/B _5315_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6295_ _6295_/I _6298_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5246_ _5258_/B2 _5343_/A2 _5389_/A2 _5255_/A2 _5246_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_114_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold38 hold38/I hold38/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold16 hold16/I hold16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold27 hold27/I hold27/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5177_ _4414_/Z _4878_/Z _5180_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_68_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold49 hold49/I hold49/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_28_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4128_ _5520_/C _3533_/Z _5513_/A3 _5839_/A3 _4136_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4059_ _6753_/Q input77/Z _4059_/S _4059_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_38__1359_ net413_53/I net613_300/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xnet613_253 net613_253/I _6972_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_118__1359_ net613_293/I net413_90/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_35_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_264 net613_264/I _6961_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet613_286 net663_324/I _6939_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_297 net613_297/I _6928_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_275 net613_281/I _6950_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold508 _7070_/Q hold508/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3430_ _7300_/Q _7283_/Q _3430_/S _7300_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold519 _5680_/Z _7033_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3361_ _7071_/Q _3361_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_171_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5100_ _5100_/A1 _5312_/A2 _5220_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6080_ hold65/I _5972_/Z _6021_/Z _6999_/Q _6085_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_3_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5031_ _5028_/Z _5354_/A1 _5202_/A3 _5035_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_3292_ _7303_/Q _3422_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6982_ _6982_/D _7260_/RN _6982_/CLK _6982_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5933_ _5913_/I _6745_/Q _7232_/Q _5934_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5864_ hold15/Z hold436/Z _5865_/S _5864_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4815_ _5414_/A2 _4764_/Z _5215_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_61_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5795_ hold113/Z hold407/Z hold7/Z _7134_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4746_ _4716_/Z _5230_/B _5231_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_147_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4677_ _4673_/Z _4892_/B _5392_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_107_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3628_ input27/Z _3954_/B1 _3925_/A2 input9/Z _3630_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6416_ hold64/I _6245_/Z _6262_/Z hold72/I _7032_/Q _6269_/Z _6417_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6347_ _7038_/Q _6275_/Z _6300_/Z _7104_/Q _6347_/C _6357_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3559_ _3523_/Z _3537_/Z _3923_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput117 wb_adr_i[2] _5051_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
Xinput106 wb_adr_i[1] _3402_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_131_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6278_ _6276_/Z _6277_/Z _6287_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_88_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput139 wb_dat_i[1] _3394_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput128 wb_dat_i[0] _3393_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_130_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5229_ _5229_/A1 _5479_/A2 _5234_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_69_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4600_ _4524_/Z _5399_/A2 _4546_/Z _5364_/B _4600_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_157_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5580_ hold64/Z hold62/Z hold23/Z _6944_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4531_ _5270_/A1 _4530_/I _5214_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_8_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold316 _7204_/Q hold316/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4462_ _4736_/A1 _4736_/A3 _4778_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold305 _5854_/Z _7187_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7250_ _7250_/D _7260_/RN _7260_/CLK _7250_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3413_ _3412_/Z _3409_/Z _6732_/Q _3413_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_172_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold338 _3493_/Z hold338/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold349 _6680_/Q hold349/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold327 _5836_/Z _7171_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6201_ _6201_/A1 _6201_/A2 _6201_/A3 _6201_/A4 _6201_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4393_ _4385_/Z _4387_/Z _4390_/Z _4489_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7181_ _7181_/D _7221_/RN _7181_/CLK _7181_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_98_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3344_ _6926_/Q _6364_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6132_ hold42/I _5994_/I _6132_/B _6133_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_86_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6063_ _6555_/C _7242_/Q _6063_/B _6064_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5014_ _4555_/C _5439_/A1 _5349_/A1 _5439_/B2 _5350_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _6965_/D _7193_/RN _6965_/CLK _6965_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xnet813_459 net813_473/I _6706_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5916_ _7228_/Q _7227_/Q _6210_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xclkbuf_leaf_21__1359_ net613_253/I _4073__47/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_35_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_101__1359_ clkbuf_4_5_0__1359_/Z net663_326/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6896_ _6896_/D _7260_/RN _6896_/CLK _6896_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_179_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5847_ hold2/Z hold377/Z _5847_/S _5847_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5778_ hold271/Z hold921/Z _5784_/S _5778_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4729_ _4765_/A1 _5302_/B _5099_/A2 _4700_/Z _4729_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_163_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold850 _6739_/Q hold850/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold872 _6823_/Q hold872/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold861 _4279_/Z _6790_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_150_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold883 _5885_/Z _7214_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold894 _7158_/Q hold894/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_130_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6750_ _6750_/D _7238_/RN _6750_/CLK _6750_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_188_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5701_ _5701_/A1 hold18/Z _5709_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_92_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3962_ _3938_/Z _3944_/Z _3949_/Z _3961_/Z _3962_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_44_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6681_ _6681_/D _7297_/RN _6681_/CLK _6681_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3893_ _7151_/Q _3916_/A2 _5536_/A1 _6907_/Q _3894_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_148_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5632_ hold86/Z hold106/Z _5637_/S _5632_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5563_ hold29/Z hold192/Z _5565_/S _5563_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7302_ _7302_/D _6654_/Z _7303_/CLK _7302_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_163_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4514_ _4414_/Z _4421_/Z _4452_/Z _4810_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_145_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold135 _3477_/Z hold135/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold113 _4102_/Z hold113/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold124 _6774_/Q hold124/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5494_ hold38/Z _3515_/Z hold6/Z hold135/Z _5496_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold102 _4114_/Z _6671_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4445_ _4853_/A1 _4501_/B _5309_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7233_ _7233_/D _7237_/RN _7258_/CLK _7233_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_132_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold168 _4249_/Z _6765_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold157 _5664_/Z _7019_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold146 _7154_/Q hold146/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4376_ _3401_/I _3402_/I _4456_/B _5051_/S _4376_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold179 _5691_/Z _7043_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7164_ _7164_/D _7221_/RN _7164_/CLK _7164_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_99_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3327_ _7232_/Q _6279_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_112_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6115_ hold43/I wire348/Z _6211_/B1 _6993_/Q _6116_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_112_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_7095_ _7095_/D _7193_/RN _7095_/CLK _7095_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XTAP_3019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6046_ _7160_/Q _7231_/Q wire348/Z _6117_/A4 _6047_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6948_ _6948_/D _7238_/RN _6948_/CLK _6948_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_179_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6879_ _6879_/D _7297_/RN _6879_/CLK _6879_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_179_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold680 _5779_/Z _7120_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_150_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold691 _6754_/Q hold691/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_103_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_76 net413_76/I _7149_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__13 net413_77/I _7212_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_65 net413_65/I _7160_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_54 net413_62/I _7171_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073__24 _4073__36/I _7201_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__46 net413_61/I _7179_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_98 net413_98/I _7127_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__35 net413_66/I _7190_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet413_87 net413_88/I _7138_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput207 _3371_/ZN mgmt_gpio_oeb[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput218 _6737_/Q mgmt_gpio_out[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_154_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput229 _6912_/Q mgmt_gpio_out[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4230_ hold257/Z _4102_/Z _4244_/S _4230_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4161_ _4161_/A1 hold18/Z _4163_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_49_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4092_ _4092_/I _4092_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6802_ _6802_/D _7243_/CLK _6802_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4994_ _5083_/C _4997_/C _4546_/Z _4422_/Z _4994_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_23_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6733_ _6733_/D _6624_/Z _7303_/CLK _6733_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3945_ _7174_/Q _3945_/A2 _3945_/B1 _7086_/Q _6682_/Q _3945_/C2 _3949_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_189_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6664_ _6664_/D _6619_/Z _7304_/CLK _6664_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_143_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5615_ hold52/Z _6975_/Q _5619_/S hold53/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3876_ _3873_/Z _3876_/A2 _3876_/A3 _3876_/A4 _3876_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6595_ _6595_/A1 _4313_/Z _6595_/B _6596_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_165_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5546_ hold15/Z hold201/Z _5547_/S _5546_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5477_ _5352_/Z _5390_/Z _5437_/Z _5476_/Z _5477_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_145_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4428_ _4427_/Z _4402_/B _4373_/Z _4428_/B2 _5337_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_160_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7216_ _7216_/D _7221_/RN _7216_/CLK _7216_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_160_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_3__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _7303_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7147_ hold46/Z _7238_/RN _7147_/CLK hold45/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_24_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4359_ _4359_/A1 hold18/Z _4361_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_48_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7078_ _7078_/D _7210_/RN _7078_/CLK _7078_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_6029_ _7103_/Q _5967_/Z _5969_/Z _7119_/Q _6030_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_46_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_151 _4073__20/I _7074_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet463_140 net613_263/I _7085_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3730_ _7071_/Q _3943_/A2 _3945_/B1 _7089_/Q _3757_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_1992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3661_ _7057_/Q _5701_/A1 _3925_/A2 input8/Z _3663_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6380_ _6380_/A1 _6380_/A2 _6380_/A3 _6380_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_5400_ _5400_/A1 _5400_/A2 _5399_/Z _4729_/Z _5401_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_86_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3592_ _3592_/A1 _3592_/A2 _3592_/A3 _3592_/A4 _3592_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_9_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5331_ _5331_/I _5482_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5262_ _5340_/A1 _5262_/A2 _5328_/A2 _5442_/A4 _5262_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_142_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7001_ _7001_/D _7238_/RN _7001_/CLK hold41/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5193_ _5193_/A1 _5193_/A2 _5437_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_114_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4213_ hold230/Z _4102_/Z _4227_/S _4213_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4144_ hold666/Z _4103_/I _4145_/S _4144_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4075_ input83/Z _4075_/I1 _7299_/Q _4075_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4977_ _5262_/A2 _5343_/A2 _4495_/Z _4497_/Z _4977_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_149_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6716_ _6716_/D _7193_/RN _6716_/CLK _6716_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_138_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3928_ _6940_/Q _5575_/A1 _3928_/B1 _6789_/Q _3928_/C1 _6822_/Q _3929_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_32_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6647_ _7237_/RN _6657_/A2 _6647_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_149_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3859_ _6933_/Q _3910_/A2 _3959_/B1 _6667_/Q _3925_/A2 input35/Z _3860_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6578_ _6578_/A1 _6578_/A2 _6602_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_165_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5529_ hold18/Z hold665/Z _6901_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_117_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_302 net663_305/I _6923_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet663_324 net663_324/I _6901_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_313 net663_313/I _6912_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_335 net813_495/I _6890_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_346 net713_358/I _6879_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_92_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4900_ _5343_/B _5255_/A2 _4900_/B _5341_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5880_ hold62/Z hold656/Z _5883_/S _5880_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4831_ _5214_/A2 _5420_/A1 _5223_/A2 _5291_/C _5276_/A1 _4840_/B1 _4834_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_61_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4762_ _5420_/A2 _5270_/A1 _4761_/I _3401_/I _4762_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_53_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6501_ _6555_/C _7257_/Q _6501_/B _6502_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4693_ _5099_/A1 _5099_/A2 _5097_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3713_ _3713_/I _3714_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6432_ _6432_/A1 _6239_/Z _6433_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3644_ _7010_/Q _3934_/A2 _3916_/A2 _7156_/Q _3645_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_161_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3575_ _7067_/Q _3927_/B1 _3592_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6363_ _6554_/A1 _6363_/A2 _6363_/A3 _6363_/A4 _6363_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_142_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5314_ _5314_/A1 _5314_/A2 _5314_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_6294_ _7142_/Q _6292_/Z _6293_/Z _7150_/Q _6295_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5245_ _4421_/Z _4510_/Z _4666_/Z _4703_/Z _5245_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_143_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold28 hold28/I hold28/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold17 hold17/I hold17/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_130_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5176_ _5175_/Z _4313_/Z _5184_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_96_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold39 hold39/I hold39/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_110_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4127_ hold2/Z hold262/Z _4127_/S _4127_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4058_ _6755_/Q input67/Z _7302_/Q _4058_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet613_254 net613_258/I _6971_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_265 net413_79/I _6960_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet613_287 net613_287/I _6938_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_298 net613_300/I _6927_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_76_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_276 net613_276/I _6949_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold509 _5722_/Z _7070_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_128_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3360_ _6701_/Q _3360_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5030_ _5471_/B2 _5376_/B2 _5002_/Z _5353_/A1 _5202_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_151_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6981_ _6981_/D _7210_/RN _6981_/CLK _6981_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_20_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5932_ _5932_/I _7231_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_179_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5863_ hold29/Z hold469/Z _5865_/S _5863_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4814_ _5414_/A2 _5287_/B _4876_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5794_ _3507_/Z _3552_/Z _5520_/C hold7/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_166_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _4700_/Z _5230_/B _4747_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4676_ _4675_/Z _4501_/B _4472_/B _4524_/Z _4892_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_179_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3627_ _7002_/Q _5638_/A1 _3959_/B1 hold97/I input32/Z _3927_/C2 _3630_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6415_ _7048_/Q _6241_/Z _6251_/Z _6984_/Q _6268_/Z hold79/I _6417_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_115_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3558_ _3515_/Z _3552_/Z _3916_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6346_ _7096_/Q _6250_/Z _6302_/Z _7088_/Q _6292_/Z _7144_/Q _6357_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_163_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput118 wb_adr_i[30] _4035_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput107 wb_adr_i[20] _4483_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_131_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6277_ _6261_/Z _6265_/Z _6268_/Z _6269_/Z _6277_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xclkbuf_leaf_44__1359_ net463_109/I net413_77/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_103_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3489_ _3489_/I _3653_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
Xclkbuf_leaf_124__1359_ _4073__15/I _4073__14/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput129 wb_dat_i[10] _6585_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5228_ _5287_/C _5302_/B _4784_/Z _5228_/B _5479_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_5159_ _4422_/Z _4568_/Z _4641_/Z _4483_/B _5160_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_99_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4530_ _4530_/I _4860_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold317 _5873_/Z _7204_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold306 _6918_/Q hold306/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4461_ _5281_/C _4481_/A2 _4469_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3412_ _3451_/I0 _7292_/Q _7293_/Q _3412_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_171_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7180_ _7180_/D _7221_/RN _7180_/CLK _7180_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_113_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6200_ _6843_/Q _5971_/Z _5981_/Z _6787_/Q _6005_/Z _6849_/Q _6201_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold328 _7162_/Q hold328/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold339 _3904_/Z hold339/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4392_ _4385_/Z _4387_/Z _4390_/Z _4392_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_113_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6131_ _6703_/Q _5965_/Z _5967_/Z _7107_/Q _7171_/Q _6006_/Z _6133_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_124_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3343_ _7136_/Q _6051_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6062_ _6053_/Z _6061_/Z _6364_/B1 _6168_/C _6555_/C _6063_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _5347_/A1 _5012_/Z _5347_/A4 _5192_/B _5013_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6964_ _6964_/D _7210_/RN _6964_/CLK _6964_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_179_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5915_ _5945_/A1 _6745_/Q _5941_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_81_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6895_ _6895_/D _7260_/RN _6895_/CLK _6895_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_34_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5846_ hold15/Z hold442/Z _5847_/S _5846_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5777_ hold113/Z hold387/Z _5784_/S _5777_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4728_ _4765_/A1 _5302_/B _5099_/A2 _4728_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_162_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4659_ _5281_/C _4436_/B _4472_/B _4501_/B _4659_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_108_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold851 _4205_/Z _6739_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_66_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold840 _6972_/Q hold840/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold873 _4325_/Z _6823_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold862 _6850_/Q hold862/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_107_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6329_ _6329_/A1 _6329_/A2 _6322_/Z _6328_/Z _6329_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold895 _5822_/Z _7158_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold884 _6719_/Q hold884/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_153_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_90__1359_ clkbuf_4_13_0__1359_/Z net763_426/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3961_ _3953_/Z _3958_/Z _3961_/A3 _3961_/A4 _3961_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_189_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5700_ hold2/Z hold142/Z _5700_/S _5700_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_177_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6680_ _6680_/D _7297_/RN _6680_/CLK _6680_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3892_ _7111_/Q _3917_/A2 _3950_/B1 _6725_/Q _3894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_31_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5631_ hold271/Z hold919/Z _5637_/S _5631_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5562_ hold62/Z hold224/Z _5565_/S _5562_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7301_ _7301_/D _6653_/Z _7304_/CLK _7301_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_157_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4513_ _4421_/Z _4506_/Z _5180_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_144_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7232_ _7232_/D _7237_/RN _4067_/I1 _7232_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xhold125 _4259_/Z _6774_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5493_ hold271/Z hold852/Z _5493_/S _5493_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold114 _5666_/Z _7020_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold103 _6966_/Q hold103/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4444_ _5288_/B _4472_/B _4868_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_132_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold158 _7035_/Q hold158/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold136 _5647_/Z _5655_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold147 _5817_/Z _7154_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4375_ _3401_/I _3402_/I _5170_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold169 _6923_/Q hold169/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7163_ _7163_/D _7297_/RN _7163_/CLK _7163_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3326_ _7233_/Q _6282_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_113_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6114_ hold49/I _5958_/Z _5969_/Z hold59/I _6133_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_7094_ _7094_/D _7193_/RN _7094_/CLK _7094_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_140_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6045_ _7088_/Q _6002_/Z _6048_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6947_ hold3/Z _7238_/RN _6947_/CLK _6947_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6878_ _6878_/D _7193_/RN _6878_/CLK _6878_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_167_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5829_ hold2/Z hold381/Z _5829_/S _5829_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold681 _6906_/Q hold681/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold670 _6724_/Q hold670/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold692 _4228_/Z _6754_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_77 net413_77/I _7148_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_66 net413_66/I _7159_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__14 _4073__14/I _7211_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_55 net413_55/I _7170_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__36 _4073__36/I _7189_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_99 net413_99/I _7126_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__47 _4073__47/I _7178_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__25 _4073__41/I _7200_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_88 net413_88/I _7137_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput208 _3370_/ZN mgmt_gpio_oeb[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput219 _6738_/Q mgmt_gpio_out[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_175_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4160_ hold271/Z hold878/Z _4160_/S _4160_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4091_ _7300_/Q input75/Z _4092_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_95_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6801_ _6801_/D _7243_/CLK _6801_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4993_ _4993_/A1 _4988_/Z _4993_/A3 _4999_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_6732_ _6732_/D _6623_/Z _7303_/CLK _6732_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_51_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3944_ _3944_/A1 _3944_/A2 _3944_/A3 _3944_/A4 _3944_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6663_ _6663_/D _6618_/Z _7303_/CLK _6663_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3875_ _7053_/Q _5701_/A1 _4188_/A1 _6727_/Q _3914_/B1 _6877_/Q _3876_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_31_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5614_ hold86/Z hold685/Z _5619_/S _5614_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6594_ _6834_/Q _6594_/A2 _6594_/B1 _6835_/Q _6836_/Q _6594_/C2 _6595_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5545_ hold29/Z hold236/Z _5547_/S _5545_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5476_ _5476_/A1 _5476_/A2 _5475_/Z _5151_/B _5476_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_117_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4427_ _4374_/Z _4427_/A2 _4427_/A3 _4481_/A1 _4427_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7215_ _7215_/D _7219_/RN _7215_/CLK _7215_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_132_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7146_ _7146_/D _7297_/RN _7146_/CLK _7146_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_99_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4358_ hold271/Z hold844/Z _4358_/S _4358_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3309_ hold9/Z hold10/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_4289_ _4289_/A1 hold18/Z _4291_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_7077_ _7077_/D _7297_/RN _7077_/CLK _7077_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6028_ _7151_/Q _5960_/Z _5965_/Z _6699_/Q _6030_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_58_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet463_141 net613_287/I _7084_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_130 net713_361/I _7095_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3660_ hold66/I _3910_/A2 _5575_/A1 _6945_/Q _3663_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_139_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3591_ _7141_/Q _3951_/A2 _3954_/B1 input28/Z _3959_/B1 hold93/I _3592_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_173_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5330_ _4936_/I _5246_/Z _5445_/B2 _5330_/B2 _5330_/C _5331_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_126_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5261_ _5261_/I _5264_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4212_ _4227_/S _4194_/Z _6652_/A2 _3519_/Z hold18/Z _4228_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_7000_ _7000_/D _7260_/RN _7000_/CLK _7000_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_48_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5192_ _5438_/C _4547_/Z _5192_/B _5192_/C _5193_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_110_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4143_ _4143_/A1 hold18/Z _4145_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_83_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4074_ input84/Z input67/Z _7300_/Q _4074_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4976_ _4421_/Z _5263_/A2 _5324_/A1 _5263_/A4 _5337_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_52_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6715_ _6715_/D _7193_/RN _6715_/CLK _6715_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_20_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3927_ _6698_/Q _3927_/A2 _3927_/B1 _7060_/Q input4/Z _3927_/C2 _3929_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6646_ _7237_/RN _6657_/A2 _6646_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3858_ _6699_/Q _3927_/A2 _3902_/A2 _6890_/Q input15/Z _3927_/C2 _3860_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_20_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6577_ _6834_/Q _6607_/A2 _6605_/A2 _6835_/Q _6577_/C _6578_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_118_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3789_ _7006_/Q _3934_/A2 _5528_/S hold88/I _3790_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_30_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5528_ hold664/Z _4102_/Z _5528_/S _5528_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_14_0__1359_ clkbuf_0__1359_/Z net663_324/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_117_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5459_ _5459_/A1 _5098_/B _5098_/C _5458_/Z _5460_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_105_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7129_ _7129_/D _7221_/RN _7129_/CLK _7129_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_115_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_8__1359_ net413_58/I net413_67/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_3_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_314 net663_316/I _6911_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_303 net663_305/I _6922_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_120_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xnet663_325 net663_326/I _6900_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_336 net813_495/I _6889_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_347 net813_471/I _6878_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_92_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4830_ _5287_/B _4586_/Z _4840_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4761_ _4761_/I _5071_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6500_ _6493_/Z _6499_/Z _6500_/B1 _6286_/Z _6555_/C _6501_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4692_ _4735_/A2 _4764_/A3 _4692_/B _4692_/C _5099_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_3712_ hold83/I _3954_/A2 _3954_/B1 input24/Z _3713_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_14_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6431_ _7131_/Q _6484_/A2 _6533_/A3 _7115_/Q _6432_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3643_ _6688_/Q _3945_/C2 _3941_/A2 _7164_/Q _3645_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6362_ _6942_/Q _6245_/Z _6273_/Z _6974_/Q _7120_/Q _6288_/Z _6363_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_155_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5313_ _5313_/A1 _5313_/A2 _5313_/A3 _5312_/Z _5314_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_3574_ _3521_/Z _3537_/Z _3927_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_143_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6293_ _7235_/Q _7234_/Q _6302_/A3 _6484_/A3 _6293_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5244_ _5324_/A1 _5324_/A2 _5324_/C _5250_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_114_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5175_ _5175_/A1 _5380_/C _5175_/A3 _5175_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_111_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold29 hold29/I hold29/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold18 hold22/Z hold18/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_60_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4126_ hold15/Z hold349/Z _4127_/S _4126_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4057_ _6756_/Q _4072_/B2 _7301_/Q _4057_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4959_ _4959_/A1 _4959_/A2 _4957_/Z _4958_/Z _4963_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xclkbuf_leaf_67__1359_ clkbuf_4_15_0__1359_/Z net613_295/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_165_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_147__1359_ net713_387/I net713_358/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_138_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6629_ _7193_/RN _6652_/A2 _6629_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_153_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet613_255 net613_255/I _6970_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet613_266 net613_297/I _6959_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_299 net613_299/I _6926_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_277 net613_285/I _6948_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_288 net613_288/I _6937_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6980_ _6980_/D _7210_/RN _6980_/CLK _6980_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5931_ _5931_/I0 _7231_/Q _5931_/S _5932_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5862_ hold62/Z hold334/Z _5865_/S _5862_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5793_ hold2/Z hold220/Z _5793_/S _5793_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4813_ _4422_/Z _4997_/C _4554_/Z _4483_/B _5167_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_178_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4744_ _5302_/B _4501_/B _4786_/A2 _5099_/A1 _5230_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_30_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4675_ _4424_/B _4026_/B _4026_/C _4402_/B _4675_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_147_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3626_ _7188_/Q _3959_/C1 _3923_/C1 _7084_/Q _3951_/C1 _7148_/Q _3646_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6414_ _7008_/Q _6243_/Z _6273_/Z hold73/I _6414_/C _6417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3557_ _3523_/Z _3529_/Z _5665_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6345_ _6345_/I _6347_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6276_ _6235_/Z _6237_/Z _6243_/Z _6266_/Z _6276_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_1_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput108 wb_adr_i[21] _4402_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_3488_ _3487_/Z _6862_/Q hold21/Z _3489_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_115_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5227_ _5227_/I _5228_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput119 wb_adr_i[31] _4035_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _5293_/A1 _5293_/B _5161_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4109_ hold51/Z _7273_/Q hold21/Z hold52/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_5089_ _4506_/Z _4666_/Z _5341_/C _5265_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_110_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_50__1359_ net463_109/I net413_80/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_31_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold307 _5551_/Z _6918_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4460_ _4454_/Z _4367_/Z _4460_/B _4736_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_116_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4391_ _4391_/A1 _4391_/A2 _4391_/A3 _4391_/A4 _4481_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3411_ _7293_/Q _7292_/Q _4042_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_172_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold318 _7131_/Q hold318/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold329 _5826_/Z _7162_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3342_ _7251_/Q _6310_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6130_ hold66/I _5981_/Z _5984_/Z _7115_/Q _6134_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_140_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6061_ _6057_/Z _6061_/A2 _6061_/A3 _6061_/A4 _6061_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5012_ _5350_/A1 _5192_/C _5009_/Z _4576_/C _5012_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6963_ hold13/Z _7260_/RN _6963_/CLK _6963_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_146_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5914_ _6745_/Q _5913_/I _7227_/Q _7227_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6894_ _6894_/D input75/Z _6894_/CLK _6894_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5845_ hold29/Z hold438/Z _5847_/S _5845_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5776_ _3521_/Z _3552_/Z _5520_/C _5784_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_21_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4727_ _4727_/A1 _5223_/C _4727_/A3 _5090_/A1 _4733_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4658_ _4887_/A1 _5315_/A2 _5172_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xclkbuf_4_2_0__1359_ clkbuf_0__1359_/Z net413_58/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_3609_ _7294_/Q _6732_/Q _3899_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold830 _5554_/Z _6921_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_123_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput90 spimemio_flash_io2_oeb input90/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4589_ _4835_/A2 _4454_/Z _5364_/B _4456_/B _4589_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_104_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold852 _6867_/Q hold852/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold841 _5612_/Z _6972_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold863 _4349_/Z _6850_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6328_ _6328_/A1 _6328_/A2 _6328_/A3 _6328_/A4 _6328_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold896 _6981_/Q hold896/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold874 _6889_/Q hold874/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold885 _4178_/Z _6719_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_153_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6259_ _6259_/A1 _6259_/A2 _6259_/A3 _6259_/A4 _6259_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_153_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_180_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3960_ _7206_/Q _3960_/A2 _3960_/B1 _6718_/Q _3960_/C _3961_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_177_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3891_ _6949_/Q _5584_/A1 _3954_/B1 input21/Z _5575_/A1 _6941_/Q _3894_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_176_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5630_ hold113/Z hold405/Z _5637_/S _5630_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5561_ hold52/Z hold624/Z _5565_/S _5561_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4512_ _4421_/Z _4452_/Z _5043_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5492_ _4103_/I hold777/Z _5493_/S _5492_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7300_ _7300_/D _6652_/Z _4075_/I1 _7300_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_160_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7231_ _7231_/D _7258_/RN _7260_/CLK _7231_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xhold104 _6775_/Q hold104/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold126 _7170_/Q hold126/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold115 _7022_/Q hold115/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4443_ _5288_/B _4380_/Z _4580_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_99_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold148 _6971_/Q hold148/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold159 _5682_/Z _7035_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold137 _5650_/Z _7006_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4374_ _5288_/B _4853_/A1 _4884_/A1 _4374_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_98_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7162_ _7162_/D _7219_/RN _7162_/CLK _7162_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3325_ _6745_/Q _5950_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
X_6113_ _7245_/Q _6113_/I1 _6558_/S _7245_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7093_ _7093_/D _7221_/RN _7093_/CLK _7093_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6044_ _6210_/A2 _7054_/Q _6048_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_58_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ hold24/Z _7238_/RN _6946_/CLK _6946_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6877_ _6877_/D _7193_/RN _6877_/CLK _6877_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_34_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5828_ hold15/Z hold418/Z _5829_/S _5828_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5759_ hold892/Z _4103_/I _5766_/S _5759_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold671 _4186_/Z _6724_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold660 _7046_/Q hold660/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold693 _6762_/Q hold693/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold682 _5537_/Z _6906_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_56 net413_56/I _7169_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_67 net413_67/I _7158_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4073__37 _4073__37/I _7188_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__48 _4073__48/I _7177_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__26 _4073__43/I _7199_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__15 _4073__15/I _7210_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet413_89 net413_89/I _7136_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_78 net413_78/I _7147_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_158_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput209 _4063_/Z mgmt_gpio_out[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_5_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4090_ _4097_/A1 _4686_/B _6827_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_67_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6800_ _6800_/D _7210_/RN _6800_/CLK _6800_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4992_ _5337_/A2 _5130_/B2 _5368_/A1 _5083_/B _5415_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_90_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6731_ _6731_/D _6622_/Z _7304_/CLK _6731_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3943_ _7068_/Q _3943_/A2 _5728_/A1 _7076_/Q _4182_/A1 _6722_/Q _3944_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_32_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6662_ _6662_/D _6617_/Z _7304_/CLK _6662_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_17_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3874_ _6884_/Q _3912_/B1 _3934_/B1 _6846_/Q _6858_/Q _4359_/A1 _3876_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_143_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5613_ hold271/Z hold978/Z _5619_/S _5613_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6593_ _6593_/I0 _7274_/Q _6602_/S _7274_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5544_ hold62/Z hold268/Z _5547_/S _5544_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5475_ _5438_/C _4604_/Z _5475_/A3 _4666_/Z _5475_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_118_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4426_ _4721_/A1 _4721_/A2 _5083_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_144_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7214_ _7214_/D _7219_/RN _7214_/CLK _7214_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_7145_ _7145_/D _7221_/RN _7145_/CLK _7145_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_98_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4357_ _4103_/I hold767/Z _4358_/S _4357_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3308_ hold36/I _5431_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4288_ _6571_/I0 _6798_/Q _4288_/S _6798_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7076_ _7076_/D _7297_/RN _7076_/CLK _7076_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_104_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6027_ _6949_/Q _5958_/Z _5994_/I _7135_/Q _6027_/C _6030_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xnet463_120 _4073__9/I _7105_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_142 net413_78/I _7083_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_131 net713_361/I _7094_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _6929_/D _7258_/RN _6929_/CLK _6929_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold490 _7219_/Q hold490/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_49_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3590_ _7019_/Q _5656_/A1 _3925_/A2 input10/Z _5665_/A1 _7027_/Q _3592_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_170_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5260_ _4700_/Z _4982_/Z _5260_/B _5261_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_141_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4211_ _4210_/Z hold582/Z _4211_/S _4211_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5191_ _4600_/Z _5190_/Z _5191_/A3 _5191_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_96_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4142_ hold271/Z hold848/Z _4142_/S _4142_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4975_ _4975_/A1 _4975_/A2 _4975_/A3 _4979_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_63_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3926_ _3926_/A1 _3926_/A2 _3926_/A3 _3926_/A4 _3926_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6714_ _6714_/D _7193_/RN _6714_/CLK _6714_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_149_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6645_ _7237_/RN _6657_/A2 _6645_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_137_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3857_ _6838_/Q _3923_/B1 _3960_/B1 _6719_/Q _3860_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6576_ _6832_/Q _6608_/I1 _6606_/A2 _6836_/Q _6578_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_164_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3788_ _7104_/Q _5758_/A1 _3947_/A2 _7096_/Q _3941_/B1 _7168_/Q _3790_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5527_ _6900_/Q hold271/Z hold34/Z _5527_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5458_ _4539_/I _4683_/Z _5302_/B _4460_/B _5458_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4409_ _4407_/Z _4390_/Z _4485_/A2 _5385_/A1 _4412_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5389_ _5389_/A1 _5389_/A2 _5389_/B _5389_/C _5390_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_161_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7128_ _7128_/D _7221_/RN _7128_/CLK _7128_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
Xclkbuf_leaf_27__1359_ clkbuf_4_8_0__1359_/Z net763_431/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_87_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_107__1359_ clkbuf_4_5_0__1359_/Z net613_276/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7059_ _7059_/D _7221_/RN _7059_/CLK _7059_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_87_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet663_315 net663_316/I _6910_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_304 net663_304/I _6921_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet663_326 net663_326/I _6899_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_348 net713_358/I _6877_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_337 net813_482/I _6888_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _5324_/A1 _4436_/B _4495_/Z _4759_/Z _4761_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_1791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4691_ _4786_/A2 _4692_/B _4692_/C _4691_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_53_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3711_ _7016_/Q _5656_/A1 _3924_/A2 hold72/I _3927_/A2 hold70/I _3715_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_186_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3642_ _3642_/A1 _3642_/A2 _3642_/A3 _3642_/A4 _3642_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6430_ _7203_/Q _6272_/Z _6275_/Z _7041_/Q _6293_/Z _7155_/Q _6434_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6361_ _7046_/Q _6241_/Z _6251_/Z _6982_/Q _6268_/Z _6950_/Q _6363_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_60_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5312_ _5312_/A1 _5312_/A2 _5376_/B2 _5312_/A4 _5312_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3573_ _3523_/Z _3552_/Z _3951_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6292_ _7235_/Q _7234_/Q _6484_/A3 _6533_/A3 _6292_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5243_ _5243_/A1 _4890_/I _5324_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_142_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5174_ _5392_/B _4893_/Z _4991_/C _5175_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_69_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold19 hold19/I hold19/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_60_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4125_ hold29/Z hold432/Z _4127_/S _4125_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4056_ _6757_/Q input58/Z _7302_/Q _4056_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4958_ _5258_/B2 _5442_/A2 _5248_/A2 _4958_/A4 _4958_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_177_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4889_ _4997_/C _4700_/Z _4890_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_138_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3909_ _7190_/Q _3909_/A2 _3915_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6628_ _7193_/RN _6652_/A2 _6628_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_165_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6559_ _6833_/D _6830_/Q _6826_/Q _6833_/Q _6559_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_134_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet613_256 net613_273/I _6969_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_267 net613_267/I _6958_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_289 net413_79/I _6936_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet613_278 net613_281/I _6947_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_10__1359_ net413_58/I net713_361/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_73__1359_ net613_299/I net613_263/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_38_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5930_ _5924_/Z _6210_/A2 _6201_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_47_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5861_ hold52/Z hold606/Z _5865_/S _5861_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5792_ hold15/Z hold434/Z _5793_/S _5792_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4812_ _4812_/A1 _4812_/A2 _5179_/B _4812_/B _5000_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_159_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4743_ _4743_/A1 _4740_/Z _4741_/Z _5111_/C _4747_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_175_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4674_ _4424_/B _4422_/Z _5172_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_147_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6413_ _6413_/I _6414_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3625_ _3625_/A1 _3625_/A2 _3625_/A3 _3866_/B _3625_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_127_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3556_ _3525_/Z _3529_/Z _5701_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6344_ _7062_/Q _6257_/Z _6299_/Z _7054_/Q _6345_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_142_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6275_ _7235_/Q _7234_/Q _6484_/A2 _6533_/A2 _6275_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_88_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput109 wb_adr_i[22] _4026_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_170_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3487_ _6658_/Q _7305_/Q _6733_/Q _3487_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5226_ _4716_/Z _5310_/A2 _5226_/B _5226_/C _5227_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_29_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5157_ _5157_/A1 _5423_/A1 _5161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5088_ _5340_/C _5417_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4108_ hold86/Z hold385/Z _4118_/S _4108_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4039_ _6730_/Q _3464_/Z _6734_/Q _4040_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_112_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold308 _7115_/Q hold308/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_8_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4390_ _4391_/A1 _4391_/A2 _4391_/A3 _4391_/A4 _4390_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3410_ _6732_/Q _3409_/Z _3991_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_172_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold319 _5791_/Z _7131_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_7_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3341_ _6925_/Q _6336_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _6974_/Q _5964_/Z _5984_/Z _7112_/Q _6061_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5011_ _5389_/C _5011_/A2 _5002_/Z _5194_/B1 _5350_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_79_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6962_ _6962_/D _7258_/RN _6962_/CLK _6962_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_53_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5913_ _5913_/I _5952_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6893_ _6893_/D input75/Z _6893_/CLK _6893_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5844_ hold62/Z hold444/Z _5847_/S _5844_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5775_ hold2/Z hold207/Z _5775_/S _5775_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4726_ _4703_/Z _5222_/A1 _5090_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4657_ _4657_/A1 _4654_/Z _4657_/A3 _4656_/Z _4664_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xinput91 spimemio_flash_io3_do input91/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3608_ _3589_/Z _3596_/Z _3607_/Z _6571_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xhold820 _6612_/Z _7296_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xnet513_200 net563_212/I _7025_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput80 spi_sck input80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_162_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4588_ _4546_/Z _5364_/B _5205_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold831 _6917_/Q hold831/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold853 _5493_/Z _6867_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6327_ _7021_/Q _6235_/Z _6262_/Z _6965_/Q _6327_/C _6328_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold864 _6825_/Q hold864/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold842 _6675_/Q hold842/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3539_ _3509_/Z _3525_/Z _3954_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold875 _5511_/Z _6889_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold897 _5622_/Z _6981_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold886 _7297_/Q hold886/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_130_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6258_ _7206_/Q _6256_/Z _6257_/Z _7060_/Q _6259_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5209_ _5438_/B _4397_/Z _5209_/A3 _4666_/Z _5209_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_76_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6189_ _6690_/Q _5985_/Z _5999_/Z _6847_/Q _6822_/Q _5964_/Z _6193_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_85_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3890_ _7135_/Q _3951_/A2 _3924_/B1 _6821_/Q _3951_/C1 _7143_/Q _3895_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_43_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5560_ hold86/Z hold779/Z _5565_/S _5560_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4511_ _5129_/A3 _5343_/B _4835_/A2 _3402_/I _4511_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_144_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5491_ _3485_/Z _5857_/A2 hold637/Z _5520_/C _5493_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4442_ _4380_/Z _4579_/A2 _4607_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_129_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7230_ _7230_/D _7258_/RN _7230_/CLK _7230_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
Xhold105 _4260_/Z _6775_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold116 _5668_/Z _7022_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold149 _7003_/Q hold149/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold138 _6882_/Q hold138/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold127 _5835_/Z _7170_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4373_ _4501_/B _5288_/C _4369_/Z _4373_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_144_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7161_ _7161_/D _7219_/RN _7161_/CLK _7161_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3324_ _6744_/Q _5957_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_140_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7092_ _7092_/D _7221_/RN _7092_/CLK _7092_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_101_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6112_ _6555_/C _6109_/Z _6112_/A3 _6112_/B _6113_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_86_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ _7022_/Q wire348/Z _6211_/B1 _6990_/Q _6051_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_152_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ hold30/Z _7238_/RN _6945_/CLK _6945_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_42_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6876_ _6876_/D _7193_/RN _6876_/CLK _6876_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_34_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5827_ hold29/Z hold324/Z _5829_/S _5827_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5758_ _5758_/A1 hold18/Z _5766_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_136_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4709_ _5459_/A1 _5098_/B _4705_/Z _4709_/A4 _4709_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_175_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5689_ hold781/Z hold29/Z _5691_/S _5689_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold672 _6710_/Q hold672/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold650 _6716_/Q hold650/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold661 _5695_/Z _7046_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold694 _4245_/Z _6762_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_103_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold683 _6851_/Q hold683/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_68 net413_68/I _7157_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_57 net413_57/I _7168_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2888 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__16 net413_72/I _7209_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__27 _4073__43/I _7198_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__38 net413_73/I _7187_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_79 net413_79/I _7146_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__49 net413_65/I _7176_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6730_ _6730_/D _6621_/Z _7303_/CLK _6730_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4991_ _5340_/A1 _5370_/B _4991_/B _4991_/C _4993_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_90_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3942_ _3907_/Z _3942_/A2 _7036_/Q _5683_/A1 _3942_/C1 _6853_/Q _3944_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6661_ _6661_/D _6616_/Z _7303_/CLK _6661_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_176_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3873_ _3873_/A1 _3873_/A2 _3873_/A3 _3873_/A4 _3873_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6592_ _6592_/A1 _4313_/Z _6592_/B _6593_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_176_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5612_ hold113/Z hold840/Z _5619_/S _5612_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5543_ hold52/Z hold596/Z _5547_/S _5543_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5474_ hold10/I _5299_/C _5466_/Z _5473_/Z _5474_/C _6864_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_4425_ _4483_/B _4373_/Z _4485_/A2 _4390_/Z _4721_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_133_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7213_ _7213_/D _7221_/RN _7213_/CLK _7213_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_117_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4356_ _3485_/Z hold630/Z _5520_/C _4358_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_7144_ _7144_/D _7258_/RN _7144_/CLK _7144_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_141_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3307_ _3307_/I hold337/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7075_ _7075_/D _7237_/RN _7075_/CLK _7075_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_140_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4287_ _6570_/I0 _6797_/Q _4288_/S _6797_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6026_ _6026_/A1 _6026_/A2 _6026_/A3 _6026_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_55_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet463_110 net513_152/I _7115_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet463_132 net413_61/I _7093_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet463_121 net613_267/I _7104_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_143 net413_89/I _7082_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6928_ _6928_/D _7258_/RN _6928_/CLK _6928_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_42_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6859_ _6859_/D _7279_/RN _7230_/CLK _6859_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold480 _5688_/Z _7040_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold491 _5890_/Z _7219_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4210_ hold95/Z hold2/Z _4210_/S _4210_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5190_ _5464_/A1 _5190_/A2 _5438_/C _5435_/A2 _5190_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_69_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4141_ _4103_/I hold789/Z _4142_/S _4141_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4072_ hold21/I _4072_/A2 _4072_/B1 _4072_/B2 _4072_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_68_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4974_ _5359_/A1 _4973_/Z _4975_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_52_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3925_ input34/Z _3925_/A2 _3925_/B1 _6824_/Q _6839_/Q _3925_/C2 _3926_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6713_ _6713_/D _7297_/RN _6713_/CLK _6713_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6644_ _7237_/RN _6656_/A2 _6644_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_149_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3856_ _7013_/Q _5656_/A1 _5638_/A1 _6997_/Q _5665_/A1 _7021_/Q _3860_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6575_ _6575_/A1 _6575_/A2 _6606_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3787_ _7192_/Q _3909_/A2 _4210_/S input45/Z _4227_/S input58/Z _3795_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_118_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5526_ _6899_/Q hold15/Z hold34/I hold16/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5457_ _5457_/A1 _5457_/A2 _5316_/Z _5457_/A4 _5457_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4408_ _4719_/A2 _4489_/A1 _4428_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5388_ _5388_/A1 _5202_/Z _5354_/Z _5388_/A4 _5388_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_160_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7127_ _7127_/D _7219_/RN _7127_/CLK _7127_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_59_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4339_ _4103_/I hold658/Z _4340_/S _4339_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7058_ _7058_/D _7258_/RN _7058_/CLK _7058_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_86_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6009_ _6009_/A1 _6009_/A2 _6009_/A3 _6008_/Z _6010_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_189_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_305 net663_305/I _6920_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet663_316 net663_316/I _6909_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet663_338 net663_341/I _6887_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_349 net713_358/I _6876_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet663_327 net763_425/I _6898_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3710_ hold73/I _3923_/A2 _3910_/A2 _6936_/Q _3956_/A2 _7122_/Q _3715_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_174_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4690_ _4736_/A1 _4736_/A3 _4690_/B _4690_/C _5099_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_53_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_33__1359_ clkbuf_4_8_0__1359_/Z _4073__48/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3641_ _6704_/Q _3927_/A2 _3924_/A2 _6970_/Q _3642_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3572_ _3529_/Z _3542_/Z _3952_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6360_ _6966_/Q _6262_/Z _6269_/Z _7030_/Q _6360_/C _6363_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xclkbuf_leaf_113__1359_ clkbuf_4_5_0__1359_/Z net413_86/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_96__1359_ clkbuf_4_5_0__1359_/Z net613_264/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_143_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5311_ _5308_/Z _5479_/A3 _5318_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_53_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6291_ _7190_/Q _6285_/Z _6290_/Z _7078_/Q _6307_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_130_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5242_ _4812_/B _5242_/A2 _5242_/A3 _4810_/B _5242_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_102_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5173_ _4424_/B _4422_/Z _5269_/A2 _4997_/C _5173_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_142_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4124_ hold62/Z hold131/Z _4127_/S _4124_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 debug_mode input1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4055_ _6766_/Q input81/Z _4055_/S _4055_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4957_ _5389_/A2 _5442_/A2 _5248_/A2 _4958_/A4 _4957_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_61_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4888_ _5263_/A2 _4700_/Z _5445_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3908_ _5821_/A3 _3533_/Z hold637/I _3942_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_165_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3839_ _3485_/Z _3680_/Z _3922_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6627_ _7193_/RN _6652_/A2 _6627_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_6558_ _7260_/Q _6558_/I1 _6558_/S _7260_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6489_ _6489_/I _6490_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5509_ hold280/Z hold29/Z _5509_/S _5509_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet613_268 net413_98/I _6957_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_76_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet613_279 net613_281/I _6946_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet613_257 net413_89/I _6968_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5860_ hold86/Z hold705/Z _5865_/S _5860_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4811_ _5094_/C _5312_/A2 _5137_/B1 _5220_/B2 _5179_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_22_806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5791_ hold29/Z hold318/Z _5793_/S _5791_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4742_ _5302_/B _4695_/Z _4703_/Z _5226_/C _5111_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_174_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4673_ _5420_/A3 _5129_/A3 _5051_/S _3402_/I _4673_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_119_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3624_ _7058_/Q _5701_/A1 _5674_/A1 _7034_/Q _3952_/A2 _7050_/Q _3625_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6412_ hold89/I _6235_/Z _6265_/Z _7000_/Q _6288_/Z _7122_/Q _6413_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_179_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3555_ _3507_/Z _3552_/Z _3951_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6343_ _7080_/Q _6290_/Z _6357_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3486_ _7305_/Q _6733_/Q _3987_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_131_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6274_ _7234_/Q _6282_/A1 _6302_/A3 _5943_/S _6274_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_0_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5225_ _4728_/Z _5310_/A2 _5225_/B _5310_/C _5229_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_5156_ _5356_/A1 _5403_/B2 _5156_/B _5423_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_97_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4107_ hold85/Z _7272_/Q hold21/Z hold86/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_5087_ _5087_/A1 _4982_/Z _5340_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4038_ _4038_/A1 _6561_/B2 _6826_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_99_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5989_ _7142_/Q _5987_/Z _5988_/Z _6980_/Q _6009_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_178_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput190 _3352_/ZN mgmt_gpio_oeb[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_opt_2_0__1359_ clkbuf_4_8_0__1359_/Z clkbuf_opt_2_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold309 _5773_/Z _7115_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _4421_/Z _5438_/C _5435_/A2 _4606_/Z _5192_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6961_ _6961_/D _7260_/RN _6961_/CLK hold58/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_47_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5912_ _6743_/Q _6745_/Q _5913_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6892_ _6892_/D _7297_/RN _6892_/CLK _6892_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_35_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5843_ hold52/Z hold543/Z _5847_/S _5843_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5774_ hold15/Z hold724/Z _5775_/S _5774_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_652 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4725_ _4510_/Z _5325_/B _4727_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4656_ _5420_/A3 _4374_/Z _5165_/A4 _5209_/A3 _4656_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_147_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4587_ _4454_/Z _5269_/A2 _5364_/B _4586_/Z _4587_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_135_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3607_ _3601_/Z _3607_/A2 _3606_/Z _3607_/A4 _3607_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xinput70 mgmt_gpio_in[7] input70/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xnet513_201 net413_78/I _7024_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold821 _7076_/Q hold821/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold810 _4147_/Z _6696_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput81 spi_sdo input81/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold832 _5550_/Z _6917_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold854 _6909_/Q hold854/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput92 spimemio_flash_io3_oeb input92/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3538_ _3505_/Z _3537_/Z _3943_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6326_ _7079_/Q _6290_/Z _6302_/Z _7087_/Q _6326_/C _6328_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold843 _4121_/Z _6675_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_66_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold898 _7190_/Q hold898/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold865 _4328_/Z _6825_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold876 _6800_/Q hold876/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold887 _6613_/Z _7297_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3469_ _3991_/A1 _3469_/A2 _7280_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6257_ _6484_/A3 _6282_/A2 _7232_/Q _6452_/A4 _6257_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5208_ _5206_/Z _4662_/B _5433_/A1 _5208_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_88_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6188_ _6857_/Q _5924_/Z _6201_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5139_ _4376_/Z _5139_/A2 _5139_/A3 _5291_/C _5139_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_72_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5490_ _5490_/A1 _5299_/C _5466_/Z _5489_/Z _5490_/C _6865_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_4510_ _5420_/A2 _4456_/B _5051_/S _3401_/I _4510_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_8_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4441_ _5420_/A3 _5315_/A1 _4884_/A1 _4441_/B _4579_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_145_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold106 _6990_/Q hold106/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold117 _7136_/Q hold117/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_176_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7160_ _7160_/D _7210_/RN _7160_/CLK _7160_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xhold139 _5502_/Z _6882_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold128 _6942_/Q hold128/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4372_ _4853_/A1 _4884_/A1 _4759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6111_ _6555_/C _7244_/Q _6112_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3323_ _6832_/Q _4096_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7091_ _7091_/D _7297_/RN _7091_/CLK _7091_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6042_ _7168_/Q _6006_/Z _6053_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6944_ _6944_/D _7238_/RN _6944_/CLK hold64/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6875_ _6875_/D _6633_/Z _4075_/I1 _6875_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_179_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5826_ hold62/Z hold328/Z _5829_/S _5826_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5757_ hold2/Z hold391/Z _5757_/S _5757_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4708_ _4708_/A1 _5312_/A2 _5312_/A1 _5094_/C _4709_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5688_ hold479/Z hold62/Z _5691_/S _5688_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4639_ _4639_/A1 _5039_/A4 _4638_/Z _4644_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_135_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold662 _7112_/Q hold662/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold640 _6841_/Q hold640/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold651 _4174_/Z _6716_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7289_ _7289_/D _6643_/Z _7304_/CLK hold14/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6309_ _6554_/A1 _6924_/Q _6310_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_104_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold673 _4165_/Z _6710_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold684 _4351_/Z _6851_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold695 _6980_/Q hold695/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_134_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet413_58 net413_58/I _7167_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2867 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__28 _4073__36/I _7197_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__17 _4073__21/I _7208_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet413_69 net413_77/I _7156_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__39 _4073__39/I _7186_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4990_ _4551_/Z _4892_/B _4991_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_64_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3941_ _7158_/Q _3941_/A2 _3941_/B1 _7166_/Q _3941_/C _3944_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6660_ _6660_/D _6615_/Z _7304_/CLK _6660_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_177_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3872_ _6675_/Q _3546_/Z _3945_/C2 _6683_/Q _3873_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6591_ _6834_/Q _6591_/A2 _6591_/B1 _6835_/Q _6836_/Q _6591_/C2 _6592_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_177_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5611_ _3509_/Z _5520_/C _5821_/A3 _5857_/A3 _5619_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_32_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5542_ hold86/Z hold602/Z _5547_/S _5542_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5473_ _5469_/Z _5489_/A2 _5472_/Z _5473_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_117_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4424_ _4374_/Z _4489_/A1 _4424_/B _4721_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_144_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7212_ _7212_/D _7221_/RN _7212_/CLK _7212_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_99_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4355_ hold271/Z hold723/Z _4355_/S _6854_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7143_ _7143_/D _7210_/RN _7143_/CLK _7143_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_7074_ _7074_/D _7221_/RN _7074_/CLK _7074_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3306_ _6860_/Q _5185_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4286_ _6569_/I0 _6796_/Q _4288_/S _6796_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6025_ _7053_/Q _5924_/Z _6002_/Z _7087_/Q _6168_/C _6026_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_2108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet463_133 net463_133/I _7092_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_111 net413_99/I _7114_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_122 net813_472/I _7103_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet463_144 _4073__30/I _7081_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6927_ _6927_/D _7219_/RN _6927_/CLK _6927_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_120_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6858_ _6858_/D _7193_/RN _6858_/CLK _6858_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_168_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5809_ hold29/Z hold45/Z _5811_/S hold46/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6789_ _6789_/D _7210_/RN _6789_/CLK _6789_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_148_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold470 _5863_/Z _7195_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold481 _7096_/Q hold481/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_8_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold492 _6676_/Q hold492/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4140_ _3485_/Z _5857_/A2 _5513_/A3 _5520_/C _4142_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_68_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4071_ _3994_/Z hold21/I _4072_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_110_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_56__1359_ net663_324/I net513_152/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_136__1359_ net563_220/I net813_489/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_52_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4973_ _5324_/A1 _5263_/A4 _4718_/B _5072_/A4 _4973_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_36_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6712_ _6712_/D _7297_/RN _6712_/CLK _6712_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3924_ _6964_/Q _3924_/A2 _3924_/B1 _6820_/Q _3926_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6643_ _7221_/RN _6656_/A2 _6643_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_60_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3855_ _3855_/A1 _3855_/A2 _3855_/A3 _3855_/A4 _3855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6574_ _6575_/A2 _6574_/A2 _6605_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3786_ _3786_/A1 _3786_/A2 _3786_/A3 _3786_/A4 _3786_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_145_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5525_ _6898_/Q hold29/Z hold34/Z hold35/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5456_ _5456_/A1 _5456_/A2 _5456_/B _5457_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_4407_ _4402_/B _4483_/B _4407_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_172_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5387_ _5387_/A1 _5387_/A2 _5387_/B _5388_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_132_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7126_ _7126_/D _7219_/RN _7126_/CLK _7126_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4338_ _3529_/Z _5520_/C hold637/Z _5857_/A2 _4340_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_75_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7057_ _7057_/D _7260_/RN _7057_/CLK _7057_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4269_ hold99/Z hold15/Z _4270_/S _4269_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6008_ _6008_/A1 _6008_/A2 _6008_/A3 _6008_/A4 _6008_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_46_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet663_306 net763_416/I _6919_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_120_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet663_317 net763_409/I _6908_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_339 net663_341/I _6886_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_328 net763_424/I _6897_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3640_ _6962_/Q _3957_/A2 _3901_/A2 _6986_/Q _3642_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_128_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3571_ _3542_/Z _3552_/Z _3941_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_155_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6290_ _6484_/A3 _5943_/S _7234_/Q _6533_/A3 _6290_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5310_ _4728_/Z _5310_/A2 _5310_/B _5310_/C _5479_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_127_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5241_ _5321_/A1 _5241_/A2 _5451_/B _5242_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_69_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5172_ _5172_/A1 _5368_/A1 _5172_/B _5172_/C _5380_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_114_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4123_ hold52/Z hold483/Z _4127_/S _4123_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4054_ _6764_/Q input78/Z _4055_/S _4054_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput2 debug_oeb input2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4956_ _5359_/A1 _4761_/I _4959_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_80_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ _4887_/A1 _5315_/A2 _4554_/Z _4675_/Z _4887_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3907_ _7300_/Q _7283_/Q _6893_/Q _3907_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_20_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3838_ _3485_/Z _3617_/Z _3920_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6626_ _7193_/RN _6652_/A2 _6626_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_153_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6557_ _6557_/I _6558_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3769_ _7038_/Q _5683_/A1 _5674_/A1 _7030_/Q _3912_/B1 _6885_/Q _3773_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5508_ hold498/Z hold62/Z _5509_/S _5508_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6488_ _7149_/Q _6292_/Z _6300_/Z _7109_/Q _6489_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_10_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _5439_/A1 _5468_/A1 _5439_/B1 _5439_/B2 _5439_/C _5440_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_121_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7109_ _7109_/D _7221_/RN _7109_/CLK _7109_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_101_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet613_258 net613_258/I _6967_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet613_269 net413_79/I _6956_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4810_ _4997_/C _4675_/Z _4683_/Z _4810_/B _4812_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_22_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5790_ hold62/Z hold488/Z _5793_/S _5790_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4741_ _4510_/Z _5302_/B _4695_/Z _5226_/C _4741_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_1590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4672_ _5269_/A2 _4530_/I _5291_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_174_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3623_ _7108_/Q _5758_/A1 _5683_/A1 _7042_/Q _6930_/Q _3935_/A2 _3625_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6411_ _6401_/Z _6408_/Z _6411_/A3 _6411_/A4 _6411_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_179_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6342_ _7070_/Q _6484_/A2 _6484_/A3 _6452_/A4 _6348_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3554_ _3505_/Z _3552_/Z _3930_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_170_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6273_ _6484_/A2 _5943_/S _7234_/Q _6533_/A2 _6273_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3485_ _3473_/Z hold11/Z hold37/Z _3484_/Z _3485_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_115_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5224_ _5224_/A1 _5224_/A2 _5401_/B _5400_/A2 _5225_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_97_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5155_ _5275_/B _5153_/Z _5157_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_57_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5086_ _5086_/A1 _5412_/A1 _5412_/A2 _5260_/B _5182_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_96_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4106_ hold271/Z hold925/Z _4118_/S _4106_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_186_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4037_ _4036_/I _6826_/Q _6561_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_37_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5988_ _7228_/Q _7227_/Q _6002_/A2 _6210_/A2 _5988_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XPHY_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4939_ _4939_/A1 _5061_/B _4937_/Z _4938_/Z _4939_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_36_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6609_ _6608_/Z _6833_/Q _6830_/Q _4313_/Z _6610_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_123_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput180 _3361_/ZN mgmt_gpio_oeb[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput191 _3351_/ZN mgmt_gpio_oeb[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_121_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6960_ _6960_/D _7297_/RN _6960_/CLK _6960_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_26_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5911_ _5911_/A1 _5901_/B _5911_/B _7226_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_98_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6891_ _6891_/D input75/Z _6891_/CLK _6891_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_179_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5842_ hold86/Z hold642/Z _5847_/S _5842_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5773_ hold29/Z hold308/Z _5775_/S _5773_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4724_ _5442_/A2 _4500_/Z _5072_/A4 _5248_/A2 _5325_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_166_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4655_ _5043_/A2 _5043_/B _4657_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_163_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput60 mgmt_gpio_in[31] input60/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4586_ _5288_/B _5281_/C _4436_/B _4472_/B _4586_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xinput71 mgmt_gpio_in[8] input71/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3606_ _3606_/A1 _3606_/A2 _3606_/A3 _3606_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xhold800 _4278_/Z _6789_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold811 _6718_/Q hold811/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput82 spi_sdoenb input82/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold855 _5541_/Z _6909_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold833 _6760_/Q hold833/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3537_ _3477_/Z hold37/Z _3484_/Z _3473_/Z _3537_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_104_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold844 _6856_/Q hold844/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6325_ _6325_/I _6326_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput93 trap _3339_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xhold822 _5729_/Z _7076_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold866 _6786_/Q hold866/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold877 _4291_/Z _6800_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold888 _7077_/Q hold888/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3468_ _7295_/Q hold4/Z _3469_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6256_ _6282_/A1 _5943_/S _7234_/Q _6533_/A3 _6256_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_103_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold899 _5858_/Z _7190_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3399_ _3399_/I _6598_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5207_ _4662_/B _5433_/A1 _5362_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_85_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6187_ _6187_/A1 _5991_/Z _6192_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5138_ _5138_/A1 _5287_/B _5148_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_85_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5069_ _4761_/I _5078_/A2 _5070_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_26_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4440_ _4436_/B _4648_/A1 _4472_/B _4604_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_157_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold107 _5632_/Z _6990_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold118 _6766_/Q hold118/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold129 _7012_/Q hold129/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4371_ _3402_/I _4456_/B _5051_/S _4460_/B _4497_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_171_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6110_ _6201_/A3 _6928_/Q _6112_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3322_ _6746_/Q _4005_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_140_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7090_ _7090_/D _7297_/RN _7090_/CLK _7090_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6041_ _7242_/Q _6041_/I1 _6558_/S _7242_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6943_ _6943_/D _7238_/RN _6943_/CLK hold65/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6874_ _6874_/D _6632_/Z _4075_/I1 _6874_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_34_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5825_ hold52/Z hold276/Z _5829_/S _5825_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5756_ hold15/Z hold456/Z _5757_/S _5756_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5687_ hold525/Z hold52/Z _5691_/S _5687_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4707_ _5420_/A3 _5269_/A2 _4708_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4638_ _4436_/B _4638_/A2 _5356_/C _5356_/A1 _4638_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold630 _3560_/Z hold630/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4569_ _5364_/B _4568_/Z _5356_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold663 _5770_/Z _7112_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap360 _7297_/RN _7210_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold641 _4336_/Z _6841_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold652 _6690_/Q hold652/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7288_ _7288_/D _6642_/Z _7304_/CLK hold28/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_103_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold674 _6998_/Q hold674/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6308_ _6554_/A1 _6307_/Z _6271_/Z _6308_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xhold685 _6974_/Q hold685/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold696 _5621_/Z _6980_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_134_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6239_ _5943_/S _6285_/A2 _7237_/Q _7234_/Q _6239_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_103_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2802 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet413_59 net413_67/I _7166_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__29 net413_80/I _7196_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4073__18 _4073__18/I _7207_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3940_ _3940_/I _3941_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_182_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3871_ _6697_/Q _4146_/A1 _3936_/B1 _6691_/Q _3873_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6590_ _6590_/I0 _7273_/Q _6602_/S _7273_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5610_ hold2/Z hold148/Z hold39/Z _6971_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5541_ hold271/Z hold854/Z _5547_/S _5541_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_16__1359_ net413_58/I net413_66/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_8_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5472_ _5472_/A1 _5472_/A2 _4841_/B _5472_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xclkbuf_leaf_79__1359_ net613_299/I _4073__41/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7211_ _7211_/D _7297_/RN _7211_/CLK _7211_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4423_ _4373_/Z _4385_/Z _4922_/A3 _4423_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_172_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7142_ _7142_/D _7210_/RN _7142_/CLK _7142_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4354_ _4103_/I _6853_/Q _4355_/S _4354_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7073_ _7073_/D _7237_/RN _7073_/CLK _7073_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3305_ _3305_/I _3500_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4285_ _6568_/I0 _6795_/Q _4288_/S _6795_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6024_ _6981_/Q _5988_/Z _6015_/Z _7005_/Q _6024_/C _6026_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_100_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet463_112 _4073__36/I _7113_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_123 net813_472/I _7102_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_134 net813_465/I _7091_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet463_145 net613_288/I _7080_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6926_ _6926_/D _7258_/RN _6926_/CLK _6926_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6857_ _6857_/D _7193_/RN _6857_/CLK _6857_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5808_ hold62/Z hold211/Z _5811_/S _5808_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6788_ _6788_/D _7193_/RN _6788_/CLK _6788_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_183_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5739_ hold2/Z hold395/Z _5739_/S _5739_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold460 _7203_/Q hold460/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold471 _6685_/Q hold471/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold482 _5752_/Z _7096_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold493 _4122_/Z _6676_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_2_2__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _7304_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_181_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4070_ _7240_/Q _6896_/Q _6900_/Q _4070_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_3__1359_ net713_387/I net763_448/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4972_ _4496_/Z _5262_/A2 _5323_/B _4495_/Z _4972_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_17_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6711_ _6711_/D input75/Z _6711_/CLK _6711_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3923_ _6972_/Q _3923_/A2 _3923_/B1 _6837_/Q _3923_/C1 _7078_/Q _3926_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_189_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6642_ _7221_/RN _6656_/A2 _6642_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3854_ _7191_/Q _3909_/A2 _4210_/S input44/Z _3854_/C _3855_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_60_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6573_ _6575_/A2 _6573_/A2 _6607_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3785_ _6934_/Q _3910_/A2 _3959_/C1 _7184_/Q _3785_/C _3786_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_173_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5524_ hold88/Z hold86/Z hold34/Z _6897_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5455_ _5455_/I _5485_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_106_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4406_ _4402_/B _4483_/B _4719_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_172_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5386_ _5386_/A1 _5432_/A1 _5386_/A3 _5434_/A1 _5386_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_7125_ _7125_/D _7258_/RN _7125_/CLK _7125_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_114_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4337_ hold271/Z hold719/Z _4337_/S _4337_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4268_ hold533/Z hold29/Z _4270_/S _4268_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7056_ _7056_/D _7210_/RN _7056_/CLK _7056_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6007_ _7036_/Q _6005_/Z _6006_/Z _7166_/Q _6008_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_39_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4199_ _4198_/Z hold856/Z _4211_/S _4199_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6909_ _6909_/D _7193_/RN _6909_/CLK _6909_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_62__1359_ clkbuf_4_15_0__1359_/Z net763_418/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_142__1359_ net563_220/I _4073__3/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_151_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold290 _7073_/Q hold290/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_78_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet663_307 net763_419/I _6918_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_318 net813_471/I _6907_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet663_329 net663_329/I _6896_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3570_ _3521_/Z _3552_/Z _3956_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_161_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5240_ _5368_/A1 _5389_/A2 _5240_/B _5451_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_142_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5171_ _5169_/Z _5170_/Z _5175_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_39_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4122_ hold86/Z hold492/Z _4127_/S _4122_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4053_ _6763_/Q input80/Z _4055_/S _4053_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput3 debug_out input3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_65_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4955_ _4419_/Z _4951_/Z _4955_/B _5068_/B _4959_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_80_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3906_ _3485_/Z _3578_/Z _3920_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4886_ _4880_/Z _4886_/A2 _4884_/Z _4885_/Z _4886_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_32_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6625_ _7237_/RN _6657_/A2 _6625_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_165_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3837_ input47/Z _4227_/S _3855_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3768_ _3527_/Z _3540_/Z _5532_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6556_ _6555_/C _7259_/Q _6556_/B _6557_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_173_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5507_ hold351/Z hold52/Z _5509_/S _5507_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6487_ _7101_/Q _6250_/Z _6299_/Z _7059_/Q _6995_/Q _6237_/Z _6492_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3699_ _6887_/Q _3912_/B1 _3916_/B1 _6882_/Q _3701_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xclkbuf_4_5_0__1359_ clkbuf_0__1359_/Z clkbuf_4_5_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_5438_ _4568_/Z _4666_/Z _5438_/B _5438_/C _5439_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_161_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput340 _6818_/Q wb_dat_o[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_126_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5369_ _5287_/B _5369_/A2 _5369_/B _5369_/C _5421_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_114_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7108_ _7108_/D _7221_/RN _7108_/CLK _7108_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_59_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7039_ _7039_/D _7221_/RN _7039_/CLK _7039_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_87_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet613_259 net663_326/I _6966_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4740_ _5302_/B _4695_/Z _4716_/Z _5226_/C _4740_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_1591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4671_ _4530_/I _5051_/S _5137_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_186_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3622_ _7180_/Q _3945_/A2 _3913_/A2 input18/Z _3941_/B1 _7172_/Q _3647_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6410_ _7146_/Q _6292_/Z _6300_/Z _7106_/Q hold68/I _6290_/Z _6411_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_174_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6341_ _6934_/Q _6263_/Z _6266_/Z _7014_/Q _6355_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_155_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3553_ _3525_/Z _3552_/Z _3945_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3484_ _4317_/A1 _3483_/Z _3484_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_143_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6272_ _6300_/A2 _6285_/A2 _7237_/Q _6452_/A4 _6272_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5223_ _5094_/B _5223_/A2 _5223_/B _5223_/C _5400_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_5154_ _4568_/Z _4624_/Z _5376_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_116_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4105_ hold270/Z hold273/Z hold21/Z _4105_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_97_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5085_ _4987_/Z _5085_/A2 _5260_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4036_ _4036_/I _4045_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5987_ _7231_/Q _7230_/Q _7229_/Q _6210_/B _5987_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XPHY_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4938_ _4998_/A2 _5389_/A2 _5056_/C _5442_/A2 _4938_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_178_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4869_ _4869_/A1 _4866_/Z _4867_/Z _4868_/Z _4872_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6608_ _6608_/I0 _6608_/I1 _6832_/Q _6608_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6539_ _6729_/Q _6247_/Z _6297_/Z _7077_/Q _6547_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_133_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput170 _4089_/Z irq[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput181 _3360_/ZN mgmt_gpio_oeb[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput192 _3350_/ZN mgmt_gpio_oeb[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5910_ _6746_/Q _4006_/Z _5910_/B _5910_/C _5911_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_35_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6890_ _6890_/D _7297_/RN _6890_/CLK _6890_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_5841_ hold271/Z hold970/Z _5847_/S _5841_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5772_ hold62/Z hold567/Z _5775_/S _5772_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4723_ _4495_/Z _4436_/B _5248_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_147_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4654_ _4467_/B _5315_/A2 _4589_/Z _4460_/B _4654_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_135_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput61 mgmt_gpio_in[32] input61/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4585_ _4887_/A1 _5399_/A2 _5276_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xinput50 mgmt_gpio_in[22] input50/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput72 mgmt_gpio_in[9] input72/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3605_ _7085_/Q _3923_/C1 _3956_/A2 _7125_/Q _3606_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold801 _6824_/Q hold801/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold812 _4177_/Z _6718_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold834 _4241_/Z _6760_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_115_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput83 spimemio_flash_clk input83/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold845 _4358_/Z _6856_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_66_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6324_ _7143_/Q _6292_/Z _6300_/Z _7103_/Q _6325_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3536_ _3533_/Z _3535_/Z _3927_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold823 _6799_/Q hold823/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput94 uart_enabled _4059_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold856 _6736_/Q hold856/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_143_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold867 _4273_/Z _6786_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold878 _6707_/Q hold878/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6255_ _7134_/Q _6253_/Z _6254_/Z _7174_/Q _6259_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold889 _5730_/Z _7077_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3467_ _3467_/I _7282_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5206_ _5189_/Z _5203_/Z _5357_/A2 _5440_/A1 _5206_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3398_ _3398_/I _6595_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6186_ _6845_/Q wire348/Z _6211_/B1 _6837_/Q _6187_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5137_ _5276_/C _5137_/A2 _5137_/B1 _5279_/A2 _5370_/B _5138_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_96_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5068_ _4700_/Z _4761_/I _5068_/B _5334_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_42_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4019_ _4006_/Z _4019_/A2 _4014_/Z _4019_/B _6745_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_16_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold108 _6950_/Q hold108/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4370_ _3402_/I _4456_/B _5051_/S _4884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_176_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold119 _4250_/Z _6766_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3321_ _7226_/Q _5911_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_99_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6040_ _6040_/I _6041_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_844 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6942_ _6942_/D _7238_/RN _6942_/CLK _6942_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_81_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6873_ _6873_/D _6631_/Z _4075_/I1 _6873_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_23_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5824_ hold86/Z hold633/Z _5829_/S _5824_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5755_ hold29/Z hold462/Z _5757_/S _5755_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4706_ _4765_/A1 _4782_/A1 _5302_/B _5218_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_5686_ hold610/Z hold86/Z _5691_/S _5686_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4637_ _4565_/Z _5293_/B _5039_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_148_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold620 _6949_/Q hold620/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_150_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4568_ _5129_/A3 _4835_/A2 _3401_/I _3402_/I _4568_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold642 _7176_/Q hold642/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap361 input75/Z _7297_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_2_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold631 _4341_/Z _4343_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold653 _4138_/Z _6690_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4499_ _4759_/A2 _4759_/A3 _4718_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7287_ _7287_/D _6641_/Z _4072_/B2 hold61/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold664 _6901_/Q hold664/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3519_ _3653_/A1 hold629/Z hold338/Z _3497_/I _3519_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_89_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold686 _5614_/Z _6974_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6307_ _6307_/A1 _6307_/A2 _6307_/A3 _6306_/Z _6307_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold675 _6720_/Q hold675/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold697 _6821_/Q hold697/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6238_ _7020_/Q _6235_/Z _6237_/Z _6988_/Q _6260_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6169_ _6169_/A1 _6169_/A2 _6169_/A3 _6169_/A4 _6169_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__19 _4073__19/I _7206_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_185_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_663 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3870_ _7103_/Q _5758_/A1 _3947_/A2 _7095_/Q _3873_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_32_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5540_ hold113/Z hold165/Z _5547_/S _5540_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5471_ _5471_/A1 _5291_/C _4555_/C _5471_/B2 _5472_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4422_ _4402_/B _4026_/B _4026_/C _4422_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_69_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7210_ _7210_/D _7210_/RN _7210_/CLK _7210_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_8_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7141_ hold8/Z _7238_/RN _7141_/CLK _7141_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4353_ _3529_/Z _5520_/C hold637/Z _5821_/A3 _4353_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3304_ _6733_/Q _4041_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_101_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4284_ _6567_/I0 _6794_/Q _4288_/S _6794_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7072_ _7072_/D _7260_/RN _7072_/CLK _7072_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_99_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6023_ _6941_/Q _5972_/Z _6021_/Z _6997_/Q _6026_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_67_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_124 net463_133/I _7101_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet463_113 net613_291/I _7112_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_102 net613_264/I _7123_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet463_135 net413_73/I _7090_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_146 net463_147/I _7079_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6925_ _6925_/D _7210_/RN _6925_/CLK _6925_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6856_ _6856_/D _7219_/RN _6856_/CLK _6856_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_167_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3999_ _3999_/I _6835_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5807_ hold52/Z hold514/Z _5811_/S _5807_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6787_ _6787_/D _7193_/RN _6787_/CLK _6787_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_22_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5738_ hold15/Z hold448/Z _5739_/S _5738_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5669_ hold264/Z hold52/Z _5673_/S _5669_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold450 _6938_/Q hold450/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold461 _5872_/Z _7203_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold472 _4132_/Z _6685_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold494 _7206_/Q hold494/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold483 _6677_/Q hold483/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_78_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_22__1359_ net613_253/I net413_98/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_102__1359_ clkbuf_4_5_0__1359_/Z net763_424/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_85__1359_ net613_299/I net613_291/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_14_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4971_ _5464_/A1 _4905_/Z _4975_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_91_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3922_ _6855_/Q _3922_/A2 _3922_/B1 _6692_/Q _3922_/C _3963_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6710_ _6710_/D input75/Z _6710_/CLK _6710_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6641_ _7221_/RN _6656_/A2 _6641_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_149_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3853_ _3853_/I _3854_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6572_ _6575_/A2 _6572_/A2 _6608_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_118_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3784_ _3784_/I _3785_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5523_ hold559/Z hold52/Z hold34/Z _6896_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5454_ _5454_/A1 _5454_/A2 _5454_/A3 _5453_/Z _5455_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_105_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5385_ _5385_/A1 _5389_/C _5439_/B1 _5393_/A1 _5385_/C _5434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4405_ _4489_/B _4483_/B _4722_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_133_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7124_ _7124_/D _7258_/RN _7124_/CLK _7124_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4336_ _4103_/I hold640/Z _4337_/S _4336_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7055_ _7055_/D _7258_/RN _7055_/CLK _7055_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4267_ hold81/Z hold62/Z _4270_/S hold82/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4198_ hold795/Z hold271/Z _4210_/S _4198_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6006_ _7231_/Q _7228_/Q _7227_/Q wire348/I _6006_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_83_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6908_ _6908_/D _7193_/RN _6908_/CLK _6908_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_70_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6839_ _6839_/D _7210_/RN _6839_/CLK _6839_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_24_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold280 _6888_/Q hold280/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold291 _5725_/Z _7073_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet663_308 net763_418/I _6917_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_319 net813_470/I _6906_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5170_ _5172_/B _5170_/A2 _5170_/A3 _5172_/C _5170_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_110_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4121_ hold271/Z hold842/Z _4127_/S _4121_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4052_ _4052_/I _4052_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 mask_rev_in[0] input4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4954_ _5464_/A1 _5324_/A1 _4759_/Z _5263_/A4 _5068_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_91_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3905_ _6894_/Q _3904_/Z _3944_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_177_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4885_ _4887_/A1 _5315_/A2 _4551_/Z _4675_/Z _4885_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_60_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6624_ _7237_/RN _6656_/A2 _6624_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_165_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3836_ _3515_/Z _3533_/Z _3914_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3767_ _6700_/Q _3927_/A2 _3786_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6555_ _6548_/Z _6554_/Z _6555_/B1 _6286_/Z _6555_/C _6556_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_118_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5506_ hold366/Z hold86/Z _5509_/S _5506_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6486_ _6486_/A1 _6486_/A2 _6486_/A3 _6486_/A4 _6486_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_106_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3698_ _7056_/Q _5701_/A1 _5674_/A1 _7032_/Q _3952_/A2 _7048_/Q _3701_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5437_ _5437_/A1 _5437_/A2 _5436_/Z _5437_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xoutput330 _7265_/Q wb_dat_o[27] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput341 _6801_/Q wb_dat_o[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5368_ _5368_/A1 _5276_/C _5368_/B _5368_/C _5369_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_4319_ _4318_/Z _6833_/Q _6832_/Q _4313_/Z _6819_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_141_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5299_ _5210_/Z _5396_/A1 _5267_/Z _5298_/Z _5299_/C _5300_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_7107_ _7107_/D _7210_/RN _7107_/CLK _7107_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_102_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7038_ _7038_/D _7258_/RN _7038_/CLK _7038_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_75_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4670_ _4670_/A1 _4667_/Z _4669_/Z _4670_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_159_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3621_ _6946_/Q _5575_/A1 _3642_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_30_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3552_ _3473_/Z _3552_/A2 _3484_/Z _3477_/Z _3552_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6340_ _7176_/Q _6254_/Z _6355_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_183_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3483_ _6662_/Q _6661_/Q _6733_/Q _3483_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6271_ _6260_/Z _6271_/A2 _6271_/A3 _6271_/A4 _6271_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_143_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5222_ _5222_/A1 _5310_/A2 _5223_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5153_ _5150_/Z _5487_/A2 _5153_/A3 _5289_/A3 _5153_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_111_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4104_ _4103_/I hold846/Z _4118_/S _4104_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5084_ _5359_/A1 _4982_/Z _5085_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4035_ _4034_/Z _4035_/A2 _4035_/A3 _4035_/A4 _4036_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_65_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ _7110_/Q _5984_/Z _5985_/Z _7060_/Q _6009_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4937_ _4998_/A2 _5328_/A1 _5056_/C _5442_/A2 _4937_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_80_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4868_ _4868_/A1 _4524_/Z _5287_/B _4683_/Z _4868_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_177_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6607_ _4900_/B _6607_/A2 _6610_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3819_ _3552_/Z hold630/Z _4182_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_165_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4799_ _4422_/Z _4534_/Z _4568_/Z _5312_/A1 _4799_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_107_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6538_ _6723_/Q _6292_/Z _6299_/Z _6858_/Q _6548_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_134_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6469_ _7010_/Q _6243_/Z _6269_/Z _7034_/Q _6469_/C _6472_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput182 _4064_/Z mgmt_gpio_oeb[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput171 _4065_/Z mgmt_gpio_oeb[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput193 _3377_/ZN mgmt_gpio_oeb[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_101_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5840_ hold113/Z hold580/Z _5847_/S _5840_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5771_ hold52/Z hold590/Z _5775_/S _5771_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4722_ _5083_/C _4722_/A2 _4923_/A2 _5083_/B _5324_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_14_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4653_ _4653_/A1 _5040_/C _4653_/A3 _5041_/B _4657_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_147_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput40 mgmt_gpio_in[13] input40/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4584_ _4584_/A1 _4584_/A2 _5349_/B _4591_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_175_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput62 mgmt_gpio_in[33] input62/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput51 mgmt_gpio_in[23] input51/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3604_ _7149_/Q _3951_/C1 _5638_/A1 _7003_/Q _3606_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xinput73 pad_flash_io0_di input73/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold802 _4327_/Z _6824_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput95 wb_adr_i[0] _3401_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_128_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3535_ hold338/Z _3617_/A1 hold629/Z _3489_/I _3535_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xinput84 spimemio_flash_csb input84/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6323_ _7095_/Q _6250_/Z _6257_/Z _7061_/Q _6275_/Z _7037_/Q _6328_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold835 _6933_/Q hold835/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold846 _6666_/Q hold846/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold824 _4290_/Z _6799_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold813 _6847_/Q hold813/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3466_ _3465_/Z hold999/Z input58/Z _3430_/S _3467_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold857 _4199_/Z _6736_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_153_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6254_ _7237_/Q _6533_/A3 _6452_/A4 _6285_/A2 _6254_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_104_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold868 _6740_/Q hold868/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold879 _4160_/Z _6707_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5205_ _5205_/A1 _5468_/A1 _5205_/B1 _5356_/C _5205_/C _5440_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_130_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3397_ _3397_/I _6592_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6185_ _7248_/Q _6185_/I1 _6558_/S _7248_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5136_ _5287_/C _4570_/Z _4598_/Z _4784_/Z _5374_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_69_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5067_ _4951_/Z _5078_/A2 _5070_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4018_ _6743_/Q _6901_/Q _4019_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_83_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5969_ _7231_/Q _6211_/B1 _6021_/A2 _7227_/Q _5969_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_12_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_172_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold109 _5587_/Z _6950_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_153_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3320_ _7224_/Q _5954_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_98_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6941_ _6941_/D _7238_/RN _6941_/CLK _6941_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_35_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6872_ _6872_/D _6630_/Z _4075_/I1 _6872_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_5823_ hold271/Z hold940/Z _5829_/S _5823_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5754_ hold62/Z hold569/Z _5757_/S _5754_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4705_ _5220_/B2 _4536_/Z _4491_/B _4705_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_5685_ hold966/Z hold271/Z _5691_/S _5685_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4636_ _4636_/A1 _5034_/B _4635_/Z _4639_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_120_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold610 _7038_/Q hold610/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold621 _5586_/Z _6949_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_162_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4567_ _5270_/A1 _4454_/Z _5389_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold643 _5842_/Z _7176_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6306_ _6306_/A1 _6306_/A2 _6306_/A3 _6306_/A4 _6306_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_1_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold654 _6726_/Q hold654/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold632 _4342_/Z _6845_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7286_ _7286_/D _6640_/Z _4072_/B2 hold51/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4498_ _4494_/Z _4496_/Z _4998_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold665 _5528_/Z hold665/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3518_ _3617_/A1 _3501_/Z _5513_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold687 _6728_/Q hold687/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold676 _4180_/Z _6720_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3449_ _7292_/Q _3449_/A2 _3450_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6237_ _7235_/Q _6533_/A2 _6533_/A3 _5942_/S _6237_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold698 _4322_/Z _6821_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6168_ _7059_/Q _5924_/Z _6015_/Z _7011_/Q _6168_/C _6169_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_76_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5119_ _4773_/Z _4874_/C _5238_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6099_ _7138_/Q _5994_/I _6015_/Z _7008_/Q hold64/I _5972_/Z _6101_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_2837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_45__1359_ net663_324/I _4073__12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_136_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5470_ _5470_/A1 _5372_/Z _5470_/A3 _5489_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_129_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4421_ _5420_/A3 _5420_/A2 _4456_/B _5051_/S _4421_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_172_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7140_ _7140_/D _7238_/RN _7140_/CLK hold25/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4352_ hold271/Z hold721/Z _4352_/S _4352_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3303_ hold21/Z _4317_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7071_ _7071_/D _7221_/RN _7071_/CLK _7071_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_113_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4283_ _6566_/I0 _6793_/Q _4288_/S _6793_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6022_ _7079_/Q _5996_/Z _6005_/Z _7037_/Q _6965_/Q _5979_/Z _6031_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_58_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet463_125 net413_97/I _7100_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_114 _4073__47/I _7111_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_103 net413_79/I _7122_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_136 net413_61/I _7089_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet463_147 net463_147/I _7078_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6924_ _6924_/D _7221_/RN _6924_/CLK _6924_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_81_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6855_ _6855_/D _7219_/RN _6855_/CLK _6855_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_50_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3998_ _6835_/Q _4097_/A1 _6829_/Q _3999_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5806_ hold86/Z hold408/Z _5811_/S _5806_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6786_ _6786_/D _7219_/RN _6786_/CLK _6786_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5737_ hold29/Z hold47/Z _5739_/S hold48/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5668_ hold115/Z hold86/Z _5673_/S _5668_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4619_ _4565_/Z _4614_/Z _5029_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_151_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5599_ hold29/Z hold58/Z hold12/Z _6961_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold451 _5573_/Z _6938_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold462 _7099_/Q hold462/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold440 _6784_/Q hold440/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7269_ _7269_/D _7269_/CLK _7269_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold473 _7054_/Q hold473/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold495 _5876_/Z _7206_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold484 _4123_/Z _6677_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_77_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4970_ _4970_/A1 _4967_/Z _4968_/Z _4969_/Z _4975_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_17_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3921_ _3921_/I _3922_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6640_ _7221_/RN _6656_/A2 _6640_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3852_ _7215_/Q _3912_/A2 _3922_/A2 _6856_/Q _3853_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_60_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6571_ _6571_/I0 _7269_/Q _6571_/S _7269_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5522_ hold566/Z hold62/Z hold34/Z _6895_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3783_ _7022_/Q _5665_/A1 _3959_/B1 _6668_/Q _3923_/C1 _7080_/Q _3784_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_157_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5453_ _5126_/I _5452_/Z _5129_/Z _5453_/A4 _5453_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4404_ _4424_/B _4402_/B _4922_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_173_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5384_ _6577_/C _5267_/Z _5382_/Z _5384_/B _6862_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_5_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7123_ hold60/Z _7260_/RN _7123_/CLK hold59/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4335_ _5520_/C _3529_/Z _5513_/A3 _5857_/A2 _4337_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_114_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4266_ hold75/Z hold52/Z _4270_/S hold76/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7054_ _7054_/D _7210_/RN _7054_/CLK _7054_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xclkbuf_leaf_91__1359_ net813_465/I net763_422/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_189_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4197_ _4196_/Z hold747/Z _4211_/S _4197_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6005_ _7230_/Q _7229_/Q _6117_/A4 _6210_/A2 _6005_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_28_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6907_ _6907_/D input75/Z _6907_/CLK _6907_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_39_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6838_ _6838_/D _7210_/RN _6838_/CLK _6838_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_168_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6769_ _6769_/D _7237_/RN _6769_/CLK _6769_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_149_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold270 _7284_/Q hold270/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold292 _6704_/Q hold292/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_105_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold281 _5509_/Z _6888_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet663_309 net763_419/I _6916_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_120_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4120_ _4103_/I hold759/Z _4127_/S _4120_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4051_ _7201_/Q input82/Z _4055_/S _4052_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput5 mask_rev_in[10] input5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4953_ _4953_/A1 _5065_/B _4953_/A3 _4955_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_149_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3904_ _3489_/I _3904_/A2 hold338/Z _3904_/A4 _3904_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_33_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6623_ _7237_/RN _6657_/A2 _6623_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_4884_ _4884_/A1 _4659_/Z _4675_/Z _3401_/I _4884_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_20_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3835_ _3485_/Z _3560_/Z _3922_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_20_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3766_ input26/Z _3927_/C2 _3794_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6554_ _6554_/A1 _6554_/A2 _6554_/A3 _6553_/Z _6554_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_146_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6485_ _7117_/Q _6240_/Z _6297_/Z _6705_/Q _6485_/C _6486_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_5505_ hold741/Z hold271/Z _5509_/S _5505_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5436_ _4576_/C _5472_/A2 _5009_/Z _5435_/Z _5436_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_161_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3697_ hold64/I _5575_/A1 _3707_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_126_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput331 _7266_/Q wb_dat_o[28] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput320 _6793_/Q wb_dat_o[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_10_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput342 _6802_/Q wb_dat_o[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5367_ _4568_/Z _4586_/Z _5368_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_120_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4318_ _4316_/Z _4318_/A2 _6833_/D _6828_/Q _4318_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5298_ _5296_/Z _5382_/A3 _5173_/Z _5464_/B _5298_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_59_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7106_ _7106_/D _7297_/RN _7106_/CLK _7106_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4249_ hold86/Z hold167/Z _4252_/S _4249_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7037_ _7037_/D _7219_/RN _7037_/CLK _7037_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_67_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3620_ hold26/I _5584_/A1 _3630_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3551_ _3525_/Z _3537_/Z _3917_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_183_892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3482_ _4041_/B1 _6662_/Q _3975_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_170_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6270_ _6948_/Q _6268_/Z _6269_/Z _7028_/Q _6271_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_102_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5221_ _5221_/I _5401_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_44_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5152_ _5364_/B _4614_/Z _4784_/Z _4624_/Z _4570_/Z _5153_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_116_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4103_ _4103_/I _5520_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5083_ _4977_/Z _4981_/Z _5083_/B _5083_/C _5337_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_110_152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4034_ _4033_/Z _4034_/A2 _4388_/A2 _4388_/A1 _4034_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_37_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5985_ _7231_/Q _6210_/C _6021_/A2 _7227_/Q _5985_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XPHY_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_162_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4936_ _4936_/I _5410_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_36_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4867_ _5269_/A2 _4530_/I _5287_/B _5293_/B _4867_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XANTENNA_10 _5538_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6606_ _4686_/B _6606_/A2 _6610_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_138_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3818_ _3535_/Z _3552_/Z _3960_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_181_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4798_ _4568_/Z _4793_/Z _5452_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6537_ _6717_/Q _6250_/Z _6290_/Z _6709_/Q _6302_/Z _6713_/Q _6548_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_119_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3749_ _7129_/Q _3930_/A2 _5758_/A1 _7105_/Q _3941_/B1 _7169_/Q _3751_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_122_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6468_ _6468_/I _6469_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5419_ _5419_/A1 _5419_/A2 _5418_/Z _5431_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_133_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6399_ _7218_/Q _6274_/Z _6285_/Z _7194_/Q _7178_/Q _6254_/Z _6401_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xnet713_390 net713_390/I _6784_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput194 _3349_/ZN mgmt_gpio_oeb[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput183 _3359_/ZN mgmt_gpio_oeb[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_115_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput172 _3369_/ZN mgmt_gpio_oeb[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_82_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_472 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ hold86/Z hold662/Z _5775_/S _5770_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4721_ _4721_/A1 _4721_/A2 _4721_/B _5323_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_159_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4652_ _4436_/B _5139_/A2 _5471_/B2 _5281_/C _5041_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3603_ _7117_/Q _3917_/A2 _5758_/A1 _7109_/Q _5674_/A1 _7035_/Q _3606_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xinput30 mask_rev_in[4] input30/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4583_ _4570_/Z _5016_/B2 _5349_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput63 mgmt_gpio_in[34] input63/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput41 mgmt_gpio_in[14] input41/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput52 mgmt_gpio_in[24] input52/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold803 _6839_/Q hold803/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput96 wb_adr_i[10] input96/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_174_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3534_ _3497_/I _3501_/Z hold637/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xinput85 spimemio_flash_io0_do input85/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6322_ _6322_/A1 _6322_/A2 _6322_/A3 _6322_/A4 _6322_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold825 _6838_/Q hold825/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold836 _5568_/Z _6933_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput74 pad_flash_io1_di _3337_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold814 _4345_/Z _6847_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3465_ _3464_/Z _3442_/B _3465_/A3 _3465_/A4 _3465_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_171_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6253_ _7236_/Q _6300_/A2 _6533_/A4 _6302_/A4 _6253_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold869 _4207_/Z _6740_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold847 _4104_/Z _6666_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold858 _6893_/Q hold858/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5204_ _5346_/A2 _5387_/A1 _5403_/B2 _5205_/A1 _5204_/C _5357_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_103_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_9__1359_ net413_58/I net813_473/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3396_ _3396_/I _6589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6184_ _6555_/C _6181_/Z _6184_/A3 _6184_/B _6185_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_5135_ _4589_/Z _4817_/Z _5287_/C _5487_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_97_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5066_ _4944_/Z _5078_/A2 _5066_/B _5481_/C _5070_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_4017_ _4006_/Z _4019_/A2 _4020_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5968_ _6014_/A2 _7229_/Q _6211_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_52_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4919_ _5343_/A1 _4496_/Z _5056_/C _5442_/A2 _4927_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5899_ _5910_/B _5899_/I1 _7223_/Q _7223_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_68__1359_ clkbuf_4_15_0__1359_/Z net763_419/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_148__1359_ net713_387/I net813_471/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_157_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6940_ _6940_/D _7238_/RN _6940_/CLK _6940_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_81_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6871_ _6871_/D _6629_/Z _4075_/I1 _6871_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_5822_ _4103_/I hold894/Z _5829_/S _5822_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5753_ hold52/Z hold300/Z _5757_/S _5753_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4704_ _4687_/Z _4704_/A2 _5255_/A2 _5092_/A1 _5098_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_148_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5684_ hold942/Z _4103_/I _5691_/S _5684_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4635_ _4868_/A1 _4524_/Z _4546_/Z _5364_/B _4635_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_136_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _4422_/Z _5278_/C _4554_/Z _4483_/B _4576_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_118_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold600 _6741_/Q hold600/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold611 _5686_/Z _7038_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_162_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xmax_cap352 _5364_/B _5287_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
Xhold644 _7217_/Q hold644/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3517_ _3489_/I _3492_/Z _5839_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold633 _7160_/Q hold633/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6305_ _7198_/Q _6272_/Z _6275_/Z _7036_/Q _6306_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold622 _7021_/Q hold622/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4497_ _4436_/B _4497_/A2 _4497_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
XFILLER_171_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7285_ _7285_/D _6639_/Z _4072_/B2 hold85/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_131_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold666 _6694_/Q hold666/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold688 _4192_/Z _6728_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold655 _4189_/Z _6726_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold677 _6857_/Q hold677/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3448_ _3448_/I _7293_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6236_ _5943_/S _7234_/Q _6533_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_131_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold699 _6932_/Q hold699/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_134_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6167_ _6947_/Q _5972_/Z _6021_/Z _7003_/Q _6169_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_58_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3379_ _6929_/Q _6447_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_5118_ _5115_/Z _5117_/Z _5118_/A3 _5215_/C _5118_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6098_ _7090_/Q _6002_/Z _6019_/Z _7048_/Q _6098_/C _6101_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_45_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5049_ _5049_/A1 _5210_/A4 _5180_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_84_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4420_ _5170_/A2 _4836_/A4 _5258_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_172_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4351_ _4103_/I hold683/Z _4352_/S _4351_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3302_ hold17/I _6608_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7070_ _7070_/D _7221_/RN _7070_/CLK _7070_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_99_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4282_ _6565_/I0 _6792_/Q _4288_/S _6792_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6021_ _6211_/B1 _6021_/A2 _6210_/A2 _7227_/Q _6021_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xnet463_104 _4073__22/I _7121_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_115 _4073__51/I _7110_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_126 _4073__22/I _7099_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet463_137 net413_57/I _7088_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_148 _4073__3/I _7077_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6923_ _6923_/D _7258_/RN _6923_/CLK _6923_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_62_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6854_ _6854_/D input75/Z _6854_/CLK _6854_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_149_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3997_ _3997_/I _6834_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6785_ _6785_/D _7219_/RN _6785_/CLK _6785_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5805_ hold271/Z hold923/Z _5811_/S _5805_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5736_ hold62/Z hold68/Z _5739_/S hold69/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_131__1359_ _4073__15/I net713_379/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_148_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5667_ hold622/Z hold271/Z _5673_/S _5667_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4618_ _4618_/A1 _5151_/B _4616_/Z _4617_/Z _4622_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_135_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5598_ hold62/Z hold215/Z hold12/Z _6960_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4549_ _5288_/B _4467_/B _4460_/B _4472_/B _4549_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_144_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold430 _7220_/Q hold430/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold452 _6768_/Q hold452/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold463 _5755_/Z _7099_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold441 _4270_/Z _6784_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_145_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7268_ _7268_/D _7269_/CLK _7268_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold474 _5704_/Z _7054_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold485 _6958_/Q hold485/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold496 _7044_/Q hold496/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6219_ _6844_/Q _5971_/Z _5981_/Z _6788_/Q _6005_/Z _6850_/Q _6220_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_131_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7199_ _7199_/D _7219_/RN _7199_/CLK _7199_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_58_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3920_ input71/Z _4244_/S _3920_/B1 _6866_/Q _6902_/Q _3920_/C2 _3921_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_44_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3851_ _7159_/Q _3941_/A2 _3912_/C1 _6707_/Q _4170_/A1 _6715_/Q _3855_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_158_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6570_ _6570_/I0 _7268_/Q _6571_/S _7268_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3782_ _7014_/Q _5656_/A1 _5638_/A1 _6998_/Q _3951_/C1 _7144_/Q _3786_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_185_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5521_ hold33/Z _5521_/A2 hold18/Z hold11/Z hold34/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_74_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5452_ _4791_/Z _5452_/A2 _5452_/A3 _4801_/Z _5452_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4403_ _4424_/B _4402_/B _4923_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5383_ _6862_/Q _6577_/C _5212_/Z _5320_/Z _5383_/C _5384_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4334_ hold271/Z hold890/Z _4334_/S _4334_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7122_ _7122_/D _7297_/RN _7122_/CLK _7122_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_119_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7053_ _7053_/D _7210_/RN _7053_/CLK _7053_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_6004_ _7086_/Q _6002_/Z _6003_/Z _7158_/Q _6008_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4265_ _6779_/Q hold86/Z _4270_/S hold87/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4196_ hold238/Z _4102_/Z _4210_/S _4196_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6906_ _6906_/D input75/Z _6906_/CLK _6906_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_42_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6837_ _6837_/D _7210_/RN _6837_/CLK _6837_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6768_ _6768_/D _7193_/RN _6768_/CLK _6768_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5719_ _5857_/A2 _5857_/A3 _3537_/Z hold6/Z _5727_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6699_ _6699_/D _7297_/RN _6699_/CLK _6699_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_137_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold271 hold274/Z hold271/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold260 _6880_/Q hold260/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_46_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold293 _4156_/Z _6704_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold282 _6930_/Q hold282/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_105_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_10_0__1359_ clkbuf_0__1359_/Z net663_304/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_2421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2498 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4050_ _4050_/I0 input90/Z _4050_/S _4050_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput6 mask_rev_in[11] input6/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4952_ _5359_/A1 _4951_/Z _4953_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_149_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4883_ _4881_/Z _4882_/Z _4886_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_51_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3903_ _3903_/A1 _5821_/A3 _5513_/A3 _3533_/Z _3903_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6622_ _7237_/RN _4064_/S _6622_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3834_ _3485_/Z _3535_/Z _3956_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_177_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3765_ _7046_/Q _3952_/A2 _3916_/B1 _6880_/Q _3790_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6553_ _6553_/A1 _6553_/A2 _6553_/A3 _6553_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6484_ _7133_/Q _6484_/A2 _6484_/A3 _6533_/A4 _6485_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5504_ hold420/Z _4103_/I _5509_/S _5504_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3696_ _7008_/Q _3934_/A2 _3701_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5435_ _5438_/C _5435_/A2 _5475_/A3 _4666_/Z _5435_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_145_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput310 _7261_/Q wb_ack_o VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_156_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput332 _7267_/Q wb_dat_o[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput321 _6794_/Q wb_dat_o[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5366_ _5366_/A1 _5366_/A2 _5365_/Z _5469_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_114_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4317_ _4317_/A1 _6826_/Q _4318_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5297_ _4882_/Z _5170_/Z _5382_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7105_ _7105_/D _7221_/RN _7105_/CLK _7105_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_114_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4248_ hold271/Z hold715/Z _4252_/S _4248_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7036_ _7036_/D _7193_/RN _7036_/CLK _7036_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_45_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4179_ _5821_/A3 hold637/Z _3537_/Z _5520_/C _4181_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_71_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet763_450 net413_71/I _6715_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3550_ _3485_/Z _3507_/Z _3955_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_128_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3481_ hold37/Z _3552_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
X_5220_ _4694_/Z _5310_/A2 _5220_/B1 _5220_/B2 _5221_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_170_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5151_ _5287_/C _5364_/B _4784_/Z _5151_/B _5487_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_96_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4102_ input58/Z hold112/Z hold21/Z _4102_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_5082_ _4980_/Z _5081_/Z _5412_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_110_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4033_ _4028_/Z _4030_/Z _4026_/B _4026_/C _4033_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_38_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5984_ _5984_/A1 _6210_/B _7231_/Q _7230_/Q _5984_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4935_ _5442_/A2 _4497_/Z _4495_/Z _5056_/C _4936_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_52_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4866_ _4868_/A1 _4524_/Z _5414_/A2 _5287_/B _4866_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XANTENNA_11 debug_oeb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6605_ _4415_/B _6605_/A2 _6610_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_159_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4797_ _4791_/Z _5452_/A2 _5453_/A4 _4797_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_3817_ _3527_/Z _3542_/Z _5536_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3748_ _6677_/Q _3546_/Z _3947_/A2 _7097_/Q _6896_/Q _5528_/S _3758_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_20_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6536_ _6691_/Q _6257_/Z _6275_/Z _6850_/Q _6300_/Z _6721_/Q _6548_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_180_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3679_ _5857_/A2 _5513_/A3 _5503_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6467_ _7026_/Q _6235_/Z _6262_/Z _6970_/Q _6265_/Z _7002_/Q _6468_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5418_ _5418_/A1 _5418_/A2 _5417_/Z _5418_/A4 _5418_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_82_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6398_ _7098_/Q _6250_/Z _6302_/Z _7090_/Q _6401_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xnet713_380 net763_447/I _6810_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5349_ _5349_/A1 _5387_/A2 _5349_/B _5350_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xoutput195 _3348_/ZN mgmt_gpio_oeb[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput184 _3358_/ZN mgmt_gpio_oeb[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput173 _3368_/ZN mgmt_gpio_oeb[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_87_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet713_391 net813_491/I _6783_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7019_ _7019_/D _7258_/RN _7019_/CLK _7019_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_46_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_28__1359_ clkbuf_opt_2_0__1359_/Z net763_409/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_108__1359_ clkbuf_4_5_0__1359_/Z net613_288/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_39_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4720_ _5083_/C _5083_/B _5259_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_1391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4651_ _4467_/B _4460_/B _4501_/B _4472_/B _4651_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3602_ _7213_/Q _3960_/A2 _3955_/A2 _7205_/Q hold91/I _5584_/A1 _3607_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xinput20 mask_rev_in[24] input20/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput31 mask_rev_in[5] input31/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4582_ _4638_/A2 _5345_/A2 _4438_/B _4467_/B _5016_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xinput64 mgmt_gpio_in[35] input64/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput42 mgmt_gpio_in[15] input42/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput53 mgmt_gpio_in[25] input53/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput97 wb_adr_i[11] input97/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_115_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3533_ hold32/Z _3477_/Z hold37/Z _3484_/Z _3533_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xinput86 spimemio_flash_io0_oeb input86/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6321_ _7069_/Q _6248_/Z _6297_/Z _6699_/Q _6321_/C _6322_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold826 _4331_/Z _6838_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold804 _4333_/Z _6839_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput75 porb input75/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
Xhold815 _6809_/Q hold815/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold837 _7005_/Q hold837/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3464_ _7283_/Q _6665_/Q _6664_/Q _6663_/Q _3464_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_66_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold848 _6693_/Q hold848/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold859 _5518_/Z _6893_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6252_ _7094_/Q _6250_/Z _6251_/Z _6980_/Q _6259_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5203_ _5199_/Z _5354_/A2 _5202_/Z _5203_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_130_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6183_ _6555_/C _7247_/Q _6184_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3395_ _3395_/I _6586_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5134_ _5293_/A1 _4624_/Z _5275_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5065_ _4699_/Z _5252_/B _5065_/B _5481_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_96_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4016_ _6744_/Q _5896_/I0 _4019_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_25_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5967_ _7231_/Q _7228_/Q _7227_/Q _6002_/A2 _5967_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_80_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4918_ _4927_/A1 _4927_/A2 _5444_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_40_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5898_ _5901_/B _5899_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4849_ _4598_/Z _4681_/Z _4849_/B _5373_/B _4852_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_20_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6519_ _6716_/Q _6250_/Z _6293_/Z _6718_/Q _6521_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_134_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6870_ _6870_/D _6628_/Z _4075_/I1 _6870_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_179_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5821_ _5520_/C _3552_/Z _5821_/A3 _5857_/A3 _5829_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_34_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5752_ hold86/Z hold481/Z _5757_/S _5752_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4703_ _5420_/A2 _5129_/A3 _4835_/A2 _3401_/I _4703_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5683_ _5683_/A1 hold18/Z _5691_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_4634_ _4868_/A1 _4524_/Z _4551_/Z _5364_/B _5034_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_163_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4565_ _5364_/B _5051_/S _4456_/B _4454_/Z _4565_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold612 _7209_/Q hold612/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold601 _4209_/Z _6741_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmax_cap353 _7221_/RN _7237_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_128_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold645 _5888_/Z _7217_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3516_ _3485_/Z _3515_/Z _3912_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold634 _5824_/Z _7160_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6304_ _7166_/Q _5948_/Z _6273_/Z _6972_/Q _6306_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold623 _5667_/Z _7021_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4496_ _4467_/B _4497_/A2 _4496_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_7284_ _7284_/D _6638_/Z _4072_/B2 _7284_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_143_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold656 _7210_/Q hold656/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold667 _4144_/Z _6694_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold678 _4360_/Z _6857_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3447_ _7293_/Q _3449_/A2 _3447_/B1 _7292_/Q _3448_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_6235_ _7235_/Q _7234_/Q _6533_/A2 _6533_/A3 _6235_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold689 _6722_/Q hold689/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_100_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6166_ _6987_/Q _5988_/Z _6019_/Z _7051_/Q _6169_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_57_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3378_ _6928_/Q _6418_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_74__1359_ net663_324/I net413_68/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5117_ _5117_/A1 _5117_/A2 _5117_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_58_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6097_ _6097_/I _6098_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5048_ _5395_/A1 _4991_/C _5210_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_111_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2806 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6999_ _6999_/D _7260_/RN _6999_/CLK _6999_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_41_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_292 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4350_ _3485_/Z _3535_/Z _5520_/C _4352_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_3301_ _6663_/Q _3971_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_141_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4281_ _6564_/I0 _6791_/Q _4288_/S _6791_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6020_ _6933_/Q _5981_/Z _6019_/Z _7045_/Q _6037_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_67_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_116 net413_68/I _7109_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet463_105 net563_251/I _7120_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_127 net413_99/I _7098_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_138 net613_253/I _7087_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_149 _4073__3/I _7076_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6922_ _6922_/D _7258_/RN _6922_/CLK _6922_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6853_ _6853_/D input75/Z _6853_/CLK _6853_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5804_ hold113/Z hold401/Z _5811_/S _5804_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3996_ _6834_/Q _4097_/A1 _6828_/Q _3997_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6784_ _6784_/D _7260_/RN _6784_/CLK _6784_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5735_ hold52/Z hold551/Z _5739_/S _5735_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5666_ _7020_/Q hold113/Z _5673_/S _5666_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4617_ _4422_/Z _4546_/Z _4614_/Z _4483_/B _4617_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_108_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5597_ hold52/Z hold259/Z hold12/Z _6959_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold420 _6883_/Q hold420/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4548_ _4441_/B _5281_/C _4436_/B _4501_/B _4555_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_144_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold431 _5891_/Z _7220_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold442 _7180_/Q hold442/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_117_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold453 _4252_/Z _6768_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xclkbuf_4_8_0__1359_ clkbuf_0__1359_/Z clkbuf_4_8_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_171_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4479_ _4786_/A1 _4786_/A2 _4786_/A3 _5094_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
Xhold464 _6962_/Q hold464/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7267_ _7267_/D _7269_/CLK _7267_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold486 _7152_/Q hold486/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold475 _6684_/Q hold475/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold497 _5693_/Z _7044_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6218_ _6790_/Q _5972_/Z _6021_/Z _6840_/Q _6220_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_86_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7198_ _7198_/D _7219_/RN _7198_/CLK _7198_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_100_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6149_ _6986_/Q _5988_/Z _5996_/Z _7084_/Q _6152_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_57_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3850_ _7069_/Q _3943_/A2 _4244_/S input72/Z _4161_/A1 _6709_/Q _3855_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3781_ _6974_/Q _3923_/A2 _3957_/A2 _6958_/Q _3956_/A2 _7120_/Q _3786_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_13_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5520_ hold339/Z _5520_/A2 _5520_/B _5520_/C hold340/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_8_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5451_ _4492_/Z _4536_/Z _5451_/B _5451_/C _5454_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_67_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4402_ _4580_/C _4489_/A1 _4402_/B _4412_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_145_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5382_ _5379_/Z _5464_/B _5382_/A3 _5382_/A4 _5382_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_126_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7121_ _7121_/D _7219_/RN _7121_/CLK _7121_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4333_ _4103_/I hold803/Z _4334_/S _4333_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7052_ _7052_/D _7210_/RN _7052_/CLK _7052_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4264_ hold763/Z hold271/Z _4270_/S _4264_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6003_ _6015_/A3 wire348/Z _7231_/Q _7228_/Q _6003_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4195_ _4210_/S _4194_/Z _6652_/A2 _3540_/Z hold18/Z _4211_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_95_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6905_ _6905_/D _7219_/RN _6905_/CLK _6905_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_70_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6836_ _6836_/D _7279_/RN _7279_/CLK _6836_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_126_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6767_ _6767_/D _7193_/RN _6767_/CLK _6767_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3979_ _3978_/Z _6661_/Q _3988_/S _6661_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5718_ hold2/Z hold190/Z _5718_/S _5718_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6698_ _6698_/D _7210_/RN _6698_/CLK _6698_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_164_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5649_ hold837/Z hold271/Z _5655_/S _7005_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold250 _6967_/Q hold250/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold261 _5500_/Z _6880_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_6_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold283 _5564_/Z _6930_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_85_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold272 _5496_/Z _6877_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold294 _7065_/Q hold294/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_46_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput7 mask_rev_in[12] input7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4951_ _4407_/Z _5259_/A1 _4759_/Z _5263_/A4 _4951_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_91_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4882_ _4367_/Z _4555_/B _5172_/B _5172_/C _4882_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3902_ _6889_/Q _3902_/A2 _3960_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_6621_ _7237_/RN _6657_/A2 _6621_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_20_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3833_ _3529_/Z _3578_/Z _3936_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_177_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3764_ _6676_/Q _3546_/Z _3776_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6552_ _6848_/Q _6269_/Z _6273_/Z _6823_/Q _6553_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_146_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6483_ _7205_/Q _6272_/Z _6296_/Z _7165_/Q _7067_/Q _6257_/Z _6486_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5503_ hold33/Z _5503_/A2 hold18/Z hold11/Z _5509_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_69_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3695_ _7106_/Q _5758_/A1 _3719_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_9_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5434_ _5434_/A1 _5434_/A2 _5432_/Z _5433_/Z _5441_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xoutput300 _3990_/I serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput322 _6812_/Q wb_dat_o[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput311 _6811_/Q wb_dat_o[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput333 _6813_/Q wb_dat_o[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5365_ _5468_/B1 _5288_/B _4441_/B _4363_/Z _5365_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_113_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7104_ _7104_/D _7258_/RN _7104_/CLK _7104_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4316_ _6830_/Q _6829_/Q _6831_/Q _4316_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_141_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5296_ _5271_/Z _5296_/A2 _5295_/Z _5467_/B _5296_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_101_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7035_ _7035_/D _7260_/RN _7035_/CLK _7035_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_75_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4247_ _4103_/I hold668/Z _4252_/S _4247_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4178_ hold271/Z hold884/Z _4178_/S _4178_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6819_ _6819_/D _7279_/RN _7279_/CLK hold21/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_143_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet763_440 net763_441/I _6725_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_451 net413_67/I _6714_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_611 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_159_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3480_ _3479_/Z hold36/Z hold21/Z hold37/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_151_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5150_ _5374_/A2 _5148_/Z _5374_/A1 _5487_/A1 _5150_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5081_ _5340_/A1 _5262_/A2 _5343_/A2 _5442_/A4 _5081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_111_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4101_ _3533_/Z _5520_/C hold637/Z _5839_/A3 _4118_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4032_ _4032_/A1 _4032_/A2 _4031_/Z _4035_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_111_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5983_ _7231_/Q _5983_/A2 _5983_/B _5983_/C _6010_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_24_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4934_ _5464_/A1 _5325_/B _5061_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_52_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4865_ _4865_/A1 _4865_/A2 _5156_/B _4869_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA_12 debug_out VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_6604_ _4316_/Z _6604_/A2 _6833_/D _6828_/Q _7278_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4796_ _4793_/Z _5394_/A2 _5453_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_119_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3816_ _3521_/Z _3527_/Z _3902_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_118_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3747_ _3747_/A1 _3747_/A2 _3747_/A3 _3747_/A4 _3747_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6535_ _6856_/Q _6256_/Z _6546_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_20_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6466_ _6466_/A1 _6466_/A2 _6466_/A3 _6465_/Z _6466_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3678_ input31/Z _3927_/C2 _3951_/A2 hold42/I _3686_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_12_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5417_ _5417_/A1 _5417_/A2 _5263_/Z _5417_/A4 _5417_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_133_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6397_ _7186_/Q _6282_/Z _6299_/Z _7056_/Q hold83/I _6237_/Z _6401_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xnet713_370 net813_489/I _6840_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_381 net763_447/I _6809_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5348_ _5348_/I _5437_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput174 _3367_/ZN mgmt_gpio_oeb[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_130_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput185 _3357_/ZN mgmt_gpio_oeb[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_114_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet713_392 net763_422/I _6782_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput196 _3732_/A1 mgmt_gpio_oeb[32] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_99_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5279_ _5288_/A1 _5279_/A2 _4555_/C _5439_/A1 _5279_/C _5284_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_88_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7018_ _7018_/D _7258_/RN _7018_/CLK _7018_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_56_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4650_ _4441_/B _5288_/B _5281_/C _4436_/B _4650_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_174_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3601_ _3601_/A1 _3601_/A2 _3601_/A3 _3601_/A4 _3601_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xinput10 mask_rev_in[15] input10/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 mask_rev_in[25] input21/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4581_ _4557_/Z _5435_/A2 _5349_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_174_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput43 mgmt_gpio_in[16] input43/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput54 mgmt_gpio_in[26] input54/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6320_ _6320_/A1 _6239_/Z _6321_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput32 mask_rev_in[6] input32/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput98 wb_adr_i[12] input98/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput65 mgmt_gpio_in[36] _7308_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput87 spimemio_flash_io1_do _7307_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3532_ hold38/Z hold135/Z _3904_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold827 _6748_/Q hold827/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold805 _6822_/Q hold805/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_7_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold816 _4302_/Z _6809_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput76 qspi_enabled _4050_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3463_ _7283_/Q _3462_/Z _3463_/S _7283_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold838 _6756_/Q hold838/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6251_ _6300_/A2 _5943_/S _7234_/Q _6533_/A2 _6251_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_116_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold849 _4142_/Z _6693_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_6_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5202_ _4626_/Z _5201_/Z _5202_/A3 _5202_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_131_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6182_ _6201_/A3 _6931_/Q _6184_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_88_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3394_ _3394_/I _6583_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5133_ _5165_/A2 _5287_/B _5288_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5064_ _5064_/A1 _5410_/B _5063_/I _5064_/A4 _5066_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_111_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4015_ _5957_/S _3990_/I _5953_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_53_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5966_ _6972_/Q _5964_/Z _5965_/Z _6698_/Q _5974_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_40_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4917_ _5328_/A1 _5056_/C _5442_/A2 _5442_/A4 _4927_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5897_ _6744_/Q _3990_/I _5901_/A1 _5950_/A1 _5901_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_33_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4848_ _4853_/A1 _5414_/A2 _5287_/B _4501_/B _5373_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_32_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_34__1359_ net463_109/I net413_72/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_114__1359_ net613_293/I net413_88/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_119_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4779_ _4700_/Z _4778_/Z _5456_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_97__1359_ clkbuf_4_5_0__1359_/Z net563_248/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_146_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6518_ _6824_/Q _6251_/Z _6256_/Z _6855_/Q _6521_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_10_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6449_ _6449_/I _6450_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5820_ hold2/Z hold232/Z _5820_/S _5820_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5751_ hold271/Z hold944/Z _5757_/S _5751_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4702_ _4884_/A1 _3401_/I _5255_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_15_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5682_ hold158/Z hold2/Z _5682_/S _5682_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4633_ _4633_/A1 _5035_/A4 _5387_/B _4636_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_129_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4564_ _4554_/Z _5364_/B _5439_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold602 _6910_/Q hold602/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7283_ _7283_/D _6637_/Z _7303_/CLK _7283_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xmax_cap343 _6657_/A2 _6656_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
Xhold635 _6860_/Q hold635/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold613 _5879_/Z _7209_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap354 _7219_/RN _7221_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold624 _6927_/Q hold624/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3515_ _3653_/A1 _3492_/Z _3497_/I _3501_/Z _3515_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6303_ _7214_/Q _6274_/Z _6302_/Z _7086_/Q _6306_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4495_ _4460_/B _4884_/A1 _4495_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
XFILLER_144_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6234_ _7233_/Q _7232_/Q _6533_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_89_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold646 _7200_/Q hold646/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold657 _5880_/Z _7210_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold679 _7120_/Q hold679/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold668 _6763_/Q hold668/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3446_ _3449_/A2 _3450_/A1 _3447_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6165_ _7019_/Q _5971_/Z _6005_/Z _7043_/Q _6169_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_69_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3377_ hold65/I _3377_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ _5117_/A1 _5117_/A2 _5316_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6096_ _7146_/Q _5987_/Z _6003_/Z _7162_/Q _6097_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5047_ _5047_/A1 _5360_/B _5049_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6998_ _6998_/D _7260_/RN _6998_/CLK _6998_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_26_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5949_ _6282_/A1 _5948_/Z _5950_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_129_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_80__1359_ _4073__15/I net613_267/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3300_ _6664_/Q _3465_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_125_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4280_ _6831_/Q _7279_/RN _4288_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_101_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet463_106 net463_147/I _7119_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_117 _4073__12/I _7108_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_128 net413_56/I _7097_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_139 net513_188/I _7086_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6921_ _6921_/D _7221_/RN _6921_/CLK _6921_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6852_ _6852_/D _7297_/RN _6852_/CLK _6852_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5803_ _3523_/Z _3552_/Z hold6/Z _5811_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_50_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3995_ _3994_/Z _3995_/A2 _4097_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_148_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6783_ _6783_/D input75/Z _6783_/CLK hold99/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5734_ hold86/Z hold144/Z _5739_/S _5734_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5665_ _5665_/A1 hold18/Z _5673_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_31_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4616_ _4422_/Z _4551_/Z _4614_/Z _4483_/B _4616_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_135_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5596_ hold86/Z hold485/Z hold12/Z _6958_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold410 _6879_/Q hold410/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_150_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4547_ _5278_/C _4878_/A2 _3401_/I _3402_/I _4547_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold443 _5846_/Z _7180_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold454 _7052_/Q hold454/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold421 _5504_/Z _6883_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold432 _6679_/Q hold432/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4478_ _4786_/A2 _4786_/A3 _4782_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7266_ _7266_/D _7269_/CLK _7266_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold487 _5815_/Z _7152_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold465 _6698_/Q hold465/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold476 _4131_/Z _6684_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3429_ _3971_/A1 _6730_/Q _6665_/Q _6664_/Q _3430_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_132_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7197_ _7197_/D _7221_/RN _7197_/CLK _7197_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold498 _6887_/Q hold498/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6217_ _6217_/A1 _6217_/A2 _6217_/A3 _6217_/A4 _6217_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6148_ _6970_/Q _5979_/Z _5999_/Z _7034_/Q _6152_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6079_ _7129_/Q _6000_/Z _6019_/Z _7047_/Q _6967_/Q _5979_/Z _6085_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_85_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3780_ _7208_/Q _3960_/A2 _3955_/A2 _7200_/Q _3796_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_185_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5450_ _5450_/I _5463_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4401_ _4412_/A1 _4399_/Z _5083_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_160_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5381_ _5381_/I _5382_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7120_ _7120_/D _7260_/RN _7120_/CLK _7120_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_5_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4332_ _3509_/Z _5839_/A3 hold637/Z _5520_/C _4334_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_114_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7051_ _7051_/D _7260_/RN _7051_/CLK _7051_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_87_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4263_ hold230/Z hold113/Z _4270_/S _4263_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6002_ _7231_/Q _6002_/A2 _6021_/A2 _7227_/Q _6002_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4194_ _4194_/A1 _3994_/Z _4194_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_94_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6904_ _6904_/D _7219_/RN _6904_/CLK _6904_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_82_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6835_ _6835_/D _7279_/RN _7230_/CLK _6835_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_51_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3978_ _3977_/Z _6660_/Q _6733_/Q _3978_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6766_ _6766_/D input75/Z _6766_/CLK _6766_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5717_ hold15/Z hold284/Z _5718_/S _5717_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_2_1__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _4072_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6697_ _6697_/D _7193_/RN _6697_/CLK _6697_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5648_ hold398/Z hold113/Z _5655_/S _7004_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5579_ hold65/Z hold52/Z hold23/Z _6943_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold251 _7007_/Q hold251/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold262 _6681_/Q hold262/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold240 _7048_/Q hold240/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold273 _7271_/Q hold273/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold284 _7066_/Q hold284/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_49_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold295 _5716_/Z _7065_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7249_ _7249_/D _7260_/RN _7260_/CLK _7249_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_120_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 mask_rev_in[13] input8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4950_ _5442_/A2 _4495_/Z _4496_/Z _4958_/A4 _5252_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_91_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4881_ _5104_/A1 _4555_/B _4650_/Z _5172_/C _4881_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3901_ _6980_/Q _3901_/A2 _3926_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_33_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6620_ _7237_/RN _6657_/A2 _6620_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3832_ _3519_/Z _3529_/Z _4359_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_158_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6551_ _6790_/Q _6245_/Z _6288_/Z _7297_/Q _6553_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3763_ input54/Z _4194_/A1 _3795_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5502_ hold138/Z hold62/Z _5502_/S _5502_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6482_ _7075_/Q _6248_/Z _6253_/Z _7141_/Q _7157_/Q _6293_/Z _6486_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3694_ _7064_/Q _3927_/B1 _3715_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_173_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5433_ _5433_/A1 _5433_/A2 _5433_/A3 _4662_/B _5433_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xoutput301 _3683_/Z serial_data_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5364_ _5414_/A2 _4551_/Z _5364_/B _5468_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_133_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput334 _7268_/Q wb_dat_o[30] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput323 _6795_/Q wb_dat_o[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput312 _6803_/Q wb_dat_o[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4315_ _6834_/Q _6835_/Q _6836_/Q _6832_/Q _5299_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_102_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7103_ _7103_/D _7219_/RN _7103_/CLK _7103_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_0_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5295_ _5295_/A1 _4501_/B _4472_/B _5315_/A1 _5295_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_141_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7034_ _7034_/D _7258_/RN _7034_/CLK _7034_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4246_ _3485_/Z _5821_/A3 _5513_/A3 _5520_/C _4252_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_95_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4177_ _4103_/I hold811/Z _4178_/S _4177_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6818_ _6818_/D _7243_/CLK _6818_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet763_430 net763_431/I _6740_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_441 net763_441/I _6724_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6749_ _6749_/D _7260_/RN _6749_/CLK _6749_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_109_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5080_ _4977_/Z _4981_/Z _5083_/B _5080_/C _5412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_4100_ hold4/Z hold17/Z hold21/Z hold22/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_110_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4031_ _4031_/A1 _4031_/A2 _4031_/A3 _4031_/A4 _4031_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_77_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5982_ _6964_/Q _5979_/Z _5981_/Z _6932_/Q _5980_/Z _7068_/Q _5983_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_4933_ _4933_/A1 _4930_/Z _4933_/A3 _4933_/A4 _4939_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_80_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_13 hold56/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4864_ _4624_/Z _4844_/Z _5156_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_61_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6603_ _5299_/C _6833_/Q _6826_/Q _6603_/A4 _6604_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_4795_ _5328_/A1 _4699_/Z _5394_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_119_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3815_ _3552_/Z _3617_/Z _4188_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_146_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3746_ _7185_/Q _3959_/C1 _3901_/A2 _6983_/Q _3747_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_20_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6534_ _6727_/Q _6253_/Z _6296_/Z _6715_/Q _6542_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6465_ _6465_/A1 _6465_/A2 _6465_/A3 _6464_/Z _6465_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5416_ _5416_/I _5417_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3677_ input49/Z _4210_/S _5521_/A2 _3904_/A2 _3947_/A2 _7099_/Q _3687_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_161_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet713_360 net713_361/I _6850_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_371 net713_385/I _6839_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6396_ _7064_/Q _6257_/Z _6408_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5347_ _5347_/A1 _5347_/A2 _5347_/A3 _5347_/A4 _5348_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xoutput175 _3366_/ZN mgmt_gpio_oeb[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput186 _3356_/ZN mgmt_gpio_oeb[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xnet713_393 net713_394/I _6781_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_382 net763_447/I _6800_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput197 _3346_/ZN mgmt_gpio_oeb[33] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5278_ _4554_/Z _4683_/Z _5364_/B _5278_/C _5279_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_87_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4229_ _4244_/S _4194_/Z _6652_/A2 _3542_/Z hold18/Z _4245_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_102_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7017_ _7017_/D _7260_/RN _7017_/CLK _7017_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_101_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_137__1359_ net563_220/I net713_385/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_28_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4580_ _4604_/A2 _4604_/A3 _4580_/B _4580_/C _5435_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_128_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3600_ _7181_/Q _3945_/A2 _3945_/B1 _7093_/Q _3601_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xinput22 mask_rev_in[26] input22/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput11 mask_rev_in[16] input11/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput44 mgmt_gpio_in[17] input44/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput55 mgmt_gpio_in[27] input55/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3531_ _3505_/Z _3529_/Z _3934_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_7_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput33 mask_rev_in[7] input33/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput66 mgmt_gpio_in[37] _7309_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_171_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput88 spimemio_flash_io1_oeb input88/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold828 _4216_/Z _6748_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold817 _6712_/Q hold817/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold806 _4324_/Z _6822_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput77 ser_tx input77/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput99 wb_adr_i[13] input99/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3462_ _3465_/A3 _6665_/Q input58/Z _3462_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_171_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6250_ _7236_/Q _6484_/A2 _6311_/A3 _6302_/A4 _6250_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold839 _4233_/Z _6756_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3393_ _3393_/I _6580_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5201_ _5464_/A1 _5438_/C _4557_/Z _4604_/Z _5201_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_143_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6181_ _6169_/Z _6181_/A2 _6181_/A3 _6180_/Z _6181_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_42_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5132_ _5205_/A1 _5132_/A2 _5293_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_97_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_816 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5063_ _5063_/I _5330_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4014_ _7237_/Q _6484_/A2 _6311_/A3 _6285_/A2 _4014_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_37_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5965_ _7231_/Q _7228_/Q _7227_/Q _6210_/C _5965_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_34_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4916_ _5324_/A1 _5263_/A4 _5056_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5896_ _5896_/I0 _6746_/Q _5957_/S _5910_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4847_ _4530_/I _5399_/A2 _5104_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_166_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4778_ _4468_/Z _4782_/A1 _5302_/B _4778_/A4 _4778_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_174_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3729_ _7201_/Q _3955_/A2 _3747_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_6517_ _6706_/Q _6254_/Z _6273_/Z _6822_/Q _6521_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_162_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6448_ _6744_/Q _7255_/Q _6448_/B _6449_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_164_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6379_ _7137_/Q _6253_/Z _6297_/Z _6701_/Q _6380_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_138_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_40__1359_ net413_53/I net413_61/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_120__1359_ net613_293/I net413_91/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_19_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5750_ _4103_/I hold900/Z _5757_/S _5750_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4701_ _4687_/Z _5097_/A1 _4699_/Z _5092_/A1 _5459_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_5681_ hold218/Z hold15/Z _5682_/S _5681_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4632_ _4441_/B _4501_/B _4460_/B _4436_/B _5293_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_30_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4563_ _4402_/B _4483_/B _4026_/B _4026_/C _5364_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold603 _5542_/Z _6910_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_118_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4494_ _5281_/C _4884_/A1 _4494_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_4
Xmax_cap344 _4064_/S _6657_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_8
X_7282_ _7282_/D _6636_/Z _7304_/CLK _7282_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_156_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6302_ _7236_/Q _6311_/A3 _6302_/A3 _6302_/A4 _6302_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold614 _7128_/Q hold614/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold636 _3496_/Z _3497_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold625 _5561_/Z _6927_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3514_ _6979_/Q _3923_/A2 _3592_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3445_ _3452_/S _7291_/Q _3450_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_171_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6233_ _7236_/Q _7237_/Q _6533_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold647 _5869_/Z _7200_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold669 _4247_/Z _6763_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold658 _6843_/Q hold658/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap355 _7193_/RN _7219_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_170_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6164_ _7027_/Q wire348/Z _6211_/B1 _6995_/Q _6176_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3376_ hold77/I _3376_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5115_ _5113_/Z _5403_/C _5233_/A1 _5156_/B _5115_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6095_ hold72/I _5979_/Z _5996_/Z hold68/I _6095_/C _6101_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_5046_ _5044_/Z _5433_/A1 _5047_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_111_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6997_ _6997_/D _7260_/RN _6997_/CLK _6997_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5948_ _7235_/Q _7234_/Q _6300_/A2 _6484_/A3 _5948_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_129_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5879_ hold52/Z hold612/Z _5883_/S _5879_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet463_107 net463_147/I _7118_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet463_129 net613_267/I _7096_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet463_118 net813_467/I _7107_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6920_ _6920_/D _7258_/RN _6920_/CLK _6920_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_90_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6851_ _6851_/D _7297_/RN _6851_/CLK _6851_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5802_ hold2/Z _7141_/Q hold7/Z hold8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3994_ _3994_/A1 _6902_/Q input67/Z _3994_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_6782_ _6782_/D _7260_/RN _6782_/CLK _6782_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5733_ hold271/Z hold908/Z _5739_/S _5733_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5664_ hold156/Z hold2/Z _5664_/S _5664_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4615_ _4422_/Z _4568_/Z _4614_/Z _4483_/B _5151_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5595_ hold271/Z hold955/Z hold12/Z _6957_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4546_ _4835_/A2 _4456_/B _3402_/I _3401_/I _4546_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_117_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold411 _5499_/Z _6879_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold400 _4112_/Z _6670_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold422 _7156_/Q hold422/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold444 _7178_/Q hold444/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold433 _4125_/Z _6679_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold477 _7062_/Q hold477/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4477_ _4692_/B _4692_/C _4786_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_89_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7265_ _7265_/D _7265_/CLK _7265_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold455 _5702_/Z _7052_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold466 _4150_/Z _6698_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3428_ _3427_/Z _6734_/Q _3428_/A3 _3428_/B _7301_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
Xhold488 _7130_/Q hold488/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7196_ _7196_/D _7221_/RN _7196_/CLK _7196_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold499 _5508_/Z _6887_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6216_ _6723_/Q _5987_/Z _6015_/Z _6842_/Q _6217_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_131_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3359_ _7081_/Q _3359_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6147_ _6147_/A1 _6147_/A2 _6147_/A3 _6147_/A4 _6147_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_58_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6078_ _6078_/A1 _6078_/A2 _6078_/A3 _6078_/A4 _6078_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_86_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5029_ _5353_/A1 _5439_/B2 _5029_/B _5354_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_2627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4400_ _4412_/A1 _4399_/Z _4491_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_157_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5380_ _4568_/Z _4892_/B _4821_/Z _4675_/Z _5380_/C _5381_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_126_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4331_ hold271/Z hold825/Z _4331_/S _4331_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7050_ _7050_/D _7258_/RN _7050_/CLK _7050_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4262_ _4227_/S _3994_/Z hold18/Z _4270_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_140_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6001_ _7028_/Q _5999_/Z _6000_/Z _7126_/Q _6008_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4193_ hold737/Z hold271/Z _4193_/S _4193_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6903_ _6903_/D _7219_/RN _6903_/CLK _6903_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_70_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6834_ _6834_/D _7279_/RN _7279_/CLK _6834_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_50_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3977_ _6661_/Q _3973_/Z _3977_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6765_ _6765_/D _7193_/RN _6765_/CLK _6765_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_11_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5716_ hold29/Z hold294/Z _5718_/S _5716_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6696_ _6696_/D _7193_/RN _6696_/CLK _6696_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_164_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5647_ _5647_/A1 hold18/Z hold33/Z hold135/Z _5647_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_163_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5578_ hold128/Z hold86/Z hold23/Z _6942_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4529_ _5420_/A2 _3401_/I _4530_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold252 _6991_/Q hold252/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold230 _6777_/Q hold230/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold241 _5697_/Z _7048_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_160_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold285 _5717_/Z _7066_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold274 _4105_/Z hold274/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold296 _7169_/Q hold296/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7248_ _7248_/D _7260_/RN _7260_/CLK _7248_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold263 _4127_/Z _6681_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_46_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7179_ _7179_/D _7221_/RN _7179_/CLK _7179_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_3103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7238__362 _7238_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_3169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 mask_rev_in[14] input9/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4880_ _4880_/A1 _4877_/Z _4879_/Z _5167_/B _4880_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3900_ _6728_/Q _4191_/A1 _3919_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_32_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3831_ _3537_/Z _3578_/Z _6611_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_32_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3762_ _3761_/Z hold991/Z _3899_/S _6871_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6550_ _6854_/Q _6241_/Z _6251_/Z _6825_/Q _6268_/Z _6800_/Q _6553_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_186_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5501_ hold110/Z hold52/Z _5502_/S _5501_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6481_ _7213_/Q _6256_/Z _6263_/Z _6939_/Q _6493_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3693_ _7000_/Q _5638_/A1 _3724_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5432_ _5432_/A1 _5189_/Z _5209_/Z _4985_/Z _5432_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_134_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5363_ _5363_/A1 _5342_/I _5363_/B1 _5396_/A1 _5383_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_127_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput335 _7269_/Q wb_dat_o[31] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput302 _3619_/Z serial_data_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput324 _6796_/Q wb_dat_o[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput313 _6804_/Q wb_dat_o[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4314_ _4313_/Z _6832_/Q _6577_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7102_ _7102_/D _7219_/RN _7102_/CLK _7102_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5294_ _5294_/A1 _5366_/A2 _5296_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_114_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4245_ _4244_/Z hold693/Z _4245_/S _4245_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7033_ _7033_/D _7260_/RN _7033_/CLK _7033_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_132_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4176_ _3535_/Z _3552_/Z _5520_/C _4178_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_28_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6817_ _6817_/D _7243_/CLK _6817_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet763_431 net763_431/I _6739_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6748_ _6748_/D _7260_/RN _6748_/CLK _6748_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet763_420 net763_426/I _6754_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet763_442 net763_443/I _6723_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_17__1359_ net413_58/I net813_472/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6679_ _6679_/D _7297_/RN _6679_/CLK _6679_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_164_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_174_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4030_ _4386_/A3 _4386_/A4 _4391_/A1 _4391_/A2 _4030_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_37_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5981_ _6210_/C _6021_/A2 _6210_/A2 _7227_/Q _5981_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4932_ _5258_/B2 _5056_/C _5442_/A2 _5248_/A2 _4933_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_80_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6602_ _6602_/I0 _7277_/Q _6602_/S _7277_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_14 user_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_4863_ _4624_/Z _4833_/Z _4865_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4794_ _4673_/Z _4793_/Z _5452_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3814_ _6729_/Q _4191_/A1 _3876_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_158_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3745_ _7209_/Q _3960_/A2 _5665_/A1 _7023_/Q _3747_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6533_ _6838_/Q _6533_/A2 _6533_/A3 _6533_/A4 _6540_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6464_ _6464_/A1 _6464_/A2 _6464_/A3 _6464_/A4 _6464_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_119_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5415_ _4703_/Z _4982_/Z _5415_/B1 _5083_/C _5416_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_133_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3676_ _7115_/Q _3917_/A2 _5683_/A1 _7041_/Q _3687_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6395_ _7254_/Q _6395_/I1 _6558_/S _7254_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet713_372 net813_485/I _6838_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_361 net713_361/I _6849_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5346_ _5393_/A2 _5346_/A2 _5346_/B _5347_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xoutput176 _3365_/ZN mgmt_gpio_oeb[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_115_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet713_394 net713_394/I _6780_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_383 net713_383/I _6799_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput198 _3345_/ZN mgmt_gpio_oeb[34] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput187 _3355_/ZN mgmt_gpio_oeb[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5277_ _5277_/I _5421_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4228_ _4227_/Z hold691/Z _4228_/S _4228_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7016_ hold63/Z _7260_/RN _7016_/CLK _7016_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_130_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4159_ _4103_/I hold791/Z _4160_/S _4159_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_4__1359_ net713_387/I net813_475/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_169_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 mask_rev_in[17] input12/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput45 mgmt_gpio_in[18] input45/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3530_ _3507_/Z _3529_/Z _5656_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xinput23 mask_rev_in[27] input23/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput34 mask_rev_in[8] input34/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold807 _6758_/Q hold807/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput56 mgmt_gpio_in[28] input56/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput89 spimemio_flash_io2_do input89/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput78 spi_csb input78/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xhold818 _4168_/Z _6712_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput67 mgmt_gpio_in[3] input67/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3461_ _6665_/Q _6663_/Q _6730_/Q _3463_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_170_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_63__1359_ clkbuf_4_15_0__1359_/Z net513_182/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold829 _6921_/Q hold829/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5200_ _5205_/A1 _5291_/B _5200_/B1 _5346_/A2 _5200_/C _5354_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_112_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6180_ _6180_/A1 _6180_/A2 _6180_/A3 _6180_/A4 _6180_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3392_ _6891_/Q _3903_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5131_ _5172_/A1 _5291_/A2 _5165_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_35_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5062_ _4699_/Z _5330_/B2 _5062_/B _5063_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_112_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4013_ _5942_/S _7235_/Q _6311_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_96_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5964_ _6117_/A4 _6014_/A2 _6210_/A2 _7229_/Q _5964_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4915_ _4496_/Z _4495_/Z _5263_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5895_ _6746_/Q _6744_/Q _5901_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_34_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4846_ _4846_/A1 _4846_/A2 _5090_/A2 _4849_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_20_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ _4782_/A1 _5099_/A1 _5456_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6516_ _6512_/Z _6516_/A2 _6516_/A3 _6516_/A4 _6516_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_146_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3728_ input46/Z _4210_/S _3739_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3659_ _7091_/Q _3945_/B1 _3927_/B1 _7065_/Q _3663_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6447_ _6440_/Z _6446_/Z _6447_/B1 _6286_/Z _6555_/C _6448_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_161_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6378_ _7071_/Q _6248_/Z _6293_/Z _7153_/Q _6380_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_115_771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5329_ _5359_/A1 _4716_/Z _5445_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_103_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4700_ _5420_/A2 _5129_/A3 _5051_/S _3401_/I _4700_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_1180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5680_ hold518/Z hold29/Z _5682_/S _5680_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4631_ _4868_/A1 _4524_/Z _5403_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_147_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4562_ _4422_/Z _4483_/B _5291_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_116_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7281_ _7281_/D _6635_/Z _7303_/CLK _7281_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
Xhold615 _5788_/Z _7128_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4493_ _4808_/A2 _4492_/Z _5240_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3513_ _3509_/Z _3512_/Z _3923_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold604 _7088_/Q hold604/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6301_ _7052_/Q _6299_/Z _6300_/Z _7102_/Q _6306_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold626 _7013_/Q hold626/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3444_ _3442_/B _3452_/S _3449_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_170_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold648 _7184_/Q hold648/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap345 _4064_/S _6652_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xhold637 hold637/I hold637/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap356 input75/Z _7193_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold659 _4339_/Z _6843_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6232_ _7250_/Q _6232_/I1 _6558_/S _7250_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6163_ _7125_/Q _5969_/Z _6176_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3375_ _6959_/Q _3375_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _4762_/Z _4867_/Z _5403_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_84_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6094_ _6094_/I _6095_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5045_ _5214_/A2 _5389_/A1 _5172_/B _5045_/C _5433_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_97_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6996_ _6996_/D _7260_/RN _6996_/CLK _6996_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_5947_ _6285_/A2 _7237_/Q _6484_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_41_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5878_ hold86/Z hold372/Z _5883_/S _5878_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4829_ _4673_/Z _4683_/Z _5276_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_21_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_13_0__1359_ clkbuf_0__1359_/Z clkbuf_4_13_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_72_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold1 hold1/I hold1/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_95_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet463_108 net513_152/I _7117_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet463_119 _4073__14/I _7106_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6850_ _6850_/D _7193_/RN _6850_/CLK _6850_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_90_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6781_ hold82/Z _7238_/RN _6781_/CLK hold81/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5801_ hold15/Z hold25/Z hold7/Z _7140_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3993_ _3994_/A1 hold773/Z input67/Z _4064_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_50_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5732_ hold113/Z hold389/Z _5739_/S _5732_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5663_ hold188/Z hold15/Z _5664_/S _5663_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4614_ _4441_/B _4467_/B _4460_/B _4501_/B _4614_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5594_ hold113/Z hold376/Z hold12/Z _6956_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4545_ _4454_/Z _4878_/A2 _5172_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_116_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold401 _7142_/Q hold401/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold434 _7132_/Q hold434/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold423 _5819_/Z _7156_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold445 _5844_/Z _7178_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold412 _7030_/Q hold412/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold478 _5713_/Z _7062_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4476_ _4853_/A1 _4481_/A2 _5288_/B _4692_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xhold456 _7100_/Q hold456/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7264_ _7264_/D _7265_/CLK _7264_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold467 _6686_/Q hold467/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3427_ _6733_/Q _6732_/Q _6730_/Q _3427_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
Xhold489 _5790_/Z _7130_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7195_ _7195_/D _7219_/RN _7195_/CLK _7195_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6215_ _6713_/Q _6002_/Z _6003_/Z _6715_/Q _6217_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3358_ _7089_/Q _3358_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6146_ _7124_/Q _5969_/Z _6146_/B _6147_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6077_ _7055_/Q _5924_/Z _5988_/Z _6983_/Q _6168_/C _6078_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_85_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5028_ _5023_/Z _5476_/A1 _5027_/I _5028_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XTAP_2617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6979_ _6979_/D _7258_/RN _6979_/CLK _6979_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_16_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold990 _6873_/Q hold990/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_135_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4330_ _4103_/I hold751/Z _4331_/S _4330_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4261_ hold2/Z hold95/Z _4261_/S hold96/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6000_ _6015_/A3 _6211_/B1 _7231_/Q _7228_/Q _6000_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_79_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4192_ hold687/Z _4103_/I _4193_/S _4192_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6902_ _6902_/D _7219_/RN _6902_/CLK _6902_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6833_ _6833_/D _7279_/RN _7279_/CLK _6833_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_36_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3976_ _3975_/Z _6662_/Q _3988_/S _6662_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ _6764_/D input75/Z _6764_/CLK _6764_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6695_ _6695_/D _7193_/RN _6695_/CLK _6695_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5715_ hold62/Z hold244/Z _5718_/S _5715_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5646_ hold149/Z hold2/Z hold19/Z _7003_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold220 _7133_/Q hold220/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_117_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5577_ hold616/Z hold271/Z hold23/Z _6941_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4528_ _5359_/A1 _4524_/Z _4472_/B _4501_/B _4528_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold242 _7213_/Q hold242/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold253 _5633_/Z _6991_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold231 _4263_/Z _6777_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4459_ _4555_/B _5270_/A1 _5281_/C _4459_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_7247_ _7247_/D _7260_/RN _7260_/CLK _7247_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_105_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold286 _7031_/Q hold286/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_85_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold264 _7023_/Q hold264/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold275 _5527_/Z _6900_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold297 _5834_/Z _7169_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7178_ _7178_/D _7219_/RN _7178_/CLK _7178_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_3104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6129_ hold54/I _5964_/Z _6014_/Z hold58/I _6000_/Z _7131_/Q _6134_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_3137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3830_ _3529_/Z _3540_/Z _3942_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3761_ _6567_/I0 _6870_/Q _3898_/S _3761_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5500_ hold260/Z hold86/Z _5502_/S _5500_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6480_ _7221_/Q _6274_/Z _6285_/Z _7197_/Q _7181_/Q _6254_/Z _6493_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3692_ _3505_/Z _3527_/Z _3916_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_145_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5431_ _5431_/A1 _5299_/C _5431_/B _5431_/C _6863_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_65_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5362_ _5362_/A1 _5362_/A2 _5362_/A3 _5363_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_126_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput314 _6805_/Q wb_dat_o[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput303 _4070_/Z serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput325 _6797_/Q wb_dat_o[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4313_ _6834_/Q _6835_/Q _6836_/Q _4313_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_154_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7101_ _7101_/D _7221_/RN _7101_/CLK _7101_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xoutput336 _6814_/Q wb_dat_o[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_142_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5293_ _5293_/A1 _5295_/A1 _5293_/B _5366_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_113_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7032_ _7032_/D _7297_/RN _7032_/CLK _7032_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4244_ hold169/Z hold2/Z _4244_/S _4244_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4175_ hold271/Z hold717/Z _4175_/S _4175_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6816_ _6816_/D _7243_/CLK _6816_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6747_ _6747_/D _7238_/RN _6747_/CLK _6747_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_177_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xnet763_432 net763_435/I _6738_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet763_421 net813_491/I _6753_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_410 net763_448/I _6764_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3959_ _7012_/Q _5656_/A1 _3959_/B1 _6666_/Q _3959_/C1 _7182_/Q _3961_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_167_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6678_ _6678_/D input75/Z _6678_/CLK _6678_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xnet763_443 net763_443/I _6722_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5629_ _3509_/Z _5520_/C _5839_/A3 _5857_/A3 _5637_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_145_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_1_0__1359_ clkbuf_0__1359_/Z net563_220/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_2299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5980_ _6015_/A3 _6210_/C _7231_/Q _7228_/Q _5980_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xclkbuf_leaf_23__1359_ net613_253/I net513_188/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_103__1359_ clkbuf_4_5_0__1359_/Z net713_394/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_24_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4931_ _5389_/A2 _5056_/C _5442_/A2 _5248_/A2 _4933_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xclkbuf_leaf_86__1359_ clkbuf_4_13_0__1359_/Z net563_230/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4862_ _4862_/A1 _4859_/Z _4861_/Z _4819_/Z _4865_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_6601_ _6601_/A1 _4313_/Z _6601_/B _6602_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_3813_ _3552_/Z _3680_/Z _4191_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_159_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4793_ _4534_/Z _5312_/A1 _4491_/B _4402_/B _4793_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XANTENNA_15 user_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_3744_ _6959_/Q _3957_/A2 _3927_/A2 _6701_/Q _3747_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6532_ _6697_/Q _6282_/Z _6542_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_174_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6463_ _6938_/Q _6263_/Z _6266_/Z _7018_/Q _6464_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3675_ _7179_/Q _3945_/A2 _5758_/A1 _7107_/Q _3687_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5414_ _4997_/B _5414_/A2 _4659_/Z _5414_/B _5418_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_134_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6394_ _6394_/I _6395_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_362 net713_383/I _6848_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5345_ _5389_/C _5345_/A2 _5356_/B _5389_/A2 _5346_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xoutput177 _3364_/ZN mgmt_gpio_oeb[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_115_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet713_373 net813_485/I _6837_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_384 net713_385/I _6790_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_395 net763_424/I _6779_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput199 _4052_/ZN mgmt_gpio_oeb[35] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_141_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput188 _3354_/ZN mgmt_gpio_oeb[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5276_ _5276_/A1 _5276_/A2 _5291_/C _5276_/C _5277_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_101_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7015_ hold57/Z _7238_/RN _7015_/CLK hold56/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_4227_ hold440/Z hold2/Z _4227_/S _4227_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4158_ _5520_/C _3552_/Z _5513_/A3 _5839_/A3 _4160_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_83_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4089_ _6907_/Q input39/Z _4089_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_43_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_466 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput13 mask_rev_in[18] input13/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput46 mgmt_gpio_in[19] input46/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput24 mask_rev_in[28] input24/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput35 mask_rev_in[9] input35/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput57 mgmt_gpio_in[29] input57/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xhold808 _4237_/Z _6758_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_128_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput68 mgmt_gpio_in[5] input68/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xhold819 _7296_/Q hold819/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xinput79 spi_enabled _4055_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_171_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3460_ hold270/Z input58/Z _3460_/S _7284_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3391_ _7222_/Q _5894_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5130_ _5240_/B _5328_/A2 _5130_/B1 _5130_/B2 _5321_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5061_ _4699_/Z _4936_/I _5061_/B _5410_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_69_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4012_ _6302_/A4 _7236_/Q _6282_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5963_ _6021_/A2 _7227_/Q _6117_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_25_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4914_ _4497_/Z _4494_/Z _5442_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_52_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5894_ _5894_/A1 _5894_/A2 _5894_/A3 _4019_/B _6746_/Q _7222_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_4845_ _4596_/Z _4817_/Z _5090_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4776_ _4703_/Z _5236_/B _5121_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3727_ _3726_/Z _6872_/Q _3899_/S _6872_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6515_ _6845_/Q _6235_/Z _6237_/Z _6837_/Q _6516_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_180_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3658_ hold45/I _3951_/C1 _3924_/A2 _6969_/Q input25/Z _3954_/B1 _3688_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6446_ _6554_/A1 _6446_/A2 _6446_/A3 _6446_/A4 _6446_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_164_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6377_ _7201_/Q _6272_/Z _6282_/Z _7185_/Q _6296_/Z _7161_/Q _6384_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_121_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3589_ _3589_/A1 _3589_/A2 _3589_/A3 _3589_/A4 _3589_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_88_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5328_ _5328_/A1 _5328_/A2 _5481_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_115_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5259_ _5259_/A1 _5259_/A2 _5337_/A2 _5449_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_130_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_823 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_855 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_285 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4630_ _4367_/Z _4555_/B _5291_/C _5387_/A1 _5387_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4561_ _4556_/Z _4561_/A2 _5003_/A2 _4561_/B _4584_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_162_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6300_ _7234_/Q _6300_/A2 _6484_/A3 _5943_/S _6300_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_7280_ _7280_/D _6634_/Z _7303_/CLK hold4/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
X_4492_ _4402_/B _4026_/B _4026_/C _5312_/A1 _4492_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_116_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3512_ _3653_/A1 _3617_/A1 _3501_/Z _3492_/Z _3512_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold605 _5743_/Z _7088_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold627 _5658_/Z _7013_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold616 _6941_/Q hold616/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3443_ _3438_/S _3440_/S _3443_/A3 _3443_/A4 _3452_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_144_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold649 _5851_/Z _7184_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap357 _7210_/RN _7258_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold638 _4353_/Z _4355_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap346 _4225_/S _4227_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
X_6231_ _6231_/I _6232_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6162_ _7247_/Q _6162_/I1 _6558_/S _7247_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5113_ _5113_/A1 _5113_/A2 _5313_/A1 _5313_/A3 _5113_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_69_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3374_ _6967_/Q _3374_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ _7000_/Q _6021_/Z _6090_/Z _5924_/Z _6094_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5044_ _5044_/A1 _5386_/A1 _5044_/A3 _5432_/A1 _5044_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_57_339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6995_ _6995_/D _7258_/RN _6995_/CLK _6995_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5946_ _5950_/B1 _5945_/B _7236_/Q _7236_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5877_ hold271/Z hold938/Z _5883_/S _5877_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4828_ _5364_/B _4586_/Z _4784_/Z _4598_/Z _5414_/A2 _5421_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_182_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4759_ _4501_/B _4759_/A2 _4759_/A3 _4759_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_182_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6429_ hold42/I _6253_/Z _6296_/Z _7163_/Q _6434_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_161_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold2 hold2/I hold2/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_181_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet463_109 net463_109/I _7116_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3992_ _7298_/Q hold4/I _3995_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6780_ hold76/Z _7238_/RN _6780_/CLK hold75/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5800_ hold29/Z hold42/Z hold7/Z _7139_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5731_ _3523_/Z _3537_/Z hold6/Z _5739_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_95_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5662_ hold555/Z hold29/Z _5664_/S _5662_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4613_ _5288_/B _5281_/C _4436_/B _4472_/B _5291_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5593_ hold6/Z _3523_/Z hold38/I hold11/Z hold12/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_163_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4544_ _4454_/Z _4456_/B _5276_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold402 _5804_/Z _7142_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_143_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold435 _5792_/Z _7132_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7263_ _7263_/D _7269_/CLK _7263_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold413 _5677_/Z _7030_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold424 _6878_/Q hold424/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4475_ _5288_/C _4454_/Z _4367_/Z _4501_/B _4692_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_116_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold457 _5756_/Z _7100_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold446 _7092_/Q hold446/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6214_ _6825_/Q _5988_/Z _6019_/Z _6854_/Q _6217_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold468 _4133_/Z _6686_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3426_ _6733_/Q _6732_/Q _6730_/Q _3434_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_98_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7194_ _7194_/D _7219_/RN _7194_/CLK _7194_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xhold479 _7040_/Q hold479/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3357_ _7097_/Q _3357_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6145_ hold26/I _5958_/Z _5994_/I hold25/I _6147_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_85_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6076_ _7089_/Q _6002_/Z _6015_/Z _7007_/Q _6076_/C _6078_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_97_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5027_ _5027_/I _5200_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6978_ _6978_/D _7258_/RN _6978_/CLK _6978_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_41_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5929_ _5925_/Z _7231_/Q _6168_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_55_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold980 _7061_/Q hold980/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold991 _6871_/Q hold991/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_88_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4260_ hold15/Z hold104/Z _4261_/S _4260_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4191_ _4191_/A1 hold18/Z _4193_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_68_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6901_ _6901_/D _7237_/RN _6901_/CLK _6901_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_82_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6832_ _6832_/D _7279_/RN _7279_/CLK _6832_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_165_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3975_ _3483_/Z _3975_/I1 _3975_/S _3975_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6763_ _6763_/D input75/Z _6763_/CLK _6763_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_176_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5714_ hold52/Z hold362/Z _5718_/S _5714_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6694_ _6694_/D _7193_/RN _6694_/CLK _6694_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_31_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5645_ _7002_/Q hold15/Z hold19/Z hold20/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5576_ hold121/Z hold113/Z hold23/Z _6940_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold210 _5781_/Z _7122_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4527_ _5359_/A1 _4997_/C _5243_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold221 _5793_/Z _7133_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold243 _5883_/Z _7213_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold232 _7157_/Q hold232/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4458_ _4467_/A1 _4555_/B _4736_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7246_ _7246_/D _7258_/RN _7260_/CLK _7246_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold287 _5678_/Z _7031_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_85_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold265 _5669_/Z _7023_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold276 _7161_/Q hold276/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold254 _6999_/Q hold254/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3409_ _6665_/Q _6664_/Q _6663_/Q _3409_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_172_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold298 _7074_/Q hold298/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7177_ _7177_/D _7219_/RN _7177_/CLK _7177_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4389_ _4427_/A2 _4427_/A3 _4485_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_58_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6128_ _7065_/Q _5985_/Z _5997_/Z _7099_/Q _6128_/C _6134_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6059_ _7030_/Q _5999_/Z _6014_/Z _6958_/Q _6000_/Z _7128_/Q _6061_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_3149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet513_190 net563_215/I _7035_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_437 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3760_ _3760_/A1 _3739_/Z _3759_/Z _6567_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_60_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5430_ _5268_/Z _5430_/A2 _5428_/Z _5429_/Z _5431_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3691_ _3690_/Z hold990/Z _3899_/S _6873_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5361_ _5361_/A1 _5209_/Z _5362_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_114_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput326 _6798_/Q wb_dat_o[23] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_58_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput315 _6806_/Q wb_dat_o[13] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput304 _4069_/Z serial_resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5292_ _5423_/A2 _5292_/A2 _5292_/A3 _5292_/A4 _5294_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xclkbuf_leaf_46__1359_ net663_324/I _4073__21/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7100_ _7100_/D _7221_/RN _7100_/CLK _7100_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xoutput337 _6815_/Q wb_dat_o[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_126__1359_ _4073__15/I net813_467/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_5_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4312_ _6571_/I0 _6818_/Q _4312_/S _6818_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4243_ _4242_/Z hold753/Z _4245_/S _4243_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7031_ _7031_/D _7260_/RN _7031_/CLK _7031_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_45_1041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4174_ _4103_/I hold650/Z _4175_/S _4174_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6815_ _6815_/D _7243_/CLK _6815_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6746_ _6746_/D _7237_/RN _4067_/I1 _6746_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_51_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet763_433 net763_435/I _6737_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_422 net763_422/I _6752_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet763_411 net763_441/I _6763_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3958_ _3958_/A1 _3958_/A2 _3958_/A3 _3958_/A4 _3958_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_176_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6677_ _6677_/D _7297_/RN _6677_/CLK _6677_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3889_ _3889_/A1 _3889_/A2 _3889_/A3 _3889_/A4 _3889_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xnet763_444 net763_445/I _6721_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5628_ hold2/Z hold140/Z _5628_/S _5628_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5559_ hold271/Z hold956/Z _5565_/S _5559_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7229_ _7229_/D _7258_/RN _7258_/CLK _7229_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_101_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_167_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4930_ _5129_/A3 _5325_/B _5051_/S _5170_/A2 _4930_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_17_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4861_ _4887_/A1 _4868_/A1 _5414_/A2 _5287_/B _4861_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_75_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6600_ _6834_/Q _6600_/A2 _6600_/B1 _6835_/Q _6836_/Q _6600_/C2 _6601_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_178_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3812_ _3552_/Z _3578_/Z _4146_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_16 hold271/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4792_ _4492_/Z _4534_/Z _5129_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_20_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3743_ _7063_/Q _3927_/B1 _3924_/A2 _6967_/Q _3743_/C _3759_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6531_ _6821_/Q _6262_/Z _6554_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_146_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6462_ _7172_/Q _5948_/Z _6261_/Z _6962_/Q _6464_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3674_ _3674_/A1 _3674_/A2 _3674_/A3 _3673_/Z _3674_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_173_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5413_ _5448_/A1 _5483_/A1 _5412_/Z _5414_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6393_ _6744_/Q _7253_/Q _6393_/B _6394_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5344_ _5438_/C _4666_/Z _5387_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_161_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet713_363 net713_383/I _6847_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_352 net413_55/I _6858_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput167 _4087_/Z debug_in VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xnet713_396 net763_426/I _6778_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_385 net713_385/I _6789_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_374 net713_385/I _6825_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput178 _3363_/ZN mgmt_gpio_oeb[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput189 _3353_/ZN mgmt_gpio_oeb[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5275_ _5376_/B2 _5468_/A2 _5275_/B _5423_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_99_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4226_ _4225_/Z hold588/Z _4228_/S _4226_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7014_ _7014_/D _7260_/RN _7014_/CLK _7014_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4157_ hold2/Z hold197/Z _4157_/S _4157_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4088_ _6906_/Q input70/Z _4088_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_37_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6729_ _6729_/D input75/Z _6729_/CLK _6729_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_165_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_92__1359_ net813_465/I net713_390/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_28_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput25 mask_rev_in[29] input25/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput14 mask_rev_in[19] input14/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput36 mgmt_gpio_in[0] input36/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_155_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput69 mgmt_gpio_in[6] input69/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput47 mgmt_gpio_in[1] input47/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput58 mgmt_gpio_in[2] input58/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xhold809 _6696_/Q hold809/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_182_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3390_ _7241_/Q _6011_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5060_ _5058_/Z _5060_/A2 _4928_/Z _5060_/A4 _5064_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_123_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4011_ _6282_/A2 _7232_/Q _6484_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_84_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5962_ _5984_/A1 _7230_/Q _6002_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_52_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4913_ _4376_/Z _5442_/A2 _4909_/Z _4927_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_5893_ _5945_/A1 _6746_/Q _5894_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4844_ _5287_/B _4456_/B _4530_/I _5051_/S _4844_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_33_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4775_ _4775_/A1 _4772_/Z _4773_/Z _4774_/Z _4781_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_158_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3726_ _4309_/I0 _6871_/Q _3898_/S _3726_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6514_ _6787_/Q _6263_/Z _6266_/Z _6843_/Q _6516_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3657_ _3657_/A1 _3657_/A2 _3657_/A3 _3657_/A4 _3657_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6445_ _7049_/Q _6241_/Z _6268_/Z hold49/I _6256_/Z _7211_/Q _6446_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6376_ _7113_/Q _6240_/Z _6376_/B _6384_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3588_ _7133_/Q _3930_/A2 _3941_/B1 _7173_/Q _3588_/C _3589_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_5327_ _4928_/Z _5326_/Z _5327_/A3 _5327_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_114_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5258_ _4890_/I _5258_/A2 _4972_/Z _5258_/B2 _5258_/C _5412_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_5189_ _5386_/A1 _5386_/A3 _5189_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_4209_ _4208_/Z hold600/Z _4211_/S _4209_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4560_ _5002_/A3 _5002_/A4 _5083_/B _5393_/B1 _4561_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_129_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4491_ _4491_/A1 _4491_/A2 _4491_/B _5312_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xhold617 _7126_/Q hold617/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold606 _7193_/Q hold606/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3511_ hold338/Z _3489_/I _5821_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3442_ _3991_/A1 _4042_/A3 _6733_/Q _3442_/B _3443_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
Xmax_cap347 _5323_/B _5442_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
Xhold628 _6859_/Q _3305_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6230_ _6555_/C _7249_/Q _6230_/B _6231_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
Xmax_cap358 _7238_/RN _7260_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
Xhold639 _4354_/Z _6853_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6161_ _6161_/I _6162_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3373_ _6975_/Q _3373_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5112_ _4614_/Z _5302_/B _4784_/Z _5230_/B _4716_/Z _5113_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XTAP_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6092_ _6092_/A1 _5991_/Z _6102_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _5385_/A1 _5043_/A2 _5043_/B _5432_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_111_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_wbbd_sck _7278_/Q clkbuf_0_wbbd_sck/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_81_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6994_ _6994_/D _7260_/RN _6994_/CLK _6994_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5945_ _5945_/A1 _6745_/Q _5945_/B _5950_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_22_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5876_ hold113/Z hold494/Z _5883_/S _5876_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4827_ _4586_/Z _4784_/Z _5223_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_119_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4758_ _5072_/A4 _4500_/Z _4958_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_175_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4689_ _4687_/Z _5092_/A1 _5302_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3709_ _7210_/Q _3960_/A2 _3955_/A2 _7202_/Q _7186_/Q _3959_/C1 _3724_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_4_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6428_ _7009_/Q _6243_/Z _6269_/Z _7033_/Q _6440_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_175_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6359_ _6359_/I _6360_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold3 hold3/I hold3/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_47_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3991_ _3991_/A1 _3412_/Z _3442_/B _3409_/Z _6730_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_62_343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5730_ hold888/Z hold271/Z _5730_/S _5730_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5661_ _7016_/Q hold62/Z _5664_/S hold63/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4612_ _4612_/A1 _4612_/A2 _5025_/B _4618_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_135_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5592_ hold91/Z hold2/Z _5592_/S hold92/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4543_ _5129_/A3 _5051_/S _4878_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_144_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold436 _7196_/Q hold436/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7262_ _7262_/D _7265_/CLK _7262_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xhold414 _6982_/Q hold414/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold403 _6688_/Q hold403/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold425 _5498_/Z _6878_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4474_ _5288_/C _4454_/Z _4367_/Z _4501_/B _4474_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_144_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold469 _7195_/Q hold469/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold447 _5747_/Z _7092_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold458 _7028_/Q hold458/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6213_ _6821_/Q _5979_/Z _5996_/Z _6709_/Q _6217_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3425_ _4041_/A3 _7302_/Q _3425_/S _7302_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7193_ _7193_/D _7193_/RN _7193_/CLK _7193_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_174_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3356_ _7105_/Q _3356_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6144_ _7066_/Q _5985_/Z _6000_/Z _7132_/Q _6144_/C _6147_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_58_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6075_ hold56/I _5971_/Z _6003_/Z _7161_/Q _6078_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xload_slew350 hold113/Z _4103_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_16
XFILLER_57_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5026_ _5471_/B2 _5291_/B _5002_/Z _5200_/B1 _5027_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2608 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6977_ hold55/Z _7260_/RN _6977_/CLK hold54/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_110_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5928_ _7231_/Q _5941_/A1 _5931_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_81_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5859_ hold271/Z hold972/Z _5865_/S _5859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold981 _5712_/Z _7061_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold970 _7175_/Q hold970/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_135_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold992 _6869_/Q hold992/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_49_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet563_250 net663_326/I _6975_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4190_ hold701/Z hold271/Z _4190_/S _4190_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6900_ _6900_/D _7238_/RN _6900_/CLK _6900_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_35_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6831_ _6831_/D _7279_/RN _7230_/CLK _6831_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_69__1359_ clkbuf_4_13_0__1359_/Z net513_194/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_62_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_149__1359_ net713_387/I net813_470/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3974_ _6661_/Q _6660_/Q _6659_/Q _3972_/Z _3975_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_165_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6762_ _6762_/D _7258_/RN _6762_/CLK _6762_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_189_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5713_ hold86/Z hold477/Z _5718_/S _5713_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6693_ _6693_/D _7219_/RN _6693_/CLK _6693_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_137_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5644_ hold41/Z hold29/Z hold19/Z _7001_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold200 _5565_/Z _6931_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5575_ _5575_/A1 hold18/Z hold23/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
Xhold211 _7146_/Q hold211/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4526_ _4472_/B _4501_/B _4460_/B _4436_/B _4997_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_145_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold233 _5820_/Z _7157_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold222 _7137_/Q hold222/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold244 _7064_/Q hold244/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold266 _6922_/Q hold266/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4457_ _4456_/B _5051_/S _4460_/B _4467_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7245_ _7245_/D _7258_/RN _7258_/CLK _7245_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold277 _5825_/Z _7161_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold255 _6876_/Q hold255/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_160_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold288 _7188_/Q hold288/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold299 _5726_/Z _7074_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3408_ _4436_/B _4467_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_12
X_7176_ _7176_/D _7210_/RN _7176_/CLK _7176_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4388_ _4388_/A1 _4388_/A2 input97/Z input96/Z _4427_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_113_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6127_ _6127_/A1 _6124_/Z _6127_/A3 _6127_/A4 _6127_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_112_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3339_ _3339_/I _3932_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6058_ _7062_/Q _5985_/Z _5997_/Z _7096_/Q _6061_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_58_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5009_ _5438_/C _5359_/A1 _5435_/A2 _5475_/A3 _5009_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_2416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet513_191 net513_191/I _7034_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_180 net513_188/I _7045_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3690_ _6569_/I0 _6872_/Q _3898_/S _3690_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5360_ _5045_/C _5393_/B1 _5360_/B _5360_/C _5361_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_127_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput305 _4086_/Z spi_sdi VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput316 _6807_/Q wb_dat_o[14] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5291_ _4542_/Z _5291_/A2 _5291_/B _5291_/C _5377_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_99_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput327 _7262_/Q wb_dat_o[24] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput338 _6816_/Q wb_dat_o[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_5_770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4311_ _6570_/I0 _6817_/Q _4312_/S _6817_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4242_ hold266/Z hold15/Z _4244_/S _4242_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7030_ _7030_/D _7258_/RN _7030_/CLK _7030_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_113_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_opt_1_0__1359_ clkbuf_4_8_0__1359_/Z clkbuf_opt_1_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_84_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4173_ _5821_/A3 _5513_/A3 _3537_/Z _5520_/C _4175_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_45_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6814_ _6814_/D _7243_/CLK _6814_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6745_ _6745_/D _7237_/RN _4067_/I1 _6745_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3957_ _6956_/Q _3957_/A2 _4289_/A1 _6799_/Q _3958_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xnet763_412 net763_413/I _6762_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_423 net763_424/I _6751_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_434 net763_435/I _6736_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6676_ _6676_/D _7297_/RN _6676_/CLK _6676_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3888_ _6989_/Q _3954_/A2 _3956_/A2 _7119_/Q _3889_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xnet763_445 net763_445/I _6720_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5627_ hold15/Z hold174/Z _5628_/S _5627_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5558_ hold113/Z hold594/Z _5565_/S _5558_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4509_ _5087_/A1 _5051_/S _5343_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_133_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5489_ _5489_/A1 _5489_/A2 _5472_/Z _5489_/A4 _5489_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_120_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7228_ _7228_/D _7258_/RN _7258_/CLK _7228_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_116_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7159_ _7159_/D _7219_/RN _7159_/CLK _7159_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_58_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_155_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_52__1359_ net663_324/I net513_159/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_183_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4860_ _5104_/A1 _4860_/A2 _5291_/C _5291_/B _5376_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_75_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3811_ _3509_/Z _3578_/Z _3925_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_177_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4791_ _5312_/A2 _5214_/A2 _5456_/A1 _5220_/B2 _4791_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XANTENNA_17 _4275_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6530_ _7259_/Q _6529_/Z _6558_/S _7259_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3742_ _3742_/I _3743_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6461_ _7220_/Q _6274_/Z _6285_/Z _7196_/Q _7180_/Q _6254_/Z _6464_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3673_ _3673_/A1 _3673_/A2 _3673_/A3 _3673_/A4 _3673_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5412_ _5412_/A1 _5412_/A2 _5412_/A3 _4984_/B _5412_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6392_ _6385_/Z _6391_/Z _6392_/B1 _6286_/Z _6744_/Q _6393_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_5343_ _5343_/A1 _5343_/A2 _5343_/B _5418_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xnet713_353 net413_71/I _6857_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput168 _6894_/Q irq[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xnet713_375 net713_385/I _6824_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_386 net763_437/I _6788_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_364 net413_55/I _6846_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput179 _3362_/ZN mgmt_gpio_oeb[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_141_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5274_ _5370_/A1 _5312_/A4 _5291_/C _5295_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_102_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet713_397 net413_88/I _6777_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7013_ _7013_/D _7260_/RN _7013_/CLK _7013_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4225_ hold99/Z hold15/Z _4225_/S _4225_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4156_ hold15/Z hold292/Z _4157_/S _4156_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4087_ input1/Z input36/Z _4087_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_36_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4989_ _5340_/A1 _5262_/A2 _5328_/A2 _5248_/A2 _4991_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_11_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6728_ _6728_/D input75/Z _6728_/CLK _6728_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_164_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6659_ _6659_/D _6614_/Z _4072_/B2 _6659_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_109_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_817 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2087 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput37 mgmt_gpio_in[10] input37/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 mask_rev_in[2] input26/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput15 mask_rev_in[1] input15/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput59 mgmt_gpio_in[30] input59/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput48 mgmt_gpio_in[20] input48/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4010_ _4010_/I _6744_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5961_ _6948_/Q _5958_/Z _5960_/Z _7150_/Q _5974_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4912_ _5464_/A1 _5443_/A1 _5193_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_179_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5892_ hold2/Z hold379/Z _5892_/S _5892_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4843_ _5287_/B _4784_/Z _5231_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_61_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4774_ _4782_/A1 _4510_/Z _5302_/B _4695_/Z _4774_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_146_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3725_ _3708_/Z _3724_/Z _3725_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_20_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6513_ _6809_/Q _6261_/Z _6268_/Z _6799_/Q _6265_/Z _6839_/Q _6516_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6444_ _7219_/Q _6274_/Z _6285_/Z _7195_/Q _7179_/Q _6254_/Z _6446_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3656_ _6679_/Q _3546_/Z _3945_/C2 _6687_/Q _3657_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_161_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6375_ _7129_/Q _6484_/A2 _6484_/A3 _6533_/A4 _6376_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_134_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3587_ _3587_/I _3588_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5326_ _5246_/Z _5442_/A4 _5442_/A2 _5056_/C _5326_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_103_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5257_ _5257_/A1 _5246_/Z _5257_/B _5257_/C _5264_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_130_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4208_ hold104/Z hold15/Z _4210_/S _4208_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5188_ _5243_/A1 _5043_/B _5205_/A1 _4650_/Z _5386_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4139_ hold271/Z hold727/Z _4139_/S _4139_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3510_ _3507_/Z _3509_/Z _5584_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_143_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4490_ _4491_/A1 _4491_/A2 _5092_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold618 _5786_/Z _7126_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold607 _5861_/Z _7193_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3441_ _6664_/Q _6663_/Q _6730_/Q _6665_/Q _3443_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_143_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold629 _3500_/Z hold629/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xmax_cap359 _7297_/RN _7238_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
X_6160_ _6555_/C _7246_/Q _6160_/B _6161_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_98_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3372_ _6983_/Q _3372_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5111_ _4614_/Z _4817_/Z _5111_/B _5111_/C _5113_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_33_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6091_ hold89/I wire348/Z _6211_/B1 hold83/I _6092_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5042_ _5385_/A1 _5389_/C _5439_/B1 _5393_/A1 _5044_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_97_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6993_ _6993_/D _7260_/RN _6993_/CLK _6993_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5944_ _6745_/Q _7235_/Q _7234_/Q _6300_/A2 _5945_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_41_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5875_ _3485_/Z _3523_/Z hold6/Z _5883_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_4826_ _4826_/A1 _5370_/B _4826_/A3 _4826_/B _4834_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_21_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4757_ _4757_/I _4766_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4688_ _5083_/B _5092_/A1 _5312_/A1 _5094_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_3708_ _3701_/Z _3708_/A2 _3708_/A3 _3707_/Z _3708_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_161_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3639_ hold25/I _3951_/A2 _5665_/A1 _7026_/Q _7018_/Q _5656_/A1 _3642_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6427_ _6945_/Q _6245_/Z _6288_/Z hold59/I _6440_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_115_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6358_ _7022_/Q _6235_/Z _6243_/Z _7006_/Q _6265_/Z _6998_/Q _6359_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5309_ _4699_/Z _5309_/A2 _5456_/A2 _5309_/B2 _5309_/C _5310_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6289_ _7182_/Q _6282_/Z _6288_/Z _7118_/Q _6307_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_130_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_166_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold4 hold4/I hold4/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_79_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3990_ _3990_/I _5896_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_23_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5660_ hold56/Z hold52/Z _5664_/S hold57/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4611_ _5287_/C _4565_/Z _5025_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_30_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5591_ hold26/Z hold15/Z _5592_/S hold27/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4542_ _5420_/A2 _5129_/A3 _5051_/S _4542_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_8_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7261_ _7261_/D _7279_/RN _7279_/CLK _7261_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_128_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold426 _7148_/Q hold426/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4473_ _4472_/B _4473_/A2 _4481_/A2 _4853_/A1 _4786_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
Xhold415 _5623_/Z _6982_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold404 _4135_/Z _6688_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3424_ _3465_/A4 _3465_/A3 _3971_/A1 _3442_/B _3425_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_171_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold437 _5864_/Z _7196_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold448 _7084_/Q hold448/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold459 _5675_/Z _7028_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6212_ _6212_/A1 _5991_/Z _6226_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_171_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_29__1359_ net663_304/I net663_316/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7192_ _7192_/D _7221_/RN _7192_/CLK _7192_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
Xclkbuf_leaf_109__1359_ clkbuf_4_5_0__1359_/Z net413_78/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3355_ _7113_/Q _3355_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6143_ _6143_/I _6144_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xload_slew351 _6744_/Q _6555_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
X_6074_ _7081_/Q _5996_/Z _6005_/Z _7039_/Q _6078_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_85_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5025_ _5439_/B2 _5200_/B1 _5025_/B _5476_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_100_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6976_ hold74/Z _7297_/RN _6976_/CLK hold73/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5927_ _5919_/Z _6014_/A2 _5941_/A1 _5925_/Z _5950_/A1 _7230_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_181_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5858_ _4103_/I hold898/Z _5865_/S _5858_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5789_ hold52/Z hold504/Z _5793_/S _5789_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4809_ _4809_/A1 _4805_/Z _4807_/Z _4808_/Z _4812_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_182_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_983 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold960 _7029_/Q hold960/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold971 _5841_/Z _7175_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold982 _7167_/Q hold982/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_115_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold993 _6868_/Q hold993/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_103_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet563_240 net663_329/I _6985_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_166_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet563_251 net563_251/I _6974_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6830_ _6833_/Q _7279_/RN _7279_/CLK _6830_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_23_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6761_ _6761_/D _7258_/RN _6761_/CLK _6761_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_189_861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3973_ _6660_/Q _6659_/Q _3972_/Z _3973_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_5712_ hold271/Z hold980/Z _5718_/S _5712_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6692_ _6692_/D _7219_/RN _6692_/CLK _6692_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_176_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5643_ hold575/Z hold62/Z hold19/Z _7000_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5574_ hold2/Z hold586/Z _5574_/S _5574_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold201 _6914_/Q hold201/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_141_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4525_ _5315_/A2 _4524_/Z _5130_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_102_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold234 _7109_/Q hold234/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold223 _7138_/Q hold223/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold212 _5808_/Z _7146_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4456_ _3401_/I _3402_/I _4456_/B _5051_/S _4481_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xhold267 _5555_/Z _6922_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold278 _7042_/Q hold278/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7244_ _7244_/D _7260_/RN _7260_/CLK _7244_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold256 _5495_/Z _6876_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold245 _5715_/Z _7064_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4387_ _4388_/A1 _4388_/A2 input97/Z input96/Z _4387_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3407_ _4460_/B _5281_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_12
Xhold289 _5855_/Z _7188_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7175_ _7175_/D _7219_/RN _7175_/CLK _7175_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3338_ _6927_/Q _6392_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_58_403 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6126_ hold47/I _5996_/Z _5999_/Z _7033_/Q _6969_/Q _5979_/Z _6127_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6057_ _6057_/A1 _6057_/A2 _6057_/A3 _6057_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_22_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5008_ _5438_/C _5359_/A1 _5439_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_2417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6959_ _6959_/D _7258_/RN _6959_/CLK _6959_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_139_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet513_170 net513_182/I _7055_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold790 _4141_/Z _6692_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet513_181 net413_70/I _7044_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_192 net663_329/I _7033_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_75__1359_ net613_299/I net613_287/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_39_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_0__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/Z _4075_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput306 _4081_/Z spimemio_flash_io0_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput317 _6808_/Q wb_dat_o[15] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5290_ _4422_/Z _4554_/Z _4614_/Z _4483_/B _5290_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4310_ _6569_/I0 _6816_/Q _4312_/S _6816_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput328 _7263_/Q wb_dat_o[25] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput339 _6817_/Q wb_dat_o[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_141_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4241_ _4240_/Z hold833/Z _4245_/S _4241_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4172_ hold711/Z hold271/Z _4172_/S _4172_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6813_ _6813_/D _7243_/CLK _6813_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6744_ _6744_/D _7258_/RN _4067_/I1 _6744_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_3956_ _7118_/Q _3956_/A2 _3956_/B1 _6712_/Q _3956_/C1 _6851_/Q _3958_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_149_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet763_402 net763_413/I _6772_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_413 net763_413/I _6761_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet763_424 net763_424/I _6750_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6675_ _6675_/D input75/Z _6675_/CLK _6675_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_164_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet763_435 net763_435/I _6735_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_446 net813_482/I _6719_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3887_ _6840_/Q _3925_/C2 _3956_/C1 _6852_/Q _3889_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5626_ hold29/Z hold516/Z _5628_/S _5626_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5557_ hold6/Z _3527_/Z _5839_/A3 _5857_/A3 _5565_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_3_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4508_ _4698_/B _5087_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_145_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _5374_/Z _5487_/Z _5489_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_117_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4439_ _4363_/Z _4369_/Z _4472_/B _4759_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_7227_ _7227_/D _7237_/RN _7258_/CLK _7227_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_104_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7158_ _7158_/D _7219_/RN _7158_/CLK _7158_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_7089_ _7089_/D _7221_/RN _7089_/CLK _7089_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XTAP_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6109_ _6101_/Z _6106_/Z _6109_/A3 _6109_/A4 _6109_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_46_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_296 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2770 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4790_ _4790_/A1 _5213_/C _4787_/Z _4789_/Z _4803_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_3810_ _3509_/Z hold630/Z _4301_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_158_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3741_ _7081_/Q _3923_/C1 _5575_/A1 hold65/I _3925_/A2 input6/Z _3742_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA_18 _7151_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_856 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6460_ _6994_/Q _6237_/Z _6247_/Z _7132_/Q _6460_/C _6465_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3672_ _7073_/Q _3943_/A2 _3941_/A2 _7163_/Q _3673_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5411_ _5248_/Z _5327_/Z _5411_/A3 _5483_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6391_ _6554_/A1 _6391_/A2 _6391_/A3 _6390_/Z _6391_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_63_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5342_ _5342_/I _5418_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet713_354 _4073__7/I _6856_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_807 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet713_376 net713_385/I _6823_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_387 net713_387/I _6787_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_365 net413_55/I _6845_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5273_ _4554_/Z _4683_/Z _5287_/B _5468_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_99_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet713_398 net763_429/I _6776_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xoutput169 _4088_/Z irq[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_7012_ _7012_/D _7260_/RN _7012_/CLK _7012_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_68_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4224_ _4223_/Z hold870/Z _4228_/S _4224_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4155_ hold29/Z hold310/Z _4157_/S _4155_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4086_ _4055_/S input63/Z _4086_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_24_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4988_ _5083_/C _4568_/Z _4659_/Z _4422_/Z _4988_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_183_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6727_ _6727_/D _7193_/RN _6727_/CLK _6727_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3939_ _6696_/Q _4146_/A1 _4359_/A1 _6857_/Q _3939_/C1 _6710_/Q _3940_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_176_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6658_ _6658_/D _4098_/Z _4072_/B2 _6658_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_180_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ hold15/Z hold173/Z hold39/Z _6970_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6589_ _6589_/A1 _4313_/Z _6589_/B _6590_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_178_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2099 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput27 mask_rev_in[30] input27/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput16 mask_rev_in[20] input16/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput38 mgmt_gpio_in[11] input38/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput49 mgmt_gpio_in[21] input49/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5960_ _7231_/Q wire348/Z _6021_/A2 _7227_/Q _5960_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_19_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4911_ _5464_/A1 _4903_/Z _5205_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5891_ hold15/Z hold430/Z _5892_/S _5891_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4842_ _5104_/A1 _4860_/A2 _4555_/C _5291_/C _4842_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_60_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4773_ _4782_/A1 _5302_/B _4695_/Z _4716_/Z _4773_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_159_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3724_ _3715_/Z _3724_/A2 _3724_/A3 _3723_/Z _3724_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6512_ _6512_/A1 _6512_/A2 _6512_/A3 _6511_/Z _6512_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_173_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3655_ _7219_/Q _3912_/A2 _3948_/C1 _7309_/I _3657_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6443_ hold43/I _6235_/Z _6261_/Z hold58/I _6443_/C _6446_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_162_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6374_ _7209_/Q _6256_/Z _6263_/Z _6935_/Q _6385_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_115_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3586_ _6931_/Q _3935_/A2 _3943_/A2 _7075_/Q _7157_/Q _3916_/A2 _3587_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5325_ _4716_/Z _5394_/A2 _5325_/B _5327_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5256_ _5262_/A2 _4902_/Z _5246_/Z _5257_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_114_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4207_ _4206_/Z hold868/Z _4211_/S _4207_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5187_ _5392_/B _5339_/A4 _5417_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_111_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4138_ _4103_/I hold652/Z _4139_/S _4138_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4069_ _7238_/Q hold88/I _6900_/Q _4069_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold608 _7168_/Q hold608/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_6_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3440_ input58/Z _3440_/I1 _3440_/S _7294_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold619 _6997_/Q hold619/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3371_ _6991_/Q _3371_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_152_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5110_ _4614_/Z _4817_/Z _5111_/C _5479_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6090_ _6210_/A2 _7056_/Q _6090_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XTAP_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ _5439_/B1 _5002_/Z _5041_/B _5386_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_98_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i clkbuf_0_wb_clk_i/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_53_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6992_ hold84/Z _7238_/RN _6992_/CLK hold83/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_179_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5943_ _5943_/I0 _5940_/Z _5943_/S _7235_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5874_ hold2/Z hold205/Z _5874_/S _5874_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4825_ _4539_/I _4683_/Z _4826_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_138_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4756_ _4510_/Z _4752_/Z _4757_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4687_ _5083_/B _4687_/A2 _4687_/A3 _4687_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_3707_ _3707_/A1 _3707_/A2 _3707_/A3 _3707_/A4 _3707_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_162_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3638_ _3638_/A1 _3638_/A2 _3638_/A3 _3638_/A4 _3638_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6426_ _6969_/Q _6262_/Z _6266_/Z _7017_/Q _6426_/C _6440_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_161_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3569_ _3515_/Z _3529_/Z _5674_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6357_ _6357_/A1 _6357_/A2 _6356_/Z _6357_/A4 _6357_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5308_ _5303_/Z _5308_/A2 _5221_/I _5480_/A1 _5308_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_88_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6288_ _7236_/Q _6302_/A3 _6533_/A4 _6302_/A4 _6288_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_103_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _5238_/Z _4801_/Z _5453_/A4 _5452_/A2 _5241_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_102_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_267 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_642 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_449 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_483 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold5 hold5/I hold5/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_90_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_194 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4610_ _5287_/C _4589_/Z _4612_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_129_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5590_ hold49/Z hold29/Z _5592_/S hold50/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4541_ _5278_/C _5279_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_4472_ _4464_/Z _4454_/Z _4472_/B _4764_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_117_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold427 _5810_/Z _7148_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold416 _6687_/Q hold416/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold405 _6988_/Q hold405/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7260_ _7260_/D _7260_/RN _7260_/CLK _7260_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3423_ _3422_/Z _7303_/Q _3988_/S _7303_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold449 _5738_/Z _7084_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold438 _7179_/Q hold438/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7191_ _7191_/D _7219_/RN _7191_/CLK _7191_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_6211_ _6846_/Q wire348/Z _6211_/B1 _6838_/Q _6212_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6142_ _6978_/Q _5964_/Z _5981_/Z _6938_/Q _6014_/Z _6962_/Q _6143_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3354_ _7121_/Q _3354_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6073_ _6073_/A1 _6073_/A2 _6073_/A3 _6073_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XTAP_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _4604_/Z _5475_/A3 _5200_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_57_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6975_ hold53/Z _7238_/RN _6975_/CLK _6975_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_41_507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5926_ _5950_/A1 _5925_/Z _5931_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_80_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5857_ _3485_/Z _5857_/A2 _5857_/A3 _5520_/C _5865_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_55_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5788_ hold86/Z hold614/Z _5793_/S _5788_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4808_ _4422_/Z _4808_/A2 _5312_/A1 _4666_/Z _4808_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_21_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4739_ _4739_/A1 _5106_/A1 _4738_/Z _4743_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_163_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6409_ _7170_/Q _5948_/Z _6261_/Z _6960_/Q _6266_/Z _7016_/Q _6411_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_122_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold972 _7191_/Q hold972/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold961 _5676_/Z _7029_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold950 _6683_/Q hold950/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold994 _6875_/Q hold994/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold983 _5832_/Z _7167_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_95_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_4_0__1359_ clkbuf_0__1359_/Z net613_293/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_leaf_35__1359_ net413_53/I _4073__30/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_115__1359_ net613_293/I net413_79/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_185_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_98__1359_ net813_465/I net663_329/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet563_230 net563_230/I _6995_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet563_241 net413_79/I _6984_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6760_ _6760_/D _7219_/RN _6760_/CLK _6760_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_91_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3972_ _7305_/Q _7304_/Q _7303_/Q _6658_/Q _3972_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_93_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5711_ hold113/Z hold393/Z _5718_/S _5711_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6691_ _6691_/D _7193_/RN _6691_/CLK _6691_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_176_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5642_ hold254/Z hold52/Z hold19/Z _6999_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5573_ hold15/Z hold450/Z _5574_/S _5573_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold202 _5546_/Z _6914_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_145_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4524_ _4460_/B _4436_/B _4524_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_116_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold235 _5766_/Z _7109_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold224 _6928_/Q hold224/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold213 _6984_/Q hold213/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4455_ _4555_/B _5270_/A1 _5170_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold268 _6912_/Q hold268/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold257 _6916_/Q hold257/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7243_ _7243_/D _7260_/RN _7243_/CLK _7243_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold246 _7032_/Q hold246/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4386_ input99/Z input98/Z _4386_/A3 _4386_/A4 _4427_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_160_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3406_ _4501_/B _5288_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
Xhold279 _5690_/Z _7042_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_113_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7174_ _7174_/D _7219_/RN _7174_/CLK _7174_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XTAP_551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6125_ _6945_/Q _5972_/Z _6021_/Z hold41/I _6127_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3337_ _3337_/I _4082_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6056_ _7070_/Q _5980_/Z _6005_/Z _7038_/Q _6057_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5007_ _5435_/A2 _5475_/A3 _5194_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2429 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6958_ _6958_/D _7258_/RN _6958_/CLK _6958_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_41_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5909_ _7226_/Q _5908_/Z _5910_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6889_ _6889_/D _7297_/RN _6889_/CLK _6889_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_14_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold780 _5560_/Z _6926_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold791 _6706_/Q hold791/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xnet513_160 net413_70/I _7065_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_182 net513_182/I _7043_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet513_171 _4073__39/I _7054_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_193 net563_221/I _7032_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2963 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput307 _4082_/ZN spimemio_flash_io1_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput329 _7264_/Q wb_dat_o[26] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_5_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput318 _6791_/Q wb_dat_o[16] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ hold829/Z hold29/Z _4244_/S _4240_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4171_ hold797/Z _4103_/I _4172_/S _4171_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6812_ _6812_/D _7265_/CLK _6812_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6743_ _6743_/D _7237_/RN _4067_/I1 _6743_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_52_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3955_ _7198_/Q _3955_/A2 _3955_/B1 _6847_/Q _3958_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_177_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet763_403 net763_413/I _6771_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_414 net413_72/I _6760_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_91_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6674_ _6674_/D input75/Z _6674_/CLK _6674_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_137_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5625_ hold62/Z hold213/Z _5628_/S _5625_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3886_ _6790_/Q _3928_/B1 _4289_/A1 _6800_/Q _6810_/Q _4301_/A1 _3889_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xnet763_447 net763_447/I _6718_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_436 net763_437/I _6729_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_425 net763_425/I _6749_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_81__1359_ _4073__15/I net413_73/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5556_ hold2/Z hold169/Z _5556_/S _5556_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5487_ _5487_/A1 _5487_/A2 _5487_/A3 _5487_/A4 _5487_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4507_ _5420_/A3 _5129_/A3 _3402_/I _4698_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_4438_ _4648_/A1 _4648_/A2 _4438_/B _4438_/C _5190_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_7226_ _7226_/D _7237_/RN _4067_/I1 _7226_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4369_ _3402_/I _4456_/B _5051_/S _4369_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_7157_ _7157_/D _7221_/RN _7157_/CLK _7157_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_113_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7088_ _7088_/D _7258_/RN _7088_/CLK _7088_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_58_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6108_ _7154_/Q _5960_/Z _5964_/Z hold73/I _5981_/Z _6936_/Q _6109_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_74_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6039_ _6555_/C _7241_/Q _6039_/B _6040_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_73_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2771 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2793 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3740_ _6935_/Q _3910_/A2 _3927_/C2 input29/Z _3954_/A2 _6991_/Q _3759_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_20_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_19 hold75/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3671_ hold54/I _3923_/A2 _5665_/A1 hold43/I _3673_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5410_ _5410_/A1 _5481_/B1 _5410_/B _5411_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6390_ _6390_/A1 _6390_/A2 _6390_/A3 _6390_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_173_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5341_ _4997_/B _4878_/Z _5341_/B _5341_/C _5342_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_126_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet713_355 _4073__7/I _6855_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_377 net813_482/I _6822_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_366 net813_475/I _6844_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5272_ _5165_/Z _5270_/Z _4877_/Z _5425_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_7011_ _7011_/D _7260_/RN _7011_/CLK _7011_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xnet713_399 net763_429/I _6775_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_388 net413_66/I _6786_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4223_ hold533/Z hold29/Z _4227_/S _4223_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4154_ hold62/Z hold70/Z _4157_/S hold71/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4085_ _4059_/S input68/Z _4085_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_102_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4987_ _4367_/Z _5340_/A1 _4555_/B _5172_/B _4987_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6726_ _6726_/D _7193_/RN _6726_/CLK _6726_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3938_ _3929_/Z _3938_/A2 _3938_/A3 _3937_/Z _3938_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_178_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6657_ _7237_/RN _6657_/A2 _6657_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_20_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3869_ _3869_/A1 _3869_/A2 _3869_/A3 _3868_/Z _3869_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6588_ _6834_/Q _6588_/A2 _6588_/B1 _6835_/Q _6836_/Q _6588_/C2 _6589_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_11_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5608_ hold29/Z _6969_/Q hold39/Z hold40/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5539_ _3485_/Z _5857_/A3 _5821_/A3 _5520_/C _5547_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_117_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7209_ _7209_/D _7221_/RN _7209_/CLK _7209_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_154_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2034 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2089 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput28 mask_rev_in[31] input28/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput17 mask_rev_in[21] input17/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput39 mgmt_gpio_in[12] input39/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_6_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_404 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_179_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4910_ _5442_/A2 _4909_/Z _5443_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5890_ hold29/Z hold490/Z _5892_/S _5890_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4841_ _5287_/B _4836_/Z _4841_/B _4841_/C _4846_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_34_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4772_ _4782_/A1 _5302_/B _4695_/Z _4700_/Z _4772_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_119_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3723_ _3719_/Z _3723_/A2 _3723_/A3 _3723_/A4 _3723_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6511_ _6511_/A1 _6511_/A2 _6511_/A3 _6511_/A4 _6511_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3654_ _3485_/Z _3653_/Z _3948_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6442_ _6442_/I _6443_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3585_ _7221_/Q _3912_/A2 _3959_/C1 _7189_/Q _3589_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6373_ _7217_/Q _6274_/Z _6285_/Z _7193_/Q _7177_/Q _6254_/Z _6385_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5324_ _5324_/A1 _5324_/A2 _5324_/B _5324_/C _5444_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_138_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5255_ _5258_/B2 _5255_/A2 _5051_/Z _5255_/B _5446_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_4206_ hold124/Z hold29/Z _4210_/S _4206_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5186_ _4506_/Z _4700_/Z _5339_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_111_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4137_ _3529_/Z _5520_/C hold637/Z _5839_/A3 _4139_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4068_ _6760_/Q _3339_/I _6905_/Q _4068_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_273 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6709_ _6709_/D _7219_/RN _6709_/CLK _6709_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_11_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_275 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1152 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold609 _5833_/Z _7168_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_183_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3370_ _6999_/Q _3370_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5040_ _5439_/B1 _5439_/B2 _5040_/B _5040_/C _5044_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6991_ _6991_/D _7260_/RN _6991_/CLK _6991_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_168_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5942_ _5943_/I0 _5936_/Z _5942_/S _7234_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5873_ hold15/Z hold316/Z _5874_/S _5873_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4824_ _4997_/C _4703_/Z _5370_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_21_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4755_ _4755_/A1 _5313_/A2 _5233_/A1 _4766_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_3706_ hold79/I _5584_/A1 _3951_/C1 _7146_/Q _3707_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_175_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_985 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4686_ _5240_/B _5214_/A2 _4686_/B _4812_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_107_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3637_ input59/Z _4194_/A1 _3917_/A2 _7116_/Q _5528_/S _3619_/Z _3638_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6425_ _6425_/I _6426_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3568_ _3512_/Z _3552_/Z _3941_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_89_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6356_ _6356_/A1 _6356_/A2 _6356_/A3 _6355_/Z _6356_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_142_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5307_ _4586_/Z _4683_/Z _5302_/B _5307_/B _5480_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_0_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3499_ _3499_/I _3500_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6287_ _6287_/A1 _6287_/A2 _6287_/A3 _6554_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_102_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5238_ _5238_/A1 _5454_/A1 _5238_/A3 _5238_/A4 _5238_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_64_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5169_ _5169_/A1 _5425_/A1 _5425_/A3 _5169_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_56_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_224 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_443 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_58__1359_ clkbuf_4_15_0__1359_/Z net763_435/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold6 hold6/I hold6/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_121_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_138__1359_ net563_220/I net813_483/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_75_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4540_ _4441_/B _4501_/B _4460_/B _4436_/B _5278_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_144_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4471_ _4853_/A1 _4481_/A2 _4735_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold417 _4134_/Z _6687_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold406 _5630_/Z _6988_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3422_ _3422_/I0 input58/Z _6733_/Q _3422_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold428 _7212_/Q hold428/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold439 _5845_/Z _7179_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7190_ _7190_/D _7219_/RN _7190_/CLK _7190_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_6210_ _6858_/Q _6210_/A2 _6210_/B _6210_/C _6220_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_172_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6141_ _6141_/A1 _5991_/Z _6146_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_48_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3353_ _7129_/Q _3353_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6072_ _7121_/Q _5969_/Z _6072_/B _6073_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XTAP_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5023_ _5019_/Z _5020_/Z _5023_/A3 _5285_/B _5023_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6974_ _6974_/D _7260_/RN _6974_/CLK _6974_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_53_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5925_ _7228_/Q _7227_/Q _7230_/Q _7229_/Q _5925_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_80_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5856_ hold2/Z hold535/Z _5856_/S _5856_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4807_ _4422_/Z _4534_/Z _5312_/A1 _5414_/A2 _4807_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_55_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5787_ hold271/Z hold976/Z _5793_/S _5787_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4738_ _4699_/Z _5309_/A2 _4738_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_5_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4669_ _4397_/Z _5209_/A3 _4997_/C _5464_/A1 _4669_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_147_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold940 _7159_/Q hold940/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6408_ _6408_/A1 _6408_/A2 _6408_/A3 _6408_/A4 _6408_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold973 _5859_/Z _7191_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold962 _7045_/Q hold962/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold951 _4130_/Z _6683_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold995 _6731_/Q hold995/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_135_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6339_ _7252_/Q _6339_/I1 _6558_/S _7252_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xhold984 _7183_/Q hold984/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet563_231 net613_255/I _6994_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_220 net563_220/I _7005_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_242 net613_258/I _6983_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_431 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3971_ _3971_/A1 _3434_/B _6663_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5710_ _3521_/Z _3537_/Z hold6/Z _5718_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_90_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6690_ _6690_/D _7193_/RN _6690_/CLK _6690_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_86_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5641_ hold674/Z hold86/Z hold19/Z _6998_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5572_ hold29/Z hold66/Z _5574_/S hold67/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4523_ _4460_/B _4436_/B _5139_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold225 _5562_/Z _6928_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold203 _7050_/Q hold203/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_102_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7242_ _7242_/D _7260_/RN _7260_/CLK _7242_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold214 _5625_/Z _6984_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold236 _6913_/Q hold236/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold269 _5544_/Z _6912_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold258 _5549_/Z _6916_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4454_ _3401_/I _3402_/I _4454_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_116_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold247 _5679_/Z _7032_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4385_ input99/Z input98/Z _4386_/A3 _4386_/A4 _4385_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3405_ _4472_/B _4441_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
X_7173_ _7173_/D _7221_/RN _7173_/CLK _7173_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3336_ _7209_/Q _4050_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6124_ _6124_/A1 _6124_/A2 _6124_/A3 _6124_/A4 _6124_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_112_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6055_ _7014_/Q _5971_/Z _5979_/Z _6966_/Q _5996_/Z _7080_/Q _6057_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5006_ _5389_/C _5170_/A2 _5170_/A3 _5130_/B2 _5347_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_100_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_41__1359_ net463_109/I _4073__45/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_66_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_121__1359_ net613_293/I net413_83/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6957_ _6957_/D _7219_/RN _6957_/CLK _6957_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_81_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5908_ _7223_/Q _7224_/Q _7225_/Q _5908_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_139_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6888_ _6888_/D _7210_/RN _6888_/CLK _6888_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_14_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5839_ hold6/Z _3552_/Z _5839_/A3 _5857_/A3 _5847_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_108_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold770 _4272_/Z _6785_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet513_161 net563_221/I _7064_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold781 _7041_/Q hold781/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xnet513_183 net413_76/I _7042_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet513_194 net513_194/I _7031_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_172 _4073__19/I _7053_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold792 _4159_/Z _6706_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_7_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2997 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput308 _7308_/Z spimemio_flash_io2_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_153_262 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput319 _6792_/Q wb_dat_o[17] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4170_ _4170_/A1 hold18/Z _4172_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_171_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_603 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6811_ _6811_/D _7265_/CLK _6811_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6742_ _6742_/D _7193_/RN _6742_/CLK _6742_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3954_ _6988_/Q _3954_/A2 _3954_/B1 input20/Z _4301_/A1 _6809_/Q _3958_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_176_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet763_404 net763_435/I _6770_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_415 net763_416/I _6759_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6673_ hold94/Z _7238_/RN _6673_/CLK hold93/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3885_ _3876_/Z _3885_/A2 _3885_/A3 _3884_/Z _3885_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5624_ hold52/Z hold248/Z _5628_/S _5624_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet763_426 net763_426/I _6748_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_437 net763_437/I _6728_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_448 net763_448/I _6717_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5555_ hold15/Z hold266/Z _5556_/S _5555_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4506_ _4997_/B _4494_/Z _4496_/Z _5263_/A2 _4506_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_133_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5486_ _4616_/Z _4855_/C _5487_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4437_ _4438_/B _4438_/C _4648_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_172_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7225_ _7225_/D _7237_/RN _4067_/I1 _7225_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
XFILLER_105_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7156_ _7156_/D _7221_/RN _7156_/CLK _7156_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4368_ _4456_/B _5051_/S _5270_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_112_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6107_ _7064_/Q _5985_/Z _5997_/Z _7098_/Q _7170_/Q _6006_/Z _6109_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3319_ _7223_/Q _5900_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4299_ _6570_/I0 _6807_/Q _4300_/S _6807_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7087_ _7087_/D _7193_/RN _7087_/CLK _7087_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XTAP_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6038_ _6031_/Z _6037_/Z _6336_/B1 _6168_/C _6555_/C _6039_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_132_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2761 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3670_ _6703_/Q _3927_/A2 _3952_/A2 _7049_/Q _3673_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_173_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5340_ _5340_/A1 _5370_/B _5340_/B _5340_/C _5363_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_127_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5271_ _5165_/Z _5270_/Z _4877_/Z _5271_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_115_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet713_378 net713_379/I _6821_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet713_356 net763_448/I _6854_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_367 net813_475/I _6843_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7010_ _7010_/D _7260_/RN _7010_/CLK _7010_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xnet713_389 net813_472/I _6785_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4222_ _4221_/Z hold547/Z _4228_/S _4222_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4153_ hold52/Z hold502/Z _4157_/S _4153_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4084_ _4084_/I0 _4084_/I1 _6732_/Q _7281_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_441 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4986_ _4986_/A1 _4980_/Z _4986_/A3 _4993_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_51_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6725_ _6725_/D input75/Z _6725_/CLK _6725_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3937_ _3937_/A1 _3937_/A2 _3937_/A3 _3903_/Z _3937_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_177_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6656_ _7237_/RN _6656_/A2 _6656_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3868_ _3868_/A1 _3868_/A2 _3868_/A3 _3868_/A4 _3868_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_20_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6587_ _6587_/I0 _7272_/Q _6602_/S _7272_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5607_ hold62/Z hold72/Z hold39/Z _6968_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3799_ _3798_/Z hold988/Z _3899_/S _6870_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5538_ hold707/Z hold271/Z _5538_/S _5538_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5469_ _5469_/A1 _5423_/Z _5469_/A3 _5469_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_7208_ _7208_/D _7221_/RN _7208_/CLK _7208_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_101_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7139_ _7139_/D _7260_/RN _7139_/CLK hold42/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_98_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1356 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 mask_rev_in[22] input18/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput29 mask_rev_in[3] input29/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_438 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4840_ _5281_/B _5132_/A2 _4840_/B1 _5214_/A2 _4841_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_2591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4771_ _4467_/B _4463_/Z _4782_/A1 _5302_/B _5236_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_20_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6510_ _6841_/Q _6243_/Z _6288_/Z _7296_/Q _6511_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_33_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3722_ _7194_/Q _3909_/A2 _3948_/C1 _7308_/I _4225_/S _4075_/I1 _3723_/A4 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3653_ _3653_/A1 _3492_/Z _3497_/I hold629/Z _3653_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6441_ _6985_/Q _6251_/Z _6273_/Z hold54/I _6265_/Z hold41/I _6442_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6372_ _7169_/Q _5948_/Z _6261_/Z _6959_/Q _6266_/Z hold56/I _6385_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5323_ _5323_/A1 _4920_/Z _5322_/Z _5323_/B _5324_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_3584_ _7197_/Q _3909_/A2 _4227_/S input70/Z _4194_/A1 input60/Z _3589_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_142_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5254_ _4761_/I _5245_/Z _5254_/B _5254_/C _5257_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_114_276 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5185_ _5185_/A1 _5185_/A2 _6577_/C _5185_/B2 _6860_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_130_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4205_ _4204_/Z hold850/Z _4211_/S _4205_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4136_ hold2/Z hold370/Z _4136_/S _4136_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4067_ _6761_/Q _4067_/I1 _6903_/Q _4067_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4969_ _4718_/B _4903_/Z _5072_/A4 _4421_/Z _4969_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_178_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6708_ _6708_/D _7219_/RN _6708_/CLK _6708_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_22_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ _7221_/RN _6656_/A2 _6639_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_138_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_805 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet613_300 net613_300/I _6925_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1164 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6990_ _6990_/D _7238_/RN _6990_/CLK _6990_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5941_ _5941_/A1 _5940_/Z _5943_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_93_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5872_ hold29/Z hold460/Z _5874_/S _5872_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4823_ _5270_/A1 _4454_/Z _4997_/C _4554_/Z _4659_/Z _4826_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_187_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4754_ _4716_/Z _4752_/Z _5233_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_105_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3705_ _6960_/Q _3957_/A2 _3959_/B1 _6670_/Q _3707_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_174_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4685_ _4685_/A1 _4685_/A2 _5180_/A3 _5211_/C _5001_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_119_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3636_ _7196_/Q _3909_/A2 _4227_/S input69/Z _3945_/B1 _7092_/Q _3638_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_88_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6424_ _7171_/Q _5948_/Z _6263_/Z hold66/I _6425_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_161_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3567_ _3512_/Z _3529_/Z _5683_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6355_ _6355_/A1 _6355_/A2 _6355_/A3 _6355_/A4 _6355_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6286_ _6287_/A1 _6287_/A2 _6287_/A3 _6286_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_5306_ _5306_/I _5307_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3498_ _7303_/Q input58/Z _6733_/Q _3499_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5237_ _5238_/A1 _5238_/A4 _5457_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_88_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5168_ _4454_/Z _4997_/C _4820_/Z _4456_/B _5425_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_111_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5099_ _5099_/A1 _5099_/A2 _4716_/Z _4784_/Z _4549_/Z _5100_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_84_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_355 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4119_ _5520_/C _3533_/Z _5839_/A3 _5857_/A3 _4127_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_71_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_1_1__f__1062_ clkbuf_0__1062_/Z _6568_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_153_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold7 hold7/I hold7/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_47_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_5__1359_ net713_387/I net413_55/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_677 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold418 _7164_/Q hold418/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4470_ _4463_/Z _4468_/Z _4765_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold407 _7134_/Q hold407/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3421_ _3421_/A1 _3421_/A2 _7304_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xhold429 _5882_/Z _7212_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3352_ _7137_/Q _3352_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6140_ _7026_/Q wire348/Z _6211_/B1 _6994_/Q _6141_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6071_ _7153_/Q _5960_/Z _5965_/Z _6701_/Q _5981_/Z _6935_/Q _6073_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_85_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _5198_/C _5023_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_4_0__1359_ net663_304/I clkbuf_opt_4_1__1359_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_85_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6973_ _6973_/D _7219_/RN _6973_/CLK _6973_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_0_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5924_ _6021_/A2 _6015_/A3 _6014_/A2 _5984_/A1 _5924_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_94_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5855_ hold15/Z hold288/Z _5856_/S _5855_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4806_ _4492_/Z _4536_/Z _5319_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_10_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5786_ hold113/Z hold617/Z _5793_/S _5786_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4737_ _5226_/C _5226_/B _5309_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_299 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4668_ _4411_/Z _5343_/A1 _5393_/A2 _5165_/A4 _5360_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xclkbuf_leaf_64__1359_ clkbuf_4_15_0__1359_/Z net413_76/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_134_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_144__1359_ net713_387/I net763_443/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_135_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold930 _6890_/Q hold930/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3619_ _7260_/Q _6899_/Q _6900_/Q _3619_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6407_ _7072_/Q _6248_/Z _6293_/Z _7154_/Q _6407_/C _6408_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4599_ _5129_/A3 _4598_/Z _5051_/S _4454_/Z _4599_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_134_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold963 _5694_/Z _7045_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold941 _5823_/Z _7159_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold952 _7068_/Q hold952/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold996 _7298_/Q _3433_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_143_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6338_ _6338_/I _6339_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold985 _5850_/Z _7183_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold974 _6709_/Q hold974/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_0_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6269_ _7235_/Q _7234_/Q _6302_/A3 _6533_/A2 _6269_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_103_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet563_210 net663_326/I _7015_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_221 net563_221/I _7004_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_243 net763_426/I _6982_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_232 net663_329/I _6993_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_962 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3970_ _3967_/Z _3970_/A2 _6664_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_189_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5640_ hold619/Z hold271/Z hold19/Z _6997_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5571_ hold62/Z hold216/Z _5574_/S _5571_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4522_ _4441_/B _5288_/B _5315_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_144_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold226 _7059_/Q hold226/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7241_ _7241_/D _7258_/RN _7258_/CLK _7241_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4453_ _3401_/I _3402_/I _4555_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_117_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold204 _5699_/Z _7050_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold215 _6960_/Q hold215/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold237 _5545_/Z _6913_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3404_ _5051_/S _4835_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_116_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold259 _6959_/Q hold259/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold248 _6983_/Q hold248/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4384_ _4376_/Z _4381_/Z _4580_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_131_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7172_ _7172_/D _7221_/RN _7172_/CLK _7172_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_98_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3335_ _7217_/Q _4049_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6123_ hold45/I _5987_/Z _6015_/Z _7009_/Q _6124_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_105_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6054_ _6934_/Q _5981_/Z _5988_/Z _6982_/Q _7046_/Q _6019_/Z _6057_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ _5043_/A2 _5389_/C _5393_/B1 _5043_/B _5347_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3340__1 _3340__1/I _6603_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_859 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6956_ _6956_/D _7297_/RN _6956_/CLK _6956_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_42_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5907_ _5906_/Z _5904_/B _7225_/Q _7225_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6887_ _6887_/D _7297_/RN _6887_/CLK _6887_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_22_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5838_ hold2/Z hold228/Z _5838_/S _5838_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5769_ hold271/Z hold968/Z _5775_/S _5769_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_625 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold771 _6757_/Q hold771/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold760 _4120_/Z _6674_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold782 _5689_/Z _7041_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xnet513_162 _4073__37/I _7063_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet513_195 net413_81/I _7030_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_173 _4073__39/I _7052_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_184 net813_465/I _7041_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold793 _6849_/Q hold793/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput309 _7309_/Z spimemio_flash_io3_di VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_142_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_442 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6810_ _6810_/D _7210_/RN _6810_/CLK _6810_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_24_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6741_ _6741_/D _7193_/RN _6741_/CLK _6741_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3953_ _3953_/A1 _3953_/A2 _3953_/A3 _3953_/A4 _3953_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_189_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet763_405 net763_435/I _6769_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6672_ hold98/Z _7238_/RN _6672_/CLK hold97/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_3884_ _3884_/A1 _3884_/A2 _3884_/A3 _3884_/A4 _3884_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_137_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet763_416 net763_416/I _6758_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5623_ hold86/Z hold414/Z _5628_/S _5623_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet763_427 net413_88/I _6747_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_438 net413_55/I _6727_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_449 net813_475/I _6716_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5554_ hold29/Z hold829/Z _5556_/S _5554_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4505_ _5340_/A1 _4495_/Z _4497_/Z _5262_/A2 _5343_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_133_937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5485_ _5480_/Z _5485_/A2 _5485_/B _5490_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_105_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4436_ _5281_/C _5464_/A1 _4436_/B _4438_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_7224_ _7224_/D _7237_/RN _4067_/I1 _7224_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_117_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4367_ _4456_/B _5051_/S _4367_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_116_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7155_ _7155_/D _7297_/RN _7155_/CLK _7155_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3318_ _6743_/Q _5945_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_6106_ _6106_/A1 _6106_/A2 _6106_/A3 _6106_/A4 _6106_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_86_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7086_ _7086_/D _7219_/RN _7086_/CLK _7086_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_58_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4298_ _6569_/I0 _6806_/Q _4300_/S _6806_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6037_ _6037_/A1 _6037_/A2 _6037_/A3 _6037_/A4 _6037_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_6_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6939_ _6939_/D _7221_/RN _6939_/CLK _6939_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_81_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_179_171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold590 _7113_/Q hold590/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2784 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5270_ _5270_/A1 _4454_/Z _4997_/C _4820_/Z _5270_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_99_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet713_368 net763_448/I _6842_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_357 net763_448/I _6853_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4221_ hold81/Z hold62/Z _4227_/S _4221_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet713_379 net713_379/I _6820_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4152_ hold86/Z hold914/Z _4157_/S _4152_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4083_ _6734_/Q _6731_/Q _4084_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_110_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4985_ _4397_/Z _5209_/A3 _4659_/Z _4703_/Z _4985_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_63_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6724_ _6724_/D input75/Z _6724_/CLK _6724_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3936_ _7028_/Q _5674_/A1 _3936_/B1 _6690_/Q _3937_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6655_ _7237_/RN _6657_/A2 _6655_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3867_ _7079_/Q _3923_/C1 _3956_/B1 _6713_/Q _3867_/C _3868_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6586_ _6586_/A1 _4313_/Z _6586_/B _6587_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_5606_ hold52/Z hold250/Z hold39/Z _6967_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3798_ _6566_/I0 _6869_/Q _3898_/S _3798_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5537_ hold681/Z _4103_/I _5538_/S _5537_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5468_ _5468_/A1 _5468_/A2 _5468_/B1 _4650_/Z _5468_/C _5469_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_127_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7207_ _7207_/D _7219_/RN _7207_/CLK _7207_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4419_ _5420_/A3 _5420_/A2 _4456_/B _4419_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_132_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5399_ _4524_/Z _5399_/A2 _4683_/Z _5302_/B _5399_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_87_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7138_ _7138_/D _7238_/RN _7138_/CLK _7138_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_143_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7069_ _7069_/D _7219_/RN _7069_/CLK _7069_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_59_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2069 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 mask_rev_in[23] input19/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_762 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2592 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_618 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ _4770_/A1 _5118_/A3 _4770_/A3 _5117_/A1 _4775_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_186_450 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3721_ _6678_/Q _3546_/Z _3916_/A2 _7154_/Q _7170_/Q _3941_/B1 _3723_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3652_ input68/Z _4227_/S _4244_/S input40/Z _3657_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6440_ _6440_/A1 _6440_/A2 _6440_/A3 _6439_/Z _6440_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_173_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6371_ _7063_/Q _6257_/Z _6299_/Z _7055_/Q _6383_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_127_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3583_ _6971_/Q _3924_/A2 _3607_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_61_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5322_ _4436_/B _4494_/Z _5328_/A2 _5056_/C _5322_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1022 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5253_ _5254_/C _5334_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5184_ _6834_/Q _5182_/Z _5184_/B _5184_/C _5185_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_4204_ hold562/Z hold62/Z _4210_/S _4204_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4135_ hold15/Z hold403/Z _4136_/S _4135_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4066_ _6762_/Q user_clock _6904_/Q _4066_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4968_ _4903_/Z _5072_/A4 _4718_/B _4666_/Z _4968_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_51_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4899_ _6577_/C _4899_/A2 _5000_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6707_ _6707_/D _7219_/RN _6707_/CLK _6707_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3919_ _3919_/A1 _3919_/A2 _3919_/A3 _3919_/A4 _3919_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6638_ _7221_/RN _6656_/A2 _6638_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_149_185 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6569_ _6569_/I0 _7267_/Q _6571_/S _7267_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_269 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_494 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet613_301 _4073__45/I _6924_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__2 _4073__2/I _7297_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_156_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_334 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5940_ _6745_/Q _7233_/Q _7232_/Q _7234_/Q _5940_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_92_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3090 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5871_ hold62/Z hold529/Z _5874_/S _5871_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4822_ _4554_/Z _4659_/Z _4820_/Z _5364_/B _4826_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_33_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4753_ _4700_/Z _4752_/Z _5313_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3704_ _7138_/Q _3951_/A2 _3901_/A2 _6984_/Q input30/Z _3927_/C2 _3707_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_175_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4684_ _4414_/Z _4452_/Z _4666_/Z _4892_/B _4683_/Z _4685_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_6423_ _7099_/Q _6250_/Z _6439_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_162_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3635_ input50/Z _4210_/S _3947_/A2 _7100_/Q _3638_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_143_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6354_ _7168_/Q _5948_/Z _6261_/Z _6958_/Q _6355_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3566_ _3507_/Z _3533_/Z _3954_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6285_ _6484_/A2 _6285_/A2 _7237_/Q _6452_/A4 _6285_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3497_ _3497_/I _3617_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
X_5305_ _4586_/Z _4673_/Z _5302_/B _5305_/B _5306_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_170_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5236_ _4510_/Z _5414_/A2 _5236_/B _5238_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_124_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5167_ _4546_/Z _4651_/Z _4675_/Z _5167_/B _5425_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_84_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1077 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5098_ _5098_/A1 _5302_/B _5098_/B _5098_/C _5101_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_4118_ hold2/Z hold93/Z _4118_/S hold94/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4049_ _4049_/I0 input92/Z _4050_/S _4049_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_24__1359_ net613_253/I _4073__18/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_56_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_104__1359_ clkbuf_4_5_0__1359_/Z net613_281/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_87__1359_ clkbuf_4_13_0__1359_/Z net413_81/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_204 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold8 hold8/I hold8/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_181_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold408 _7144_/Q hold408/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_172_979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3420_ _3988_/S _3422_/I0 _3421_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_128_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold419 _5828_/Z _7164_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_87_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3351_ _7145_/Q _3351_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6070_ hold77/I _5958_/Z _5967_/Z _7105_/Q _7137_/Q _5994_/I _6073_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_79_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5021_ _4604_/Z _4606_/Z _5003_/Z _5021_/B _5198_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_79_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6972_ _6972_/D _7193_/RN _6972_/CLK _6972_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_19_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_581 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5923_ _7230_/Q _7229_/Q _6210_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_94_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5854_ hold29/Z hold304/Z _5856_/S _5854_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4805_ _4835_/A2 _4492_/Z _4534_/Z _4681_/Z _4805_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_21_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5785_ _5520_/C _3552_/Z _5857_/A3 _5857_/A2 _5793_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_181_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4736_ _4736_/A1 _5302_/B _4736_/A3 _4467_/B _5226_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_175_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4667_ _4414_/Z _5038_/A1 _4557_/Z _4666_/Z _4667_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_163_935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3618_ _3527_/Z _3617_/Z _5528_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold920 _5631_/Z _6989_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold931 _5512_/Z _6890_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6406_ _6406_/I _6407_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_150_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6337_ _6744_/Q _7251_/Q _6337_/B _6338_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_122_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4598_ _5287_/B _4460_/B _5399_/A2 _4436_/B _4598_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold964 _7069_/Q hold964/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold942 _7036_/Q hold942/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold953 _5720_/Z _7068_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold997 _7295_/Q hold997/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3549_ _3485_/Z _3512_/Z _4194_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_88_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold986 _7087_/Q hold986/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold975 _4163_/Z _6709_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6268_ _7233_/Q _7232_/Q _6533_/A2 _6452_/A4 _6268_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_103_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5219_ _5303_/A1 _5303_/A3 _5224_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_9_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6199_ _6789_/Q _5972_/Z _6021_/Z _6839_/Q _6201_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_57_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_222 net563_246/I _7003_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_211 net813_465/I _7014_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet563_233 net613_276/I _6992_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet563_244 net413_90/I _6981_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_158_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_70__1359_ clkbuf_4_13_0__1359_/Z net563_215/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_679 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_150__1359_ net713_387/I net813_491/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_31_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5570_ hold52/Z hold598/Z _5574_/S _5570_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_184_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4521_ _4472_/B _4501_/B _5139_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_129_475 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4452_ _5038_/A1 _4648_/B _4638_/A2 _4452_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_172_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7240_ _7240_/D _7258_/RN _4067_/I1 _7240_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold205 _7205_/Q hold205/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_117_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold216 _6936_/Q hold216/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold238 _6769_/Q hold238/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_160_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold227 _5709_/Z _7059_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3403_ _4456_/B _5129_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
Xhold249 _5624_/Z _6983_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4383_ _5464_/A1 _4383_/A2 _5385_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_171_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7171_ _7171_/D _7297_/RN _7171_/CLK _7171_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3334_ _3334_/I _4029_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6122_ _7091_/Q _6002_/Z _6003_/Z _7163_/Q _6124_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_140_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6053_ _6053_/A1 _6053_/A2 _6053_/A3 _6053_/A4 _6053_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5004_ _5368_/A1 _5420_/A1 _5002_/Z _5389_/B _5191_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_100_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_465 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6955_ hold92/Z _7238_/RN _6955_/CLK hold91/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5906_ _7223_/Q _7224_/Q _5910_/B _5906_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_41_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6886_ _6886_/D _7297_/RN _6886_/CLK _6886_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_34_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5837_ hold15/Z hold729/Z _5838_/S _5837_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5768_ hold113/Z hold573/Z _5775_/S _5768_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4719_ _5083_/B _4719_/A2 _4721_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_175_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5699_ hold15/Z hold203/Z _5700_/S _5699_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet513_152 net513_152/I _7073_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold772 _4235_/Z _6757_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold761 _6891_/Q hold761/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold750 _4181_/Z _6721_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_150_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet513_163 _4073__37/I _7062_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet513_174 net613_258/I _7051_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_185 net513_185/I _7040_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold783 _7091_/Q hold783/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold794 _4348_/Z _6849_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_162_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet513_196 _4073__43/I _7029_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1058 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6740_ _6740_/D _7193_/RN _6740_/CLK _6740_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3952_ _7044_/Q _3952_/A2 _5638_/A1 _6996_/Q _6948_/Q _5584_/A1 _3953_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_149_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet763_406 net763_431/I _6768_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_91_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3883_ input53/Z _4194_/A1 _3948_/C1 input62/Z _3941_/B1 _7167_/Q _3884_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6671_ _6671_/D _7238_/RN _6671_/CLK _6671_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_31_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet763_417 net763_419/I _6757_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_428 net763_429/I _6742_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5622_ hold271/Z hold896/Z _5628_/S _5622_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet763_439 net413_55/I _6726_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_367 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5553_ hold62/Z hold330/Z _5556_/S _5553_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4504_ _4759_/A2 _4759_/A3 _4504_/B _4504_/C _5263_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_145_721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5484_ _5483_/Z _5450_/I _5477_/Z _5441_/B _5485_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_160_713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4435_ _5281_/C _5270_/A1 _5170_/A2 _4436_/B _4438_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7223_ _7223_/D _7237_/RN _4067_/I1 _7223_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4366_ _4472_/B _4460_/B _4436_/B _4853_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_116_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7154_ _7154_/D _7193_/RN _7154_/CLK _7154_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3317_ _6836_/Q _4686_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_141_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6105_ _7114_/Q _5984_/Z _6000_/Z _7130_/Q _6106_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_7085_ _7085_/D _7221_/RN _7085_/CLK _7085_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_86_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4297_ _4309_/I0 _6805_/Q _4300_/S _6805_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _6973_/Q _5964_/Z _5984_/Z _7111_/Q _6036_/C _6037_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6938_ _6938_/D _7221_/RN _6938_/CLK _6938_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XPHY_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6869_ _6869_/D _6627_/Z _4075_/I1 _6869_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_50_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_827 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_378 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold580 _7174_/Q hold580/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold591 _5771_/Z _7113_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2796 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet713_358 net713_358/I _6852_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet713_369 net763_448/I _6841_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4220_ _4219_/Z hold541/Z _4228_/S _4220_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4151_ hold271/Z hold916/Z _4157_/S _4151_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4082_ _4082_/A1 _7299_/Q _4082_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_37_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4984_ _4700_/Z _4982_/Z _4984_/B _4986_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_177_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6723_ _6723_/D _7297_/RN _6723_/CLK _6723_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3935_ _6924_/Q _3935_/A2 _3935_/B1 _6849_/Q _3937_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_189_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6654_ _7237_/RN _6657_/A2 _6654_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_32_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3866_ _3866_/A1 _3537_/Z _3617_/Z _3866_/B _3867_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_5605_ hold86/Z hold103/Z hold39/Z _6966_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6585_ _6834_/Q _6585_/A2 _6585_/B1 _6835_/Q _6836_/Q _6585_/C2 _6586_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_178_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3797_ _3776_/Z _3797_/A2 _3797_/A3 _3796_/Z _6566_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_145_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5536_ _5536_/A1 hold18/Z _5538_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_5467_ _4570_/Z _4651_/Z _5467_/B _5467_/C _5468_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_117_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4418_ _5170_/A2 _4456_/B _5343_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_133_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7206_ _7206_/D _7210_/RN _7206_/CLK _7206_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_5398_ _5391_/Z _5398_/A2 _5419_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_114_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4349_ hold271/Z hold862/Z _4349_/S _4349_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7137_ _7137_/D _7238_/RN _7137_/CLK _7137_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_7068_ _7068_/D _7193_/RN _7068_/CLK _7068_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_6019_ _7228_/Q _7227_/Q wire348/Z _6210_/A2 _6019_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_2015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_410 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2571 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_3720_ _7114_/Q _3917_/A2 _3947_/A2 _7098_/Q _3945_/A2 _7178_/Q _3723_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_187_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_665 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3651_ _7187_/Q _3959_/C1 _3960_/A2 _7211_/Q _3657_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6370_ _6991_/Q _6237_/Z _6380_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3582_ _3509_/Z _3515_/Z _3924_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_161_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5321_ _5321_/A1 _5212_/Z _5454_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_54_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1045 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5252_ _5343_/A1 _5343_/A2 _5255_/A2 _5252_/B _5254_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_142_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4203_ _4202_/Z hold775/Z _4211_/S _4203_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5183_ _5181_/Z _4686_/B _5299_/C _5184_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_87_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_866 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4134_ hold29/Z hold416/Z _4136_/S _4134_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4065_ _6392_/B1 input2/Z input1/Z _4065_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1046 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4967_ _4903_/Z _5072_/A4 _4718_/B _5359_/A1 _4967_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_33_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_974 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4898_ _3401_/I _4893_/Z _4898_/B _4898_/C _4899_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_6706_ _6706_/D _7219_/RN _6706_/CLK _6706_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3918_ input36/Z _4225_/S _4143_/A1 _6694_/Q _3919_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6637_ _7237_/RN _6656_/A2 _6637_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
X_3849_ _7175_/Q _3945_/A2 _3939_/C1 _6711_/Q _3897_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_180_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6568_ _6568_/I0 _7266_/Q _6571_/S _7266_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_47__1359_ net463_109/I net413_96/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_127__1359_ _4073__15/I _4073__19/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5519_ _6894_/Q hold339/Z _5520_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_105_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6499_ _6554_/A1 _6499_/A2 _6499_/A3 _6498_/Z _6499_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_87_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_674 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__3 _4073__3/I _7296_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_7_0__1359_ clkbuf_0__1359_/Z net813_465/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_11_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3091 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5870_ hold52/Z hold592/Z _5874_/S _5870_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4821_ _4554_/Z _4472_/B _4887_/A1 _4501_/B _4821_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_2390 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_760 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4752_ _5302_/B _4436_/B _4463_/Z _5226_/C _4752_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_175_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4683_ _5420_/A3 _4835_/A2 _4456_/B _3402_/I _4683_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_105_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3703_ input48/Z _4210_/S _4244_/S input39/Z _3708_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_162_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3634_ _7220_/Q _3912_/A2 _4244_/S input41/Z _3930_/A2 _7132_/Q _3638_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_88_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6422_ _7065_/Q _6257_/Z _6434_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_134_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6353_ _7208_/Q _6256_/Z _6285_/Z _7192_/Q _6274_/Z _7216_/Q _6355_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_115_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3565_ _3509_/Z _3542_/Z _3901_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_142_362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3496_ _3495_/Z hold635/Z hold21/Z _3496_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_6284_ _6281_/Z _6283_/Z _6251_/Z _6273_/Z _6287_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_103_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5304_ _4683_/Z _5302_/B _5456_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5235_ _5316_/A2 _5234_/Z _5238_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_69_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5166_ _5166_/A1 _5467_/B _5166_/A3 _5165_/Z _5169_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_96_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_836 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4117_ hold1/Z _7277_/Q hold21/I hold2/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_151_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5097_ _5097_/A1 _5328_/A2 _5368_/B _3401_/I _5098_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_112_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4048_ _6767_/Q input89/Z _4050_/S _4048_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_216 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5999_ wire348/Z _6021_/A2 _6210_/A2 _7227_/Q _5999_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_138_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_782 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput290 _6685_/Q pll_trim[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold9 hold9/I hold9/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_59_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_281 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold409 _5806_/Z _7144_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_174_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_30__1359_ clkbuf_opt_3_0__1359_/Z net663_313/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3350_ _7153_/Q _3350_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_110__1359_ _4073__15/I net413_70/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_152_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_93__1359_ net813_465/I net563_225/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5020_ _5438_/C _5359_/A1 _4604_/Z _4606_/Z _5020_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6971_ _6971_/D _7260_/RN _6971_/CLK _6971_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_0_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5922_ _5922_/I _7229_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5853_ hold62/Z hold343/Z _5856_/S _5853_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4804_ _4681_/Z _4793_/Z _5319_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5784_ hold2/Z hold163/Z _5784_/S _5784_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4735_ _4501_/B _4735_/A2 _4764_/A3 _5226_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_9_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_487 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4666_ _5420_/A3 _5420_/A2 _4835_/A2 _4456_/B _4666_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4597_ _5287_/B _4596_/Z _5420_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3617_ _3617_/A1 hold629/Z _3489_/I _3492_/Z _3617_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold921 _7119_/Q hold921/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6405_ _7138_/Q _6253_/Z _6297_/Z hold70/I _6406_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold910 _7150_/Q hold910/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3548_ _3519_/Z _3533_/Z _3945_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6336_ _6329_/Z _6335_/Z _6336_/B1 _6286_/Z _6555_/C _6337_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold954 _6965_/Q hold954/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold943 _5684_/Z _7036_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold932 _7103_/Q hold932/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold998 _6731_/Q _3312_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold976 _7127_/Q hold976/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold965 _5721_/Z _7069_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold987 _5742_/Z _7087_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3479_ _6659_/Q _6658_/Q _6733_/Q _3479_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6267_ _6996_/Q _6265_/Z _6266_/Z _7012_/Q _6271_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5218_ _4673_/Z _4700_/Z _5218_/B _5303_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_88_268 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6198_ _6198_/A1 _6198_/A2 _6198_/A3 _6198_/A4 _6198_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5149_ _5165_/A2 _4598_/Z _5374_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xnet563_212 net563_212/I _7013_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_234 net613_255/I _6991_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_223 net613_281/I _7002_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_245 net613_293/I _6980_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_446 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_485 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_833 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1000 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ _4835_/A2 _4456_/B _3402_/I _3401_/I _5359_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_116_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4451_ _4604_/A2 _4604_/A3 _4451_/B _4451_/C _5038_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_144_435 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold206 _5874_/Z _7205_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold217 _5571_/Z _6936_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_7_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold239 _4254_/Z _6769_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3402_ _3402_/I _5420_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
Xhold228 _7173_/Q hold228/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7170_ _7170_/D _7193_/RN _7170_/CLK _7170_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4382_ _4472_/B _4501_/B _4460_/B _4436_/B _4383_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_153_980 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6121_ _6985_/Q _5988_/Z _6019_/Z _7049_/Q _6124_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3333_ _4483_/B _4424_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_112_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6052_ _6950_/Q _5958_/Z _5967_/Z _7104_/Q _6052_/C _6053_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _5165_/A4 _5003_/A2 _4421_/Z _4491_/B _5003_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_79_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0__1062_ _3725_/ZN clkbuf_0__1062_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6954_ hold27/Z _7238_/RN _6954_/CLK hold26/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5905_ _5905_/I _7224_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6885_ _6885_/D _7297_/RN _6885_/CLK _6885_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_14_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5836_ hold29/Z hold326/Z _5838_/S _5836_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5767_ _5857_/A3 _5839_/A3 _3537_/Z _5520_/C _5775_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4718_ _4504_/B _4504_/C _4718_/B _5056_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_135_402 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_627 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5698_ hold29/Z hold506/Z _5700_/S _5698_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4649_ _4570_/Z _5438_/B _4653_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_107_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold773 _6902_/Q hold773/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold740 _4214_/Z _6747_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold751 _6837_/Q hold751/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold762 _5514_/Z _6891_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold795 _6770_/Q hold795/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7299_ _7299_/D _6651_/Z _7304_/CLK _7299_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
Xnet513_186 net413_80/I _7039_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet513_175 net513_194/I _7050_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6319_ _7127_/Q _6484_/A2 _6533_/A3 _7111_/Q _6320_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xnet513_164 net413_57/I _7061_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold784 _5746_/Z _7091_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xnet513_153 net563_251/I _7072_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet513_197 _4073__39/I _7028_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_452 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2945 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2923 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3951_ _7134_/Q _3951_/A2 _5665_/A1 _7020_/Q _3951_/C1 _7142_/Q _3953_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_63_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3882_ _6925_/Q _3935_/A2 _3933_/B1 _6786_/Q _3942_/C1 _6854_/Q _3884_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6670_ _6670_/D _7238_/RN _6670_/CLK _6670_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_31_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet763_418 net763_418/I _6756_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet763_407 net763_431/I _6767_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_91_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet763_429 net763_429/I _6741_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ hold113/Z hold695/Z _5628_/S _5621_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_560 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5552_ hold52/Z hold347/Z _5556_/S _5552_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4503_ _4718_/B _5072_/A4 _5262_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_145_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5483_ _5483_/A1 _5483_/A2 _5483_/A3 _5483_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_144_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_457 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7222_ _7222_/D _7237_/RN _4067_/I1 _7222_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4434_ _4467_/B _4460_/B _4887_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_132_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4365_ _4472_/B _4460_/B _4436_/B _5288_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_160_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7153_ _7153_/D _7221_/RN _7153_/CLK _7153_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_113_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3316_ _6835_/Q _4415_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_7084_ _7084_/D _7221_/RN _7084_/CLK _7084_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6104_ _7106_/Q _5967_/Z _5980_/Z _7072_/Q _5969_/Z _7122_/Q _6106_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_101_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6035_ _6035_/I _6036_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4296_ _6567_/I0 _6804_/Q _4300_/S _6804_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_978 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1518 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1507 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6937_ hold67/Z _7238_/RN _6937_/CLK hold66/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XPHY_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6868_ _6868_/D _6626_/Z _4075_/I1 _6868_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
XFILLER_167_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5819_ hold15/Z hold422/Z _5820_/S _5819_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6799_ _6799_/D _7210_/RN _6799_/CLK _6799_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_182_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold570 _5754_/Z _7098_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold581 _5840_/Z _7174_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold592 _7201_/Q hold592/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_278 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2764 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet713_359 net763_443/I _6851_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4150_ hold113/Z hold465/Z _4157_/S _4150_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4081_ _4081_/A1 input73/Z _4081_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_83_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4983_ _5083_/C _4659_/Z _4703_/Z _4422_/Z _4984_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_51_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6722_ _6722_/D _7297_/RN _6722_/CLK _6722_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3934_ _7004_/Q _3934_/A2 _3934_/B1 _6845_/Q _5532_/A1 _6905_/Q _3937_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6653_ _7237_/RN _4064_/S _6653_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_20_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3865_ _6900_/Q _5528_/S _6611_/A1 _7297_/Q _3868_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_149_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5604_ hold271/Z hold954/Z hold39/Z _6965_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6584_ _6584_/I0 _7271_/Q _6602_/S _7271_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3796_ _3796_/A1 _3796_/A2 _3786_/Z _3795_/Z _3796_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_20_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5535_ hold537/Z hold113/Z _5535_/S _5535_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5466_ _5425_/Z _5428_/Z _5429_/Z _5465_/Z _5466_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4417_ _5129_/A3 _4835_/A2 _4836_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7205_ _7205_/D _7237_/RN _7205_/CLK _7205_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5397_ _5433_/A2 _5433_/A3 _5434_/A2 _5209_/Z _5398_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_120_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7136_ _7136_/D _7238_/RN _7136_/CLK _7136_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
X_4348_ _4103_/I hold793/Z _4349_/S _4348_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7067_ _7067_/D _7237_/RN _7067_/CLK _7067_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4279_ hold271/Z hold860/Z _4279_/S _4279_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_688 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6018_ _7143_/Q _7231_/Q _6210_/B wire348/Z _6024_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_2016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2005 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_183_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_170_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2594 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_187 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3650_ _7195_/Q _3909_/A2 _4194_/A1 input57/Z _3955_/A2 _7203_/Q _3689_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_174_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3581_ _3523_/Z _3533_/Z _3925_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_170_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5320_ _5320_/A1 _5319_/Z _5452_/A2 _5453_/A4 _5320_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5251_ _5330_/B2 _5246_/Z _5251_/B _5254_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_114_213 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4202_ hold332/Z hold52/Z _4210_/S _4202_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5182_ _5182_/A1 _5340_/C _5265_/A4 _4511_/Z _5182_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_123_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4133_ hold62/Z hold467/Z _4136_/S _4133_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4064_ _6392_/B1 _7281_/Q _4064_/S _4064_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4966_ _4966_/A1 _4966_/A2 _5073_/B _4970_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_149_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6705_ _6705_/D _7237_/RN _6705_/CLK _6705_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_149_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4897_ _6834_/Q _6835_/Q _6836_/Q _4897_/A4 _4898_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3917_ _7110_/Q _3917_/A2 _6611_/A1 _7296_/Q _3919_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_177_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6636_ _7237_/RN _6657_/A2 _6636_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_165_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3848_ _7127_/Q _3930_/A2 _3920_/B1 _6867_/Q _3922_/B1 _6693_/Q _3897_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_22_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3779_ _6982_/Q _3901_/A2 _3927_/B1 _7062_/Q _3796_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6567_ _6567_/I0 _7265_/Q _6571_/S _7265_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5518_ _4103_/I hold858/Z _5518_/S _5518_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6498_ _6498_/A1 _6498_/A2 _6498_/A3 _6498_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_172_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5449_ _5449_/A1 _5342_/I _5416_/I _5449_/A4 _5450_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_133_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7119_ _7119_/D _7210_/RN _7119_/CLK _7119_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_86_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1123 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/Z _4072_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_151_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_931 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4073__4 _4073__9/I _7221_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_956 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3092 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3081 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3070 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4820_ _4489_/B _4483_/B _4026_/B _4026_/C _4820_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_2380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_227 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_53__1359_ net663_324/I _4073__37/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2391 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1690 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4751_ _4751_/A1 _4748_/Z _4750_/Z _4755_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_15_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4682_ _4530_/I _4878_/A2 _5312_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3702_ _7218_/Q _3912_/A2 _4194_/A1 input56/Z _3941_/A2 _7162_/Q _3708_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_30_984 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6421_ _7255_/Q _6421_/I1 _6558_/S _7255_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3633_ _6978_/Q _3923_/A2 _3960_/A2 _7212_/Q _3633_/C _3646_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_146_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3564_ _3515_/Z _3537_/Z _3945_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6352_ _6990_/Q _6237_/Z _6240_/Z _7112_/Q _6352_/C _6356_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3495_ _7304_/Q _7303_/Q _6733_/Q _3495_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6283_ _6241_/Z _6275_/Z _6282_/Z _6283_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_5303_ _5303_/A1 _5303_/A2 _5303_/A3 _5303_/A4 _5303_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_170_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5234_ _5234_/A1 _5314_/A1 _5404_/A1 _5234_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_5165_ _5209_/A3 _5165_/A2 _4651_/Z _5165_/A4 _5165_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_124_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4116_ hold15/Z hold97/Z _4118_/S hold98/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5096_ _4539_/I _5287_/B _4673_/Z _4460_/B _5098_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4047_ _6768_/Q input91/Z _4050_/S _4047_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5998_ _7078_/Q _5996_/Z _5997_/Z _7094_/Q _6008_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_185_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4949_ _5464_/A1 _4944_/Z _5065_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_166_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6619_ _7237_/RN _6657_/A2 _6619_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_177_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_606 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_800 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput280 _6668_/Q pll_trim[18] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_94_409 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput291 _6686_/Q pll_trim[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_48_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_488 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_988 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_639 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1010 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6970_ _6970_/D _7260_/RN _6970_/CLK _6970_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_65_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ _5920_/Z _6745_/Q _7229_/Q _5913_/I _5922_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5852_ hold52/Z hold520/Z _5856_/S _5852_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4803_ _4803_/A1 _4797_/Z _4803_/B _4809_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_5783_ hold15/Z hold180/Z _5784_/S _5783_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4734_ _4703_/Z _4728_/Z _5106_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_147_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_809 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4665_ _5170_/A2 _4878_/A2 _5389_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_147_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4596_ _5288_/B _4460_/B _4436_/B _4472_/B _4596_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_3616_ _5857_/A2 hold637/I _5521_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6404_ _7202_/Q _6272_/Z _6275_/Z _7040_/Q _6296_/Z _7162_/Q _6408_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold922 _5778_/Z _7119_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold900 _7094_/Q hold900/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold911 _5813_/Z _7150_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3547_ _3485_/Z _3523_/Z _3960_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold955 _6957_/Q hold955/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6335_ _6554_/A1 _6335_/A2 _6335_/A3 _6335_/A4 _6335_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold933 _5760_/Z _7103_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold944 _7095_/Q hold944/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_834 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold977 _5787_/Z _7127_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold966 _7037_/Q hold966/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold988 _6870_/Q hold988/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_0_107 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold999 _7282_/Q hold999/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3478_ _3478_/I0 hold10/Z hold21/I hold11/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_6266_ _6300_/A2 _6533_/A4 _6285_/A2 _6302_/A4 _6266_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_88_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5217_ _5460_/A1 _5460_/A4 _5224_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6197_ _6722_/Q _5987_/Z _6015_/Z _6841_/Q _6198_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5148_ _5147_/Z _5139_/Z _5148_/A3 _5470_/A3 _5148_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5079_ _5079_/A1 _5258_/C _5086_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_85_987 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet563_202 net563_246/I _7023_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_213 net563_248/I _7012_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_181_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_246 net563_246/I _6979_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_235 net613_281/I _6990_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_224 net613_285/I _7001_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_181_745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_797 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_206 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_453 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_467 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4450_ _4607_/A1 _4451_/B _4451_/C _5356_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_145_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold207 _7117_/Q hold207/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_129_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4381_ _4472_/B _4501_/B _4460_/B _4436_/B _4381_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3401_ _3401_/I _5420_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_8
Xhold229 _5838_/Z _7173_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold218 _7034_/Q hold218/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_153_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3332_ _4402_/B _4489_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_125_683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6120_ _7017_/Q _5971_/Z _6005_/Z _7041_/Q _6124_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_98_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ _6051_/A1 _6051_/A2 _6051_/B1 _5991_/Z _6052_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_5002_ _4411_/Z _5258_/B2 _5002_/A3 _5002_/A4 _5002_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_112_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_612 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_751 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_188 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6953_ hold50/Z _7238_/RN _6953_/CLK hold49/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5904_ _7224_/Q _5903_/Z _5904_/B _5905_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_6884_ _6884_/D _7297_/RN _6884_/CLK _6884_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_35_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5835_ hold62/Z hold126/Z _5838_/S _5835_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5766_ hold234/Z hold2/Z _5766_/S _5766_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4717_ _5222_/A1 _4716_/Z _5223_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5697_ hold62/Z hold240/Z _5700_/S _5697_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4648_ _4648_/A1 _4648_/A2 _4648_/B _5356_/C _5438_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_163_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold730 _5837_/Z _7172_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_107_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4579_ _4380_/Z _4579_/A2 _4451_/B _4451_/C _5345_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_162_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold763 _6778_/Q hold763/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold752 _4330_/Z _6837_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold741 _6884_/Q hold741/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7298_ _7298_/D _6650_/Z _7303_/CLK _7298_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold796 _4255_/Z _6770_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xnet513_154 net513_159/I _7071_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6318_ _7199_/Q _6272_/Z _6293_/Z _7151_/Q _6318_/C _6322_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold774 _5531_/Z _6902_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold785 _6708_/Q hold785/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xnet513_165 net563_221/I _7060_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_176 net663_329/I _7049_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet513_198 net413_81/I _7027_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_187 net413_57/I _7038_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6249_ _7126_/Q _6247_/Z _6248_/Z _7068_/Q _6259_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_130_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2979 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_572 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_417 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_913 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_486 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold90 hold90/I hold90/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_75_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3950_ _6726_/Q _4188_/A1 _3950_/B1 _6724_/Q _3950_/C1 _6843_/Q _3953_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_72_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3881_ _7037_/Q _5683_/A1 _5674_/A1 _7029_/Q _3881_/C _3884_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_176_347 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet763_419 net763_419/I _6755_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5620_ hold6/Z _3542_/Z hold38/Z hold11/Z _5628_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xnet763_408 net763_441/I _6766_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5551_ hold86/Z hold306/Z _5556_/S _5551_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4502_ _4504_/B _4504_/C _5072_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_145_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5482_ _5482_/A1 _5482_/A2 _5483_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7221_ _7221_/D _7221_/RN _7221_/CLK _7221_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4433_ _4648_/A1 _4648_/A2 _4638_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_104_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4364_ _4460_/B _4436_/B _5315_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_99_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_331 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7152_ _7152_/D _7297_/RN _7152_/CLK _7152_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_3315_ _6834_/Q _4900_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_98_364 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7083_ hold48/Z _7260_/RN _7083_/CLK hold47/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6103_ hold70/I _5965_/Z _6014_/Z _6960_/Q _6106_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4295_ _6566_/I0 _6803_/Q _4300_/S _6803_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6034_ _7029_/Q _5999_/Z _6014_/Z _6957_/Q _6000_/Z _7127_/Q _6035_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_6_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_795 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_412 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1508 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6936_ _6936_/D _7297_/RN _6936_/CLK _6936_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XPHY_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6867_ _6867_/D _7219_/RN _6867_/CLK _6867_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6798_ _6798_/D _7265_/CLK _6798_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5818_ hold29/Z hold302/Z _5820_/S _5818_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5749_ _5857_/A3 _5821_/A3 _3537_/Z _5520_/C _5757_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_22_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold560 _6767_/Q hold560/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold571 _7072_/Q hold571/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold593 _5870_/Z _7201_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_103_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_130 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold582 _6742_/Q hold582/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_181_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_401 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2721 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_426 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_448 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_380 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_225 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4080_ input85/Z input58/Z _7300_/Q _4080_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4982_ _4997_/B _4495_/Z _5263_/A2 _4436_/B _4982_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_63_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3933_ _7222_/Q _5528_/S _3933_/B1 _6785_/Q _3933_/C _3938_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_6721_ _6721_/D input75/Z _6721_/CLK _6721_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_23_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3864_ _6723_/Q _4182_/A1 _3946_/A2 _6721_/Q input12/Z _3913_/A2 _3868_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_32_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6652_ _7193_/RN _6652_/A2 _6652_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_176_155 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5603_ hold113/Z hold397/Z hold39/Z _6964_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6583_ _6583_/A1 _4313_/Z _6583_/B _6584_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_176_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3795_ _3795_/A1 _3790_/Z _3794_/Z _3795_/A4 _3795_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5534_ hold946/Z hold271/Z _5535_/S _5534_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5465_ _5465_/A1 _5170_/Z _4882_/Z _4881_/Z _5465_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_117_255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7204_ _7204_/D _7221_/RN _7204_/CLK _7204_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4416_ _4456_/B _5051_/S _5104_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_105_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5396_ _5396_/A1 _5395_/Z _5434_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_132_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7135_ _7135_/D _7210_/RN _7135_/CLK _7135_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_28_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4347_ _5520_/C _3529_/Z _5513_/A3 _5821_/A3 _4349_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7066_ _7066_/D _7237_/RN _7066_/CLK _7066_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_140_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_645 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4278_ _4103_/I hold799/Z _4279_/S _4278_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_678 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6017_ _7167_/Q _6006_/Z _6030_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_2006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/Z _3340__1/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6919_ _6919_/D _7258_/RN _6919_/CLK _6919_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_74_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1349 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_604 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_637 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_501 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold390 _5732_/Z _7078_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_150 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3252 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_634 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1872 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3580_ _3505_/Z _3509_/Z _5575_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_182_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5250_ _5250_/A1 _5247_/Z _5248_/Z _5250_/A4 _5251_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_154_394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_883 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4201_ _4200_/Z hold765/Z _4211_/S _4201_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_13__1359_ net413_58/I net413_56/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5181_ _5127_/Z _5181_/A2 _5321_/A1 _5242_/A3 _5181_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_68_301 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_868 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4132_ hold52/Z hold471/Z _4136_/S _4132_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4063_ _6747_/Q input3/Z input1/Z _4063_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_1023 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4965_ _5464_/A1 _4908_/Z _5073_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_145_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6704_ _6704_/D _7221_/RN _6704_/CLK _6704_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3916_ _7150_/Q _3916_/A2 _3916_/B1 _6878_/Q _4274_/A1 _6787_/Q _3919_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_33_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_291 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4896_ _4554_/Z _4892_/B _4897_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_138_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6635_ _7237_/RN _4064_/S _6635_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_149_177 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3847_ _3552_/Z _3653_/Z _4170_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3778_ input37/Z _4244_/S _3948_/C1 input63/Z _3797_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6566_ _6566_/I0 _7264_/Q _6571_/S _7264_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5517_ _5821_/A3 _3533_/Z hold637/Z _5520_/C _5518_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_105_203 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6497_ _7035_/Q _6269_/Z _6273_/Z _6979_/Q _6498_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_161_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5448_ _5448_/A1 _5483_/A2 _5448_/A3 _5463_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_154_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5379_ _5469_/A1 _5379_/A2 _5377_/Z _5379_/A4 _5379_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_120_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_792 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7118_ _7118_/D _7210_/RN _7118_/CLK _7118_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_102_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7049_ _7049_/D _7260_/RN _7049_/CLK _7049_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_86_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4073__5 _4073__9/I _7220_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1157 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_418 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_397 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3082 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3071 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3093 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_982 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1680 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ _5302_/B _5099_/A1 _4703_/Z _5226_/C _4750_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xclkbuf_leaf_0__1359_ net713_387/I net763_441/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_186_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4681_ _5420_/A3 _3402_/I _4456_/B _4681_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_3701_ _3701_/A1 _3701_/A2 _3701_/A3 _3701_/A4 _3701_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_186_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6420_ _6420_/I _6421_/I1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_1057 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3632_ _3632_/I _3633_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_607 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6351_ _6351_/I _6352_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5302_ _4536_/Z _5283_/B _5302_/B _5303_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_3563_ _3537_/Z _3542_/Z _5758_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_143_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6282_ _6282_/A1 _6282_/A2 _7232_/Q _6452_/A4 _6282_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3494_ _3653_/A1 hold338/Z _5857_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_143_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_386 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5233_ _5233_/A1 _4757_/I _5156_/B _5233_/A4 _5404_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5164_ _5315_/A1 _5315_/A2 _5287_/B _4784_/Z _5467_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_64_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4115_ hold14/Z _7276_/Q hold21/I hold15/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
XFILLER_151_1033 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5095_ _5278_/C _5302_/B _4784_/Z _4716_/Z _4697_/Z _5460_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_69_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_315 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4046_ _4046_/I _6832_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_294 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_167 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_229 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ _7231_/Q _6117_/A4 _6014_/A2 _7229_/Q _5997_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4948_ _4948_/A1 _4945_/Z _4946_/Z _4947_/Z _4953_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_177_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4879_ _5315_/A2 _4524_/Z _4546_/Z _4820_/Z _4879_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_71_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6618_ _7237_/RN _6656_/A2 _6618_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_71_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6549_ _6846_/Q _6235_/Z _6243_/Z _6842_/Q _6265_/Z _6840_/Q _6554_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_133_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput270 _6885_/Q pll_sel[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_88_941 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput292 _6687_/Q pll_trim[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput281 _6669_/Q pll_trim[19] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_87_462 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_348 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_743 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_705 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_860 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5920_ _7229_/Q _6210_/B _5920_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_111_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_1004 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5851_ hold86/Z hold648/Z _5856_/S _5851_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4802_ _5453_/A4 _5420_/A3 _5456_/A1 _5130_/B1 _5129_/A2 _5389_/A1 _4803_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_21_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5782_ hold29/Z hold59/Z _5784_/S hold60/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4733_ _4733_/A1 _4729_/Z _4731_/Z _4732_/Z _4739_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_175_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4664_ _4664_/A1 _4664_/A2 _4663_/Z _4670_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6403_ _7114_/Q _6240_/Z _6403_/B _6408_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_31_1040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4595_ _5190_/A2 _5364_/B _4568_/Z _5435_/A2 _4595_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_135_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3615_ _5857_/A2 _5857_/A3 hold38/I _3477_/Z _3866_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold912 _6682_/Q hold912/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold901 _5750_/Z _7094_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3546_ _3489_/I _3492_/Z _3904_/A4 _3904_/A2 _3546_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold934 _7215_/Q hold934/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6334_ _7045_/Q _6241_/Z _6268_/Z _6949_/Q _6274_/Z _7215_/Q _6335_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold923 _7143_/Q hold923/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold945 _5751_/Z _7095_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6265_ _6302_/A3 _6533_/A4 _6285_/A2 _6302_/A4 _6265_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold956 _6925_/Q hold956/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold978 _6973_/Q hold978/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold989 _6874_/Q hold989/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold967 _5685_/Z _7037_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3477_ hold134/Z hold9/Z hold21/Z _3477_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_5216_ _4697_/Z _5310_/A2 _5460_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_131_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6196_ _6712_/Q _6002_/Z _6003_/Z _6714_/Q _6198_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5147_ _4842_/Z _5147_/A2 _5147_/A3 _5147_/A4 _5147_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_130_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_624 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5078_ _5324_/A1 _5078_/A2 _5263_/A4 _5263_/A2 _5337_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_72_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4029_ _4029_/A1 _4029_/A2 _4391_/A3 _4391_/A4 _4031_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_38_893 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_649 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet563_203 net763_425/I _7022_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_154_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet563_214 net563_215/I _7011_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_247 net413_81/I _6978_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_225 net563_225/I _7000_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_236 net813_485/I _6989_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold208 _5775_/Z _7117_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_8_786 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3400_ _3400_/I _6601_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4380_ _4853_/A1 _5270_/A1 _5170_/A2 _4380_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_171_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold219 _5681_/Z _7034_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3331_ _7237_/Q _6302_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XTAP_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6050_ _7152_/Q _5960_/Z _5965_/Z _6700_/Q _5969_/Z _7120_/Q _6053_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XTAP_557 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5001_ _5000_/Z _5001_/A2 _5001_/B _6859_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_100_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_568 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_579 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6952_ hold80/Z _7260_/RN _6952_/CLK hold79/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5903_ _5901_/B _5902_/Z _7223_/Q _5903_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_6883_ _6883_/D _7297_/RN _6883_/CLK _6883_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5834_ hold52/Z hold296/Z _5838_/S _5834_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5765_ hold341/Z hold15/Z _5766_/S _5765_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_754 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4716_ _5420_/A2 _4835_/A2 _4456_/B _3401_/I _4716_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5696_ hold52/Z hold345/Z _5700_/S _5696_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4647_ _5038_/A1 _5475_/A3 _5439_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_148_798 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold720 _4337_/Z _6842_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4578_ _5464_/A1 _5438_/C _5346_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold753 _6761_/Q hold753/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_144_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_824 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6317_ _7135_/Q _6253_/Z _6296_/Z _7159_/Q _6322_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold764 _4264_/Z _6778_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold742 _5505_/Z _6884_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold731 _6723_/Q hold731/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold775 _6738_/Q hold775/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_143_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet513_155 _4073__20/I _7070_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_166 _4073__21/I _7059_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3529_ hold11/Z _3552_/A2 _3484_/Z hold32/Z _3529_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold786 _4162_/Z _6708_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7297_ _7297_/D _7297_/RN _7297_/CLK _7297_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
Xnet513_177 net563_221/I _7048_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold797 _6714_/Q hold797/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6248_ _7236_/Q _6484_/A2 _6452_/A4 _6302_/A4 _6248_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_77_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet513_199 net563_246/I _7026_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_188 net513_188/I _7037_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6179_ _7117_/Q _5984_/Z _5997_/Z _7101_/Q _7075_/Q _5980_/Z _6180_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_76_218 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_240 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_785 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2936 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2947 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_529 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_584 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_461 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold80 hold80/I hold80/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_36_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold91 hold91/I hold91/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_21_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_698 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3880_ _3880_/I _3881_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_43_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet763_409 net763_409/I _6765_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5550_ hold271/Z hold831/Z _5556_/S _5550_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4501_ _4853_/A1 _4884_/A1 _4501_/B _4504_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_5481_ _4944_/Z _5245_/Z _5481_/B1 _4951_/Z _5481_/C _5482_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_129_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4432_ _4460_/B _4376_/Z _4648_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7220_ _7220_/D _7221_/RN _7220_/CLK _7220_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_126_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4363_ _4460_/B _4436_/B _4363_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_116_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7151_ _7151_/D _7219_/RN _7151_/CLK _7151_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_112_142 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3314_ _6950_/Q _3994_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
X_7082_ hold69/Z _7238_/RN _7082_/CLK hold68/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6102_ hold79/I _5958_/Z _5999_/Z _7032_/Q _6102_/C _6106_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4294_ _6565_/I0 _6802_/Q _4300_/S _6802_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_495 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6033_ _7061_/Q _5985_/Z _5997_/Z _7095_/Q _6037_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_100_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6935_ _6935_/D _7221_/RN _6935_/CLK _6935_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_81_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_298 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6866_ _6866_/D _7219_/RN _6866_/CLK _6866_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_22_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_197 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6797_ _6797_/D _7265_/CLK _6797_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5817_ hold62/Z hold146/Z _5820_/S _5817_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5748_ hold2/Z hold374/Z _5748_/S _5748_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_509 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5679_ hold246/Z hold62/Z _5682_/S _5679_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold550 _5533_/Z _6903_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold561 _4251_/Z _6767_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold572 _5724_/Z _7072_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_9_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold594 _6924_/Q hold594/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold583 _4211_/Z _6742_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2711 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_134 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_284 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4981_ _5262_/A2 _5255_/A2 _4495_/Z _4497_/Z _4981_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_177_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3932_ _3932_/A1 _3533_/Z _3542_/Z _3932_/B _3933_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_16_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6720_ _6720_/D input75/Z _6720_/CLK _6720_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6651_ _7237_/RN _6657_/A2 _6651_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
Xclkbuf_leaf_36__1359_ clkbuf_4_8_0__1359_/Z _4073__8/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3863_ _6973_/Q _3923_/A2 _3959_/C1 _7183_/Q _3869_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xclkbuf_leaf_116__1359_ net613_293/I net813_495/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6582_ _6834_/Q _6582_/A2 _6582_/B1 _6835_/Q _6836_/Q _6582_/C2 _6583_/B VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_165_819 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5602_ hold6/Z _3515_/Z hold38/Z hold11/Z hold39/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xclkbuf_leaf_99__1359_ clkbuf_4_5_0__1359_/Z net763_425/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_164_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5533_ hold549/Z hold86/Z _5535_/S _5533_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3794_ _3794_/A1 _3794_/A2 _3794_/A3 _3794_/A4 _3794_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_118_735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5464_ _5464_/A1 _4659_/Z _4675_/Z _5464_/B _5465_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
X_4415_ _5385_/A1 _5045_/C _4415_/B _5211_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5395_ _5395_/A1 _4991_/C _5428_/A2 _5395_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_132_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7203_ _7203_/D _7219_/RN _7203_/CLK _7203_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_154_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7134_ _7134_/D _7297_/RN _7134_/CLK _7134_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4346_ hold271/Z hold904/Z _4346_/S _4346_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_1042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4277_ _3509_/Z _5520_/C _5513_/A3 _5857_/A2 _4279_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_7065_ _7065_/D _7297_/RN _7065_/CLK _7065_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_6016_ _7013_/Q _5971_/Z _6031_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_2007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2029 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6918_ _6918_/D _7258_/RN _6918_/CLK _6918_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_74_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6849_ _6849_/D _7193_/RN _6849_/CLK _6849_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_168_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_178 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_381 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_328 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold380 _5892_/Z _7221_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_89_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold391 _7101_/Q hold391/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_105_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_184 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3253 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet813_490 net813_491/I _6675_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_187_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1884 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1895 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1026 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4200_ hold312/Z hold86/Z _4210_/S _4200_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5180_ _5180_/A1 _5180_/A2 _5180_/A3 _5211_/C _5185_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_111_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_12_0__1359_ clkbuf_0__1359_/Z net613_299/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4131_ hold86/Z hold475/Z _4136_/S _4131_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4062_ _4061_/Z _3337_/I _7299_/Q _4062_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_1021 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_582 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4964_ _4421_/Z _4908_/Z _4966_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_52_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6703_ _6703_/D _7237_/RN _6703_/CLK _6703_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3915_ _3915_/A1 _3915_/A2 _3915_/A3 _3915_/A4 _3915_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4895_ _4886_/Z _4887_/Z _4891_/Z _4895_/A4 _4898_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6634_ _7237_/RN _6657_/A2 _6634_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_165_616 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_189 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3846_ _3540_/Z _3552_/Z _3939_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_644 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3777_ _7176_/Q _3945_/A2 _5532_/A1 _6903_/Q _3797_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6565_ _6565_/I0 _7263_/Q _6571_/S _7263_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6496_ _6947_/Q _6245_/Z _6288_/Z _7125_/Q _6498_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5516_ _4103_/I hold757/Z _5516_/S _5516_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5447_ _5447_/A1 _5447_/A2 _5448_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_160_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_259 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5378_ _5425_/A2 _5425_/A3 _5379_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_87_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7117_ _7117_/D _7237_/RN _7117_/CLK _7117_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_102_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4329_ _3509_/Z _5839_/A3 _5513_/A3 _5520_/C _4331_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_59_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7048_ _7048_/D _7297_/RN _7048_/CLK _7048_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_47_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4073__6 _4073__8/I _7219_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_808 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_118 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_270 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3083 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3061 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3050 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_777 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_585 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3094 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2393 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3700_ _6686_/Q _3945_/C2 _5683_/A1 _7040_/Q _3701_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_175_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4680_ _4414_/Z _4452_/Z _4666_/Z _5395_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_147_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3631_ _6938_/Q _3910_/A2 _3954_/A2 _6994_/Q _7204_/Q _3955_/A2 _3632_/I VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_174_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6350_ _7128_/Q _6247_/Z _6297_/Z _6700_/Q _6351_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3562_ _3507_/Z _3537_/Z _3927_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_155_682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5301_ _5301_/I _6861_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_681 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3493_ _3493_/I0 hold337/Z hold21/Z _3493_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_6281_ _6484_/A3 _6256_/Z _6272_/Z _6274_/Z _6281_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_170_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_207 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5232_ _5414_/A2 _4752_/Z _5233_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_88_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5163_ _5356_/A1 _4650_/Z _5231_/A2 _5468_/A1 _5166_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_112_1007 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4114_ hold29/Z hold101/Z _4118_/S _4114_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_1048 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5094_ _5328_/A1 _5389_/A1 _5094_/B _5094_/C _5347_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_83_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4045_ _6832_/Q _4097_/A1 _4045_/B1 _6826_/Q _4046_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_84_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ _7231_/Q _6210_/B _6014_/A2 _7229_/Q _5996_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_80_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4947_ _5072_/A4 _4903_/Z _4421_/Z _4500_/Z _4947_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_71_1024 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_791 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4878_ _4997_/C _4878_/A2 _3401_/I _3402_/I _4878_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_138_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6617_ _7237_/RN _6656_/A2 _6617_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_137_115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3829_ _3537_/Z hold630/Z _4161_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_986 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6548_ _6548_/A1 _6548_/A2 _6548_/A3 _6547_/Z _6548_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_161_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6479_ _7189_/Q _6282_/Z _6492_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_121_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput260 _6891_/Q pll_bypass VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput271 _6682_/Q pll_trim[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_160_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_835 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput282 _6683_/Q pll_trim[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput293 _6688_/Q pll_trim[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_741 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_474 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_628 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_722 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_969 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_468 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_994 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_205 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_183 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_901 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_975 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_477 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5850_ hold271/Z hold984/Z _5856_/S _5850_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4801_ _5312_/A2 _5312_/A4 _5456_/A1 _5220_/B2 _4801_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_62_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5781_ hold62/Z hold209/Z _5784_/S _5781_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4732_ _4765_/A1 _4510_/Z _5302_/B _5099_/A2 _4732_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_174_221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4663_ _4411_/Z _5214_/A2 _5172_/B _5165_/A4 _4663_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_147_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6402_ _7130_/Q _6484_/A2 _6484_/A3 _6533_/A4 _6403_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3614_ _3505_/Z _3533_/Z _3770_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4594_ _5190_/A2 _5435_/A2 _5389_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold913 _4129_/Z _6682_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold902 _7166_/Q hold902/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_143_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold946 _6904_/Q hold946/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3545_ _3485_/Z _3521_/Z _3959_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold935 _5886_/Z _7215_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6333_ _7207_/Q _6256_/Z _6261_/Z _6957_/Q _6285_/Z _7191_/Q _6335_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold924 _5805_/Z _7143_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_685 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3476_ _3476_/I _3478_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold957 _5559_/Z _6925_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold979 _5613_/Z _6973_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold968 _7111_/Q hold968/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_0_109 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6264_ _6956_/Q _6261_/Z _6263_/Z _6932_/Q _6262_/Z _6964_/Q _6271_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_115_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5215_ _4698_/B _5403_/A2 _5215_/B _5215_/C _5316_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_9_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6195_ _6824_/Q _5988_/Z _6019_/Z _6853_/Q _6198_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5146_ _4546_/Z _5364_/B _4586_/Z _4598_/Z _4568_/Z _5147_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_97_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_636 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5077_ _4973_/Z _5078_/A2 _5258_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_111_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4028_ input97/Z input96/Z input99/Z input98/Z _4028_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_56_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5979_ _6002_/A2 _6021_/A2 _6210_/A2 _7227_/Q _5979_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_139_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_204 net563_212/I _7021_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet563_215 net563_215/I _7010_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_226 net613_255/I _6999_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_237 net413_91/I _6988_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_153_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet563_248 net563_248/I _6977_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_630 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_632 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_803 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_825 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_814 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_313 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_469 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_732 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1055 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold209 _7122_/Q hold209/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_152_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3330_ _7236_/Q _6285_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_4_971 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _5000_/A1 _5000_/A2 _5000_/A3 _5000_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_112_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_558 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_0_0__1359_ clkbuf_0__1359_/Z net713_387/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_85_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_411 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_569 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6951_ hold78/Z _7238_/RN _6951_/CLK hold77/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
X_5902_ _5911_/A1 _6746_/Q _7225_/Q _5902_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_6882_ _6882_/D _7193_/RN _6882_/CLK _6882_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5833_ hold86/Z hold608/Z _5838_/S _5833_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5764_ hold314/Z hold29/Z _5766_/S _5764_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4715_ _4835_/A2 _5087_/A1 _5328_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5695_ hold86/Z hold660/Z _5700_/S _5695_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4646_ _4648_/A1 _4648_/A2 _4648_/B _5475_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_4577_ _5002_/A3 _5002_/A4 _5083_/B _5003_/A2 _5043_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_162_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold721 _6852_/Q hold721/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold710 _4148_/Z _6697_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold754 _4243_/Z _6761_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_150_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1002 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6316_ _7167_/Q _5948_/Z _6245_/Z _6941_/Q _6263_/Z _6933_/Q _6329_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xhold732 _4184_/Z _6723_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold743 _6725_/Q hold743/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold765 _6737_/Q hold765/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold776 _4203_/Z _6738_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold787 _6759_/Q hold787/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_118_1035 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_696 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_173 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet513_167 net613_297/I _7058_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_302 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3528_ _3525_/Z _3527_/Z _3935_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xnet513_156 _4073__51/I _7069_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7296_ _7296_/D _7297_/RN _7296_/CLK _7296_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3459_ hold85/Z hold270/Z _3460_/S _7285_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6247_ _7236_/Q _6484_/A2 _6533_/A4 _6302_/A4 _6247_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xnet513_178 net763_419/I _7047_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_335 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet513_189 _4073__51/I _7036_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold798 _4171_/Z _6714_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_130_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6178_ _7157_/Q _5960_/Z _5965_/Z _6705_/Q _6006_/Z _7173_/Q _6180_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_29_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5129_ _5420_/A2 _5129_/A2 _5129_/A3 _3401_/I _5129_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_69_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2904 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2937 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2959 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1015 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_580 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_230 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold81 hold81/I hold81/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold92 hold92/I hold92/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold70 hold70/I hold70/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_90_222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4500_ _4759_/A2 _4759_/A3 _4500_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_129_265 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5480_ _5480_/A1 _5480_/A2 _5480_/A3 _5479_/Z _5480_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4431_ _4414_/Z _4421_/Z _5393_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_1 _4124_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4362_ _5299_/C _6859_/Q _5001_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_125_482 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7150_ _7150_/D _7193_/RN _7150_/CLK _7150_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_3313_ _6830_/Q _4038_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7081_ _7081_/D _7219_/RN _7081_/CLK _7081_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4293_ _6564_/I0 _6801_/Q _4300_/S _6801_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6101_ _6101_/A1 _6101_/A2 _6101_/A3 _6101_/A4 _6101_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xclkbuf_leaf_59__1359_ clkbuf_4_15_0__1359_/Z net763_413/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_140_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_316 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6032_ _7069_/Q _5980_/Z _6003_/Z _7159_/Q _6037_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xclkbuf_leaf_139__1359_ net563_220/I net813_482/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6934_ _6934_/D _7258_/RN _6934_/CLK _6934_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_54_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6865_ _6865_/D _7279_/RN _7230_/CLK hold31/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5816_ hold52/Z hold539/Z _5820_/S _5816_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6796_ _6796_/D _7265_/CLK _6796_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5747_ hold15/Z hold446/Z _5748_/S _5747_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_388 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_235 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5678_ hold286/Z hold52/Z _5682_/S _5678_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4629_ _5190_/A2 _4604_/Z _5387_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_163_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_279 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold540 _5816_/Z _7153_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold551 _7081_/Q hold551/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold562 _6773_/Q hold562/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_1_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7279_ _7279_/D _7279_/RN _7279_/CLK hold17/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_132_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold595 _5558_/Z _6924_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_666 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold573 _7110_/Q hold573/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold584 _7086_/Q hold584/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_106_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_561 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2745 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2756 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_828 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2789 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_731 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput160 wb_rstn_i _7279_/RN VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_91_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_458 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4980_ _4998_/A2 _5262_/A2 _5255_/A2 _5442_/A2 _4980_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xnet413_100 net513_191/I _7125_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3931_ _7052_/Q _5701_/A1 _5536_/A1 _6906_/Q _3932_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_177_647 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6650_ _7237_/RN _6657_/A2 _6650_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_149_338 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_305 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3862_ _6957_/Q _3957_/A2 _3928_/C1 _6823_/Q _3925_/B1 _6825_/Q _3869_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_31_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6581_ _6581_/I0 _7270_/Q _6602_/S _7270_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5601_ hold2/Z _6963_/Q hold12/Z hold13/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_894 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5532_ _5532_/A1 hold18/Z _5535_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_9_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3793_ _7136_/Q _3951_/A2 _3924_/A2 _6966_/Q _3794_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_118_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_717 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5463_ _5463_/A1 _5463_/A2 _5485_/A2 _5463_/B2 _5463_/C _5474_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_8_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4414_ _4397_/Z _4491_/B _5003_/A2 _4414_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_5394_ _4892_/B _5394_/A2 _5428_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_105_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7202_ _7202_/D _7210_/RN _7202_/CLK _7202_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_7133_ _7133_/D _7237_/RN _7133_/CLK _7133_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_114_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4345_ _4103_/I hold813/Z _4346_/S _4345_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_675 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7064_ _7064_/D _7297_/RN _7064_/CLK _7064_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4276_ hold733/Z hold271/Z _4276_/S _4276_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6015_ _7228_/Q _6211_/B1 _6015_/A3 _6210_/A2 _6015_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_100_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_274 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2019 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_609 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1307 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6917_ _6917_/D _7258_/RN _6917_/CLK _6917_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_161_1003 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_973 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6848_ _6848_/D _7210_/RN _6848_/CLK _6848_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_168_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1047 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6779_ hold87/Z _7238_/RN _6779_/CLK _6779_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_6_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_513 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1072 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold381 _7165_/Q hold381/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_105_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold370 _6689_/Q hold370/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_131_260 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold392 _5757_/Z _7101_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_42__1359_ net413_53/I net413_97/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_306 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_122__1359_ net613_293/I net563_221/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3221 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3210 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_491 net813_491/I _6674_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_480 net813_483/I _6685_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1874 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1016 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_896 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4130_ hold271/Z hold950/Z _4136_/S _4130_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_591 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4061_ _4060_/Z input38/Z _7301_/Q _4061_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4963_ _4963_/A1 _4960_/Z _4961_/Z _4962_/Z _4966_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_145_1009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6702_ hold71/Z _7238_/RN _6702_/CLK hold70/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3914_ _7102_/Q _5758_/A1 _3914_/B1 _6876_/Q _3915_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_189_293 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4894_ _4894_/A1 _4893_/Z _4895_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6633_ _7219_/RN _6652_/A2 _6633_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_164_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3845_ _7061_/Q _3927_/B1 _3955_/B1 _6848_/Q _3895_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_177_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3776_ _3773_/Z _3776_/A2 _3776_/A3 _3776_/A4 _3776_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6564_ _6564_/I0 _7262_/Q _6571_/S _7262_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_801 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6495_ _7051_/Q _6241_/Z _6251_/Z _6987_/Q _6268_/Z hold91/I _6498_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_5515_ _3485_/Z _5857_/A3 _5839_/A3 _5520_/C _5516_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5446_ _5446_/A1 _5446_/A2 _5447_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_161_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5377_ _5377_/A1 _5290_/Z _5377_/A3 _5377_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
X_7116_ _7116_/D _7221_/RN _7116_/CLK _7116_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_113_271 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4328_ hold271/Z hold864/Z _4328_/S _4328_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7047_ _7047_/D _7258_/RN _7047_/CLK _7047_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_101_444 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4259_ hold29/Z hold124/Z _4261_/S _4259_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_369 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1115 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4073__7 _4073__7/I _7218_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1148 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_122 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_436 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_311 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_626 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3040 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3062 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3084 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3095 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_219 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2394 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_781 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_447 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3630_ _3630_/A1 _3630_/A2 _3630_/A3 _3630_/A4 _3630_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_30_976 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3561_ _3533_/Z _3560_/Z _3913_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_183_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5300_ _5242_/Z _5266_/Z _5300_/A3 _5299_/C _6861_/Q _5301_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_3492_ _3491_/I _3307_/I hold21/Z _3492_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_6280_ _6245_/Z _6262_/Z _6263_/Z _6279_/Z _6287_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_5_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5231_ _5291_/B _5231_/A2 _5231_/B _5231_/C _5314_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_97_910 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5162_ _5165_/A2 _5287_/B _5315_/A2 _5315_/A1 _5467_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_111_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_943 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4113_ hold28/Z _7275_/Q hold21/Z hold29/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_5093_ _5359_/A1 _4568_/Z _5218_/B _5303_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_151_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4044_ _4044_/I _6732_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_169 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_862 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_512 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5995_ _7052_/Q _5924_/Z _5994_/I _7134_/Q _5995_/C _6009_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_4946_ _4500_/Z _4903_/Z _5072_/A4 _4666_/Z _4946_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_178_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_921 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_263 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_926 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4877_ _4651_/Z _4483_/B _4422_/Z _4683_/Z _4877_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6616_ _7237_/RN _6656_/A2 _6616_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_165_414 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3828_ _3535_/Z _3537_/Z _3956_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6547_ _6547_/A1 _6547_/A2 _6542_/Z _6546_/Z _6547_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_20_497 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_812 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3759_ _3759_/A1 _3759_/A2 _3747_/Z _3758_/Z _3759_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6478_ _7043_/Q _6275_/Z _6486_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_3_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5429_ _4898_/C _4991_/C _5392_/B _4893_/Z _5429_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_134_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput261 _6877_/Q pll_dco_ena VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput250 _4092_/ZN pad_flash_csb_oe VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput294 _6689_/Q pll_trim[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput272 _6676_/Q pll_trim[10] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput283 _6670_/Q pll_trim[20] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_59_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_915 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_954 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_464 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_653 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_366 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1068 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_196 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xload_slew349 hold6/Z _5520_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_93_423 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_840 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_575 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_1006 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4800_ _4675_/Z _4683_/Z _5130_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5780_ hold52/Z hold545/Z _5784_/S _5780_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4731_ _4765_/A1 _5302_/B _5099_/A2 _4716_/Z _4731_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XTAP_1490 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4662_ _5464_/A1 _4414_/Z _4659_/Z _4662_/B _4664_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_147_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_767 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3613_ _7074_/Q _3943_/A2 _3647_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_70_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6401_ _6401_/A1 _6401_/A2 _6401_/A3 _6401_/A4 _6401_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_174_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4593_ _4593_/A1 _5018_/B _4601_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_134_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold903 _5831_/Z _7166_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_31_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3544_ input51/Z _4210_/S _4244_/S input42/Z _3589_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold936 _7151_/Q hold936/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold914 _6700_/Q hold914/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6332_ _6981_/Q _6251_/Z _6254_/Z _7175_/Q _6332_/C _6335_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
Xhold925 _6667_/Q hold925/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3475_ _6660_/Q hold133/Z _6733_/Q _3476_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6263_ _7232_/Q _6533_/A2 _6452_/A4 _6282_/A2 _6263_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_116_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold947 _5534_/Z _6904_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold969 _5769_/Z _7111_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold958 _7199_/Q hold958/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_5214_ _5343_/A2 _5214_/A2 _5310_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_9_1043 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6194_ _6820_/Q _5979_/Z _5996_/Z _6708_/Q _6198_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_5145_ _4570_/Z _5145_/A2 _4878_/Z _5364_/B _4820_/Z _4821_/Z _5147_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai222_4
XFILLER_96_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5076_ _5464_/A1 _4905_/Z _4973_/Z _4700_/Z _5076_/C _5079_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_84_434 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4027_ _4027_/A1 _4027_/A2 _4031_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_38_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5978_ _5924_/Z _5975_/Z _5976_/Z _5977_/Z _5983_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_166_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4929_ _4929_/A1 _4928_/Z _4929_/A3 _4933_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_60_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_773 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_238 net613_258/I _6987_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_227 net763_422/I _6998_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_205 net763_425/I _7020_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_216 net663_329/I _7009_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_300 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xnet563_249 net413_89/I _6976_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_697 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_239 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_837 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_981 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_504 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_548 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_559 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_231 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_659 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_456 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6950_ _6950_/D _7238_/RN _6950_/CLK _6950_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_5901_ _5901_/A1 _5951_/A3 _5901_/B _5904_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_93_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6881_ _6881_/D _7193_/RN _6881_/CLK _6881_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_35_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5832_ hold271/Z hold982/Z _5838_/S _5832_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5763_ hold368/Z hold62/Z _5766_/S _5763_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4714_ _4709_/Z _4711_/Z _5305_/B _4714_/A4 _4727_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xclkbuf_leaf_19__1359_ net613_253/I net513_185/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_50_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5694_ hold271/Z hold962/Z _5700_/S _5694_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4645_ _4565_/Z _4641_/Z _5040_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_147_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4576_ _4549_/Z _4570_/Z _5192_/B _4576_/C _4584_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
Xhold700 _5567_/Z _6932_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold711 _6715_/Q hold711/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_162_258 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold755 _6755_/Q hold755/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3527_ _3552_/A2 _3484_/Z hold32/Z _3477_/Z _3527_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6315_ _7183_/Q _6282_/Z _6322_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_2_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold722 _4352_/Z _6852_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold733 _6788_/Q hold733/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold744 _4187_/Z _6725_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7295_ _7295_/D _6649_/Z _7304_/CLK _7295_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold766 _4201_/Z _6737_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold788 _4239_/Z _6759_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold777 _6866_/Q hold777/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xnet513_168 net713_390/I _7057_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet513_157 net513_185/I _7068_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3458_ hold51/Z hold85/Z _3460_/S _7286_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xnet513_179 net763_422/I _7046_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold799 _6789_/Q hold799/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_6246_ _7004_/Q _6243_/Z _6245_/Z _6940_/Q _6260_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_130_166 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3389_ _7229_/Q _5984_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_97_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6177_ _7109_/Q _5967_/Z _6177_/B _6180_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5128_ _5453_/A4 _5319_/A3 _5181_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2916 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5059_ _4700_/Z _5325_/B _5060_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_297 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_670 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2949 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_620 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_202 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_174 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold82 hold82/I hold82/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_48_478 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold71 hold71/I hold71/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold60 hold60/I hold60/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_75_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold93 hold93/I hold93/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_72_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_323 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_857 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_277 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4430_ _4402_/B _4026_/B _4026_/C _5083_/C _4997_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_145_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_2 _4130_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_995 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4361_ hold703/Z hold271/Z _4361_/S _4361_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6100_ _7016_/Q _5971_/Z _5988_/Z _6984_/Q _6005_/Z _7040_/Q _6101_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_3312_ _3312_/I _3428_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_879 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4292_ _6828_/Q _7279_/RN _4300_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_7080_ _7080_/D _7238_/RN _7080_/CLK _7080_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_141_998 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6031_ _6031_/A1 _6026_/Z _6030_/Z _6031_/A4 _6031_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_6_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_6__1359_ net713_387/I net413_71/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_66_242 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_264 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6933_ _6933_/D _7210_/RN _6933_/CLK _6933_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XPHY_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6864_ _6864_/D _7279_/RN _7230_/CLK hold9/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_133 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5815_ hold86/Z hold486/Z _5820_/S _5815_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6795_ _6795_/D _7269_/CLK _6795_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1051 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5746_ hold29/Z hold783/Z _5748_/S _5746_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5677_ hold412/Z hold86/Z _5682_/S _5677_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4628_ _4565_/Z _4624_/Z _5035_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xhold530 _5871_/Z _7202_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4559_ _5464_/A1 _4997_/C _5393_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold552 _5735_/Z _7081_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold563 _4258_/Z _6773_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold541 _6750_/Q hold541/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7278_ _7278_/D _7279_/RN _7279_/CLK _7278_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold596 _6911_/Q hold596/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_132_965 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold574 _5768_/Z _7110_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold585 _5741_/Z _7086_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xclkbuf_opt_4_1__1359_ clkbuf_opt_4_1__1359_/I net663_310/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_103_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6229_ _6220_/Z _6228_/Z _6555_/B1 _6168_/C _6555_/C _6230_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_103_199 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_540 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_990 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2746 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_919 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2757 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2768 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_289 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_317 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_523 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_145__1359_ net563_220/I _4073__2/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_154_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_940 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput161 wb_sel_i[0] _6572_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput150 wb_dat_i[2] _3395_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_562 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet413_101 net563_230/I _7124_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3930_ _7126_/Q _3930_/A2 _3930_/B1 _6841_/Q _4170_/A1 _6714_/Q _3938_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_45_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3861_ _7207_/Q _3960_/A2 _3955_/A2 _7199_/Q _3924_/A2 _6965_/Q _3869_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_32_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6580_ _6580_/A1 _4313_/Z _6580_/B _6581_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_158_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5600_ hold15/Z hold464/Z hold12/Z _6962_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3792_ _6990_/Q _3954_/A2 _3954_/B1 input22/Z _3794_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_157_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5531_ _4103_/I hold773/Z _5531_/S _5531_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7201_ _7201_/D _7221_/RN _7201_/CLK _7201_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_117_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5462_ _5404_/Z _5457_/Z _5461_/I _5463_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_5393_ _5393_/A1 _5393_/A2 _5393_/B1 _5045_/C _5433_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_4413_ _5209_/A3 _4397_/Z _5045_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_7132_ _7132_/D _7221_/RN _7132_/CLK _7132_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_28_1025 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4344_ _3529_/Z _3535_/Z _5520_/C _4346_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
X_7063_ _7063_/D _7221_/RN _7063_/CLK _7063_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_140_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6014_ _6210_/B _6014_/A2 _6210_/A2 _7229_/Q _6014_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_98_175 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_337 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4275_ hold927/Z _4103_/I _4276_/S _4275_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_158 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_595 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2009 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1319 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6916_ _6916_/D _7258_/RN _6916_/CLK _6916_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_6847_ _6847_/D _7210_/RN _6847_/CLK _6847_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_168_648 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6778_ _6778_/D _7260_/RN _6778_/CLK _6778_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_51_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_629 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5729_ hold821/Z _4103_/I _5730_/S _5729_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_320 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_236 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold360 _7055_/Q hold360/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_420 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold371 _4136_/Z _6689_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_117_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold382 _5829_/Z _7165_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold393 _7060_/Q hold393/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_120_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3222 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3211 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3200 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3255 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3244 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3233 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2510 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_692 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2554 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet813_492 net413_86/I _6673_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_481 net813_482/I _6684_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_470 net813_470/I _6695_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_489 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_567 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_707 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_1044 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1039 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_280 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_902 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4060_ _6748_/Q _6875_/Q _4064_/S _4060_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_407 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4962_ _4500_/Z _4906_/Z _5072_/A4 _4666_/Z _4962_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_64_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_261 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4893_ _5139_/A2 _5139_/A3 _4542_/Z _5172_/C _4893_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6701_ _6701_/D _7221_/RN _6701_/CLK _6701_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3913_ input11/Z _3913_/A2 _3913_/B1 _6892_/Q _3915_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_32_451 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_968 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_946 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6632_ _7193_/RN _6652_/A2 _6632_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_20_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3844_ _3529_/Z _3535_/Z _3955_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6563_ _6833_/D _7279_/RN _6571_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3775_ _7112_/Q _3917_/A2 _3913_/A2 input13/Z _3916_/A2 _7152_/Q _3776_/A3 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_118_534 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6494_ _7027_/Q _6235_/Z _6243_/Z _7011_/Q _6265_/Z _7003_/Q _6499_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_9_691 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5514_ _4103_/I hold761/Z _5514_/S _5514_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5445_ _4376_/Z _5255_/B _4972_/Z _5445_/B2 _5056_/B _5445_/C2 _5446_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_7115_ _7115_/D _7237_/RN _7115_/CLK _7115_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_5376_ _5291_/C _5376_/A2 _5468_/B1 _5376_/B2 _5376_/C _5377_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_99_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_283 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4327_ _4103_/I hold801/Z _4328_/S _4327_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4258_ hold62/Z hold562/Z _4261_/S _4258_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_957 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7046_ _7046_/D _7260_/RN _7046_/CLK _7046_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_170_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4189_ hold654/Z _4103_/I _4190_/S _4189_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_716 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4073__8 _4073__8/I _7217_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_635 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_415 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_813 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_375 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_209 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_740 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold190 _7067_/Q hold190/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_272 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_250 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_702 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3030 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3063 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3041 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3085 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3074 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2395 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_220 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1683 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_900 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1049 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_459 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3560_ hold338/Z _3496_/Z hold629/Z _3489_/I _3560_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_183_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3491_ _3491_/I _3493_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5230_ _4510_/Z _5414_/A2 _5230_/B _5231_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_170_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_687 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5161_ _5161_/A1 _5161_/A2 _5366_/A1 _5166_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_123_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5092_ _5092_/A1 _4705_/Z _5218_/B _4784_/Z _5303_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_84_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_646 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1066 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4112_ hold62/Z hold399/Z _4118_/S _4112_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4043_ _4043_/A1 _6732_/Q _6733_/Q _3409_/Z _4044_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_111_776 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_159 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5994_ _5994_/I _6051_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4945_ _4500_/Z _4903_/Z _5072_/A4 _5359_/A1 _4945_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4876_ _4650_/Z _4876_/A2 _4876_/B _4876_/C _4880_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_6615_ _7237_/RN _6656_/A2 _6615_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_177_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3827_ _3537_/Z _3540_/Z _3946_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_174_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3758_ _3758_/A1 _3751_/Z _3757_/Z _3758_/A4 _3758_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6546_ _6546_/A1 _6546_/A2 _6546_/A3 _6546_/A4 _6546_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_146_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_161 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_353 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6477_ _6971_/Q _6262_/Z _6499_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_3689_ _3689_/A1 _3657_/Z _3688_/Z _6569_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_5428_ _5381_/I _5428_/A2 _6577_/C _5428_/A4 _5428_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_0_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput240 _6750_/Q mgmt_gpio_out[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput251 _4080_/Z pad_flash_io0_do VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput262 _6878_/Q pll_div[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5359_ _5359_/A1 _4892_/B _5360_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_87_421 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput295 _6674_/Q pll_trim[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput273 _6677_/Q pll_trim[11] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput284 _6671_/Q pll_trim[21] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_58_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7029_ _7029_/D _7219_/RN _7029_/CLK _7029_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_59_156 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_938 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_621 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_172 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_903 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_977 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_671 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_524 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2192 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_905 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4730_ _4716_/Z _4728_/Z _5105_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_1491 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1480 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4661_ _4414_/Z _5038_/A1 _5359_/A1 _4557_/Z _4662_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_159_286 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_779 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6400_ _7210_/Q _6256_/Z _6263_/Z _6936_/Q _6401_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_3612_ _6680_/Q _3546_/Z _3625_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_4592_ _4565_/Z _4586_/Z _5018_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_156_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6331_ _6331_/I _6332_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xhold904 _6848_/Q hold904/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_846 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3543_ _3485_/Z _3542_/Z _4244_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold937 _5814_/Z _7151_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold915 _4152_/Z _6700_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold926 _4106_/Z _6667_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3474_ _4041_/B1 _6660_/Q _3981_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_142_153 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6262_ _6302_/A3 _5943_/S _7234_/Q _6533_/A2 _6262_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xhold959 _5868_/Z _7199_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold948 _7053_/Q hold948/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_838 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5213_ _4673_/Z _5124_/B _5213_/B _5213_/C _5454_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_6193_ _6193_/A1 _6193_/A2 _6193_/A3 _6193_/A4 _6193_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5144_ _4555_/C _5276_/C _5145_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_130_359 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_752 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_476 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5075_ _5255_/B _5051_/Z _5075_/B _5076_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_85_958 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4026_ _4402_/B _4483_/B _4026_/B _4026_/C _4412_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_65_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5977_ _6996_/Q _6211_/B1 _6021_/A2 _7227_/Q _5977_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4928_ _4376_/Z _5056_/C _5442_/A2 _5442_/A4 _4928_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_100_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_927 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4859_ _4614_/Z _5051_/S _5287_/B _4681_/Z _4859_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xnet563_206 net563_230/I _7019_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_228 net413_78/I _6997_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_217 net413_70/I _7008_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_239 net613_255/I _6986_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6529_ _6529_/I0 _7258_/Q _6555_/C _6529_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_131 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_186 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_304 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_774 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_863 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_849 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1073 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1038 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_960 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_295 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_266 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_120 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_602 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_730 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1014 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5900_ _5900_/A1 _5954_/A3 _5951_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_75_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6880_ _6880_/D _7297_/RN _6880_/CLK _6880_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_34_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_326 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_162 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5831_ _4103_/I hold902/Z _5838_/S _5831_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_505 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5762_ hold527/Z hold52/Z _5766_/S _5762_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_882 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4713_ _4713_/A1 _5094_/B _4691_/Z _4699_/Z _5305_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_147_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_908 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5693_ hold113/Z hold496/Z _5700_/S _5693_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4644_ _4644_/A1 _5038_/B _4643_/Z _4653_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_162_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_790 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4575_ _5281_/C _4539_/I _4551_/Z _5364_/B _5192_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_144_930 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_610 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold701 _6727_/Q hold701/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold712 _4172_/Z _6715_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7294_ _7294_/D _6648_/Z _7303_/CLK _7294_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3526_ _3552_/A2 _3484_/Z hold32/Z hold33/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_6314_ _7053_/Q _6299_/Z _6328_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xhold745 _6711_/Q hold745/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold734 _4276_/Z _6788_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold723 _6854_/Q hold723/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_157_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xnet513_158 net513_159/I _7067_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6245_ _7233_/Q _6533_/A2 _6452_/A4 _6279_/A3 _6245_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_116_676 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold756 _4231_/Z _6755_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold767 _6855_/Q hold767/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold778 _5492_/Z _6866_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3457_ hold61/Z hold51/Z _3460_/S _7287_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_112 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold789 _6692_/Q hold789/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xnet513_169 net813_467/I _7056_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_871 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3388_ _7230_/Q _6014_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_85_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6176_ _5991_/Z _6176_/A2 _6176_/B _6176_/C _6177_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_5127_ _5127_/A1 _5457_/A1 _5213_/B _5127_/A4 _5127_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5058_ _5058_/A1 _5055_/Z _5193_/A2 _5058_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_85_766 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2928 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2917 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2906 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4009_ _4009_/A1 _6744_/Q _6745_/Q _4010_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_84_287 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2939 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_310 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1076 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_516 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_370 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_749 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_932 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_999 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_700 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold50 hold50/I hold50/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold61 hold61/I hold61/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_152_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_392 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_25__1359_ clkbuf_4_8_0__1359_/Z net413_99/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_76_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_105__1359_ clkbuf_4_5_0__1359_/Z net613_285/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold72 hold72/I hold72/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_21_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold83 hold83/I hold83/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xclkbuf_leaf_88__1359_ clkbuf_4_13_0__1359_/Z net563_246/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_60_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold94 hold94/I hold94/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_91_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_181 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_657 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_176_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_371 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_3 _4165_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_952 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_440 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4360_ hold677/Z _4103_/I _4361_/S _4360_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3311_ _6730_/Q _3442_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_141_911 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_484 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_955 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4291_ hold876/Z hold271/Z _4291_/S _4291_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6030_ _6030_/A1 _6030_/A2 _6030_/A3 _6030_/A4 _6030_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_100_329 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_424 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1013 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_6932_ _6932_/D _7297_/RN _6932_/CLK _6932_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_35_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6863_ _6863_/D _7279_/RN _7230_/CLK hold36/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_63_961 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5814_ hold271/Z hold936/Z _5820_/S _5814_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_318 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6794_ _6794_/D _7265_/CLK _6794_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5745_ hold62/Z hold353/Z _5748_/S _5745_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_565 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5676_ hold960/Z hold271/Z _5682_/S _5676_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4627_ _4627_/A1 _4625_/Z _4626_/Z _4633_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_136_727 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xhold520 _7185_/Q hold520/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4558_ _5038_/A1 _4557_/Z _5393_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xhold531 _7197_/Q hold531/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_117_996 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_613 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xhold542 _4220_/Z _6750_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_718 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold553 _7057_/Q hold553/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7277_ _7277_/D _7279_/RN _7279_/CLK _7277_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold597 _5543_/Z _6911_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4489_ _4489_/A1 _4692_/B _4489_/B _4491_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai21_4
Xhold586 _6939_/Q hold586/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3509_ hold11/Z hold37/Z _3484_/Z hold32/Z _3509_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold564 _6934_/Q hold564/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold575 _7000_/Q hold575/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_104_668 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ _6228_/A1 _6228_/A2 _6228_/A3 _6227_/Z _6228_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_44_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1012 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6159_ _6147_/Z _6158_/Z _6473_/B1 _6168_/C _6555_/C _6160_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_98_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_880 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_254 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_885 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2736 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2725 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_340 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_598 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1079 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_877 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_237 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_545 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_365 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_473 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_398 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_590 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput162 wb_sel_i[1] _6574_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput151 wb_dat_i[30] _6597_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput140 wb_dat_i[20] _6591_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_232 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_416 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_622 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_964 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3860_ _3860_/A1 _3860_/A2 _3860_/A3 _3860_/A4 _3860_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_177_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3791_ _6950_/Q _5584_/A1 _5575_/A1 _6942_/Q _3925_/A2 input5/Z _3794_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XPHY_190 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_5530_ _3485_/Z _5839_/A3 hold637/Z _5520_/C _5531_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_9_851 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_822 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_215 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5461_ _5461_/I _5480_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4412_ _4412_/A1 _4399_/Z _4412_/B _4412_/C _5209_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_172_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7200_ _7200_/D _7258_/RN _7200_/CLK _7200_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
XFILLER_68_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5392_ _5051_/S _5360_/B _5392_/B _5433_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_67_1020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7131_ _7131_/D _7237_/RN _7131_/CLK _7131_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_114_933 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_432 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_633 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4343_ hold271/Z hold726/Z _4343_/S _6846_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7062_ _7062_/D _7221_/RN _7062_/CLK _7062_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_141_763 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_966 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_132 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4274_ _4274_/A1 hold18/Z _4276_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_101_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6013_ _6013_/A1 _5991_/Z _6027_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_100_137 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_360 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_405 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6915_ _6915_/D _7193_/RN _6915_/CLK _6915_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xclkbuf_leaf_71__1359_ clkbuf_4_13_0__1359_/Z net613_258/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1309 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_246 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_605 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6846_ _6846_/D input75/Z _6846_/CLK _6846_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_50_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6777_ _6777_/D _7238_/RN _6777_/CLK _6777_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3989_ _7239_/Q _6895_/Q _6900_/Q _3990_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_5728_ _5728_/A1 hold18/Z _5730_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_182_129 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_693 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_708 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5659_ hold918/Z hold86/Z _5664_/S _7014_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_899 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_549 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold361 _5705_/Z _7055_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_7_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold350 _4126_/Z _6680_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold372 _7208_/Q hold372/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_120_914 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold383 _6669_/Q hold383/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold394 _5711_/Z _7060_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_77_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_530 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3201 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3256 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3245 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3234 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3223 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet813_460 _4073__37/I _6705_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2533 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xnet813_482 net813_482/I _6683_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_493 net413_86/I _6672_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet813_471 net813_471/I _6694_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_186_413 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_638 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1898 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_170 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_811 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_384 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_342 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_570 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_168 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_842 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1027 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1008 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4961_ _4500_/Z _4906_/Z _5072_/A4 _5359_/A1 _4961_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_92_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4892_ _4551_/Z _4716_/Z _4892_/B _4894_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_6700_ _6700_/D _7258_/RN _6700_/CLK _6700_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_3912_ _7214_/Q _3912_/A2 _3912_/B1 _6883_/Q _3912_/C1 _6706_/Q _3915_/A1 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_6631_ _7193_/RN _6652_/A2 _6631_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_32_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3843_ _3529_/Z _3617_/Z _3950_/C1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_32_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6562_ _6562_/I _7261_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_502 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3774_ _6926_/Q _3935_/A2 _3945_/C2 _6684_/Q _5701_/A1 _7054_/Q _3776_/A2 VDD VSS
+ gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_173_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6493_ _6493_/A1 _6493_/A2 _6486_/Z _6492_/Z _6493_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_5513_ _5520_/C _3533_/Z _5513_/A3 _5821_/A3 _5514_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_5444_ _5444_/A1 _5444_/A2 _5442_/Z _5444_/A4 _5483_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_145_376 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_379 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5375_ _5421_/A2 _5470_/A1 _5372_/Z _5374_/Z _5379_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7114_ _7114_/D _7219_/RN _7114_/CLK _7114_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_99_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4326_ _3509_/Z _5821_/A3 hold637/Z _5520_/C _4328_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4257_ hold52/Z hold332/Z _4261_/S _4257_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_146 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7045_ _7045_/D _7219_/RN _7045_/CLK _7045_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_86_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4188_ _4188_/A1 hold18/Z _4190_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_55_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1128 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_920 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1106 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_925 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1139 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6829_ _6829_/D _7279_/RN _7279_/CLK _6829_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_144_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4073__9 _4073__9/I _7216_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_479 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_619 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_387 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold180 _7124_/Q hold180/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold191 _5718_/Z _7067_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_2_389 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3020 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_820 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3053 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_769 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3086 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1052 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_953 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1060 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1684 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1036 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1695 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_934 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_600 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3490_ _7305_/Q _7304_/Q _6733_/Q _3491_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_140 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_673 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_346 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_519 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5160_ _5287_/B _5293_/B _4784_/Z _5160_/B _5366_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_68_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4111_ hold61/Z _7274_/Q hold21/Z hold62/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_4
X_5091_ _4586_/Z _5302_/B _4784_/Z _4716_/Z _5222_/A1 _5103_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai32_4
XFILLER_64_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4042_ _7291_/Q _3409_/Z _4042_/A3 _4043_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_83_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_511 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_330 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_672 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5993_ _7231_/Q _7228_/Q _7227_/Q _6211_/B1 _5994_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_4944_ _4467_/B _4495_/Z _5324_/A1 _4759_/Z _4944_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_64_396 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_290 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_744 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4875_ _4651_/Z _4817_/Z _4876_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_178_788 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6614_ _7221_/RN _6656_/A2 _6614_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_159_991 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3826_ _3529_/Z _3560_/Z _3934_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_118_321 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3757_ _3757_/A1 _3757_/A2 _3757_/A3 _3757_/A4 _3757_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_6545_ _6788_/Q _6263_/Z _6266_/Z _6844_/Q _6546_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_180_419 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6476_ _7257_/Q _6476_/I1 _6558_/S _7257_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_538 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3688_ _3688_/A1 _3663_/Z _3674_/Z _3687_/Z _3688_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
Xoutput230 _6913_/Q mgmt_gpio_out[29] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5427_ _5427_/A1 _5425_/Z _5426_/Z _4881_/Z _5430_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_134_869 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput252 _4079_/ZN pad_flash_io0_ie VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput241 _6751_/Q mgmt_gpio_out[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5358_ _5432_/A1 _5189_/Z _5355_/Z _5357_/Z _5362_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xoutput274 _6678_/Q pll_trim[12] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput285 hold97/I pll_trim[22] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
Xoutput263 _6879_/Q pll_div[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_593 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_733 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4309_ _4309_/I0 _6815_/Q _4312_/S _6815_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput296 _6675_/Q pll_trim[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5289_ _5029_/B _5289_/A2 _5289_/A3 _5292_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_74_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7028_ _7028_/D _7210_/RN _7028_/CLK _7028_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
XFILLER_87_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_694 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_514 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1028 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_755 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_243 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_799 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_427 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_967 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_354 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_858 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_847 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_643 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_891 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_563 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_617 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_864 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2171 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2160 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2193 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1492 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_720 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4660_ _4376_/Z _4411_/Z _5172_/B _5165_/A4 _5385_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
X_3611_ _3610_/Z hold994/Z _3899_/S _6875_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_1011 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4591_ _4591_/A1 _4587_/Z _4590_/Z _4593_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_156_972 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6330_ _7005_/Q _6243_/Z _6269_/Z _7029_/Q _7119_/Q _6288_/Z _6331_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_142_110 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3542_ _3653_/A1 hold338/Z _3497_/I _3501_/Z _3542_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_50_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_993 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold916 _6699_/Q hold916/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold927 _6787_/Q hold927/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold905 _4346_/Z _6848_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_430 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_655 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_121 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3473_ _3471_/I _5490_/A1 hold21/Z _3473_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6261_ _7234_/Q _6533_/A2 _6533_/A3 _5943_/S _6261_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_115_357 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold938 _7207_/Q hold938/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold949 _5703_/Z _7053_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5212_ _5242_/A3 _4810_/B _4812_/B _5212_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_9_1001 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6192_ _6718_/Q _5960_/Z _6192_/B _6193_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_5143_ _4820_/Z _4821_/Z _4878_/Z _5364_/B _5372_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_9_1078 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1067 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5074_ _5074_/A1 _5408_/C _5072_/Z _5335_/C _5075_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_69_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_116 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4025_ _4489_/B _4424_/B _4034_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_38_853 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_385 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5976_ _6015_/A3 _6211_/B1 _7004_/Q _7228_/Q _5976_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_13_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4927_ _4927_/A1 _4927_/A2 _4927_/A3 _4929_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_4858_ _4858_/A1 _4858_/A2 _5289_/A2 _4862_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_166_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_909 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xnet563_218 net613_258/I _7007_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xnet563_207 net563_230/I _7018_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3809_ _3509_/Z _3617_/Z _4289_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xnet563_229 net763_425/I _6996_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_181_728 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_641 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4789_ _5270_/A1 _4808_/A2 _4530_/I _5302_/B _4789_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_146_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6528_ _6516_/Z _6527_/Z _6528_/B1 _6286_/Z _6529_/I0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_6459_ _6459_/I _6460_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_195 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_327 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_596 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_439 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_352 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_897 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_631 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_839 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_742 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_758 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_775 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_566 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_950 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_780 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_942 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_471 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_48__1359_ net463_109/I _4073__9/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_128__1359_ _4073__15/I _4073__39/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_171_249 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_154 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_506 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_241 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_948 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_138 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_951 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5830_ _3542_/Z _3552_/Z _5520_/C _5838_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_61_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_804 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_377 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5761_ hold500/Z hold86/Z _5766_/S _5761_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4712_ _4687_/Z _5092_/A1 _4713_/A1 _4691_/Z _5222_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_148_747 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5692_ _3529_/Z _3542_/Z hold6/Z _5700_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_30_583 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4643_ _5315_/A1 _5315_/A2 _4546_/Z _5364_/B _4643_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_4574_ _5278_/C _4551_/Z _5370_/C VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_128_460 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold702 _4190_/Z _6727_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7293_ _7293_/D _6647_/Z _7304_/CLK _7293_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xhold724 _7116_/Q hold724/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3525_ _3653_/A1 hold338/Z _3617_/A1 _3501_/Z _3525_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
X_6313_ _6997_/Q _6265_/Z _6266_/Z _7013_/Q _6329_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xhold746 _4166_/Z _6711_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold713 _6695_/Q hold713/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold735 _6844_/Q hold735/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_171_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_1054 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xnet513_159 net513_159/I _7066_/CLK VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6244_ _7235_/Q _7234_/Q _6452_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_115_165 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold779 _6926_/Q hold779/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold768 _4357_/Z _6855_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold757 _6892_/Q hold757/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_170_282 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3456_ hold28/Z hold61/Z _3460_/S _7288_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_198 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_669 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6175_ hold91/I _5958_/Z _5994_/I _7141_/Q _6176_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_85_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3387_ _7227_/Q _6015_/A3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_130_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5126_ _5126_/I _5127_/A4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5057_ _5078_/A2 _5443_/A1 _5057_/B _5324_/C _5058_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_85_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_149 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2918 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2907 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_4008_ _4008_/I _4009_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_992 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_344 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5959_ _6014_/A2 _5984_/A1 wire348/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_40_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_503 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_706 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_408 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_238 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_493 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_658 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_176 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_850 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold40 hold40/I hold40/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_48_425 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold51 hold51/I hold51/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold62 hold62/I hold62/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold73 hold73/I hold73/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_29_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold95 hold95/I hold95/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_75_288 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_406 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_970 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xhold84 hold84/I hold84/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_17_845 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_614 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_826 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_361 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_350 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_372 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_363 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_739 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_4 _4186_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_400 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3310_ hold31/Z _5490_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_98_314 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_794 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4290_ hold823/Z _4103_/I _4291_/S _4290_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_455 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_308 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_550 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_701 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_179 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_15_0__1359_ clkbuf_0__1359_/Z clkbuf_4_15_0__1359_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_94_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_597 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_929 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_119 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6931_ _6931_/D _7258_/RN _6931_/CLK _6931_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_179_113 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6862_ _6862_/D _7279_/RN _7230_/CLK _6862_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_601 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_303 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_848 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5813_ _4103_/I hold910/Z _5820_/S _5813_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6793_ _6793_/D _7265_/CLK _6793_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_656 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_667 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1031 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5744_ hold52/Z hold512/Z _5748_/S _5744_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5675_ hold458/Z hold113/Z _5682_/S _5675_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4626_ _4887_/A1 _4868_/A1 _4546_/Z _5364_/B _4626_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
XFILLER_148_599 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_547 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xhold510 _6993_/Q hold510/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_4557_ _4436_/B _4648_/A1 _4648_/A2 _4557_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
Xhold521 _5852_/Z _7185_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold532 _5865_/Z _7197_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold543 _7177_/Q hold543/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_116_463 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_94__1359_ net813_465/I net563_251/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xhold554 _5707_/Z _7057_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_7276_ _7276_/D _7279_/RN _7279_/CLK _7276_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_4488_ _4392_/Z _4474_/Z _4722_/A2 _4923_/A2 _4491_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
Xhold587 _5574_/Z _6939_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3508_ hold32/Z hold37/Z _3484_/Z hold38/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or3_4
XFILLER_103_124 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_325 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xhold576 _7182_/Q hold576/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
Xhold565 _5569_/Z _6934_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
X_3439_ _3971_/A1 _3442_/B _6665_/Q _6664_/Q _3440_/S VDD VSS gf180mcu_fd_sc_mcu7t5v0__or4_4
Xhold598 _6935_/Q hold598/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlyc_2
XFILLER_106_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6227_ _6227_/A1 _6227_/A2 _6227_/A3 _6227_/A4 _6227_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_131_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6158_ _6152_/Z _6155_/Z _6158_/A3 _6158_/A4 _6158_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XTAP_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_5109_ _5108_/Z _4853_/Z _4740_/Z _5111_/B VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_85_542 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_881 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_6089_ _7244_/Q _6089_/I1 _6558_/S _7244_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2737 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2715 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_214 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_428 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2759 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2748 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_247 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_664 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_163 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_686 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_333 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_889 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_208 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_912 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_496 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_989 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_712 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_251 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput163 wb_sel_i[2] _6573_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput152 wb_dat_i[31] _6600_/C2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput141 wb_dat_i[21] _6594_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput130 wb_dat_i[11] _6588_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_531 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_778 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_578 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_556 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_422 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1080 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1075 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1064 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1059 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3790_ _3790_/A1 _3790_/A2 _3790_/A3 _3790_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_13_870 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_818 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_144 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_689 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_191 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_180 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_886 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5460_ _5460_/A1 _5303_/Z _5460_/A3 _5460_/A4 _5461_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_8_373 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _5083_/B _4412_/B _4412_/C _4411_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and3_4
XFILLER_145_536 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_709 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5391_ _5388_/Z _4985_/Z _5386_/Z _5390_/Z _5391_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_126_772 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7130_ _7130_/D _7221_/RN _7130_/CLK _7130_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_4342_ _4103_/I _6845_/Q _4343_/S _4342_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7061_ _7061_/D _7210_/RN _7061_/CLK _7061_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
X_4273_ hold271/Z hold866/Z _4273_/S _4273_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_499 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6012_ _7021_/Q wire348/Z _6211_/B1 _6989_/Q _6013_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__aoi22_4
.ends

