magic
tech gf180mcuC
magscale 1 10
timestamp 1655307388
<< error_p >>
rect -275 -24 -229 72
rect 229 -24 275 72
<< nwell >>
rect -518 -336 518 336
<< mvpmos >>
rect -200 -26 200 74
<< mvpdiff >>
rect -288 61 -200 74
rect -288 -13 -275 61
rect -229 -13 -200 61
rect -288 -26 -200 -13
rect 200 61 288 74
rect 200 -13 229 61
rect 275 -13 288 61
rect 200 -26 288 -13
<< mvpdiffc >>
rect -275 -13 -229 61
rect 229 -13 275 61
<< mvnsubdiff >>
rect -432 237 432 250
rect -432 191 -316 237
rect 316 191 432 237
rect -432 178 432 191
rect -432 134 -360 178
rect -432 -134 -419 134
rect -373 -134 -360 134
rect 360 134 432 178
rect -432 -178 -360 -134
rect 360 -134 373 134
rect 419 -134 432 134
rect 360 -178 432 -134
rect -432 -250 432 -178
<< mvnsubdiffcont >>
rect -316 191 316 237
rect -419 -134 -373 134
rect 373 -134 419 134
<< polysilicon >>
rect -200 74 200 118
rect -200 -59 200 -26
rect -200 -105 -187 -59
rect 187 -105 200 -59
rect -200 -118 200 -105
<< polycontact >>
rect -187 -105 187 -59
<< metal1 >>
rect -419 191 -316 237
rect 316 191 419 237
rect -419 134 -373 191
rect 373 134 419 191
rect -275 61 -229 72
rect -275 -24 -229 -13
rect 229 61 275 72
rect 229 -24 275 -13
rect -198 -105 -187 -59
rect 187 -105 198 -59
rect -419 -191 -373 -134
rect 373 -191 419 -134
rect -419 -237 419 -191
<< properties >>
string FIXED_BBOX -396 -214 396 214
string gencell pmos_6p0
string library gf180mcu
string parameters w 0.5 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.5 wmin 0.3 full_metal 1 compatible {pmos_3p3 pmos_6p0}
<< end >>
