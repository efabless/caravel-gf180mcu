magic
tech gf180mcuC
magscale 1 5
timestamp 1655473103
<< obsm1 >>
rect 560 267 16408 9438
<< metal2 >>
rect 588 9600 644 10000
rect 1876 9600 1932 10000
rect 3164 9600 3220 10000
rect 4508 9600 4564 10000
rect 5796 9600 5852 10000
rect 7084 9600 7140 10000
rect 8428 9600 8484 10000
rect 9716 9600 9772 10000
rect 11060 9600 11116 10000
rect 12348 9600 12404 10000
rect 13636 9600 13692 10000
rect 14980 9600 15036 10000
rect 16268 9600 16324 10000
rect 4228 0 4284 400
rect 12740 0 12796 400
<< obsm2 >>
rect 434 9570 558 9600
rect 674 9570 1846 9600
rect 1962 9570 3134 9600
rect 3250 9570 4478 9600
rect 4594 9570 5766 9600
rect 5882 9570 7054 9600
rect 7170 9570 8398 9600
rect 8514 9570 9686 9600
rect 9802 9570 11030 9600
rect 11146 9570 12318 9600
rect 12434 9570 13606 9600
rect 13722 9570 14950 9600
rect 15066 9570 16238 9600
rect 434 430 16310 9570
rect 434 261 4198 430
rect 4314 261 12710 430
rect 12826 261 16310 430
<< metal3 >>
rect 0 9604 400 9660
rect 16600 9100 17000 9156
rect 0 8988 400 9044
rect 0 8372 400 8428
rect 0 7756 400 7812
rect 16600 7420 17000 7476
rect 0 7140 400 7196
rect 0 6524 400 6580
rect 0 5908 400 5964
rect 16600 5796 17000 5852
rect 0 5292 400 5348
rect 0 4620 400 4676
rect 16600 4116 17000 4172
rect 0 4004 400 4060
rect 0 3388 400 3444
rect 0 2772 400 2828
rect 16600 2436 17000 2492
rect 0 2156 400 2212
rect 0 1540 400 1596
rect 0 924 400 980
rect 16600 812 17000 868
rect 0 308 400 364
<< obsm3 >>
rect 430 9574 16600 9646
rect 400 9186 16600 9574
rect 400 9074 16570 9186
rect 430 9070 16570 9074
rect 430 8958 16600 9070
rect 400 8458 16600 8958
rect 430 8342 16600 8458
rect 400 7842 16600 8342
rect 430 7726 16600 7842
rect 400 7506 16600 7726
rect 400 7390 16570 7506
rect 400 7226 16600 7390
rect 430 7110 16600 7226
rect 400 6610 16600 7110
rect 430 6494 16600 6610
rect 400 5994 16600 6494
rect 430 5882 16600 5994
rect 430 5878 16570 5882
rect 400 5766 16570 5878
rect 400 5378 16600 5766
rect 430 5262 16600 5378
rect 400 4706 16600 5262
rect 430 4590 16600 4706
rect 400 4202 16600 4590
rect 400 4090 16570 4202
rect 430 4086 16570 4090
rect 430 3974 16600 4086
rect 400 3474 16600 3974
rect 430 3358 16600 3474
rect 400 2858 16600 3358
rect 430 2742 16600 2858
rect 400 2522 16600 2742
rect 400 2406 16570 2522
rect 400 2242 16600 2406
rect 430 2126 16600 2242
rect 400 1626 16600 2126
rect 430 1510 16600 1626
rect 400 1010 16600 1510
rect 430 898 16600 1010
rect 430 894 16570 898
rect 400 782 16570 894
rect 400 394 16600 782
rect 430 322 16600 394
<< metal4 >>
rect 2465 362 2625 9438
rect 4450 362 4610 9438
rect 6435 362 6595 9438
rect 8420 362 8580 9438
rect 10405 362 10565 9438
rect 12390 362 12550 9438
rect 14375 362 14535 9438
<< obsm4 >>
rect 602 485 2435 9203
rect 2655 485 4420 9203
rect 4640 485 6405 9203
rect 6625 485 8390 9203
rect 8610 485 10375 9203
rect 10595 485 12360 9203
rect 12580 485 13846 9203
<< metal5 >>
rect 530 8376 16438 8536
rect 530 7224 16438 7384
rect 530 6072 16438 6232
rect 530 4920 16438 5080
rect 530 3768 16438 3928
rect 530 2616 16438 2776
rect 530 1464 16438 1624
<< obsm5 >>
rect 762 8586 13854 9202
rect 762 7434 13854 8326
rect 762 6282 13854 7174
rect 762 5130 13854 6022
rect 762 3978 13854 4870
rect 762 2826 13854 3718
rect 762 1688 13854 2566
<< labels >>
rlabel metal4 s 2465 362 2625 9438 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 6435 362 6595 9438 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 10405 362 10565 9438 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 14375 362 14535 9438 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 530 1464 16438 1624 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 530 3768 16438 3928 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 530 6072 16438 6232 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 530 8376 16438 8536 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 4450 362 4610 9438 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 8420 362 8580 9438 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 12390 362 12550 9438 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 530 2616 16438 2776 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 530 4920 16438 5080 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 530 7224 16438 7384 6 VSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 308 400 364 6 clockp[0]
port 3 nsew signal output
rlabel metal3 s 0 924 400 980 6 clockp[1]
port 4 nsew signal output
rlabel metal3 s 0 5292 400 5348 6 dco
port 5 nsew signal input
rlabel metal3 s 0 1540 400 1596 6 div[0]
port 6 nsew signal input
rlabel metal3 s 0 2156 400 2212 6 div[1]
port 7 nsew signal input
rlabel metal3 s 0 2772 400 2828 6 div[2]
port 8 nsew signal input
rlabel metal3 s 0 3388 400 3444 6 div[3]
port 9 nsew signal input
rlabel metal3 s 0 4004 400 4060 6 div[4]
port 10 nsew signal input
rlabel metal3 s 0 4620 400 4676 6 enable
port 11 nsew signal input
rlabel metal3 s 0 5908 400 5964 6 ext_trim[0]
port 12 nsew signal input
rlabel metal2 s 4508 9600 4564 10000 6 ext_trim[10]
port 13 nsew signal input
rlabel metal2 s 5796 9600 5852 10000 6 ext_trim[11]
port 14 nsew signal input
rlabel metal2 s 7084 9600 7140 10000 6 ext_trim[12]
port 15 nsew signal input
rlabel metal2 s 8428 9600 8484 10000 6 ext_trim[13]
port 16 nsew signal input
rlabel metal2 s 9716 9600 9772 10000 6 ext_trim[14]
port 17 nsew signal input
rlabel metal2 s 11060 9600 11116 10000 6 ext_trim[15]
port 18 nsew signal input
rlabel metal2 s 12348 9600 12404 10000 6 ext_trim[16]
port 19 nsew signal input
rlabel metal2 s 13636 9600 13692 10000 6 ext_trim[17]
port 20 nsew signal input
rlabel metal2 s 14980 9600 15036 10000 6 ext_trim[18]
port 21 nsew signal input
rlabel metal2 s 16268 9600 16324 10000 6 ext_trim[19]
port 22 nsew signal input
rlabel metal3 s 0 6524 400 6580 6 ext_trim[1]
port 23 nsew signal input
rlabel metal3 s 16600 9100 17000 9156 6 ext_trim[20]
port 24 nsew signal input
rlabel metal3 s 16600 7420 17000 7476 6 ext_trim[21]
port 25 nsew signal input
rlabel metal3 s 16600 5796 17000 5852 6 ext_trim[22]
port 26 nsew signal input
rlabel metal3 s 16600 4116 17000 4172 6 ext_trim[23]
port 27 nsew signal input
rlabel metal3 s 16600 2436 17000 2492 6 ext_trim[24]
port 28 nsew signal input
rlabel metal3 s 16600 812 17000 868 6 ext_trim[25]
port 29 nsew signal input
rlabel metal3 s 0 7140 400 7196 6 ext_trim[2]
port 30 nsew signal input
rlabel metal3 s 0 7756 400 7812 6 ext_trim[3]
port 31 nsew signal input
rlabel metal3 s 0 8372 400 8428 6 ext_trim[4]
port 32 nsew signal input
rlabel metal3 s 0 8988 400 9044 6 ext_trim[5]
port 33 nsew signal input
rlabel metal3 s 0 9604 400 9660 6 ext_trim[6]
port 34 nsew signal input
rlabel metal2 s 588 9600 644 10000 6 ext_trim[7]
port 35 nsew signal input
rlabel metal2 s 1876 9600 1932 10000 6 ext_trim[8]
port 36 nsew signal input
rlabel metal2 s 3164 9600 3220 10000 6 ext_trim[9]
port 37 nsew signal input
rlabel metal2 s 12740 0 12796 400 6 osc
port 38 nsew signal input
rlabel metal2 s 4228 0 4284 400 6 resetb
port 39 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 17000 10000
string GDS_END 936528
string GDS_FILE ../gds/digital_pll.gds.gz
string GDS_START 207956
string LEFclass BLOCK
string LEFview TRUE
<< end >>
