// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

// `default_nettype none
module chip_io_alt #(
	parameter ANALOG_PADS_1 = 5,
	parameter ANALOG_PADS_2 = 6
) (
`ifdef USE_POWER_PINS
	// Power buses
	inout  vss,	// Common padframe/ESD 5.0V ground
	inout  vdd,	// Management padframe/ESD 5.0V supply
`endif

	inout  gpio,
	input  clock,
	input  resetb,
	output flash_csb,
	output flash_clk,
	inout  flash_io0,
	inout  flash_io1,

	// Chip Core Interface
	output resetb_core,
	output clock_core,
	output gpio_in_core,
	input  gpio_out_core,
	input  gpio_outen_core,
	input  gpio_inen_core,
	input  gpio_pu_select,
	input  gpio_pd_select,
	input  gpio_schmitt_select,
	input  gpio_slew_select,
	input  [1:0] gpio_drive_select_core,
	input  flash_csb_core,
	input  flash_clk_core,
	input  flash_csb_oe_core,
	input  flash_clk_oe_core,
	input  flash_io0_oe_core,
	input  flash_io1_oe_core,
	input  flash_io0_ie_core,
	input  flash_io1_ie_core,
	input  flash_io0_do_core,
	input  flash_io1_do_core,
	output flash_io0_di_core,
	output flash_io1_di_core,

	// Constant value inputs for fixed GPIO configuration
	input [5:0] const_zero,
	input [1:0] const_one,

	// User project IOs
	inout [`MPRJ_IO_PADS-1:0] mprj_io,
	// The section below is for the digital pads only
	input [`MPRJ_IO_PADS-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_out,
	input [`MPRJ_IO_PADS-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_outen,
	input [`MPRJ_IO_PADS-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_inen,
	input [`MPRJ_IO_PADS-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_schmitt_select,
	input [`MPRJ_IO_PADS-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_slew_select,
	input [`MPRJ_IO_PADS-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_pu_select,
	input [`MPRJ_IO_PADS-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_pd_select,
	input [(`MPRJ_IO_PADS-ANALOG_PADS_1-ANALOG_PADS_2)*2-1:0] mprj_io_drive_sel,
	output [`MPRJ_IO_PADS-ANALOG_PADS_1-ANALOG_PADS_2-1:0] mprj_io_in
);

	// Instantiate power and ground pads for management domain
	// 12 pads:  vddio, vssio, vdda, vssa, vccd, vssd correspond
	// to names used with sky130, with multiple voltages for each
	// domain.  The instance names reflect where these pads
	// match the position of corresponding pads on the sky130
	// caravel, but note that there is actually only one
	// 5V supply, VDD and one common ground, VSS.

	// NOTE:  Global Foundries only supplies two pads, DVDD and
	// DVSS for 5V.  Only 5V digital cells are available for this
	// process.  Therefore, all power supplies are on the 5V
	// domain.  The VDD breaker cell divides VDD domains;
	// however, all VSS domains are tied together.

    	gf180mcu_fd_io__dvdd mgmt_vddio_pad_0 (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

	// lies in user area---Does not belong to management domain
	// like it does on the Sky130 version.
    	gf180mcu_fd_io__dvdd mgmt_vddio_pad_1 (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

    	gf180mcu_fd_io__dvdd mgmt_vdda_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

    	gf180mcu_fd_io__dvdd mgmt_vccd_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

    	gf180mcu_fd_io__dvss mgmt_vssio_pad_0 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);

    	gf180mcu_fd_io__dvss mgmt_vssio_pad_1 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);

    	gf180mcu_fd_io__dvss mgmt_vssa_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);

    	gf180mcu_fd_io__dvss mgmt_vssd_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);

	// Instantiate power and ground pads for user 1 domain
	// 8 pads:  vdda, vssa, vccd, vssd;  One each HV and LV clamp.

    	gf180mcu_fd_io__dvdd user1_vdda_pad_0 (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

		gf180mcu_fd_io__dvdd user1_vdda_pad_1 (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

    	gf180mcu_fd_io__dvdd user1_vccd_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

    	gf180mcu_fd_io__dvss user1_vssa_pad_0 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);


    	gf180mcu_fd_io__dvss user1_vssa_pad_1 (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);

    	gf180mcu_fd_io__dvss user1_vssd_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);

	// Instantiate power and ground pads for user 2 domain
	// 8 pads:  vdda, vssa, vccd, vssd;  One each HV and LV clamp.

    	gf180mcu_fd_io__dvdd user2_vdda_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

    	gf180mcu_fd_io__dvdd user2_vccd_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VSS(vss)
    	);

    	gf180mcu_fd_io__dvss user2_vssa_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);

    	gf180mcu_fd_io__dvss user2_vssd_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd)
    	);

	// Management clock input pad
	gf180mcu_fd_io__in_c mgmt_clock_input_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PU(const_zero[4]),
		.PD(const_zero[4]),
		.PAD(clock),
		.Y(clock_core)
	);

	// Management GPIO pad
	gf180mcu_fd_io__bi_t mgmt_gpio_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(gpio),
		.CS(gpio_schmitt_select),
		.SL(gpio_slew_select),
		.IE(gpio_inen_core),
		.OE(gpio_outen_core),
		.PU(gpio_pu_select),
		.PD(gpio_pd_select),
		.PDRV0(gpio_drive_select_core[0]),
		.PDRV1(gpio_drive_select_core[1]),
		.A(gpio_out_core),
		.Y(gpio_in_core)
	);

	// Management Flash SPI pads
	gf180mcu_fd_io__bi_t flash_io0_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(flash_io0),
		.CS(const_zero[1]),
		.SL(const_zero[1]),
		.IE(flash_io0_ie_core),
		.OE(flash_io0_oe_core),
		.PU(const_zero[1]),
		.PD(const_zero[1]),
		.PDRV0(const_zero[1]),
		.PDRV1(const_zero[1]),
		.A(flash_io0_do_core),
		.Y(flash_io0_di_core)
	);
	
	gf180mcu_fd_io__bi_t flash_io1_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(flash_io1),
		.CS(const_zero[0]),
		.SL(const_zero[0]),
		.IE(flash_io1_ie_core),
		.OE(flash_io1_oe_core),
		.PU(const_zero[0]),
		.PD(const_zero[0]),
		.PDRV0(const_zero[0]),
		.PDRV1(const_zero[0]),
		.A(flash_io1_do_core),
		.Y(flash_io1_di_core)
	);

	gf180mcu_fd_io__bi_t flash_csb_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(flash_csb),
		.CS(const_zero[3]),
		.SL(const_zero[3]),
		.IE(const_zero[3]),
		.OE(flash_csb_oe_core),
		.PU(const_one[1]),
		.PD(const_zero[3]),
		.PDRV0(const_zero[3]),
		.PDRV1(const_zero[3]),
		.A(flash_csb_core),
		.Y()
	);

	gf180mcu_fd_io__bi_t flash_clk_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PAD(flash_clk),
		.CS(const_zero[2]),
		.SL(const_zero[2]),
		.IE(const_zero[2]),
		.OE(flash_clk_oe_core),
		.PU(const_zero[2]),
		.PD(const_zero[2]),
		.PDRV0(const_zero[2]),
		.PDRV1(const_zero[2]),
		.A(flash_clk_core),
		.Y()
	);

	// NOTE:  Resetb is active low and is configured as a pull-up

	gf180mcu_fd_io__in_s resetb_pad (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
		.PU(const_one[0]),
		.PD(const_zero[5]),
		.PAD(resetb),
		.Y(resetb_core)
	);

	// Corner cells (These are overlay cells;  it is not clear what is normally
    	// supposed to go under them.)

	gf180mcu_fd_io__cor mgmt_corner [1:0] (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	);

	gf180mcu_fd_io__cor user1_corner (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
    	);

	gf180mcu_fd_io__cor user2_corner (
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
    	);

	// generated by running ./scripts/update_chip_io_rtl.py then copying
	// ./scripts/chip_io.txt and pasting here;  edited to remove pads
	// replaced by analog pads on caravan (15 through 25)

	gf180mcu_fd_io__bi_t \mprj_pads[0]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[0]),
		.CS(mprj_io_schmitt_select[0]),
		.SL(mprj_io_slew_select[0]),
		.IE(mprj_io_inen[0]),
		.OE(mprj_io_outen[0]),
		.PU(mprj_io_pu_select[0]),
		.PD(mprj_io_pd_select[0]),
		.PDRV0(mprj_io_drive_sel[0]),
		.PDRV1(mprj_io_drive_sel[1]),
		.A(mprj_io_out[0]),
		.Y(mprj_io_in[0])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[1]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[1]),
		.CS(mprj_io_schmitt_select[1]),
		.SL(mprj_io_slew_select[1]),
		.IE(mprj_io_inen[1]),
		.OE(mprj_io_outen[1]),
		.PU(mprj_io_pu_select[1]),
		.PD(mprj_io_pd_select[1]),
		.PDRV0(mprj_io_drive_sel[2]),
		.PDRV1(mprj_io_drive_sel[3]),
		.A(mprj_io_out[1]),
		.Y(mprj_io_in[1])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[2]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[2]),
		.CS(mprj_io_schmitt_select[2]),
		.SL(mprj_io_slew_select[2]),
		.IE(mprj_io_inen[2]),
		.OE(mprj_io_outen[2]),
		.PU(mprj_io_pu_select[2]),
		.PD(mprj_io_pd_select[2]),
		.PDRV0(mprj_io_drive_sel[4]),
		.PDRV1(mprj_io_drive_sel[5]),
		.A(mprj_io_out[2]),
		.Y(mprj_io_in[2])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[3]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[3]),
		.CS(mprj_io_schmitt_select[3]),
		.SL(mprj_io_slew_select[3]),
		.IE(mprj_io_inen[3]),
		.OE(mprj_io_outen[3]),
		.PU(mprj_io_pu_select[3]),
		.PD(mprj_io_pd_select[3]),
		.PDRV0(mprj_io_drive_sel[6]),
		.PDRV1(mprj_io_drive_sel[7]),
		.A(mprj_io_out[3]),
		.Y(mprj_io_in[3])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[4]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[4]),
		.CS(mprj_io_schmitt_select[4]),
		.SL(mprj_io_slew_select[4]),
		.IE(mprj_io_inen[4]),
		.OE(mprj_io_outen[4]),
		.PU(mprj_io_pu_select[4]),
		.PD(mprj_io_pd_select[4]),
		.PDRV0(mprj_io_drive_sel[8]),
		.PDRV1(mprj_io_drive_sel[9]),
		.A(mprj_io_out[4]),
		.Y(mprj_io_in[4])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[5]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[5]),
		.CS(mprj_io_schmitt_select[5]),
		.SL(mprj_io_slew_select[5]),
		.IE(mprj_io_inen[5]),
		.OE(mprj_io_outen[5]),
		.PU(mprj_io_pu_select[5]),
		.PD(mprj_io_pd_select[5]),
		.PDRV0(mprj_io_drive_sel[10]),
		.PDRV1(mprj_io_drive_sel[11]),
		.A(mprj_io_out[5]),
		.Y(mprj_io_in[5])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[6]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[6]),
		.CS(mprj_io_schmitt_select[6]),
		.SL(mprj_io_slew_select[6]),
		.IE(mprj_io_inen[6]),
		.OE(mprj_io_outen[6]),
		.PU(mprj_io_pu_select[6]),
		.PD(mprj_io_pd_select[6]),
		.PDRV0(mprj_io_drive_sel[12]),
		.PDRV1(mprj_io_drive_sel[13]),
		.A(mprj_io_out[6]),
		.Y(mprj_io_in[6])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[7]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[7]),
		.CS(mprj_io_schmitt_select[7]),
		.SL(mprj_io_slew_select[7]),
		.IE(mprj_io_inen[7]),
		.OE(mprj_io_outen[7]),
		.PU(mprj_io_pu_select[7]),
		.PD(mprj_io_pd_select[7]),
		.PDRV0(mprj_io_drive_sel[14]),
		.PDRV1(mprj_io_drive_sel[15]),
		.A(mprj_io_out[7]),
		.Y(mprj_io_in[7])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[8]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[8]),
		.CS(mprj_io_schmitt_select[8]),
		.SL(mprj_io_slew_select[8]),
		.IE(mprj_io_inen[8]),
		.OE(mprj_io_outen[8]),
		.PU(mprj_io_pu_select[8]),
		.PD(mprj_io_pd_select[8]),
		.PDRV0(mprj_io_drive_sel[16]),
		.PDRV1(mprj_io_drive_sel[17]),
		.A(mprj_io_out[8]),
		.Y(mprj_io_in[8])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[9]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[9]),
		.CS(mprj_io_schmitt_select[9]),
		.SL(mprj_io_slew_select[9]),
		.IE(mprj_io_inen[9]),
		.OE(mprj_io_outen[9]),
		.PU(mprj_io_pu_select[9]),
		.PD(mprj_io_pd_select[9]),
		.PDRV0(mprj_io_drive_sel[18]),
		.PDRV1(mprj_io_drive_sel[19]),
		.A(mprj_io_out[9]),
		.Y(mprj_io_in[9])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[10]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[10]),
		.CS(mprj_io_schmitt_select[10]),
		.SL(mprj_io_slew_select[10]),
		.IE(mprj_io_inen[10]),
		.OE(mprj_io_outen[10]),
		.PU(mprj_io_pu_select[10]),
		.PD(mprj_io_pd_select[10]),
		.PDRV0(mprj_io_drive_sel[20]),
		.PDRV1(mprj_io_drive_sel[21]),
		.A(mprj_io_out[10]),
		.Y(mprj_io_in[10])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[11]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[11]),
		.CS(mprj_io_schmitt_select[11]),
		.SL(mprj_io_slew_select[11]),
		.IE(mprj_io_inen[11]),
		.OE(mprj_io_outen[11]),
		.PU(mprj_io_pu_select[11]),
		.PD(mprj_io_pd_select[11]),
		.PDRV0(mprj_io_drive_sel[22]),
		.PDRV1(mprj_io_drive_sel[23]),
		.A(mprj_io_out[11]),
		.Y(mprj_io_in[11])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[12]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[12]),
		.CS(mprj_io_schmitt_select[12]),
		.SL(mprj_io_slew_select[12]),
		.IE(mprj_io_inen[12]),
		.OE(mprj_io_outen[12]),
		.PU(mprj_io_pu_select[12]),
		.PD(mprj_io_pd_select[12]),
		.PDRV0(mprj_io_drive_sel[24]),
		.PDRV1(mprj_io_drive_sel[25]),
		.A(mprj_io_out[12]),
		.Y(mprj_io_in[12])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[13]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[13]),
		.CS(mprj_io_schmitt_select[13]),
		.SL(mprj_io_slew_select[13]),
		.IE(mprj_io_inen[13]),
		.OE(mprj_io_outen[13]),
		.PU(mprj_io_pu_select[13]),
		.PD(mprj_io_pd_select[13]),
		.PDRV0(mprj_io_drive_sel[26]),
		.PDRV1(mprj_io_drive_sel[27]),
		.A(mprj_io_out[13]),
		.Y(mprj_io_in[13])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[25]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[14]),
		.CS(mprj_io_schmitt_select[14]),
		.SL(mprj_io_slew_select[14]),
		.IE(mprj_io_inen[14]),
		.OE(mprj_io_outen[14]),
		.PU(mprj_io_pu_select[14]),
		.PD(mprj_io_pd_select[14]),
		.PDRV0(mprj_io_drive_sel[28]),
		.PDRV1(mprj_io_drive_sel[29]),
		.A(mprj_io_out[14]),
		.Y(mprj_io_in[14])
	);

	gf180mcu_fd_io__bi_t \mprj_pads[26]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[15]),
		.CS(mprj_io_schmitt_select[15]),
		.SL(mprj_io_slew_select[15]),
		.IE(mprj_io_inen[15]),
		.OE(mprj_io_outen[15]),
		.PU(mprj_io_pu_select[15]),
		.PD(mprj_io_pd_select[15]),
		.PDRV0(mprj_io_drive_sel[30]),
		.PDRV1(mprj_io_drive_sel[31]),
		.A(mprj_io_out[15]),
		.Y(mprj_io_in[15])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[27]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[16]),
		.CS(mprj_io_schmitt_select[16]),
		.SL(mprj_io_slew_select[16]),
		.IE(mprj_io_inen[16]),
		.OE(mprj_io_outen[16]),
		.PU(mprj_io_pu_select[16]),
		.PD(mprj_io_pd_select[16]),
		.PDRV0(mprj_io_drive_sel[32]),
		.PDRV1(mprj_io_drive_sel[33]),
		.A(mprj_io_out[16]),
		.Y(mprj_io_in[16])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[28]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[17]),
		.CS(mprj_io_schmitt_select[17]),
		.SL(mprj_io_slew_select[17]),
		.IE(mprj_io_inen[17]),
		.OE(mprj_io_outen[17]),
		.PU(mprj_io_pu_select[17]),
		.PD(mprj_io_pd_select[17]),
		.PDRV0(mprj_io_drive_sel[34]),
		.PDRV1(mprj_io_drive_sel[35]),
		.A(mprj_io_out[17]),
		.Y(mprj_io_in[17])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[29]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[18]),
		.CS(mprj_io_schmitt_select[18]),
		.SL(mprj_io_slew_select[18]),
		.IE(mprj_io_inen[18]),
		.OE(mprj_io_outen[18]),
		.PU(mprj_io_pu_select[18]),
		.PD(mprj_io_pd_select[18]),
		.PDRV0(mprj_io_drive_sel[36]),
		.PDRV1(mprj_io_drive_sel[37]),
		.A(mprj_io_out[18]),
		.Y(mprj_io_in[18])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[30]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[19]),
		.CS(mprj_io_schmitt_select[19]),
		.SL(mprj_io_slew_select[19]),
		.IE(mprj_io_inen[19]),
		.OE(mprj_io_outen[19]),
		.PU(mprj_io_pu_select[19]),
		.PD(mprj_io_pd_select[19]),
		.PDRV0(mprj_io_drive_sel[38]),
		.PDRV1(mprj_io_drive_sel[39]),
		.A(mprj_io_out[19]),
		.Y(mprj_io_in[19])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[31]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[20]),
		.CS(mprj_io_schmitt_select[20]),
		.SL(mprj_io_slew_select[20]),
		.IE(mprj_io_inen[20]),
		.OE(mprj_io_outen[20]),
		.PU(mprj_io_pu_select[20]),
		.PD(mprj_io_pd_select[20]),
		.PDRV0(mprj_io_drive_sel[40]),
		.PDRV1(mprj_io_drive_sel[41]),
		.A(mprj_io_out[20]),
		.Y(mprj_io_in[20])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[32]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[21]),
		.CS(mprj_io_schmitt_select[21]),
		.SL(mprj_io_slew_select[21]),
		.IE(mprj_io_inen[21]),
		.OE(mprj_io_outen[21]),
		.PU(mprj_io_pu_select[21]),
		.PD(mprj_io_pd_select[21]),
		.PDRV0(mprj_io_drive_sel[42]),
		.PDRV1(mprj_io_drive_sel[43]),
		.A(mprj_io_out[21]),
		.Y(mprj_io_in[21])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[33]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[22]),
		.CS(mprj_io_schmitt_select[22]),
		.SL(mprj_io_slew_select[22]),
		.IE(mprj_io_inen[22]),
		.OE(mprj_io_outen[22]),
		.PU(mprj_io_pu_select[22]),
		.PD(mprj_io_pd_select[22]),
		.PDRV0(mprj_io_drive_sel[44]),
		.PDRV1(mprj_io_drive_sel[45]),
		.A(mprj_io_out[22]),
		.Y(mprj_io_in[22])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[34]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[23]),
		.CS(mprj_io_schmitt_select[23]),
		.SL(mprj_io_slew_select[23]),
		.IE(mprj_io_inen[23]),
		.OE(mprj_io_outen[23]),
		.PU(mprj_io_pu_select[23]),
		.PD(mprj_io_pd_select[23]),
		.PDRV0(mprj_io_drive_sel[46]),
		.PDRV1(mprj_io_drive_sel[47]),
		.A(mprj_io_out[23]),
		.Y(mprj_io_in[23])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[35]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[24]),
		.CS(mprj_io_schmitt_select[24]),
		.SL(mprj_io_slew_select[24]),
		.IE(mprj_io_inen[24]),
		.OE(mprj_io_outen[24]),
		.PU(mprj_io_pu_select[24]),
		.PD(mprj_io_pd_select[24]),
		.PDRV0(mprj_io_drive_sel[48]),
		.PDRV1(mprj_io_drive_sel[49]),
		.A(mprj_io_out[24]),
		.Y(mprj_io_in[24])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[36]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[25]),
		.CS(mprj_io_schmitt_select[25]),
		.SL(mprj_io_slew_select[25]),
		.IE(mprj_io_inen[25]),
		.OE(mprj_io_outen[25]),
		.PU(mprj_io_pu_select[25]),
		.PD(mprj_io_pd_select[25]),
		.PDRV0(mprj_io_drive_sel[50]),
		.PDRV1(mprj_io_drive_sel[51]),
		.A(mprj_io_out[25]),
		.Y(mprj_io_in[25])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[37]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.PAD(mprj_io[26]),
		.CS(mprj_io_schmitt_select[26]),
		.SL(mprj_io_slew_select[26]),
		.IE(mprj_io_inen[26]),
		.OE(mprj_io_outen[26]),
		.PU(mprj_io_pu_select[26]),
		.PD(mprj_io_pd_select[26]),
		.PDRV0(mprj_io_drive_sel[52]),
		.PDRV1(mprj_io_drive_sel[53]),
		.A(mprj_io_out[26]),
		.Y(mprj_io_in[26])
	);

	gf180mcu_fd_io__asig_5p0 \mprj_pads[14]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.ASIG5V(mprj_io[14])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[15]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.ASIG5V(mprj_io[15])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[16]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.ASIG5V(mprj_io[16])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[17]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.ASIG5V(mprj_io[17])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[18]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.ASIG5V(mprj_io[18])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[19]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.ASIG5V(mprj_io[19])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[20]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.ASIG5V(mprj_io[20])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[21]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.ASIG5V(mprj_io[21])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[22]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.ASIG5V(mprj_io[22])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[23]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.ASIG5V(mprj_io[23])
	);
	gf180mcu_fd_io__bi_t \mprj_pads[24]  (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss),
	`endif
		.ASIG5V(mprj_io[24])
	);
	gf180mcu_fd_io__fill5 gf180mcu_fd_io__fill5_0 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill5 gf180mcu_fd_io__fill5_1 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill5 gf180mcu_fd_io__fill5_2 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_2 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_3 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_4 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_5 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_6 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_7 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_8 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_9 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_10 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_11 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_12 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_13 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_14 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_15 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_16 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_17 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_18 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_19 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_20 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_21 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_22 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_23 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_24 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_25 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_26 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_27 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_28 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_29 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_30 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_31 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_32 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_33 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_34 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_35 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_36 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_37 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_38 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_39 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_40 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_41 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_42 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_43 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_44 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_45 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_46 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_47 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_48 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_49 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_50 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_51 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_52 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_53 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_54 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_55 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_56 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_57 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_58 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_59 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_60 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_61 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_62 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_63 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_64 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_65 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_66 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_67 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_68 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_69 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_70 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_71 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_72 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_73 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_74 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_75 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_76 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_77 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_78 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_79 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_80 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_81 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_82 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_83 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_84 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_85 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_86 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_87 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_88 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_89 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_90 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_91 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_92 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_93 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_94 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_95 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_96 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_97 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_98 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_99 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_100 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_101 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_102 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_103 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_104 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_105 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_106 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_107 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_108 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_109 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_110 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_111 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_112 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_113 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_114 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_115 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_116 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_117 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_118 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_119 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_120 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_121 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_122 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_123 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_124 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_125 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_126 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_127 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_128 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_129 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_130 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_131 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_132 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_133 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_134 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_135 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_136 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_137 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_138 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_139 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_140 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_141 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_142 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_143 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_144 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_145 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_146 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_147 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_148 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_149 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_150 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_151 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_152 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_153 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_154 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_155 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_156 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_157 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_158 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_159 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_160 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_161 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_162 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_163 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_164 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_165 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_166 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_167 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_168 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_169 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_170 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_171 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_172 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_173 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_174 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_175 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_176 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_177 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_178 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_179 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_180 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_181 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_182 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_183 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_184 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_185 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_186 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_187 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_188 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_189 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_190 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_191 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_192 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_193 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_194 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_195 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_196 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_197 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_198 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_199 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_200 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_201 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_202 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_203 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_204 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_205 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_206 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_207 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_208 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_209 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_210 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_211 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_212 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_213 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_214 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_215 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_216 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_217 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_218 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_219 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_220 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_221 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_222 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_223 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_224 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_225 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_226 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_227 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_228 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_229 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_230 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_231 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_232 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_233 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_234 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_238 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_239 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_240 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_241 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_242 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_243 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_244 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_245 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_246 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_247 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_248 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_249 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_250 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_251 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_252 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_253 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_254 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_255 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_256 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_257 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_258 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_259 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_260 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_261 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_262 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_263 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_264 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_265 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_266 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_267 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_268 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_269 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_270 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_271 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_272 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_273 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_274 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_275 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_276 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_277 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_278 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_279 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_280 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_281 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_282 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_283 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_284 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_285 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_286 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_287 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_288 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_289 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_290 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_291 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_292 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_293 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_294 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_295 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_296 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_297 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_298 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_299 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_300 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_301 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_302 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_303 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_304 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_305 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_306 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_307 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_308 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_309 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_310 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_311 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_312 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_313 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_314 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_315 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_316 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_317 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_318 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_319 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_320 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_321 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_322 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_323 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_324 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_325 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_326 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_327 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_328 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_329 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_330 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_331 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_332 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_333 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_334 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_335 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_336 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_337 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_338 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_339 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_340 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_341 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_342 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_343 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_344 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_345 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_346 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_347 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_348 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_349 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_350 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_351 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_352 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_353 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_354 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_355 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_356 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_357 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_358 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_359 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_360 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_361 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_362 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_363 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_364 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_365 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_366 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_367 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_368 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_369 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_370 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_371 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_372 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_373 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_374 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_375 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_376 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_377 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_378 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_379 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_380 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_381 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_382 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_383 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_384 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_385 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_386 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_387 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_388 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_389 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_390 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_391 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_392 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_393 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_394 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_395 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_396 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_397 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_398 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_399 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_400 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_401 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_402 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_403 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_404 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_405 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_406 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_407 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_408 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_409 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_410 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_411 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_412 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_413 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_414 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_415 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_416 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_417 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_418 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_419 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_420 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_421 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_422 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_423 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_424 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_425 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_426 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_427 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_428 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_429 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_430 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_431 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_432 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_433 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_434 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_435 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_436 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_437 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_438 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_439 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_440 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_441 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_442 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_443 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_444 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_445 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_446 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_447 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_448 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_449 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_450 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_451 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_452 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_453 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_454 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_455 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_456 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_457 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_458 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_459 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_460 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_461 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_462 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_463 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_464 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_465 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_466 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_467 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_468 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_469 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_470 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_471 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_472 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_473 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_474 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_475 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_476 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_477 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_478 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_479 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_480 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_481 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_482 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_483 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_484 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_485 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_486 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_487 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_488 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_489 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_490 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_491 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_492 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_493 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_494 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_495 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_496 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_497 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_498 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_499 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_500 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_501 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_502 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_503 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_504 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_505 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_506 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_507 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_508 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_509 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_510 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_511 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_512 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_513 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_514 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_515 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_516 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_517 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_518 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_519 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_520 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_521 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_522 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_523 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_524 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_525 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_526 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_527 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_528 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_529 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_530 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_531 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_532 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_533 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_534 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_535 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_536 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_537 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_538 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_539 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_540 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_541 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_542 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_543 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_544 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_545 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_546 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_547 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_548 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_549 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_550 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_551 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_552 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_553 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_554 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_555 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_556 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_557 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_558 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_559 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_560 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_561 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_562 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_563 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_564 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_565 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_566 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_567 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_568 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_569 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_570 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_571 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_572 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_573 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_574 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_575 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_576 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_577 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_578 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_579 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_580 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_581 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_582 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_583 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_584 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_585 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_586 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_587 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_588 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_589 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_590 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_591 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_592 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_593 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_594 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_595 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_596 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_597 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_598 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_599 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_600 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_601 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_602 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_603 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_604 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_605 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_606 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_607 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_608 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_609 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_610 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_611 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_612 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_613 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_614 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_615 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_616 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_617 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_618 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_619 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_620 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_621 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_622 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_623 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_624 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_625 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_626 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_627 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_628 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_629 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_630 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_631 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_632 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_633 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_634 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_635 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_636 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_637 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_638 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_639 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_640 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_641 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_642 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_643 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_644 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_645 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_646 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_647 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_648 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_649 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_650 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_651 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_652 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_653 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_654 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_655 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_656 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_657 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_658 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_659 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_660 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_661 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_662 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_663 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_664 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_665 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_666 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_667 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_668 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_669 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_670 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_671 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_672 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_673 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_674 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_675 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_676 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_677 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_678 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_679 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_680 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_681 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_682 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_683 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_684 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_685 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_686 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_687 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_688 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_689 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_690 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_691 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_692 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_693 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_694 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_695 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_696 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_697 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_698 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_699 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_700 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_701 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_702 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_703 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_704 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_705 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_706 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_707 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_708 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_709 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_710 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_711 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_712 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_713 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_714 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_715 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_716 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_717 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_718 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_719 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_720 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_721 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_722 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_723 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_724 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_725 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_726 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_727 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_728 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_729 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_730 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_731 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_732 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_733 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_734 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_735 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_736 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_737 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_738 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_739 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_740 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_741 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_742 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_743 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_744 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_745 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_746 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_747 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_748 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_749 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_750 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_751 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_752 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_753 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_754 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_755 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_756 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_757 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_759 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_760 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_761 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_762 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_763 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_764 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_765 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_766 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_767 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_768 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_769 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_770 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_771 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_772 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_773 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_774 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_775 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_776 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_777 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_778 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_779 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_780 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_781 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_782 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_783 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_784 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_785 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_786 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_787 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_788 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_789 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_790 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_791 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_792 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_793 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_794 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_795 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_796 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_797 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_798 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_799 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_800 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_801 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_802 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_803 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_804 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_805 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_806 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_807 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_808 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_809 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_810 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_811 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_812 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_813 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_814 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_815 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_816 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_817 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_818 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_819 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_820 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_821 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_822 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_823 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_824 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_825 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_826 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_827 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_828 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_829 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_830 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_831 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_832 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_833 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_834 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_835 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_836 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_837 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_838 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_839 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_840 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_841 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_842 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_843 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_844 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_845 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_846 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_847 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_848 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_849 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_850 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_851 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_852 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_853 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_854 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_855 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_856 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_857 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_858 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_859 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_860 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_861 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_862 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_863 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_864 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_865 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_866 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_867 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_868 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_869 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_870 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_871 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_872 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_873 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_874 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_875 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_876 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_877 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_878 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_879 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_880 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_881 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_882 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_883 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_884 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_885 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_886 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_887 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_888 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_889 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_890 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_891 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_892 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_893 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_894 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_895 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_896 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_897 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_898 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_899 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_900 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_901 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_902 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_903 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_904 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_905 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_906 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_907 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_908 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_909 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_910 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_911 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_912 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_913 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_914 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_915 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_916 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_917 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_918 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_919 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_920 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_921 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_922 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_923 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_924 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_925 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_926 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_927 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_928 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_929 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_930 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_931 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_932 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_933 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_934 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_935 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_936 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_937 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_938 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_940 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_941 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_942 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_943 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_944 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_945 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_946 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_947 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_948 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_949 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_950 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_951 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_952 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_953 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_955 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_956 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_957 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_958 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_959 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_960 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_961 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_962 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_963 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_964 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_965 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_966 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_967 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_968 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_970 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_971 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_972 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_973 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_974 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_975 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_976 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_977 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_978 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_979 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_980 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_981 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_982 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_983 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_985 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_986 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_987 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_988 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_989 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_990 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_991 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_992 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_993 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_994 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_995 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_996 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_997 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_999 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1000 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1001 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1002 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1003 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1004 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1005 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1006 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1007 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1008 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1009 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1010 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1011 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1013 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1014 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1015 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1016 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1017 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1018 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1019 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1020 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1021 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1022 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1024 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1025 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1026 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1027 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1028 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1029 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1030 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1031 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1032 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1033 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1034 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1035 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1036 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1038 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1039 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1040 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1041 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1042 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1043 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);
	gf180mcu_fd_io__fill10 gf180mcu_fd_io__fill10_1044 (
	`ifdef USE_POWER_PINS
		.DVDD(vdd),
		.DVSS(vss),
		.VDD(vdd),
		.VSS(vss)
	`endif
	);

endmodule
// `default_nettype wire
