magic
tech gf180mcuC
magscale 1 10
timestamp 1670499160
<< checkpaint >>
rect 68000 68000 708000 946000
<< metal2 >>
rect 379272 941655 381172 944000
rect 379272 941599 379326 941655
rect 379382 941599 379450 941655
rect 379506 941599 379574 941655
rect 379630 941599 379698 941655
rect 379754 941599 379822 941655
rect 379878 941599 379946 941655
rect 380002 941599 381172 941655
rect 379272 941531 381172 941599
rect 379272 941475 379326 941531
rect 379382 941475 379450 941531
rect 379506 941475 379574 941531
rect 379630 941475 379698 941531
rect 379754 941475 379822 941531
rect 379878 941475 379946 941531
rect 380002 941475 381172 941531
rect 379272 941407 381172 941475
rect 379272 941351 379326 941407
rect 379382 941351 379450 941407
rect 379506 941351 379574 941407
rect 379630 941351 379698 941407
rect 379754 941351 379822 941407
rect 379878 941351 379946 941407
rect 380002 941351 381172 941407
rect 379272 941283 381172 941351
rect 379272 941227 379326 941283
rect 379382 941227 379450 941283
rect 379506 941227 379574 941283
rect 379630 941227 379698 941283
rect 379754 941227 379822 941283
rect 379878 941227 379946 941283
rect 380002 941227 381172 941283
rect 379272 941159 381172 941227
rect 379272 941103 379326 941159
rect 379382 941103 379450 941159
rect 379506 941103 379574 941159
rect 379630 941103 379698 941159
rect 379754 941103 379822 941159
rect 379878 941103 379946 941159
rect 380002 941103 381172 941159
rect 379272 941035 381172 941103
rect 379272 940979 379326 941035
rect 379382 940979 379450 941035
rect 379506 940979 379574 941035
rect 379630 940979 379698 941035
rect 379754 940979 379822 941035
rect 379878 940979 379946 941035
rect 380002 940979 381172 941035
rect 379272 940911 381172 940979
rect 379272 940855 379326 940911
rect 379382 940855 379450 940911
rect 379506 940855 379574 940911
rect 379630 940855 379698 940911
rect 379754 940855 379822 940911
rect 379878 940855 379946 940911
rect 380002 940855 381172 940911
rect 379272 940787 381172 940855
rect 379272 940731 379326 940787
rect 379382 940731 379450 940787
rect 379506 940731 379574 940787
rect 379630 940731 379698 940787
rect 379754 940731 379822 940787
rect 379878 940731 379946 940787
rect 380002 940731 381172 940787
rect 379272 940663 381172 940731
rect 379272 940607 379326 940663
rect 379382 940607 379450 940663
rect 379506 940607 379574 940663
rect 379630 940607 379698 940663
rect 379754 940607 379822 940663
rect 379878 940607 379946 940663
rect 380002 940607 381172 940663
rect 379272 940539 381172 940607
rect 379272 940483 379326 940539
rect 379382 940483 379450 940539
rect 379506 940483 379574 940539
rect 379630 940483 379698 940539
rect 379754 940483 379822 940539
rect 379878 940483 379946 940539
rect 380002 940483 381172 940539
rect 379272 940415 381172 940483
rect 379272 940359 379326 940415
rect 379382 940359 379450 940415
rect 379506 940359 379574 940415
rect 379630 940359 379698 940415
rect 379754 940359 379822 940415
rect 379878 940359 379946 940415
rect 380002 940359 381172 940415
rect 379272 940291 381172 940359
rect 379272 940235 379326 940291
rect 379382 940235 379450 940291
rect 379506 940235 379574 940291
rect 379630 940235 379698 940291
rect 379754 940235 379822 940291
rect 379878 940235 379946 940291
rect 380002 940235 381172 940291
rect 379272 940167 381172 940235
rect 379272 940111 379326 940167
rect 379382 940111 379450 940167
rect 379506 940111 379574 940167
rect 379630 940111 379698 940167
rect 379754 940111 379822 940167
rect 379878 940111 379946 940167
rect 380002 940111 381172 940167
rect 379272 940043 381172 940111
rect 379272 939987 379326 940043
rect 379382 939987 379450 940043
rect 379506 939987 379574 940043
rect 379630 939987 379698 940043
rect 379754 939987 379822 940043
rect 379878 939987 379946 940043
rect 380002 939987 381172 940043
rect 379272 939919 381172 939987
rect 379272 939863 379326 939919
rect 379382 939863 379450 939919
rect 379506 939863 379574 939919
rect 379630 939863 379698 939919
rect 379754 939863 379822 939919
rect 379878 939863 379946 939919
rect 380002 939863 381172 939919
rect 379272 939720 381172 939863
rect 381752 941655 383802 944000
rect 381752 941599 381832 941655
rect 381888 941599 381956 941655
rect 382012 941599 382080 941655
rect 382136 941599 382204 941655
rect 382260 941599 382328 941655
rect 382384 941599 382452 941655
rect 382508 941599 382576 941655
rect 382632 941599 382700 941655
rect 382756 941599 382824 941655
rect 382880 941599 382948 941655
rect 383004 941599 383072 941655
rect 383128 941599 383196 941655
rect 383252 941599 383320 941655
rect 383376 941599 383444 941655
rect 383500 941599 383568 941655
rect 383624 941599 383692 941655
rect 383748 941599 383802 941655
rect 381752 941531 383802 941599
rect 381752 941475 381832 941531
rect 381888 941475 381956 941531
rect 382012 941475 382080 941531
rect 382136 941475 382204 941531
rect 382260 941475 382328 941531
rect 382384 941475 382452 941531
rect 382508 941475 382576 941531
rect 382632 941475 382700 941531
rect 382756 941475 382824 941531
rect 382880 941475 382948 941531
rect 383004 941475 383072 941531
rect 383128 941475 383196 941531
rect 383252 941475 383320 941531
rect 383376 941475 383444 941531
rect 383500 941475 383568 941531
rect 383624 941475 383692 941531
rect 383748 941475 383802 941531
rect 381752 941407 383802 941475
rect 381752 941351 381832 941407
rect 381888 941351 381956 941407
rect 382012 941351 382080 941407
rect 382136 941351 382204 941407
rect 382260 941351 382328 941407
rect 382384 941351 382452 941407
rect 382508 941351 382576 941407
rect 382632 941351 382700 941407
rect 382756 941351 382824 941407
rect 382880 941351 382948 941407
rect 383004 941351 383072 941407
rect 383128 941351 383196 941407
rect 383252 941351 383320 941407
rect 383376 941351 383444 941407
rect 383500 941351 383568 941407
rect 383624 941351 383692 941407
rect 383748 941351 383802 941407
rect 381752 941283 383802 941351
rect 381752 941227 381832 941283
rect 381888 941227 381956 941283
rect 382012 941227 382080 941283
rect 382136 941227 382204 941283
rect 382260 941227 382328 941283
rect 382384 941227 382452 941283
rect 382508 941227 382576 941283
rect 382632 941227 382700 941283
rect 382756 941227 382824 941283
rect 382880 941227 382948 941283
rect 383004 941227 383072 941283
rect 383128 941227 383196 941283
rect 383252 941227 383320 941283
rect 383376 941227 383444 941283
rect 383500 941227 383568 941283
rect 383624 941227 383692 941283
rect 383748 941227 383802 941283
rect 381752 941159 383802 941227
rect 381752 941103 381832 941159
rect 381888 941103 381956 941159
rect 382012 941103 382080 941159
rect 382136 941103 382204 941159
rect 382260 941103 382328 941159
rect 382384 941103 382452 941159
rect 382508 941103 382576 941159
rect 382632 941103 382700 941159
rect 382756 941103 382824 941159
rect 382880 941103 382948 941159
rect 383004 941103 383072 941159
rect 383128 941103 383196 941159
rect 383252 941103 383320 941159
rect 383376 941103 383444 941159
rect 383500 941103 383568 941159
rect 383624 941103 383692 941159
rect 383748 941103 383802 941159
rect 381752 941035 383802 941103
rect 381752 940979 381832 941035
rect 381888 940979 381956 941035
rect 382012 940979 382080 941035
rect 382136 940979 382204 941035
rect 382260 940979 382328 941035
rect 382384 940979 382452 941035
rect 382508 940979 382576 941035
rect 382632 940979 382700 941035
rect 382756 940979 382824 941035
rect 382880 940979 382948 941035
rect 383004 940979 383072 941035
rect 383128 940979 383196 941035
rect 383252 940979 383320 941035
rect 383376 940979 383444 941035
rect 383500 940979 383568 941035
rect 383624 940979 383692 941035
rect 383748 940979 383802 941035
rect 381752 940911 383802 940979
rect 381752 940855 381832 940911
rect 381888 940855 381956 940911
rect 382012 940855 382080 940911
rect 382136 940855 382204 940911
rect 382260 940855 382328 940911
rect 382384 940855 382452 940911
rect 382508 940855 382576 940911
rect 382632 940855 382700 940911
rect 382756 940855 382824 940911
rect 382880 940855 382948 940911
rect 383004 940855 383072 940911
rect 383128 940855 383196 940911
rect 383252 940855 383320 940911
rect 383376 940855 383444 940911
rect 383500 940855 383568 940911
rect 383624 940855 383692 940911
rect 383748 940855 383802 940911
rect 381752 940787 383802 940855
rect 381752 940731 381832 940787
rect 381888 940731 381956 940787
rect 382012 940731 382080 940787
rect 382136 940731 382204 940787
rect 382260 940731 382328 940787
rect 382384 940731 382452 940787
rect 382508 940731 382576 940787
rect 382632 940731 382700 940787
rect 382756 940731 382824 940787
rect 382880 940731 382948 940787
rect 383004 940731 383072 940787
rect 383128 940731 383196 940787
rect 383252 940731 383320 940787
rect 383376 940731 383444 940787
rect 383500 940731 383568 940787
rect 383624 940731 383692 940787
rect 383748 940731 383802 940787
rect 381752 940663 383802 940731
rect 381752 940607 381832 940663
rect 381888 940607 381956 940663
rect 382012 940607 382080 940663
rect 382136 940607 382204 940663
rect 382260 940607 382328 940663
rect 382384 940607 382452 940663
rect 382508 940607 382576 940663
rect 382632 940607 382700 940663
rect 382756 940607 382824 940663
rect 382880 940607 382948 940663
rect 383004 940607 383072 940663
rect 383128 940607 383196 940663
rect 383252 940607 383320 940663
rect 383376 940607 383444 940663
rect 383500 940607 383568 940663
rect 383624 940607 383692 940663
rect 383748 940607 383802 940663
rect 381752 940539 383802 940607
rect 381752 940483 381832 940539
rect 381888 940483 381956 940539
rect 382012 940483 382080 940539
rect 382136 940483 382204 940539
rect 382260 940483 382328 940539
rect 382384 940483 382452 940539
rect 382508 940483 382576 940539
rect 382632 940483 382700 940539
rect 382756 940483 382824 940539
rect 382880 940483 382948 940539
rect 383004 940483 383072 940539
rect 383128 940483 383196 940539
rect 383252 940483 383320 940539
rect 383376 940483 383444 940539
rect 383500 940483 383568 940539
rect 383624 940483 383692 940539
rect 383748 940483 383802 940539
rect 381752 940415 383802 940483
rect 381752 940359 381832 940415
rect 381888 940359 381956 940415
rect 382012 940359 382080 940415
rect 382136 940359 382204 940415
rect 382260 940359 382328 940415
rect 382384 940359 382452 940415
rect 382508 940359 382576 940415
rect 382632 940359 382700 940415
rect 382756 940359 382824 940415
rect 382880 940359 382948 940415
rect 383004 940359 383072 940415
rect 383128 940359 383196 940415
rect 383252 940359 383320 940415
rect 383376 940359 383444 940415
rect 383500 940359 383568 940415
rect 383624 940359 383692 940415
rect 383748 940359 383802 940415
rect 381752 940291 383802 940359
rect 381752 940235 381832 940291
rect 381888 940235 381956 940291
rect 382012 940235 382080 940291
rect 382136 940235 382204 940291
rect 382260 940235 382328 940291
rect 382384 940235 382452 940291
rect 382508 940235 382576 940291
rect 382632 940235 382700 940291
rect 382756 940235 382824 940291
rect 382880 940235 382948 940291
rect 383004 940235 383072 940291
rect 383128 940235 383196 940291
rect 383252 940235 383320 940291
rect 383376 940235 383444 940291
rect 383500 940235 383568 940291
rect 383624 940235 383692 940291
rect 383748 940235 383802 940291
rect 381752 940167 383802 940235
rect 381752 940111 381832 940167
rect 381888 940111 381956 940167
rect 382012 940111 382080 940167
rect 382136 940111 382204 940167
rect 382260 940111 382328 940167
rect 382384 940111 382452 940167
rect 382508 940111 382576 940167
rect 382632 940111 382700 940167
rect 382756 940111 382824 940167
rect 382880 940111 382948 940167
rect 383004 940111 383072 940167
rect 383128 940111 383196 940167
rect 383252 940111 383320 940167
rect 383376 940111 383444 940167
rect 383500 940111 383568 940167
rect 383624 940111 383692 940167
rect 383748 940111 383802 940167
rect 381752 940043 383802 940111
rect 381752 939987 381832 940043
rect 381888 939987 381956 940043
rect 382012 939987 382080 940043
rect 382136 939987 382204 940043
rect 382260 939987 382328 940043
rect 382384 939987 382452 940043
rect 382508 939987 382576 940043
rect 382632 939987 382700 940043
rect 382756 939987 382824 940043
rect 382880 939987 382948 940043
rect 383004 939987 383072 940043
rect 383128 939987 383196 940043
rect 383252 939987 383320 940043
rect 383376 939987 383444 940043
rect 383500 939987 383568 940043
rect 383624 939987 383692 940043
rect 383748 939987 383802 940043
rect 381752 939919 383802 939987
rect 381752 939863 381832 939919
rect 381888 939863 381956 939919
rect 382012 939863 382080 939919
rect 382136 939863 382204 939919
rect 382260 939863 382328 939919
rect 382384 939863 382452 939919
rect 382508 939863 382576 939919
rect 382632 939863 382700 939919
rect 382756 939863 382824 939919
rect 382880 939863 382948 939919
rect 383004 939863 383072 939919
rect 383128 939863 383196 939919
rect 383252 939863 383320 939919
rect 383376 939863 383444 939919
rect 383500 939863 383568 939919
rect 383624 939863 383692 939919
rect 383748 939863 383802 939919
rect 381752 939720 383802 939863
rect 384122 941655 386172 944000
rect 384122 941599 384202 941655
rect 384258 941599 384326 941655
rect 384382 941599 384450 941655
rect 384506 941599 384574 941655
rect 384630 941599 384698 941655
rect 384754 941599 384822 941655
rect 384878 941599 384946 941655
rect 385002 941599 385070 941655
rect 385126 941599 385194 941655
rect 385250 941599 385318 941655
rect 385374 941599 385442 941655
rect 385498 941599 385566 941655
rect 385622 941599 385690 941655
rect 385746 941599 385814 941655
rect 385870 941599 385938 941655
rect 385994 941599 386062 941655
rect 386118 941599 386172 941655
rect 384122 941531 386172 941599
rect 384122 941475 384202 941531
rect 384258 941475 384326 941531
rect 384382 941475 384450 941531
rect 384506 941475 384574 941531
rect 384630 941475 384698 941531
rect 384754 941475 384822 941531
rect 384878 941475 384946 941531
rect 385002 941475 385070 941531
rect 385126 941475 385194 941531
rect 385250 941475 385318 941531
rect 385374 941475 385442 941531
rect 385498 941475 385566 941531
rect 385622 941475 385690 941531
rect 385746 941475 385814 941531
rect 385870 941475 385938 941531
rect 385994 941475 386062 941531
rect 386118 941475 386172 941531
rect 384122 941407 386172 941475
rect 384122 941351 384202 941407
rect 384258 941351 384326 941407
rect 384382 941351 384450 941407
rect 384506 941351 384574 941407
rect 384630 941351 384698 941407
rect 384754 941351 384822 941407
rect 384878 941351 384946 941407
rect 385002 941351 385070 941407
rect 385126 941351 385194 941407
rect 385250 941351 385318 941407
rect 385374 941351 385442 941407
rect 385498 941351 385566 941407
rect 385622 941351 385690 941407
rect 385746 941351 385814 941407
rect 385870 941351 385938 941407
rect 385994 941351 386062 941407
rect 386118 941351 386172 941407
rect 384122 941283 386172 941351
rect 384122 941227 384202 941283
rect 384258 941227 384326 941283
rect 384382 941227 384450 941283
rect 384506 941227 384574 941283
rect 384630 941227 384698 941283
rect 384754 941227 384822 941283
rect 384878 941227 384946 941283
rect 385002 941227 385070 941283
rect 385126 941227 385194 941283
rect 385250 941227 385318 941283
rect 385374 941227 385442 941283
rect 385498 941227 385566 941283
rect 385622 941227 385690 941283
rect 385746 941227 385814 941283
rect 385870 941227 385938 941283
rect 385994 941227 386062 941283
rect 386118 941227 386172 941283
rect 384122 941159 386172 941227
rect 384122 941103 384202 941159
rect 384258 941103 384326 941159
rect 384382 941103 384450 941159
rect 384506 941103 384574 941159
rect 384630 941103 384698 941159
rect 384754 941103 384822 941159
rect 384878 941103 384946 941159
rect 385002 941103 385070 941159
rect 385126 941103 385194 941159
rect 385250 941103 385318 941159
rect 385374 941103 385442 941159
rect 385498 941103 385566 941159
rect 385622 941103 385690 941159
rect 385746 941103 385814 941159
rect 385870 941103 385938 941159
rect 385994 941103 386062 941159
rect 386118 941103 386172 941159
rect 384122 941035 386172 941103
rect 384122 940979 384202 941035
rect 384258 940979 384326 941035
rect 384382 940979 384450 941035
rect 384506 940979 384574 941035
rect 384630 940979 384698 941035
rect 384754 940979 384822 941035
rect 384878 940979 384946 941035
rect 385002 940979 385070 941035
rect 385126 940979 385194 941035
rect 385250 940979 385318 941035
rect 385374 940979 385442 941035
rect 385498 940979 385566 941035
rect 385622 940979 385690 941035
rect 385746 940979 385814 941035
rect 385870 940979 385938 941035
rect 385994 940979 386062 941035
rect 386118 940979 386172 941035
rect 384122 940911 386172 940979
rect 384122 940855 384202 940911
rect 384258 940855 384326 940911
rect 384382 940855 384450 940911
rect 384506 940855 384574 940911
rect 384630 940855 384698 940911
rect 384754 940855 384822 940911
rect 384878 940855 384946 940911
rect 385002 940855 385070 940911
rect 385126 940855 385194 940911
rect 385250 940855 385318 940911
rect 385374 940855 385442 940911
rect 385498 940855 385566 940911
rect 385622 940855 385690 940911
rect 385746 940855 385814 940911
rect 385870 940855 385938 940911
rect 385994 940855 386062 940911
rect 386118 940855 386172 940911
rect 384122 940787 386172 940855
rect 384122 940731 384202 940787
rect 384258 940731 384326 940787
rect 384382 940731 384450 940787
rect 384506 940731 384574 940787
rect 384630 940731 384698 940787
rect 384754 940731 384822 940787
rect 384878 940731 384946 940787
rect 385002 940731 385070 940787
rect 385126 940731 385194 940787
rect 385250 940731 385318 940787
rect 385374 940731 385442 940787
rect 385498 940731 385566 940787
rect 385622 940731 385690 940787
rect 385746 940731 385814 940787
rect 385870 940731 385938 940787
rect 385994 940731 386062 940787
rect 386118 940731 386172 940787
rect 384122 940663 386172 940731
rect 384122 940607 384202 940663
rect 384258 940607 384326 940663
rect 384382 940607 384450 940663
rect 384506 940607 384574 940663
rect 384630 940607 384698 940663
rect 384754 940607 384822 940663
rect 384878 940607 384946 940663
rect 385002 940607 385070 940663
rect 385126 940607 385194 940663
rect 385250 940607 385318 940663
rect 385374 940607 385442 940663
rect 385498 940607 385566 940663
rect 385622 940607 385690 940663
rect 385746 940607 385814 940663
rect 385870 940607 385938 940663
rect 385994 940607 386062 940663
rect 386118 940607 386172 940663
rect 384122 940539 386172 940607
rect 384122 940483 384202 940539
rect 384258 940483 384326 940539
rect 384382 940483 384450 940539
rect 384506 940483 384574 940539
rect 384630 940483 384698 940539
rect 384754 940483 384822 940539
rect 384878 940483 384946 940539
rect 385002 940483 385070 940539
rect 385126 940483 385194 940539
rect 385250 940483 385318 940539
rect 385374 940483 385442 940539
rect 385498 940483 385566 940539
rect 385622 940483 385690 940539
rect 385746 940483 385814 940539
rect 385870 940483 385938 940539
rect 385994 940483 386062 940539
rect 386118 940483 386172 940539
rect 384122 940415 386172 940483
rect 384122 940359 384202 940415
rect 384258 940359 384326 940415
rect 384382 940359 384450 940415
rect 384506 940359 384574 940415
rect 384630 940359 384698 940415
rect 384754 940359 384822 940415
rect 384878 940359 384946 940415
rect 385002 940359 385070 940415
rect 385126 940359 385194 940415
rect 385250 940359 385318 940415
rect 385374 940359 385442 940415
rect 385498 940359 385566 940415
rect 385622 940359 385690 940415
rect 385746 940359 385814 940415
rect 385870 940359 385938 940415
rect 385994 940359 386062 940415
rect 386118 940359 386172 940415
rect 384122 940291 386172 940359
rect 384122 940235 384202 940291
rect 384258 940235 384326 940291
rect 384382 940235 384450 940291
rect 384506 940235 384574 940291
rect 384630 940235 384698 940291
rect 384754 940235 384822 940291
rect 384878 940235 384946 940291
rect 385002 940235 385070 940291
rect 385126 940235 385194 940291
rect 385250 940235 385318 940291
rect 385374 940235 385442 940291
rect 385498 940235 385566 940291
rect 385622 940235 385690 940291
rect 385746 940235 385814 940291
rect 385870 940235 385938 940291
rect 385994 940235 386062 940291
rect 386118 940235 386172 940291
rect 384122 940167 386172 940235
rect 384122 940111 384202 940167
rect 384258 940111 384326 940167
rect 384382 940111 384450 940167
rect 384506 940111 384574 940167
rect 384630 940111 384698 940167
rect 384754 940111 384822 940167
rect 384878 940111 384946 940167
rect 385002 940111 385070 940167
rect 385126 940111 385194 940167
rect 385250 940111 385318 940167
rect 385374 940111 385442 940167
rect 385498 940111 385566 940167
rect 385622 940111 385690 940167
rect 385746 940111 385814 940167
rect 385870 940111 385938 940167
rect 385994 940111 386062 940167
rect 386118 940111 386172 940167
rect 384122 940043 386172 940111
rect 384122 939987 384202 940043
rect 384258 939987 384326 940043
rect 384382 939987 384450 940043
rect 384506 939987 384574 940043
rect 384630 939987 384698 940043
rect 384754 939987 384822 940043
rect 384878 939987 384946 940043
rect 385002 939987 385070 940043
rect 385126 939987 385194 940043
rect 385250 939987 385318 940043
rect 385374 939987 385442 940043
rect 385498 939987 385566 940043
rect 385622 939987 385690 940043
rect 385746 939987 385814 940043
rect 385870 939987 385938 940043
rect 385994 939987 386062 940043
rect 386118 939987 386172 940043
rect 384122 939919 386172 939987
rect 384122 939863 384202 939919
rect 384258 939863 384326 939919
rect 384382 939863 384450 939919
rect 384506 939863 384574 939919
rect 384630 939863 384698 939919
rect 384754 939863 384822 939919
rect 384878 939863 384946 939919
rect 385002 939863 385070 939919
rect 385126 939863 385194 939919
rect 385250 939863 385318 939919
rect 385374 939863 385442 939919
rect 385498 939863 385566 939919
rect 385622 939863 385690 939919
rect 385746 939863 385814 939919
rect 385870 939863 385938 939919
rect 385994 939863 386062 939919
rect 386118 939863 386172 939919
rect 384122 939720 386172 939863
rect 386828 941655 388878 944000
rect 386828 941599 386908 941655
rect 386964 941599 387032 941655
rect 387088 941599 387156 941655
rect 387212 941599 387280 941655
rect 387336 941599 387404 941655
rect 387460 941599 387528 941655
rect 387584 941599 387652 941655
rect 387708 941599 387776 941655
rect 387832 941599 387900 941655
rect 387956 941599 388024 941655
rect 388080 941599 388148 941655
rect 388204 941599 388272 941655
rect 388328 941599 388396 941655
rect 388452 941599 388520 941655
rect 388576 941599 388644 941655
rect 388700 941599 388768 941655
rect 388824 941599 388878 941655
rect 386828 941531 388878 941599
rect 386828 941475 386908 941531
rect 386964 941475 387032 941531
rect 387088 941475 387156 941531
rect 387212 941475 387280 941531
rect 387336 941475 387404 941531
rect 387460 941475 387528 941531
rect 387584 941475 387652 941531
rect 387708 941475 387776 941531
rect 387832 941475 387900 941531
rect 387956 941475 388024 941531
rect 388080 941475 388148 941531
rect 388204 941475 388272 941531
rect 388328 941475 388396 941531
rect 388452 941475 388520 941531
rect 388576 941475 388644 941531
rect 388700 941475 388768 941531
rect 388824 941475 388878 941531
rect 386828 941407 388878 941475
rect 386828 941351 386908 941407
rect 386964 941351 387032 941407
rect 387088 941351 387156 941407
rect 387212 941351 387280 941407
rect 387336 941351 387404 941407
rect 387460 941351 387528 941407
rect 387584 941351 387652 941407
rect 387708 941351 387776 941407
rect 387832 941351 387900 941407
rect 387956 941351 388024 941407
rect 388080 941351 388148 941407
rect 388204 941351 388272 941407
rect 388328 941351 388396 941407
rect 388452 941351 388520 941407
rect 388576 941351 388644 941407
rect 388700 941351 388768 941407
rect 388824 941351 388878 941407
rect 386828 941283 388878 941351
rect 386828 941227 386908 941283
rect 386964 941227 387032 941283
rect 387088 941227 387156 941283
rect 387212 941227 387280 941283
rect 387336 941227 387404 941283
rect 387460 941227 387528 941283
rect 387584 941227 387652 941283
rect 387708 941227 387776 941283
rect 387832 941227 387900 941283
rect 387956 941227 388024 941283
rect 388080 941227 388148 941283
rect 388204 941227 388272 941283
rect 388328 941227 388396 941283
rect 388452 941227 388520 941283
rect 388576 941227 388644 941283
rect 388700 941227 388768 941283
rect 388824 941227 388878 941283
rect 386828 941159 388878 941227
rect 386828 941103 386908 941159
rect 386964 941103 387032 941159
rect 387088 941103 387156 941159
rect 387212 941103 387280 941159
rect 387336 941103 387404 941159
rect 387460 941103 387528 941159
rect 387584 941103 387652 941159
rect 387708 941103 387776 941159
rect 387832 941103 387900 941159
rect 387956 941103 388024 941159
rect 388080 941103 388148 941159
rect 388204 941103 388272 941159
rect 388328 941103 388396 941159
rect 388452 941103 388520 941159
rect 388576 941103 388644 941159
rect 388700 941103 388768 941159
rect 388824 941103 388878 941159
rect 386828 941035 388878 941103
rect 386828 940979 386908 941035
rect 386964 940979 387032 941035
rect 387088 940979 387156 941035
rect 387212 940979 387280 941035
rect 387336 940979 387404 941035
rect 387460 940979 387528 941035
rect 387584 940979 387652 941035
rect 387708 940979 387776 941035
rect 387832 940979 387900 941035
rect 387956 940979 388024 941035
rect 388080 940979 388148 941035
rect 388204 940979 388272 941035
rect 388328 940979 388396 941035
rect 388452 940979 388520 941035
rect 388576 940979 388644 941035
rect 388700 940979 388768 941035
rect 388824 940979 388878 941035
rect 386828 940911 388878 940979
rect 386828 940855 386908 940911
rect 386964 940855 387032 940911
rect 387088 940855 387156 940911
rect 387212 940855 387280 940911
rect 387336 940855 387404 940911
rect 387460 940855 387528 940911
rect 387584 940855 387652 940911
rect 387708 940855 387776 940911
rect 387832 940855 387900 940911
rect 387956 940855 388024 940911
rect 388080 940855 388148 940911
rect 388204 940855 388272 940911
rect 388328 940855 388396 940911
rect 388452 940855 388520 940911
rect 388576 940855 388644 940911
rect 388700 940855 388768 940911
rect 388824 940855 388878 940911
rect 386828 940787 388878 940855
rect 386828 940731 386908 940787
rect 386964 940731 387032 940787
rect 387088 940731 387156 940787
rect 387212 940731 387280 940787
rect 387336 940731 387404 940787
rect 387460 940731 387528 940787
rect 387584 940731 387652 940787
rect 387708 940731 387776 940787
rect 387832 940731 387900 940787
rect 387956 940731 388024 940787
rect 388080 940731 388148 940787
rect 388204 940731 388272 940787
rect 388328 940731 388396 940787
rect 388452 940731 388520 940787
rect 388576 940731 388644 940787
rect 388700 940731 388768 940787
rect 388824 940731 388878 940787
rect 386828 940663 388878 940731
rect 386828 940607 386908 940663
rect 386964 940607 387032 940663
rect 387088 940607 387156 940663
rect 387212 940607 387280 940663
rect 387336 940607 387404 940663
rect 387460 940607 387528 940663
rect 387584 940607 387652 940663
rect 387708 940607 387776 940663
rect 387832 940607 387900 940663
rect 387956 940607 388024 940663
rect 388080 940607 388148 940663
rect 388204 940607 388272 940663
rect 388328 940607 388396 940663
rect 388452 940607 388520 940663
rect 388576 940607 388644 940663
rect 388700 940607 388768 940663
rect 388824 940607 388878 940663
rect 386828 940539 388878 940607
rect 386828 940483 386908 940539
rect 386964 940483 387032 940539
rect 387088 940483 387156 940539
rect 387212 940483 387280 940539
rect 387336 940483 387404 940539
rect 387460 940483 387528 940539
rect 387584 940483 387652 940539
rect 387708 940483 387776 940539
rect 387832 940483 387900 940539
rect 387956 940483 388024 940539
rect 388080 940483 388148 940539
rect 388204 940483 388272 940539
rect 388328 940483 388396 940539
rect 388452 940483 388520 940539
rect 388576 940483 388644 940539
rect 388700 940483 388768 940539
rect 388824 940483 388878 940539
rect 386828 940415 388878 940483
rect 386828 940359 386908 940415
rect 386964 940359 387032 940415
rect 387088 940359 387156 940415
rect 387212 940359 387280 940415
rect 387336 940359 387404 940415
rect 387460 940359 387528 940415
rect 387584 940359 387652 940415
rect 387708 940359 387776 940415
rect 387832 940359 387900 940415
rect 387956 940359 388024 940415
rect 388080 940359 388148 940415
rect 388204 940359 388272 940415
rect 388328 940359 388396 940415
rect 388452 940359 388520 940415
rect 388576 940359 388644 940415
rect 388700 940359 388768 940415
rect 388824 940359 388878 940415
rect 386828 940291 388878 940359
rect 386828 940235 386908 940291
rect 386964 940235 387032 940291
rect 387088 940235 387156 940291
rect 387212 940235 387280 940291
rect 387336 940235 387404 940291
rect 387460 940235 387528 940291
rect 387584 940235 387652 940291
rect 387708 940235 387776 940291
rect 387832 940235 387900 940291
rect 387956 940235 388024 940291
rect 388080 940235 388148 940291
rect 388204 940235 388272 940291
rect 388328 940235 388396 940291
rect 388452 940235 388520 940291
rect 388576 940235 388644 940291
rect 388700 940235 388768 940291
rect 388824 940235 388878 940291
rect 386828 940167 388878 940235
rect 386828 940111 386908 940167
rect 386964 940111 387032 940167
rect 387088 940111 387156 940167
rect 387212 940111 387280 940167
rect 387336 940111 387404 940167
rect 387460 940111 387528 940167
rect 387584 940111 387652 940167
rect 387708 940111 387776 940167
rect 387832 940111 387900 940167
rect 387956 940111 388024 940167
rect 388080 940111 388148 940167
rect 388204 940111 388272 940167
rect 388328 940111 388396 940167
rect 388452 940111 388520 940167
rect 388576 940111 388644 940167
rect 388700 940111 388768 940167
rect 388824 940111 388878 940167
rect 386828 940043 388878 940111
rect 386828 939987 386908 940043
rect 386964 939987 387032 940043
rect 387088 939987 387156 940043
rect 387212 939987 387280 940043
rect 387336 939987 387404 940043
rect 387460 939987 387528 940043
rect 387584 939987 387652 940043
rect 387708 939987 387776 940043
rect 387832 939987 387900 940043
rect 387956 939987 388024 940043
rect 388080 939987 388148 940043
rect 388204 939987 388272 940043
rect 388328 939987 388396 940043
rect 388452 939987 388520 940043
rect 388576 939987 388644 940043
rect 388700 939987 388768 940043
rect 388824 939987 388878 940043
rect 386828 939919 388878 939987
rect 386828 939863 386908 939919
rect 386964 939863 387032 939919
rect 387088 939863 387156 939919
rect 387212 939863 387280 939919
rect 387336 939863 387404 939919
rect 387460 939863 387528 939919
rect 387584 939863 387652 939919
rect 387708 939863 387776 939919
rect 387832 939863 387900 939919
rect 387956 939863 388024 939919
rect 388080 939863 388148 939919
rect 388204 939863 388272 939919
rect 388328 939863 388396 939919
rect 388452 939863 388520 939919
rect 388576 939863 388644 939919
rect 388700 939863 388768 939919
rect 388824 939863 388878 939919
rect 386828 939720 388878 939863
rect 389198 941655 391248 944000
rect 389198 941599 389278 941655
rect 389334 941599 389402 941655
rect 389458 941599 389526 941655
rect 389582 941599 389650 941655
rect 389706 941599 389774 941655
rect 389830 941599 389898 941655
rect 389954 941599 390022 941655
rect 390078 941599 390146 941655
rect 390202 941599 390270 941655
rect 390326 941599 390394 941655
rect 390450 941599 390518 941655
rect 390574 941599 390642 941655
rect 390698 941599 390766 941655
rect 390822 941599 390890 941655
rect 390946 941599 391014 941655
rect 391070 941599 391138 941655
rect 391194 941599 391248 941655
rect 389198 941531 391248 941599
rect 389198 941475 389278 941531
rect 389334 941475 389402 941531
rect 389458 941475 389526 941531
rect 389582 941475 389650 941531
rect 389706 941475 389774 941531
rect 389830 941475 389898 941531
rect 389954 941475 390022 941531
rect 390078 941475 390146 941531
rect 390202 941475 390270 941531
rect 390326 941475 390394 941531
rect 390450 941475 390518 941531
rect 390574 941475 390642 941531
rect 390698 941475 390766 941531
rect 390822 941475 390890 941531
rect 390946 941475 391014 941531
rect 391070 941475 391138 941531
rect 391194 941475 391248 941531
rect 389198 941407 391248 941475
rect 389198 941351 389278 941407
rect 389334 941351 389402 941407
rect 389458 941351 389526 941407
rect 389582 941351 389650 941407
rect 389706 941351 389774 941407
rect 389830 941351 389898 941407
rect 389954 941351 390022 941407
rect 390078 941351 390146 941407
rect 390202 941351 390270 941407
rect 390326 941351 390394 941407
rect 390450 941351 390518 941407
rect 390574 941351 390642 941407
rect 390698 941351 390766 941407
rect 390822 941351 390890 941407
rect 390946 941351 391014 941407
rect 391070 941351 391138 941407
rect 391194 941351 391248 941407
rect 389198 941283 391248 941351
rect 389198 941227 389278 941283
rect 389334 941227 389402 941283
rect 389458 941227 389526 941283
rect 389582 941227 389650 941283
rect 389706 941227 389774 941283
rect 389830 941227 389898 941283
rect 389954 941227 390022 941283
rect 390078 941227 390146 941283
rect 390202 941227 390270 941283
rect 390326 941227 390394 941283
rect 390450 941227 390518 941283
rect 390574 941227 390642 941283
rect 390698 941227 390766 941283
rect 390822 941227 390890 941283
rect 390946 941227 391014 941283
rect 391070 941227 391138 941283
rect 391194 941227 391248 941283
rect 389198 941159 391248 941227
rect 389198 941103 389278 941159
rect 389334 941103 389402 941159
rect 389458 941103 389526 941159
rect 389582 941103 389650 941159
rect 389706 941103 389774 941159
rect 389830 941103 389898 941159
rect 389954 941103 390022 941159
rect 390078 941103 390146 941159
rect 390202 941103 390270 941159
rect 390326 941103 390394 941159
rect 390450 941103 390518 941159
rect 390574 941103 390642 941159
rect 390698 941103 390766 941159
rect 390822 941103 390890 941159
rect 390946 941103 391014 941159
rect 391070 941103 391138 941159
rect 391194 941103 391248 941159
rect 389198 941035 391248 941103
rect 389198 940979 389278 941035
rect 389334 940979 389402 941035
rect 389458 940979 389526 941035
rect 389582 940979 389650 941035
rect 389706 940979 389774 941035
rect 389830 940979 389898 941035
rect 389954 940979 390022 941035
rect 390078 940979 390146 941035
rect 390202 940979 390270 941035
rect 390326 940979 390394 941035
rect 390450 940979 390518 941035
rect 390574 940979 390642 941035
rect 390698 940979 390766 941035
rect 390822 940979 390890 941035
rect 390946 940979 391014 941035
rect 391070 940979 391138 941035
rect 391194 940979 391248 941035
rect 389198 940911 391248 940979
rect 389198 940855 389278 940911
rect 389334 940855 389402 940911
rect 389458 940855 389526 940911
rect 389582 940855 389650 940911
rect 389706 940855 389774 940911
rect 389830 940855 389898 940911
rect 389954 940855 390022 940911
rect 390078 940855 390146 940911
rect 390202 940855 390270 940911
rect 390326 940855 390394 940911
rect 390450 940855 390518 940911
rect 390574 940855 390642 940911
rect 390698 940855 390766 940911
rect 390822 940855 390890 940911
rect 390946 940855 391014 940911
rect 391070 940855 391138 940911
rect 391194 940855 391248 940911
rect 389198 940787 391248 940855
rect 389198 940731 389278 940787
rect 389334 940731 389402 940787
rect 389458 940731 389526 940787
rect 389582 940731 389650 940787
rect 389706 940731 389774 940787
rect 389830 940731 389898 940787
rect 389954 940731 390022 940787
rect 390078 940731 390146 940787
rect 390202 940731 390270 940787
rect 390326 940731 390394 940787
rect 390450 940731 390518 940787
rect 390574 940731 390642 940787
rect 390698 940731 390766 940787
rect 390822 940731 390890 940787
rect 390946 940731 391014 940787
rect 391070 940731 391138 940787
rect 391194 940731 391248 940787
rect 389198 940663 391248 940731
rect 389198 940607 389278 940663
rect 389334 940607 389402 940663
rect 389458 940607 389526 940663
rect 389582 940607 389650 940663
rect 389706 940607 389774 940663
rect 389830 940607 389898 940663
rect 389954 940607 390022 940663
rect 390078 940607 390146 940663
rect 390202 940607 390270 940663
rect 390326 940607 390394 940663
rect 390450 940607 390518 940663
rect 390574 940607 390642 940663
rect 390698 940607 390766 940663
rect 390822 940607 390890 940663
rect 390946 940607 391014 940663
rect 391070 940607 391138 940663
rect 391194 940607 391248 940663
rect 389198 940539 391248 940607
rect 389198 940483 389278 940539
rect 389334 940483 389402 940539
rect 389458 940483 389526 940539
rect 389582 940483 389650 940539
rect 389706 940483 389774 940539
rect 389830 940483 389898 940539
rect 389954 940483 390022 940539
rect 390078 940483 390146 940539
rect 390202 940483 390270 940539
rect 390326 940483 390394 940539
rect 390450 940483 390518 940539
rect 390574 940483 390642 940539
rect 390698 940483 390766 940539
rect 390822 940483 390890 940539
rect 390946 940483 391014 940539
rect 391070 940483 391138 940539
rect 391194 940483 391248 940539
rect 389198 940415 391248 940483
rect 389198 940359 389278 940415
rect 389334 940359 389402 940415
rect 389458 940359 389526 940415
rect 389582 940359 389650 940415
rect 389706 940359 389774 940415
rect 389830 940359 389898 940415
rect 389954 940359 390022 940415
rect 390078 940359 390146 940415
rect 390202 940359 390270 940415
rect 390326 940359 390394 940415
rect 390450 940359 390518 940415
rect 390574 940359 390642 940415
rect 390698 940359 390766 940415
rect 390822 940359 390890 940415
rect 390946 940359 391014 940415
rect 391070 940359 391138 940415
rect 391194 940359 391248 940415
rect 389198 940291 391248 940359
rect 389198 940235 389278 940291
rect 389334 940235 389402 940291
rect 389458 940235 389526 940291
rect 389582 940235 389650 940291
rect 389706 940235 389774 940291
rect 389830 940235 389898 940291
rect 389954 940235 390022 940291
rect 390078 940235 390146 940291
rect 390202 940235 390270 940291
rect 390326 940235 390394 940291
rect 390450 940235 390518 940291
rect 390574 940235 390642 940291
rect 390698 940235 390766 940291
rect 390822 940235 390890 940291
rect 390946 940235 391014 940291
rect 391070 940235 391138 940291
rect 391194 940235 391248 940291
rect 389198 940167 391248 940235
rect 389198 940111 389278 940167
rect 389334 940111 389402 940167
rect 389458 940111 389526 940167
rect 389582 940111 389650 940167
rect 389706 940111 389774 940167
rect 389830 940111 389898 940167
rect 389954 940111 390022 940167
rect 390078 940111 390146 940167
rect 390202 940111 390270 940167
rect 390326 940111 390394 940167
rect 390450 940111 390518 940167
rect 390574 940111 390642 940167
rect 390698 940111 390766 940167
rect 390822 940111 390890 940167
rect 390946 940111 391014 940167
rect 391070 940111 391138 940167
rect 391194 940111 391248 940167
rect 389198 940043 391248 940111
rect 389198 939987 389278 940043
rect 389334 939987 389402 940043
rect 389458 939987 389526 940043
rect 389582 939987 389650 940043
rect 389706 939987 389774 940043
rect 389830 939987 389898 940043
rect 389954 939987 390022 940043
rect 390078 939987 390146 940043
rect 390202 939987 390270 940043
rect 390326 939987 390394 940043
rect 390450 939987 390518 940043
rect 390574 939987 390642 940043
rect 390698 939987 390766 940043
rect 390822 939987 390890 940043
rect 390946 939987 391014 940043
rect 391070 939987 391138 940043
rect 391194 939987 391248 940043
rect 389198 939919 391248 939987
rect 389198 939863 389278 939919
rect 389334 939863 389402 939919
rect 389458 939863 389526 939919
rect 389582 939863 389650 939919
rect 389706 939863 389774 939919
rect 389830 939863 389898 939919
rect 389954 939863 390022 939919
rect 390078 939863 390146 939919
rect 390202 939863 390270 939919
rect 390326 939863 390394 939919
rect 390450 939863 390518 939919
rect 390574 939863 390642 939919
rect 390698 939863 390766 939919
rect 390822 939863 390890 939919
rect 390946 939863 391014 939919
rect 391070 939863 391138 939919
rect 391194 939863 391248 939919
rect 389198 939720 391248 939863
rect 391828 941655 393728 944000
rect 391828 941599 391882 941655
rect 391938 941599 392006 941655
rect 392062 941599 392130 941655
rect 392186 941599 392254 941655
rect 392310 941599 392378 941655
rect 392434 941599 392502 941655
rect 392558 941599 392626 941655
rect 392682 941599 392750 941655
rect 392806 941599 392874 941655
rect 392930 941599 392998 941655
rect 393054 941599 393122 941655
rect 393178 941599 393246 941655
rect 393302 941599 393370 941655
rect 393426 941599 393494 941655
rect 393550 941599 393618 941655
rect 393674 941599 393728 941655
rect 391828 941531 393728 941599
rect 391828 941475 391882 941531
rect 391938 941475 392006 941531
rect 392062 941475 392130 941531
rect 392186 941475 392254 941531
rect 392310 941475 392378 941531
rect 392434 941475 392502 941531
rect 392558 941475 392626 941531
rect 392682 941475 392750 941531
rect 392806 941475 392874 941531
rect 392930 941475 392998 941531
rect 393054 941475 393122 941531
rect 393178 941475 393246 941531
rect 393302 941475 393370 941531
rect 393426 941475 393494 941531
rect 393550 941475 393618 941531
rect 393674 941475 393728 941531
rect 391828 941407 393728 941475
rect 391828 941351 391882 941407
rect 391938 941351 392006 941407
rect 392062 941351 392130 941407
rect 392186 941351 392254 941407
rect 392310 941351 392378 941407
rect 392434 941351 392502 941407
rect 392558 941351 392626 941407
rect 392682 941351 392750 941407
rect 392806 941351 392874 941407
rect 392930 941351 392998 941407
rect 393054 941351 393122 941407
rect 393178 941351 393246 941407
rect 393302 941351 393370 941407
rect 393426 941351 393494 941407
rect 393550 941351 393618 941407
rect 393674 941351 393728 941407
rect 391828 941283 393728 941351
rect 391828 941227 391882 941283
rect 391938 941227 392006 941283
rect 392062 941227 392130 941283
rect 392186 941227 392254 941283
rect 392310 941227 392378 941283
rect 392434 941227 392502 941283
rect 392558 941227 392626 941283
rect 392682 941227 392750 941283
rect 392806 941227 392874 941283
rect 392930 941227 392998 941283
rect 393054 941227 393122 941283
rect 393178 941227 393246 941283
rect 393302 941227 393370 941283
rect 393426 941227 393494 941283
rect 393550 941227 393618 941283
rect 393674 941227 393728 941283
rect 391828 941159 393728 941227
rect 391828 941103 391882 941159
rect 391938 941103 392006 941159
rect 392062 941103 392130 941159
rect 392186 941103 392254 941159
rect 392310 941103 392378 941159
rect 392434 941103 392502 941159
rect 392558 941103 392626 941159
rect 392682 941103 392750 941159
rect 392806 941103 392874 941159
rect 392930 941103 392998 941159
rect 393054 941103 393122 941159
rect 393178 941103 393246 941159
rect 393302 941103 393370 941159
rect 393426 941103 393494 941159
rect 393550 941103 393618 941159
rect 393674 941103 393728 941159
rect 391828 941035 393728 941103
rect 391828 940979 391882 941035
rect 391938 940979 392006 941035
rect 392062 940979 392130 941035
rect 392186 940979 392254 941035
rect 392310 940979 392378 941035
rect 392434 940979 392502 941035
rect 392558 940979 392626 941035
rect 392682 940979 392750 941035
rect 392806 940979 392874 941035
rect 392930 940979 392998 941035
rect 393054 940979 393122 941035
rect 393178 940979 393246 941035
rect 393302 940979 393370 941035
rect 393426 940979 393494 941035
rect 393550 940979 393618 941035
rect 393674 940979 393728 941035
rect 391828 940911 393728 940979
rect 391828 940855 391882 940911
rect 391938 940855 392006 940911
rect 392062 940855 392130 940911
rect 392186 940855 392254 940911
rect 392310 940855 392378 940911
rect 392434 940855 392502 940911
rect 392558 940855 392626 940911
rect 392682 940855 392750 940911
rect 392806 940855 392874 940911
rect 392930 940855 392998 940911
rect 393054 940855 393122 940911
rect 393178 940855 393246 940911
rect 393302 940855 393370 940911
rect 393426 940855 393494 940911
rect 393550 940855 393618 940911
rect 393674 940855 393728 940911
rect 391828 940787 393728 940855
rect 391828 940731 391882 940787
rect 391938 940731 392006 940787
rect 392062 940731 392130 940787
rect 392186 940731 392254 940787
rect 392310 940731 392378 940787
rect 392434 940731 392502 940787
rect 392558 940731 392626 940787
rect 392682 940731 392750 940787
rect 392806 940731 392874 940787
rect 392930 940731 392998 940787
rect 393054 940731 393122 940787
rect 393178 940731 393246 940787
rect 393302 940731 393370 940787
rect 393426 940731 393494 940787
rect 393550 940731 393618 940787
rect 393674 940731 393728 940787
rect 391828 940663 393728 940731
rect 391828 940607 391882 940663
rect 391938 940607 392006 940663
rect 392062 940607 392130 940663
rect 392186 940607 392254 940663
rect 392310 940607 392378 940663
rect 392434 940607 392502 940663
rect 392558 940607 392626 940663
rect 392682 940607 392750 940663
rect 392806 940607 392874 940663
rect 392930 940607 392998 940663
rect 393054 940607 393122 940663
rect 393178 940607 393246 940663
rect 393302 940607 393370 940663
rect 393426 940607 393494 940663
rect 393550 940607 393618 940663
rect 393674 940607 393728 940663
rect 391828 940539 393728 940607
rect 391828 940483 391882 940539
rect 391938 940483 392006 940539
rect 392062 940483 392130 940539
rect 392186 940483 392254 940539
rect 392310 940483 392378 940539
rect 392434 940483 392502 940539
rect 392558 940483 392626 940539
rect 392682 940483 392750 940539
rect 392806 940483 392874 940539
rect 392930 940483 392998 940539
rect 393054 940483 393122 940539
rect 393178 940483 393246 940539
rect 393302 940483 393370 940539
rect 393426 940483 393494 940539
rect 393550 940483 393618 940539
rect 393674 940483 393728 940539
rect 391828 940415 393728 940483
rect 391828 940359 391882 940415
rect 391938 940359 392006 940415
rect 392062 940359 392130 940415
rect 392186 940359 392254 940415
rect 392310 940359 392378 940415
rect 392434 940359 392502 940415
rect 392558 940359 392626 940415
rect 392682 940359 392750 940415
rect 392806 940359 392874 940415
rect 392930 940359 392998 940415
rect 393054 940359 393122 940415
rect 393178 940359 393246 940415
rect 393302 940359 393370 940415
rect 393426 940359 393494 940415
rect 393550 940359 393618 940415
rect 393674 940359 393728 940415
rect 391828 940291 393728 940359
rect 391828 940235 391882 940291
rect 391938 940235 392006 940291
rect 392062 940235 392130 940291
rect 392186 940235 392254 940291
rect 392310 940235 392378 940291
rect 392434 940235 392502 940291
rect 392558 940235 392626 940291
rect 392682 940235 392750 940291
rect 392806 940235 392874 940291
rect 392930 940235 392998 940291
rect 393054 940235 393122 940291
rect 393178 940235 393246 940291
rect 393302 940235 393370 940291
rect 393426 940235 393494 940291
rect 393550 940235 393618 940291
rect 393674 940235 393728 940291
rect 391828 940167 393728 940235
rect 391828 940111 391882 940167
rect 391938 940111 392006 940167
rect 392062 940111 392130 940167
rect 392186 940111 392254 940167
rect 392310 940111 392378 940167
rect 392434 940111 392502 940167
rect 392558 940111 392626 940167
rect 392682 940111 392750 940167
rect 392806 940111 392874 940167
rect 392930 940111 392998 940167
rect 393054 940111 393122 940167
rect 393178 940111 393246 940167
rect 393302 940111 393370 940167
rect 393426 940111 393494 940167
rect 393550 940111 393618 940167
rect 393674 940111 393728 940167
rect 391828 940043 393728 940111
rect 391828 939987 391882 940043
rect 391938 939987 392006 940043
rect 392062 939987 392130 940043
rect 392186 939987 392254 940043
rect 392310 939987 392378 940043
rect 392434 939987 392502 940043
rect 392558 939987 392626 940043
rect 392682 939987 392750 940043
rect 392806 939987 392874 940043
rect 392930 939987 392998 940043
rect 393054 939987 393122 940043
rect 393178 939987 393246 940043
rect 393302 939987 393370 940043
rect 393426 939987 393494 940043
rect 393550 939987 393618 940043
rect 393674 939987 393728 940043
rect 391828 939919 393728 939987
rect 391828 939863 391882 939919
rect 391938 939863 392006 939919
rect 392062 939863 392130 939919
rect 392186 939863 392254 939919
rect 392310 939863 392378 939919
rect 392434 939863 392502 939919
rect 392558 939863 392626 939919
rect 392682 939863 392750 939919
rect 392806 939863 392874 939919
rect 392930 939863 392998 939919
rect 393054 939863 393122 939919
rect 393178 939863 393246 939919
rect 393302 939863 393370 939919
rect 393426 939863 393494 939919
rect 393550 939863 393618 939919
rect 393674 939863 393728 939919
rect 391828 939720 393728 939863
rect 599272 941655 601172 944000
rect 599272 941599 599326 941655
rect 599382 941599 599450 941655
rect 599506 941599 599574 941655
rect 599630 941599 599698 941655
rect 599754 941599 599822 941655
rect 599878 941599 599946 941655
rect 600002 941599 600070 941655
rect 600126 941599 600194 941655
rect 600250 941599 600318 941655
rect 600374 941599 600442 941655
rect 600498 941599 600566 941655
rect 600622 941599 600690 941655
rect 600746 941599 600814 941655
rect 600870 941599 600938 941655
rect 600994 941599 601062 941655
rect 601118 941599 601172 941655
rect 599272 941531 601172 941599
rect 599272 941475 599326 941531
rect 599382 941475 599450 941531
rect 599506 941475 599574 941531
rect 599630 941475 599698 941531
rect 599754 941475 599822 941531
rect 599878 941475 599946 941531
rect 600002 941475 600070 941531
rect 600126 941475 600194 941531
rect 600250 941475 600318 941531
rect 600374 941475 600442 941531
rect 600498 941475 600566 941531
rect 600622 941475 600690 941531
rect 600746 941475 600814 941531
rect 600870 941475 600938 941531
rect 600994 941475 601062 941531
rect 601118 941475 601172 941531
rect 599272 941407 601172 941475
rect 599272 941351 599326 941407
rect 599382 941351 599450 941407
rect 599506 941351 599574 941407
rect 599630 941351 599698 941407
rect 599754 941351 599822 941407
rect 599878 941351 599946 941407
rect 600002 941351 600070 941407
rect 600126 941351 600194 941407
rect 600250 941351 600318 941407
rect 600374 941351 600442 941407
rect 600498 941351 600566 941407
rect 600622 941351 600690 941407
rect 600746 941351 600814 941407
rect 600870 941351 600938 941407
rect 600994 941351 601062 941407
rect 601118 941351 601172 941407
rect 599272 941283 601172 941351
rect 599272 941227 599326 941283
rect 599382 941227 599450 941283
rect 599506 941227 599574 941283
rect 599630 941227 599698 941283
rect 599754 941227 599822 941283
rect 599878 941227 599946 941283
rect 600002 941227 600070 941283
rect 600126 941227 600194 941283
rect 600250 941227 600318 941283
rect 600374 941227 600442 941283
rect 600498 941227 600566 941283
rect 600622 941227 600690 941283
rect 600746 941227 600814 941283
rect 600870 941227 600938 941283
rect 600994 941227 601062 941283
rect 601118 941227 601172 941283
rect 599272 941159 601172 941227
rect 599272 941103 599326 941159
rect 599382 941103 599450 941159
rect 599506 941103 599574 941159
rect 599630 941103 599698 941159
rect 599754 941103 599822 941159
rect 599878 941103 599946 941159
rect 600002 941103 600070 941159
rect 600126 941103 600194 941159
rect 600250 941103 600318 941159
rect 600374 941103 600442 941159
rect 600498 941103 600566 941159
rect 600622 941103 600690 941159
rect 600746 941103 600814 941159
rect 600870 941103 600938 941159
rect 600994 941103 601062 941159
rect 601118 941103 601172 941159
rect 599272 941035 601172 941103
rect 599272 940979 599326 941035
rect 599382 940979 599450 941035
rect 599506 940979 599574 941035
rect 599630 940979 599698 941035
rect 599754 940979 599822 941035
rect 599878 940979 599946 941035
rect 600002 940979 600070 941035
rect 600126 940979 600194 941035
rect 600250 940979 600318 941035
rect 600374 940979 600442 941035
rect 600498 940979 600566 941035
rect 600622 940979 600690 941035
rect 600746 940979 600814 941035
rect 600870 940979 600938 941035
rect 600994 940979 601062 941035
rect 601118 940979 601172 941035
rect 599272 940911 601172 940979
rect 599272 940855 599326 940911
rect 599382 940855 599450 940911
rect 599506 940855 599574 940911
rect 599630 940855 599698 940911
rect 599754 940855 599822 940911
rect 599878 940855 599946 940911
rect 600002 940855 600070 940911
rect 600126 940855 600194 940911
rect 600250 940855 600318 940911
rect 600374 940855 600442 940911
rect 600498 940855 600566 940911
rect 600622 940855 600690 940911
rect 600746 940855 600814 940911
rect 600870 940855 600938 940911
rect 600994 940855 601062 940911
rect 601118 940855 601172 940911
rect 599272 940787 601172 940855
rect 599272 940731 599326 940787
rect 599382 940731 599450 940787
rect 599506 940731 599574 940787
rect 599630 940731 599698 940787
rect 599754 940731 599822 940787
rect 599878 940731 599946 940787
rect 600002 940731 600070 940787
rect 600126 940731 600194 940787
rect 600250 940731 600318 940787
rect 600374 940731 600442 940787
rect 600498 940731 600566 940787
rect 600622 940731 600690 940787
rect 600746 940731 600814 940787
rect 600870 940731 600938 940787
rect 600994 940731 601062 940787
rect 601118 940731 601172 940787
rect 599272 940663 601172 940731
rect 599272 940607 599326 940663
rect 599382 940607 599450 940663
rect 599506 940607 599574 940663
rect 599630 940607 599698 940663
rect 599754 940607 599822 940663
rect 599878 940607 599946 940663
rect 600002 940607 600070 940663
rect 600126 940607 600194 940663
rect 600250 940607 600318 940663
rect 600374 940607 600442 940663
rect 600498 940607 600566 940663
rect 600622 940607 600690 940663
rect 600746 940607 600814 940663
rect 600870 940607 600938 940663
rect 600994 940607 601062 940663
rect 601118 940607 601172 940663
rect 599272 940539 601172 940607
rect 599272 940483 599326 940539
rect 599382 940483 599450 940539
rect 599506 940483 599574 940539
rect 599630 940483 599698 940539
rect 599754 940483 599822 940539
rect 599878 940483 599946 940539
rect 600002 940483 600070 940539
rect 600126 940483 600194 940539
rect 600250 940483 600318 940539
rect 600374 940483 600442 940539
rect 600498 940483 600566 940539
rect 600622 940483 600690 940539
rect 600746 940483 600814 940539
rect 600870 940483 600938 940539
rect 600994 940483 601062 940539
rect 601118 940483 601172 940539
rect 599272 940415 601172 940483
rect 599272 940359 599326 940415
rect 599382 940359 599450 940415
rect 599506 940359 599574 940415
rect 599630 940359 599698 940415
rect 599754 940359 599822 940415
rect 599878 940359 599946 940415
rect 600002 940359 600070 940415
rect 600126 940359 600194 940415
rect 600250 940359 600318 940415
rect 600374 940359 600442 940415
rect 600498 940359 600566 940415
rect 600622 940359 600690 940415
rect 600746 940359 600814 940415
rect 600870 940359 600938 940415
rect 600994 940359 601062 940415
rect 601118 940359 601172 940415
rect 599272 940291 601172 940359
rect 599272 940235 599326 940291
rect 599382 940235 599450 940291
rect 599506 940235 599574 940291
rect 599630 940235 599698 940291
rect 599754 940235 599822 940291
rect 599878 940235 599946 940291
rect 600002 940235 600070 940291
rect 600126 940235 600194 940291
rect 600250 940235 600318 940291
rect 600374 940235 600442 940291
rect 600498 940235 600566 940291
rect 600622 940235 600690 940291
rect 600746 940235 600814 940291
rect 600870 940235 600938 940291
rect 600994 940235 601062 940291
rect 601118 940235 601172 940291
rect 599272 940167 601172 940235
rect 599272 940111 599326 940167
rect 599382 940111 599450 940167
rect 599506 940111 599574 940167
rect 599630 940111 599698 940167
rect 599754 940111 599822 940167
rect 599878 940111 599946 940167
rect 600002 940111 600070 940167
rect 600126 940111 600194 940167
rect 600250 940111 600318 940167
rect 600374 940111 600442 940167
rect 600498 940111 600566 940167
rect 600622 940111 600690 940167
rect 600746 940111 600814 940167
rect 600870 940111 600938 940167
rect 600994 940111 601062 940167
rect 601118 940111 601172 940167
rect 599272 940043 601172 940111
rect 599272 939987 599326 940043
rect 599382 939987 599450 940043
rect 599506 939987 599574 940043
rect 599630 939987 599698 940043
rect 599754 939987 599822 940043
rect 599878 939987 599946 940043
rect 600002 939987 600070 940043
rect 600126 939987 600194 940043
rect 600250 939987 600318 940043
rect 600374 939987 600442 940043
rect 600498 939987 600566 940043
rect 600622 939987 600690 940043
rect 600746 939987 600814 940043
rect 600870 939987 600938 940043
rect 600994 939987 601062 940043
rect 601118 939987 601172 940043
rect 599272 939919 601172 939987
rect 599272 939863 599326 939919
rect 599382 939863 599450 939919
rect 599506 939863 599574 939919
rect 599630 939863 599698 939919
rect 599754 939863 599822 939919
rect 599878 939863 599946 939919
rect 600002 939863 600070 939919
rect 600126 939863 600194 939919
rect 600250 939863 600318 939919
rect 600374 939863 600442 939919
rect 600498 939863 600566 939919
rect 600622 939863 600690 939919
rect 600746 939863 600814 939919
rect 600870 939863 600938 939919
rect 600994 939863 601062 939919
rect 601118 939863 601172 939919
rect 599272 939720 601172 939863
rect 601752 941655 603802 944000
rect 601752 941599 601832 941655
rect 601888 941599 601956 941655
rect 602012 941599 602080 941655
rect 602136 941599 602204 941655
rect 602260 941599 602328 941655
rect 602384 941599 602452 941655
rect 602508 941599 602576 941655
rect 602632 941599 602700 941655
rect 602756 941599 602824 941655
rect 602880 941599 602948 941655
rect 603004 941599 603072 941655
rect 603128 941599 603196 941655
rect 603252 941599 603320 941655
rect 603376 941599 603444 941655
rect 603500 941599 603568 941655
rect 603624 941599 603692 941655
rect 603748 941599 603802 941655
rect 601752 941531 603802 941599
rect 601752 941475 601832 941531
rect 601888 941475 601956 941531
rect 602012 941475 602080 941531
rect 602136 941475 602204 941531
rect 602260 941475 602328 941531
rect 602384 941475 602452 941531
rect 602508 941475 602576 941531
rect 602632 941475 602700 941531
rect 602756 941475 602824 941531
rect 602880 941475 602948 941531
rect 603004 941475 603072 941531
rect 603128 941475 603196 941531
rect 603252 941475 603320 941531
rect 603376 941475 603444 941531
rect 603500 941475 603568 941531
rect 603624 941475 603692 941531
rect 603748 941475 603802 941531
rect 601752 941407 603802 941475
rect 601752 941351 601832 941407
rect 601888 941351 601956 941407
rect 602012 941351 602080 941407
rect 602136 941351 602204 941407
rect 602260 941351 602328 941407
rect 602384 941351 602452 941407
rect 602508 941351 602576 941407
rect 602632 941351 602700 941407
rect 602756 941351 602824 941407
rect 602880 941351 602948 941407
rect 603004 941351 603072 941407
rect 603128 941351 603196 941407
rect 603252 941351 603320 941407
rect 603376 941351 603444 941407
rect 603500 941351 603568 941407
rect 603624 941351 603692 941407
rect 603748 941351 603802 941407
rect 601752 941283 603802 941351
rect 601752 941227 601832 941283
rect 601888 941227 601956 941283
rect 602012 941227 602080 941283
rect 602136 941227 602204 941283
rect 602260 941227 602328 941283
rect 602384 941227 602452 941283
rect 602508 941227 602576 941283
rect 602632 941227 602700 941283
rect 602756 941227 602824 941283
rect 602880 941227 602948 941283
rect 603004 941227 603072 941283
rect 603128 941227 603196 941283
rect 603252 941227 603320 941283
rect 603376 941227 603444 941283
rect 603500 941227 603568 941283
rect 603624 941227 603692 941283
rect 603748 941227 603802 941283
rect 601752 941159 603802 941227
rect 601752 941103 601832 941159
rect 601888 941103 601956 941159
rect 602012 941103 602080 941159
rect 602136 941103 602204 941159
rect 602260 941103 602328 941159
rect 602384 941103 602452 941159
rect 602508 941103 602576 941159
rect 602632 941103 602700 941159
rect 602756 941103 602824 941159
rect 602880 941103 602948 941159
rect 603004 941103 603072 941159
rect 603128 941103 603196 941159
rect 603252 941103 603320 941159
rect 603376 941103 603444 941159
rect 603500 941103 603568 941159
rect 603624 941103 603692 941159
rect 603748 941103 603802 941159
rect 601752 941035 603802 941103
rect 601752 940979 601832 941035
rect 601888 940979 601956 941035
rect 602012 940979 602080 941035
rect 602136 940979 602204 941035
rect 602260 940979 602328 941035
rect 602384 940979 602452 941035
rect 602508 940979 602576 941035
rect 602632 940979 602700 941035
rect 602756 940979 602824 941035
rect 602880 940979 602948 941035
rect 603004 940979 603072 941035
rect 603128 940979 603196 941035
rect 603252 940979 603320 941035
rect 603376 940979 603444 941035
rect 603500 940979 603568 941035
rect 603624 940979 603692 941035
rect 603748 940979 603802 941035
rect 601752 940911 603802 940979
rect 601752 940855 601832 940911
rect 601888 940855 601956 940911
rect 602012 940855 602080 940911
rect 602136 940855 602204 940911
rect 602260 940855 602328 940911
rect 602384 940855 602452 940911
rect 602508 940855 602576 940911
rect 602632 940855 602700 940911
rect 602756 940855 602824 940911
rect 602880 940855 602948 940911
rect 603004 940855 603072 940911
rect 603128 940855 603196 940911
rect 603252 940855 603320 940911
rect 603376 940855 603444 940911
rect 603500 940855 603568 940911
rect 603624 940855 603692 940911
rect 603748 940855 603802 940911
rect 601752 940787 603802 940855
rect 601752 940731 601832 940787
rect 601888 940731 601956 940787
rect 602012 940731 602080 940787
rect 602136 940731 602204 940787
rect 602260 940731 602328 940787
rect 602384 940731 602452 940787
rect 602508 940731 602576 940787
rect 602632 940731 602700 940787
rect 602756 940731 602824 940787
rect 602880 940731 602948 940787
rect 603004 940731 603072 940787
rect 603128 940731 603196 940787
rect 603252 940731 603320 940787
rect 603376 940731 603444 940787
rect 603500 940731 603568 940787
rect 603624 940731 603692 940787
rect 603748 940731 603802 940787
rect 601752 940663 603802 940731
rect 601752 940607 601832 940663
rect 601888 940607 601956 940663
rect 602012 940607 602080 940663
rect 602136 940607 602204 940663
rect 602260 940607 602328 940663
rect 602384 940607 602452 940663
rect 602508 940607 602576 940663
rect 602632 940607 602700 940663
rect 602756 940607 602824 940663
rect 602880 940607 602948 940663
rect 603004 940607 603072 940663
rect 603128 940607 603196 940663
rect 603252 940607 603320 940663
rect 603376 940607 603444 940663
rect 603500 940607 603568 940663
rect 603624 940607 603692 940663
rect 603748 940607 603802 940663
rect 601752 940539 603802 940607
rect 601752 940483 601832 940539
rect 601888 940483 601956 940539
rect 602012 940483 602080 940539
rect 602136 940483 602204 940539
rect 602260 940483 602328 940539
rect 602384 940483 602452 940539
rect 602508 940483 602576 940539
rect 602632 940483 602700 940539
rect 602756 940483 602824 940539
rect 602880 940483 602948 940539
rect 603004 940483 603072 940539
rect 603128 940483 603196 940539
rect 603252 940483 603320 940539
rect 603376 940483 603444 940539
rect 603500 940483 603568 940539
rect 603624 940483 603692 940539
rect 603748 940483 603802 940539
rect 601752 940415 603802 940483
rect 601752 940359 601832 940415
rect 601888 940359 601956 940415
rect 602012 940359 602080 940415
rect 602136 940359 602204 940415
rect 602260 940359 602328 940415
rect 602384 940359 602452 940415
rect 602508 940359 602576 940415
rect 602632 940359 602700 940415
rect 602756 940359 602824 940415
rect 602880 940359 602948 940415
rect 603004 940359 603072 940415
rect 603128 940359 603196 940415
rect 603252 940359 603320 940415
rect 603376 940359 603444 940415
rect 603500 940359 603568 940415
rect 603624 940359 603692 940415
rect 603748 940359 603802 940415
rect 601752 940291 603802 940359
rect 601752 940235 601832 940291
rect 601888 940235 601956 940291
rect 602012 940235 602080 940291
rect 602136 940235 602204 940291
rect 602260 940235 602328 940291
rect 602384 940235 602452 940291
rect 602508 940235 602576 940291
rect 602632 940235 602700 940291
rect 602756 940235 602824 940291
rect 602880 940235 602948 940291
rect 603004 940235 603072 940291
rect 603128 940235 603196 940291
rect 603252 940235 603320 940291
rect 603376 940235 603444 940291
rect 603500 940235 603568 940291
rect 603624 940235 603692 940291
rect 603748 940235 603802 940291
rect 601752 940167 603802 940235
rect 601752 940111 601832 940167
rect 601888 940111 601956 940167
rect 602012 940111 602080 940167
rect 602136 940111 602204 940167
rect 602260 940111 602328 940167
rect 602384 940111 602452 940167
rect 602508 940111 602576 940167
rect 602632 940111 602700 940167
rect 602756 940111 602824 940167
rect 602880 940111 602948 940167
rect 603004 940111 603072 940167
rect 603128 940111 603196 940167
rect 603252 940111 603320 940167
rect 603376 940111 603444 940167
rect 603500 940111 603568 940167
rect 603624 940111 603692 940167
rect 603748 940111 603802 940167
rect 601752 940043 603802 940111
rect 601752 939987 601832 940043
rect 601888 939987 601956 940043
rect 602012 939987 602080 940043
rect 602136 939987 602204 940043
rect 602260 939987 602328 940043
rect 602384 939987 602452 940043
rect 602508 939987 602576 940043
rect 602632 939987 602700 940043
rect 602756 939987 602824 940043
rect 602880 939987 602948 940043
rect 603004 939987 603072 940043
rect 603128 939987 603196 940043
rect 603252 939987 603320 940043
rect 603376 939987 603444 940043
rect 603500 939987 603568 940043
rect 603624 939987 603692 940043
rect 603748 939987 603802 940043
rect 601752 939919 603802 939987
rect 601752 939863 601832 939919
rect 601888 939863 601956 939919
rect 602012 939863 602080 939919
rect 602136 939863 602204 939919
rect 602260 939863 602328 939919
rect 602384 939863 602452 939919
rect 602508 939863 602576 939919
rect 602632 939863 602700 939919
rect 602756 939863 602824 939919
rect 602880 939863 602948 939919
rect 603004 939863 603072 939919
rect 603128 939863 603196 939919
rect 603252 939863 603320 939919
rect 603376 939863 603444 939919
rect 603500 939863 603568 939919
rect 603624 939863 603692 939919
rect 603748 939863 603802 939919
rect 601752 939720 603802 939863
rect 604122 941655 606172 944000
rect 604122 941599 605070 941655
rect 605126 941599 605194 941655
rect 605250 941599 605318 941655
rect 605374 941599 605442 941655
rect 605498 941599 605566 941655
rect 605622 941599 605690 941655
rect 605746 941599 605814 941655
rect 605870 941599 605938 941655
rect 605994 941599 606062 941655
rect 606118 941599 606172 941655
rect 604122 941531 606172 941599
rect 604122 941475 605070 941531
rect 605126 941475 605194 941531
rect 605250 941475 605318 941531
rect 605374 941475 605442 941531
rect 605498 941475 605566 941531
rect 605622 941475 605690 941531
rect 605746 941475 605814 941531
rect 605870 941475 605938 941531
rect 605994 941475 606062 941531
rect 606118 941475 606172 941531
rect 604122 941407 606172 941475
rect 604122 941351 605070 941407
rect 605126 941351 605194 941407
rect 605250 941351 605318 941407
rect 605374 941351 605442 941407
rect 605498 941351 605566 941407
rect 605622 941351 605690 941407
rect 605746 941351 605814 941407
rect 605870 941351 605938 941407
rect 605994 941351 606062 941407
rect 606118 941351 606172 941407
rect 604122 941283 606172 941351
rect 604122 941227 605070 941283
rect 605126 941227 605194 941283
rect 605250 941227 605318 941283
rect 605374 941227 605442 941283
rect 605498 941227 605566 941283
rect 605622 941227 605690 941283
rect 605746 941227 605814 941283
rect 605870 941227 605938 941283
rect 605994 941227 606062 941283
rect 606118 941227 606172 941283
rect 604122 941159 606172 941227
rect 604122 941103 605070 941159
rect 605126 941103 605194 941159
rect 605250 941103 605318 941159
rect 605374 941103 605442 941159
rect 605498 941103 605566 941159
rect 605622 941103 605690 941159
rect 605746 941103 605814 941159
rect 605870 941103 605938 941159
rect 605994 941103 606062 941159
rect 606118 941103 606172 941159
rect 604122 941035 606172 941103
rect 604122 940979 605070 941035
rect 605126 940979 605194 941035
rect 605250 940979 605318 941035
rect 605374 940979 605442 941035
rect 605498 940979 605566 941035
rect 605622 940979 605690 941035
rect 605746 940979 605814 941035
rect 605870 940979 605938 941035
rect 605994 940979 606062 941035
rect 606118 940979 606172 941035
rect 604122 940911 606172 940979
rect 604122 940855 605070 940911
rect 605126 940855 605194 940911
rect 605250 940855 605318 940911
rect 605374 940855 605442 940911
rect 605498 940855 605566 940911
rect 605622 940855 605690 940911
rect 605746 940855 605814 940911
rect 605870 940855 605938 940911
rect 605994 940855 606062 940911
rect 606118 940855 606172 940911
rect 604122 940787 606172 940855
rect 604122 940731 605070 940787
rect 605126 940731 605194 940787
rect 605250 940731 605318 940787
rect 605374 940731 605442 940787
rect 605498 940731 605566 940787
rect 605622 940731 605690 940787
rect 605746 940731 605814 940787
rect 605870 940731 605938 940787
rect 605994 940731 606062 940787
rect 606118 940731 606172 940787
rect 604122 940663 606172 940731
rect 604122 940607 605070 940663
rect 605126 940607 605194 940663
rect 605250 940607 605318 940663
rect 605374 940607 605442 940663
rect 605498 940607 605566 940663
rect 605622 940607 605690 940663
rect 605746 940607 605814 940663
rect 605870 940607 605938 940663
rect 605994 940607 606062 940663
rect 606118 940607 606172 940663
rect 604122 940539 606172 940607
rect 604122 940483 605070 940539
rect 605126 940483 605194 940539
rect 605250 940483 605318 940539
rect 605374 940483 605442 940539
rect 605498 940483 605566 940539
rect 605622 940483 605690 940539
rect 605746 940483 605814 940539
rect 605870 940483 605938 940539
rect 605994 940483 606062 940539
rect 606118 940483 606172 940539
rect 604122 940415 606172 940483
rect 604122 940359 605070 940415
rect 605126 940359 605194 940415
rect 605250 940359 605318 940415
rect 605374 940359 605442 940415
rect 605498 940359 605566 940415
rect 605622 940359 605690 940415
rect 605746 940359 605814 940415
rect 605870 940359 605938 940415
rect 605994 940359 606062 940415
rect 606118 940359 606172 940415
rect 604122 940291 606172 940359
rect 604122 940235 605070 940291
rect 605126 940235 605194 940291
rect 605250 940235 605318 940291
rect 605374 940235 605442 940291
rect 605498 940235 605566 940291
rect 605622 940235 605690 940291
rect 605746 940235 605814 940291
rect 605870 940235 605938 940291
rect 605994 940235 606062 940291
rect 606118 940235 606172 940291
rect 604122 940167 606172 940235
rect 604122 940111 605070 940167
rect 605126 940111 605194 940167
rect 605250 940111 605318 940167
rect 605374 940111 605442 940167
rect 605498 940111 605566 940167
rect 605622 940111 605690 940167
rect 605746 940111 605814 940167
rect 605870 940111 605938 940167
rect 605994 940111 606062 940167
rect 606118 940111 606172 940167
rect 604122 940043 606172 940111
rect 604122 939987 605070 940043
rect 605126 939987 605194 940043
rect 605250 939987 605318 940043
rect 605374 939987 605442 940043
rect 605498 939987 605566 940043
rect 605622 939987 605690 940043
rect 605746 939987 605814 940043
rect 605870 939987 605938 940043
rect 605994 939987 606062 940043
rect 606118 939987 606172 940043
rect 604122 939919 606172 939987
rect 604122 939863 605070 939919
rect 605126 939863 605194 939919
rect 605250 939863 605318 939919
rect 605374 939863 605442 939919
rect 605498 939863 605566 939919
rect 605622 939863 605690 939919
rect 605746 939863 605814 939919
rect 605870 939863 605938 939919
rect 605994 939863 606062 939919
rect 606118 939863 606172 939919
rect 604122 939720 606172 939863
rect 606828 941655 608878 944000
rect 606828 941599 606908 941655
rect 606964 941599 607032 941655
rect 607088 941599 607156 941655
rect 607212 941599 607280 941655
rect 607336 941599 607404 941655
rect 607460 941599 607528 941655
rect 607584 941599 607652 941655
rect 607708 941599 607776 941655
rect 607832 941599 607900 941655
rect 607956 941599 608024 941655
rect 608080 941599 608148 941655
rect 608204 941599 608272 941655
rect 608328 941599 608396 941655
rect 608452 941599 608520 941655
rect 608576 941599 608644 941655
rect 608700 941599 608768 941655
rect 608824 941599 608878 941655
rect 606828 941531 608878 941599
rect 606828 941475 606908 941531
rect 606964 941475 607032 941531
rect 607088 941475 607156 941531
rect 607212 941475 607280 941531
rect 607336 941475 607404 941531
rect 607460 941475 607528 941531
rect 607584 941475 607652 941531
rect 607708 941475 607776 941531
rect 607832 941475 607900 941531
rect 607956 941475 608024 941531
rect 608080 941475 608148 941531
rect 608204 941475 608272 941531
rect 608328 941475 608396 941531
rect 608452 941475 608520 941531
rect 608576 941475 608644 941531
rect 608700 941475 608768 941531
rect 608824 941475 608878 941531
rect 606828 941407 608878 941475
rect 606828 941351 606908 941407
rect 606964 941351 607032 941407
rect 607088 941351 607156 941407
rect 607212 941351 607280 941407
rect 607336 941351 607404 941407
rect 607460 941351 607528 941407
rect 607584 941351 607652 941407
rect 607708 941351 607776 941407
rect 607832 941351 607900 941407
rect 607956 941351 608024 941407
rect 608080 941351 608148 941407
rect 608204 941351 608272 941407
rect 608328 941351 608396 941407
rect 608452 941351 608520 941407
rect 608576 941351 608644 941407
rect 608700 941351 608768 941407
rect 608824 941351 608878 941407
rect 606828 941283 608878 941351
rect 606828 941227 606908 941283
rect 606964 941227 607032 941283
rect 607088 941227 607156 941283
rect 607212 941227 607280 941283
rect 607336 941227 607404 941283
rect 607460 941227 607528 941283
rect 607584 941227 607652 941283
rect 607708 941227 607776 941283
rect 607832 941227 607900 941283
rect 607956 941227 608024 941283
rect 608080 941227 608148 941283
rect 608204 941227 608272 941283
rect 608328 941227 608396 941283
rect 608452 941227 608520 941283
rect 608576 941227 608644 941283
rect 608700 941227 608768 941283
rect 608824 941227 608878 941283
rect 606828 941159 608878 941227
rect 606828 941103 606908 941159
rect 606964 941103 607032 941159
rect 607088 941103 607156 941159
rect 607212 941103 607280 941159
rect 607336 941103 607404 941159
rect 607460 941103 607528 941159
rect 607584 941103 607652 941159
rect 607708 941103 607776 941159
rect 607832 941103 607900 941159
rect 607956 941103 608024 941159
rect 608080 941103 608148 941159
rect 608204 941103 608272 941159
rect 608328 941103 608396 941159
rect 608452 941103 608520 941159
rect 608576 941103 608644 941159
rect 608700 941103 608768 941159
rect 608824 941103 608878 941159
rect 606828 941035 608878 941103
rect 606828 940979 606908 941035
rect 606964 940979 607032 941035
rect 607088 940979 607156 941035
rect 607212 940979 607280 941035
rect 607336 940979 607404 941035
rect 607460 940979 607528 941035
rect 607584 940979 607652 941035
rect 607708 940979 607776 941035
rect 607832 940979 607900 941035
rect 607956 940979 608024 941035
rect 608080 940979 608148 941035
rect 608204 940979 608272 941035
rect 608328 940979 608396 941035
rect 608452 940979 608520 941035
rect 608576 940979 608644 941035
rect 608700 940979 608768 941035
rect 608824 940979 608878 941035
rect 606828 940911 608878 940979
rect 606828 940855 606908 940911
rect 606964 940855 607032 940911
rect 607088 940855 607156 940911
rect 607212 940855 607280 940911
rect 607336 940855 607404 940911
rect 607460 940855 607528 940911
rect 607584 940855 607652 940911
rect 607708 940855 607776 940911
rect 607832 940855 607900 940911
rect 607956 940855 608024 940911
rect 608080 940855 608148 940911
rect 608204 940855 608272 940911
rect 608328 940855 608396 940911
rect 608452 940855 608520 940911
rect 608576 940855 608644 940911
rect 608700 940855 608768 940911
rect 608824 940855 608878 940911
rect 606828 940787 608878 940855
rect 606828 940731 606908 940787
rect 606964 940731 607032 940787
rect 607088 940731 607156 940787
rect 607212 940731 607280 940787
rect 607336 940731 607404 940787
rect 607460 940731 607528 940787
rect 607584 940731 607652 940787
rect 607708 940731 607776 940787
rect 607832 940731 607900 940787
rect 607956 940731 608024 940787
rect 608080 940731 608148 940787
rect 608204 940731 608272 940787
rect 608328 940731 608396 940787
rect 608452 940731 608520 940787
rect 608576 940731 608644 940787
rect 608700 940731 608768 940787
rect 608824 940731 608878 940787
rect 606828 940663 608878 940731
rect 606828 940607 606908 940663
rect 606964 940607 607032 940663
rect 607088 940607 607156 940663
rect 607212 940607 607280 940663
rect 607336 940607 607404 940663
rect 607460 940607 607528 940663
rect 607584 940607 607652 940663
rect 607708 940607 607776 940663
rect 607832 940607 607900 940663
rect 607956 940607 608024 940663
rect 608080 940607 608148 940663
rect 608204 940607 608272 940663
rect 608328 940607 608396 940663
rect 608452 940607 608520 940663
rect 608576 940607 608644 940663
rect 608700 940607 608768 940663
rect 608824 940607 608878 940663
rect 606828 940539 608878 940607
rect 606828 940483 606908 940539
rect 606964 940483 607032 940539
rect 607088 940483 607156 940539
rect 607212 940483 607280 940539
rect 607336 940483 607404 940539
rect 607460 940483 607528 940539
rect 607584 940483 607652 940539
rect 607708 940483 607776 940539
rect 607832 940483 607900 940539
rect 607956 940483 608024 940539
rect 608080 940483 608148 940539
rect 608204 940483 608272 940539
rect 608328 940483 608396 940539
rect 608452 940483 608520 940539
rect 608576 940483 608644 940539
rect 608700 940483 608768 940539
rect 608824 940483 608878 940539
rect 606828 940415 608878 940483
rect 606828 940359 606908 940415
rect 606964 940359 607032 940415
rect 607088 940359 607156 940415
rect 607212 940359 607280 940415
rect 607336 940359 607404 940415
rect 607460 940359 607528 940415
rect 607584 940359 607652 940415
rect 607708 940359 607776 940415
rect 607832 940359 607900 940415
rect 607956 940359 608024 940415
rect 608080 940359 608148 940415
rect 608204 940359 608272 940415
rect 608328 940359 608396 940415
rect 608452 940359 608520 940415
rect 608576 940359 608644 940415
rect 608700 940359 608768 940415
rect 608824 940359 608878 940415
rect 606828 940291 608878 940359
rect 606828 940235 606908 940291
rect 606964 940235 607032 940291
rect 607088 940235 607156 940291
rect 607212 940235 607280 940291
rect 607336 940235 607404 940291
rect 607460 940235 607528 940291
rect 607584 940235 607652 940291
rect 607708 940235 607776 940291
rect 607832 940235 607900 940291
rect 607956 940235 608024 940291
rect 608080 940235 608148 940291
rect 608204 940235 608272 940291
rect 608328 940235 608396 940291
rect 608452 940235 608520 940291
rect 608576 940235 608644 940291
rect 608700 940235 608768 940291
rect 608824 940235 608878 940291
rect 606828 940167 608878 940235
rect 606828 940111 606908 940167
rect 606964 940111 607032 940167
rect 607088 940111 607156 940167
rect 607212 940111 607280 940167
rect 607336 940111 607404 940167
rect 607460 940111 607528 940167
rect 607584 940111 607652 940167
rect 607708 940111 607776 940167
rect 607832 940111 607900 940167
rect 607956 940111 608024 940167
rect 608080 940111 608148 940167
rect 608204 940111 608272 940167
rect 608328 940111 608396 940167
rect 608452 940111 608520 940167
rect 608576 940111 608644 940167
rect 608700 940111 608768 940167
rect 608824 940111 608878 940167
rect 606828 940043 608878 940111
rect 606828 939987 606908 940043
rect 606964 939987 607032 940043
rect 607088 939987 607156 940043
rect 607212 939987 607280 940043
rect 607336 939987 607404 940043
rect 607460 939987 607528 940043
rect 607584 939987 607652 940043
rect 607708 939987 607776 940043
rect 607832 939987 607900 940043
rect 607956 939987 608024 940043
rect 608080 939987 608148 940043
rect 608204 939987 608272 940043
rect 608328 939987 608396 940043
rect 608452 939987 608520 940043
rect 608576 939987 608644 940043
rect 608700 939987 608768 940043
rect 608824 939987 608878 940043
rect 606828 939919 608878 939987
rect 606828 939863 606908 939919
rect 606964 939863 607032 939919
rect 607088 939863 607156 939919
rect 607212 939863 607280 939919
rect 607336 939863 607404 939919
rect 607460 939863 607528 939919
rect 607584 939863 607652 939919
rect 607708 939863 607776 939919
rect 607832 939863 607900 939919
rect 607956 939863 608024 939919
rect 608080 939863 608148 939919
rect 608204 939863 608272 939919
rect 608328 939863 608396 939919
rect 608452 939863 608520 939919
rect 608576 939863 608644 939919
rect 608700 939863 608768 939919
rect 608824 939863 608878 939919
rect 606828 939720 608878 939863
rect 609198 941655 611248 944000
rect 609198 941599 609278 941655
rect 609334 941599 609402 941655
rect 609458 941599 609526 941655
rect 609582 941599 609650 941655
rect 609706 941599 609774 941655
rect 609830 941599 609898 941655
rect 609954 941599 610022 941655
rect 610078 941599 610146 941655
rect 610202 941599 610270 941655
rect 610326 941599 610394 941655
rect 610450 941599 610518 941655
rect 610574 941599 610642 941655
rect 610698 941599 610766 941655
rect 610822 941599 610890 941655
rect 610946 941599 611014 941655
rect 611070 941599 611138 941655
rect 611194 941599 611248 941655
rect 609198 941531 611248 941599
rect 609198 941475 609278 941531
rect 609334 941475 609402 941531
rect 609458 941475 609526 941531
rect 609582 941475 609650 941531
rect 609706 941475 609774 941531
rect 609830 941475 609898 941531
rect 609954 941475 610022 941531
rect 610078 941475 610146 941531
rect 610202 941475 610270 941531
rect 610326 941475 610394 941531
rect 610450 941475 610518 941531
rect 610574 941475 610642 941531
rect 610698 941475 610766 941531
rect 610822 941475 610890 941531
rect 610946 941475 611014 941531
rect 611070 941475 611138 941531
rect 611194 941475 611248 941531
rect 609198 941407 611248 941475
rect 609198 941351 609278 941407
rect 609334 941351 609402 941407
rect 609458 941351 609526 941407
rect 609582 941351 609650 941407
rect 609706 941351 609774 941407
rect 609830 941351 609898 941407
rect 609954 941351 610022 941407
rect 610078 941351 610146 941407
rect 610202 941351 610270 941407
rect 610326 941351 610394 941407
rect 610450 941351 610518 941407
rect 610574 941351 610642 941407
rect 610698 941351 610766 941407
rect 610822 941351 610890 941407
rect 610946 941351 611014 941407
rect 611070 941351 611138 941407
rect 611194 941351 611248 941407
rect 609198 941283 611248 941351
rect 609198 941227 609278 941283
rect 609334 941227 609402 941283
rect 609458 941227 609526 941283
rect 609582 941227 609650 941283
rect 609706 941227 609774 941283
rect 609830 941227 609898 941283
rect 609954 941227 610022 941283
rect 610078 941227 610146 941283
rect 610202 941227 610270 941283
rect 610326 941227 610394 941283
rect 610450 941227 610518 941283
rect 610574 941227 610642 941283
rect 610698 941227 610766 941283
rect 610822 941227 610890 941283
rect 610946 941227 611014 941283
rect 611070 941227 611138 941283
rect 611194 941227 611248 941283
rect 609198 941159 611248 941227
rect 609198 941103 609278 941159
rect 609334 941103 609402 941159
rect 609458 941103 609526 941159
rect 609582 941103 609650 941159
rect 609706 941103 609774 941159
rect 609830 941103 609898 941159
rect 609954 941103 610022 941159
rect 610078 941103 610146 941159
rect 610202 941103 610270 941159
rect 610326 941103 610394 941159
rect 610450 941103 610518 941159
rect 610574 941103 610642 941159
rect 610698 941103 610766 941159
rect 610822 941103 610890 941159
rect 610946 941103 611014 941159
rect 611070 941103 611138 941159
rect 611194 941103 611248 941159
rect 609198 941035 611248 941103
rect 609198 940979 609278 941035
rect 609334 940979 609402 941035
rect 609458 940979 609526 941035
rect 609582 940979 609650 941035
rect 609706 940979 609774 941035
rect 609830 940979 609898 941035
rect 609954 940979 610022 941035
rect 610078 940979 610146 941035
rect 610202 940979 610270 941035
rect 610326 940979 610394 941035
rect 610450 940979 610518 941035
rect 610574 940979 610642 941035
rect 610698 940979 610766 941035
rect 610822 940979 610890 941035
rect 610946 940979 611014 941035
rect 611070 940979 611138 941035
rect 611194 940979 611248 941035
rect 609198 940911 611248 940979
rect 609198 940855 609278 940911
rect 609334 940855 609402 940911
rect 609458 940855 609526 940911
rect 609582 940855 609650 940911
rect 609706 940855 609774 940911
rect 609830 940855 609898 940911
rect 609954 940855 610022 940911
rect 610078 940855 610146 940911
rect 610202 940855 610270 940911
rect 610326 940855 610394 940911
rect 610450 940855 610518 940911
rect 610574 940855 610642 940911
rect 610698 940855 610766 940911
rect 610822 940855 610890 940911
rect 610946 940855 611014 940911
rect 611070 940855 611138 940911
rect 611194 940855 611248 940911
rect 609198 940787 611248 940855
rect 609198 940731 609278 940787
rect 609334 940731 609402 940787
rect 609458 940731 609526 940787
rect 609582 940731 609650 940787
rect 609706 940731 609774 940787
rect 609830 940731 609898 940787
rect 609954 940731 610022 940787
rect 610078 940731 610146 940787
rect 610202 940731 610270 940787
rect 610326 940731 610394 940787
rect 610450 940731 610518 940787
rect 610574 940731 610642 940787
rect 610698 940731 610766 940787
rect 610822 940731 610890 940787
rect 610946 940731 611014 940787
rect 611070 940731 611138 940787
rect 611194 940731 611248 940787
rect 609198 940663 611248 940731
rect 609198 940607 609278 940663
rect 609334 940607 609402 940663
rect 609458 940607 609526 940663
rect 609582 940607 609650 940663
rect 609706 940607 609774 940663
rect 609830 940607 609898 940663
rect 609954 940607 610022 940663
rect 610078 940607 610146 940663
rect 610202 940607 610270 940663
rect 610326 940607 610394 940663
rect 610450 940607 610518 940663
rect 610574 940607 610642 940663
rect 610698 940607 610766 940663
rect 610822 940607 610890 940663
rect 610946 940607 611014 940663
rect 611070 940607 611138 940663
rect 611194 940607 611248 940663
rect 609198 940539 611248 940607
rect 609198 940483 609278 940539
rect 609334 940483 609402 940539
rect 609458 940483 609526 940539
rect 609582 940483 609650 940539
rect 609706 940483 609774 940539
rect 609830 940483 609898 940539
rect 609954 940483 610022 940539
rect 610078 940483 610146 940539
rect 610202 940483 610270 940539
rect 610326 940483 610394 940539
rect 610450 940483 610518 940539
rect 610574 940483 610642 940539
rect 610698 940483 610766 940539
rect 610822 940483 610890 940539
rect 610946 940483 611014 940539
rect 611070 940483 611138 940539
rect 611194 940483 611248 940539
rect 609198 940415 611248 940483
rect 609198 940359 609278 940415
rect 609334 940359 609402 940415
rect 609458 940359 609526 940415
rect 609582 940359 609650 940415
rect 609706 940359 609774 940415
rect 609830 940359 609898 940415
rect 609954 940359 610022 940415
rect 610078 940359 610146 940415
rect 610202 940359 610270 940415
rect 610326 940359 610394 940415
rect 610450 940359 610518 940415
rect 610574 940359 610642 940415
rect 610698 940359 610766 940415
rect 610822 940359 610890 940415
rect 610946 940359 611014 940415
rect 611070 940359 611138 940415
rect 611194 940359 611248 940415
rect 609198 940291 611248 940359
rect 609198 940235 609278 940291
rect 609334 940235 609402 940291
rect 609458 940235 609526 940291
rect 609582 940235 609650 940291
rect 609706 940235 609774 940291
rect 609830 940235 609898 940291
rect 609954 940235 610022 940291
rect 610078 940235 610146 940291
rect 610202 940235 610270 940291
rect 610326 940235 610394 940291
rect 610450 940235 610518 940291
rect 610574 940235 610642 940291
rect 610698 940235 610766 940291
rect 610822 940235 610890 940291
rect 610946 940235 611014 940291
rect 611070 940235 611138 940291
rect 611194 940235 611248 940291
rect 609198 940167 611248 940235
rect 609198 940111 609278 940167
rect 609334 940111 609402 940167
rect 609458 940111 609526 940167
rect 609582 940111 609650 940167
rect 609706 940111 609774 940167
rect 609830 940111 609898 940167
rect 609954 940111 610022 940167
rect 610078 940111 610146 940167
rect 610202 940111 610270 940167
rect 610326 940111 610394 940167
rect 610450 940111 610518 940167
rect 610574 940111 610642 940167
rect 610698 940111 610766 940167
rect 610822 940111 610890 940167
rect 610946 940111 611014 940167
rect 611070 940111 611138 940167
rect 611194 940111 611248 940167
rect 609198 940043 611248 940111
rect 609198 939987 609278 940043
rect 609334 939987 609402 940043
rect 609458 939987 609526 940043
rect 609582 939987 609650 940043
rect 609706 939987 609774 940043
rect 609830 939987 609898 940043
rect 609954 939987 610022 940043
rect 610078 939987 610146 940043
rect 610202 939987 610270 940043
rect 610326 939987 610394 940043
rect 610450 939987 610518 940043
rect 610574 939987 610642 940043
rect 610698 939987 610766 940043
rect 610822 939987 610890 940043
rect 610946 939987 611014 940043
rect 611070 939987 611138 940043
rect 611194 939987 611248 940043
rect 609198 939919 611248 939987
rect 609198 939863 609278 939919
rect 609334 939863 609402 939919
rect 609458 939863 609526 939919
rect 609582 939863 609650 939919
rect 609706 939863 609774 939919
rect 609830 939863 609898 939919
rect 609954 939863 610022 939919
rect 610078 939863 610146 939919
rect 610202 939863 610270 939919
rect 610326 939863 610394 939919
rect 610450 939863 610518 939919
rect 610574 939863 610642 939919
rect 610698 939863 610766 939919
rect 610822 939863 610890 939919
rect 610946 939863 611014 939919
rect 611070 939863 611138 939919
rect 611194 939863 611248 939919
rect 609198 939720 611248 939863
rect 611828 941655 613728 944000
rect 611828 941599 611882 941655
rect 611938 941599 612006 941655
rect 612062 941599 612130 941655
rect 612186 941599 612254 941655
rect 612310 941599 612378 941655
rect 612434 941599 612502 941655
rect 612558 941599 612626 941655
rect 612682 941599 612750 941655
rect 612806 941599 612874 941655
rect 612930 941599 612998 941655
rect 613054 941599 613122 941655
rect 613178 941599 613246 941655
rect 613302 941599 613370 941655
rect 613426 941599 613494 941655
rect 613550 941599 613618 941655
rect 613674 941599 613728 941655
rect 611828 941531 613728 941599
rect 611828 941475 611882 941531
rect 611938 941475 612006 941531
rect 612062 941475 612130 941531
rect 612186 941475 612254 941531
rect 612310 941475 612378 941531
rect 612434 941475 612502 941531
rect 612558 941475 612626 941531
rect 612682 941475 612750 941531
rect 612806 941475 612874 941531
rect 612930 941475 612998 941531
rect 613054 941475 613122 941531
rect 613178 941475 613246 941531
rect 613302 941475 613370 941531
rect 613426 941475 613494 941531
rect 613550 941475 613618 941531
rect 613674 941475 613728 941531
rect 611828 941407 613728 941475
rect 611828 941351 611882 941407
rect 611938 941351 612006 941407
rect 612062 941351 612130 941407
rect 612186 941351 612254 941407
rect 612310 941351 612378 941407
rect 612434 941351 612502 941407
rect 612558 941351 612626 941407
rect 612682 941351 612750 941407
rect 612806 941351 612874 941407
rect 612930 941351 612998 941407
rect 613054 941351 613122 941407
rect 613178 941351 613246 941407
rect 613302 941351 613370 941407
rect 613426 941351 613494 941407
rect 613550 941351 613618 941407
rect 613674 941351 613728 941407
rect 611828 941283 613728 941351
rect 611828 941227 611882 941283
rect 611938 941227 612006 941283
rect 612062 941227 612130 941283
rect 612186 941227 612254 941283
rect 612310 941227 612378 941283
rect 612434 941227 612502 941283
rect 612558 941227 612626 941283
rect 612682 941227 612750 941283
rect 612806 941227 612874 941283
rect 612930 941227 612998 941283
rect 613054 941227 613122 941283
rect 613178 941227 613246 941283
rect 613302 941227 613370 941283
rect 613426 941227 613494 941283
rect 613550 941227 613618 941283
rect 613674 941227 613728 941283
rect 611828 941159 613728 941227
rect 611828 941103 611882 941159
rect 611938 941103 612006 941159
rect 612062 941103 612130 941159
rect 612186 941103 612254 941159
rect 612310 941103 612378 941159
rect 612434 941103 612502 941159
rect 612558 941103 612626 941159
rect 612682 941103 612750 941159
rect 612806 941103 612874 941159
rect 612930 941103 612998 941159
rect 613054 941103 613122 941159
rect 613178 941103 613246 941159
rect 613302 941103 613370 941159
rect 613426 941103 613494 941159
rect 613550 941103 613618 941159
rect 613674 941103 613728 941159
rect 611828 941035 613728 941103
rect 611828 940979 611882 941035
rect 611938 940979 612006 941035
rect 612062 940979 612130 941035
rect 612186 940979 612254 941035
rect 612310 940979 612378 941035
rect 612434 940979 612502 941035
rect 612558 940979 612626 941035
rect 612682 940979 612750 941035
rect 612806 940979 612874 941035
rect 612930 940979 612998 941035
rect 613054 940979 613122 941035
rect 613178 940979 613246 941035
rect 613302 940979 613370 941035
rect 613426 940979 613494 941035
rect 613550 940979 613618 941035
rect 613674 940979 613728 941035
rect 611828 940911 613728 940979
rect 611828 940855 611882 940911
rect 611938 940855 612006 940911
rect 612062 940855 612130 940911
rect 612186 940855 612254 940911
rect 612310 940855 612378 940911
rect 612434 940855 612502 940911
rect 612558 940855 612626 940911
rect 612682 940855 612750 940911
rect 612806 940855 612874 940911
rect 612930 940855 612998 940911
rect 613054 940855 613122 940911
rect 613178 940855 613246 940911
rect 613302 940855 613370 940911
rect 613426 940855 613494 940911
rect 613550 940855 613618 940911
rect 613674 940855 613728 940911
rect 611828 940787 613728 940855
rect 611828 940731 611882 940787
rect 611938 940731 612006 940787
rect 612062 940731 612130 940787
rect 612186 940731 612254 940787
rect 612310 940731 612378 940787
rect 612434 940731 612502 940787
rect 612558 940731 612626 940787
rect 612682 940731 612750 940787
rect 612806 940731 612874 940787
rect 612930 940731 612998 940787
rect 613054 940731 613122 940787
rect 613178 940731 613246 940787
rect 613302 940731 613370 940787
rect 613426 940731 613494 940787
rect 613550 940731 613618 940787
rect 613674 940731 613728 940787
rect 611828 940663 613728 940731
rect 611828 940607 611882 940663
rect 611938 940607 612006 940663
rect 612062 940607 612130 940663
rect 612186 940607 612254 940663
rect 612310 940607 612378 940663
rect 612434 940607 612502 940663
rect 612558 940607 612626 940663
rect 612682 940607 612750 940663
rect 612806 940607 612874 940663
rect 612930 940607 612998 940663
rect 613054 940607 613122 940663
rect 613178 940607 613246 940663
rect 613302 940607 613370 940663
rect 613426 940607 613494 940663
rect 613550 940607 613618 940663
rect 613674 940607 613728 940663
rect 611828 940539 613728 940607
rect 611828 940483 611882 940539
rect 611938 940483 612006 940539
rect 612062 940483 612130 940539
rect 612186 940483 612254 940539
rect 612310 940483 612378 940539
rect 612434 940483 612502 940539
rect 612558 940483 612626 940539
rect 612682 940483 612750 940539
rect 612806 940483 612874 940539
rect 612930 940483 612998 940539
rect 613054 940483 613122 940539
rect 613178 940483 613246 940539
rect 613302 940483 613370 940539
rect 613426 940483 613494 940539
rect 613550 940483 613618 940539
rect 613674 940483 613728 940539
rect 611828 940415 613728 940483
rect 611828 940359 611882 940415
rect 611938 940359 612006 940415
rect 612062 940359 612130 940415
rect 612186 940359 612254 940415
rect 612310 940359 612378 940415
rect 612434 940359 612502 940415
rect 612558 940359 612626 940415
rect 612682 940359 612750 940415
rect 612806 940359 612874 940415
rect 612930 940359 612998 940415
rect 613054 940359 613122 940415
rect 613178 940359 613246 940415
rect 613302 940359 613370 940415
rect 613426 940359 613494 940415
rect 613550 940359 613618 940415
rect 613674 940359 613728 940415
rect 611828 940291 613728 940359
rect 611828 940235 611882 940291
rect 611938 940235 612006 940291
rect 612062 940235 612130 940291
rect 612186 940235 612254 940291
rect 612310 940235 612378 940291
rect 612434 940235 612502 940291
rect 612558 940235 612626 940291
rect 612682 940235 612750 940291
rect 612806 940235 612874 940291
rect 612930 940235 612998 940291
rect 613054 940235 613122 940291
rect 613178 940235 613246 940291
rect 613302 940235 613370 940291
rect 613426 940235 613494 940291
rect 613550 940235 613618 940291
rect 613674 940235 613728 940291
rect 611828 940167 613728 940235
rect 611828 940111 611882 940167
rect 611938 940111 612006 940167
rect 612062 940111 612130 940167
rect 612186 940111 612254 940167
rect 612310 940111 612378 940167
rect 612434 940111 612502 940167
rect 612558 940111 612626 940167
rect 612682 940111 612750 940167
rect 612806 940111 612874 940167
rect 612930 940111 612998 940167
rect 613054 940111 613122 940167
rect 613178 940111 613246 940167
rect 613302 940111 613370 940167
rect 613426 940111 613494 940167
rect 613550 940111 613618 940167
rect 613674 940111 613728 940167
rect 611828 940043 613728 940111
rect 611828 939987 611882 940043
rect 611938 939987 612006 940043
rect 612062 939987 612130 940043
rect 612186 939987 612254 940043
rect 612310 939987 612378 940043
rect 612434 939987 612502 940043
rect 612558 939987 612626 940043
rect 612682 939987 612750 940043
rect 612806 939987 612874 940043
rect 612930 939987 612998 940043
rect 613054 939987 613122 940043
rect 613178 939987 613246 940043
rect 613302 939987 613370 940043
rect 613426 939987 613494 940043
rect 613550 939987 613618 940043
rect 613674 939987 613728 940043
rect 611828 939919 613728 939987
rect 611828 939863 611882 939919
rect 611938 939863 612006 939919
rect 612062 939863 612130 939919
rect 612186 939863 612254 939919
rect 612310 939863 612378 939919
rect 612434 939863 612502 939919
rect 612558 939863 612626 939919
rect 612682 939863 612750 939919
rect 612806 939863 612874 939919
rect 612930 939863 612998 939919
rect 613054 939863 613122 939919
rect 613178 939863 613246 939919
rect 613302 939863 613370 939919
rect 613426 939863 613494 939919
rect 613550 939863 613618 939919
rect 613674 939863 613728 939919
rect 611828 939720 613728 939863
rect 70000 878661 70488 878728
rect 70000 878605 70047 878661
rect 70103 878605 70171 878661
rect 70227 878605 70295 878661
rect 70351 878605 70419 878661
rect 70475 878605 70488 878661
rect 70000 878537 70488 878605
rect 70000 878481 70047 878537
rect 70103 878481 70171 878537
rect 70227 878481 70295 878537
rect 70351 878481 70419 878537
rect 70475 878481 70488 878537
rect 70000 878413 70488 878481
rect 70000 878357 70047 878413
rect 70103 878357 70171 878413
rect 70227 878357 70295 878413
rect 70351 878357 70419 878413
rect 70475 878357 70488 878413
rect 70000 878289 70488 878357
rect 70000 878233 70047 878289
rect 70103 878233 70171 878289
rect 70227 878233 70295 878289
rect 70351 878233 70419 878289
rect 70475 878233 70488 878289
rect 70000 878165 70488 878233
rect 70000 878109 70047 878165
rect 70103 878109 70171 878165
rect 70227 878109 70295 878165
rect 70351 878109 70419 878165
rect 70475 878109 70488 878165
rect 70000 878041 70488 878109
rect 70000 877985 70047 878041
rect 70103 877985 70171 878041
rect 70227 877985 70295 878041
rect 70351 877985 70419 878041
rect 70475 877985 70488 878041
rect 70000 877917 70488 877985
rect 70000 877861 70047 877917
rect 70103 877861 70171 877917
rect 70227 877861 70295 877917
rect 70351 877861 70419 877917
rect 70475 877861 70488 877917
rect 70000 877793 70488 877861
rect 70000 877737 70047 877793
rect 70103 877737 70171 877793
rect 70227 877737 70295 877793
rect 70351 877737 70419 877793
rect 70475 877737 70488 877793
rect 70000 877669 70488 877737
rect 70000 877613 70047 877669
rect 70103 877613 70171 877669
rect 70227 877613 70295 877669
rect 70351 877613 70419 877669
rect 70475 877613 70488 877669
rect 70000 877545 70488 877613
rect 70000 877489 70047 877545
rect 70103 877489 70171 877545
rect 70227 877489 70295 877545
rect 70351 877489 70419 877545
rect 70475 877489 70488 877545
rect 70000 877421 70488 877489
rect 70000 877365 70047 877421
rect 70103 877365 70171 877421
rect 70227 877365 70295 877421
rect 70351 877365 70419 877421
rect 70475 877365 70488 877421
rect 70000 877297 70488 877365
rect 70000 877241 70047 877297
rect 70103 877241 70171 877297
rect 70227 877241 70295 877297
rect 70351 877241 70419 877297
rect 70475 877241 70488 877297
rect 70000 877173 70488 877241
rect 70000 877117 70047 877173
rect 70103 877117 70171 877173
rect 70227 877117 70295 877173
rect 70351 877117 70419 877173
rect 70475 877117 70488 877173
rect 70000 877049 70488 877117
rect 70000 876993 70047 877049
rect 70103 876993 70171 877049
rect 70227 876993 70295 877049
rect 70351 876993 70419 877049
rect 70475 876993 70488 877049
rect 70000 876925 70488 876993
rect 70000 876869 70047 876925
rect 70103 876869 70171 876925
rect 70227 876869 70295 876925
rect 70351 876869 70419 876925
rect 70475 876869 70488 876925
rect 70000 876828 70488 876869
rect 705512 877687 706000 877728
rect 705512 877631 705525 877687
rect 705581 877631 705649 877687
rect 705705 877631 705773 877687
rect 705829 877631 705897 877687
rect 705953 877631 706000 877687
rect 705512 877563 706000 877631
rect 705512 877507 705525 877563
rect 705581 877507 705649 877563
rect 705705 877507 705773 877563
rect 705829 877507 705897 877563
rect 705953 877507 706000 877563
rect 705512 877439 706000 877507
rect 705512 877383 705525 877439
rect 705581 877383 705649 877439
rect 705705 877383 705773 877439
rect 705829 877383 705897 877439
rect 705953 877383 706000 877439
rect 705512 877315 706000 877383
rect 705512 877259 705525 877315
rect 705581 877259 705649 877315
rect 705705 877259 705773 877315
rect 705829 877259 705897 877315
rect 705953 877259 706000 877315
rect 705512 877191 706000 877259
rect 705512 877135 705525 877191
rect 705581 877135 705649 877191
rect 705705 877135 705773 877191
rect 705829 877135 705897 877191
rect 705953 877135 706000 877191
rect 705512 877067 706000 877135
rect 705512 877011 705525 877067
rect 705581 877011 705649 877067
rect 705705 877011 705773 877067
rect 705829 877011 705897 877067
rect 705953 877011 706000 877067
rect 705512 876943 706000 877011
rect 705512 876887 705525 876943
rect 705581 876887 705649 876943
rect 705705 876887 705773 876943
rect 705829 876887 705897 876943
rect 705953 876887 706000 876943
rect 705512 876819 706000 876887
rect 705512 876763 705525 876819
rect 705581 876763 705649 876819
rect 705705 876763 705773 876819
rect 705829 876763 705897 876819
rect 705953 876763 706000 876819
rect 705512 876695 706000 876763
rect 705512 876639 705525 876695
rect 705581 876639 705649 876695
rect 705705 876639 705773 876695
rect 705829 876639 705897 876695
rect 705953 876639 706000 876695
rect 705512 876571 706000 876639
rect 705512 876515 705525 876571
rect 705581 876515 705649 876571
rect 705705 876515 705773 876571
rect 705829 876515 705897 876571
rect 705953 876515 706000 876571
rect 705512 876447 706000 876515
rect 705512 876391 705525 876447
rect 705581 876391 705649 876447
rect 705705 876391 705773 876447
rect 705829 876391 705897 876447
rect 705953 876391 706000 876447
rect 705512 876323 706000 876391
rect 705512 876267 705525 876323
rect 705581 876267 705649 876323
rect 705705 876267 705773 876323
rect 705829 876267 705897 876323
rect 705953 876267 706000 876323
rect 70000 876181 70488 876248
rect 70000 876125 70047 876181
rect 70103 876125 70171 876181
rect 70227 876125 70295 876181
rect 70351 876125 70419 876181
rect 70475 876125 70488 876181
rect 70000 876057 70488 876125
rect 70000 876001 70047 876057
rect 70103 876001 70171 876057
rect 70227 876001 70295 876057
rect 70351 876001 70419 876057
rect 70475 876001 70488 876057
rect 70000 875933 70488 876001
rect 70000 875877 70047 875933
rect 70103 875877 70171 875933
rect 70227 875877 70295 875933
rect 70351 875877 70419 875933
rect 70475 875877 70488 875933
rect 70000 875809 70488 875877
rect 705512 876199 706000 876267
rect 705512 876143 705525 876199
rect 705581 876143 705649 876199
rect 705705 876143 705773 876199
rect 705829 876143 705897 876199
rect 705953 876143 706000 876199
rect 705512 876075 706000 876143
rect 705512 876019 705525 876075
rect 705581 876019 705649 876075
rect 705705 876019 705773 876075
rect 705829 876019 705897 876075
rect 705953 876019 706000 876075
rect 705512 875951 706000 876019
rect 705512 875895 705525 875951
rect 705581 875895 705649 875951
rect 705705 875895 705773 875951
rect 705829 875895 705897 875951
rect 705953 875895 706000 875951
rect 705512 875828 706000 875895
rect 70000 875753 70047 875809
rect 70103 875753 70171 875809
rect 70227 875753 70295 875809
rect 70351 875753 70419 875809
rect 70475 875753 70488 875809
rect 70000 875685 70488 875753
rect 70000 875629 70047 875685
rect 70103 875629 70171 875685
rect 70227 875629 70295 875685
rect 70351 875629 70419 875685
rect 70475 875629 70488 875685
rect 70000 875561 70488 875629
rect 70000 875505 70047 875561
rect 70103 875505 70171 875561
rect 70227 875505 70295 875561
rect 70351 875505 70419 875561
rect 70475 875505 70488 875561
rect 70000 875437 70488 875505
rect 70000 875381 70047 875437
rect 70103 875381 70171 875437
rect 70227 875381 70295 875437
rect 70351 875381 70419 875437
rect 70475 875381 70488 875437
rect 70000 875313 70488 875381
rect 70000 875257 70047 875313
rect 70103 875257 70171 875313
rect 70227 875257 70295 875313
rect 70351 875257 70419 875313
rect 70475 875257 70488 875313
rect 70000 875189 70488 875257
rect 70000 875133 70047 875189
rect 70103 875133 70171 875189
rect 70227 875133 70295 875189
rect 70351 875133 70419 875189
rect 70475 875133 70488 875189
rect 70000 875065 70488 875133
rect 70000 875009 70047 875065
rect 70103 875009 70171 875065
rect 70227 875009 70295 875065
rect 70351 875009 70419 875065
rect 70475 875009 70488 875065
rect 70000 874941 70488 875009
rect 70000 874885 70047 874941
rect 70103 874885 70171 874941
rect 70227 874885 70295 874941
rect 70351 874885 70419 874941
rect 70475 874885 70488 874941
rect 70000 874817 70488 874885
rect 70000 874761 70047 874817
rect 70103 874761 70171 874817
rect 70227 874761 70295 874817
rect 70351 874761 70419 874817
rect 70475 874761 70488 874817
rect 70000 874693 70488 874761
rect 70000 874637 70047 874693
rect 70103 874637 70171 874693
rect 70227 874637 70295 874693
rect 70351 874637 70419 874693
rect 70475 874637 70488 874693
rect 70000 874569 70488 874637
rect 70000 874513 70047 874569
rect 70103 874513 70171 874569
rect 70227 874513 70295 874569
rect 70351 874513 70419 874569
rect 70475 874513 70488 874569
rect 70000 874445 70488 874513
rect 70000 874389 70047 874445
rect 70103 874389 70171 874445
rect 70227 874389 70295 874445
rect 70351 874389 70419 874445
rect 70475 874389 70488 874445
rect 70000 874321 70488 874389
rect 70000 874265 70047 874321
rect 70103 874265 70171 874321
rect 70227 874265 70295 874321
rect 70351 874265 70419 874321
rect 70475 874265 70488 874321
rect 70000 874198 70488 874265
rect 705512 875181 706000 875248
rect 705512 875125 705525 875181
rect 705581 875125 705649 875181
rect 705705 875125 705773 875181
rect 705829 875125 705897 875181
rect 705953 875125 706000 875181
rect 705512 875057 706000 875125
rect 705512 875001 705525 875057
rect 705581 875001 705649 875057
rect 705705 875001 705773 875057
rect 705829 875001 705897 875057
rect 705953 875001 706000 875057
rect 705512 874933 706000 875001
rect 705512 874877 705525 874933
rect 705581 874877 705649 874933
rect 705705 874877 705773 874933
rect 705829 874877 705897 874933
rect 705953 874877 706000 874933
rect 705512 874809 706000 874877
rect 705512 874753 705525 874809
rect 705581 874753 705649 874809
rect 705705 874753 705773 874809
rect 705829 874753 705897 874809
rect 705953 874753 706000 874809
rect 705512 874685 706000 874753
rect 705512 874629 705525 874685
rect 705581 874629 705649 874685
rect 705705 874629 705773 874685
rect 705829 874629 705897 874685
rect 705953 874629 706000 874685
rect 705512 874561 706000 874629
rect 705512 874505 705525 874561
rect 705581 874505 705649 874561
rect 705705 874505 705773 874561
rect 705829 874505 705897 874561
rect 705953 874505 706000 874561
rect 705512 874437 706000 874505
rect 705512 874381 705525 874437
rect 705581 874381 705649 874437
rect 705705 874381 705773 874437
rect 705829 874381 705897 874437
rect 705953 874381 706000 874437
rect 705512 874313 706000 874381
rect 705512 874257 705525 874313
rect 705581 874257 705649 874313
rect 705705 874257 705773 874313
rect 705829 874257 705897 874313
rect 705953 874257 706000 874313
rect 705512 874189 706000 874257
rect 705512 874133 705525 874189
rect 705581 874133 705649 874189
rect 705705 874133 705773 874189
rect 705829 874133 705897 874189
rect 705953 874133 706000 874189
rect 705512 874065 706000 874133
rect 705512 874009 705525 874065
rect 705581 874009 705649 874065
rect 705705 874009 705773 874065
rect 705829 874009 705897 874065
rect 705953 874009 706000 874065
rect 705512 873941 706000 874009
rect 705512 873885 705525 873941
rect 705581 873885 705649 873941
rect 705705 873885 705773 873941
rect 705829 873885 705897 873941
rect 705953 873885 706000 873941
rect 70000 873811 70488 873878
rect 70000 873755 70047 873811
rect 70103 873755 70171 873811
rect 70227 873755 70295 873811
rect 70351 873755 70419 873811
rect 70475 873755 70488 873811
rect 70000 873687 70488 873755
rect 70000 873631 70047 873687
rect 70103 873631 70171 873687
rect 70227 873631 70295 873687
rect 70351 873631 70419 873687
rect 70475 873631 70488 873687
rect 70000 873563 70488 873631
rect 70000 873507 70047 873563
rect 70103 873507 70171 873563
rect 70227 873507 70295 873563
rect 70351 873507 70419 873563
rect 70475 873507 70488 873563
rect 70000 873439 70488 873507
rect 70000 873383 70047 873439
rect 70103 873383 70171 873439
rect 70227 873383 70295 873439
rect 70351 873383 70419 873439
rect 70475 873383 70488 873439
rect 70000 873315 70488 873383
rect 70000 873259 70047 873315
rect 70103 873259 70171 873315
rect 70227 873259 70295 873315
rect 70351 873259 70419 873315
rect 70475 873259 70488 873315
rect 70000 873191 70488 873259
rect 705512 873817 706000 873885
rect 705512 873761 705525 873817
rect 705581 873761 705649 873817
rect 705705 873761 705773 873817
rect 705829 873761 705897 873817
rect 705953 873761 706000 873817
rect 705512 873693 706000 873761
rect 705512 873637 705525 873693
rect 705581 873637 705649 873693
rect 705705 873637 705773 873693
rect 705829 873637 705897 873693
rect 705953 873637 706000 873693
rect 705512 873569 706000 873637
rect 705512 873513 705525 873569
rect 705581 873513 705649 873569
rect 705705 873513 705773 873569
rect 705829 873513 705897 873569
rect 705953 873513 706000 873569
rect 705512 873445 706000 873513
rect 705512 873389 705525 873445
rect 705581 873389 705649 873445
rect 705705 873389 705773 873445
rect 705829 873389 705897 873445
rect 705953 873389 706000 873445
rect 705512 873321 706000 873389
rect 705512 873265 705525 873321
rect 705581 873265 705649 873321
rect 705705 873265 705773 873321
rect 705829 873265 705897 873321
rect 705953 873265 706000 873321
rect 705512 873198 706000 873265
rect 70000 873135 70047 873191
rect 70103 873135 70171 873191
rect 70227 873135 70295 873191
rect 70351 873135 70419 873191
rect 70475 873135 70488 873191
rect 70000 873067 70488 873135
rect 70000 873011 70047 873067
rect 70103 873011 70171 873067
rect 70227 873011 70295 873067
rect 70351 873011 70419 873067
rect 70475 873011 70488 873067
rect 70000 872943 70488 873011
rect 70000 872887 70047 872943
rect 70103 872887 70171 872943
rect 70227 872887 70295 872943
rect 70351 872887 70419 872943
rect 70475 872887 70488 872943
rect 70000 872819 70488 872887
rect 70000 872763 70047 872819
rect 70103 872763 70171 872819
rect 70227 872763 70295 872819
rect 70351 872763 70419 872819
rect 70475 872763 70488 872819
rect 70000 872695 70488 872763
rect 70000 872639 70047 872695
rect 70103 872639 70171 872695
rect 70227 872639 70295 872695
rect 70351 872639 70419 872695
rect 70475 872639 70488 872695
rect 70000 872571 70488 872639
rect 70000 872515 70047 872571
rect 70103 872515 70171 872571
rect 70227 872515 70295 872571
rect 70351 872515 70419 872571
rect 70475 872515 70488 872571
rect 70000 872447 70488 872515
rect 70000 872391 70047 872447
rect 70103 872391 70171 872447
rect 70227 872391 70295 872447
rect 70351 872391 70419 872447
rect 70475 872391 70488 872447
rect 70000 872323 70488 872391
rect 70000 872267 70047 872323
rect 70103 872267 70171 872323
rect 70227 872267 70295 872323
rect 70351 872267 70419 872323
rect 70475 872267 70488 872323
rect 70000 872199 70488 872267
rect 70000 872143 70047 872199
rect 70103 872143 70171 872199
rect 70227 872143 70295 872199
rect 70351 872143 70419 872199
rect 70475 872143 70488 872199
rect 70000 872075 70488 872143
rect 70000 872019 70047 872075
rect 70103 872019 70171 872075
rect 70227 872019 70295 872075
rect 70351 872019 70419 872075
rect 70475 872019 70488 872075
rect 70000 871951 70488 872019
rect 70000 871895 70047 871951
rect 70103 871895 70171 871951
rect 70227 871895 70295 871951
rect 70351 871895 70419 871951
rect 70475 871895 70488 871951
rect 70000 871828 70488 871895
rect 705512 872811 706000 872878
rect 705512 872755 705525 872811
rect 705581 872755 705649 872811
rect 705705 872755 705773 872811
rect 705829 872755 705897 872811
rect 705953 872755 706000 872811
rect 705512 872687 706000 872755
rect 705512 872631 705525 872687
rect 705581 872631 705649 872687
rect 705705 872631 705773 872687
rect 705829 872631 705897 872687
rect 705953 872631 706000 872687
rect 705512 872563 706000 872631
rect 705512 872507 705525 872563
rect 705581 872507 705649 872563
rect 705705 872507 705773 872563
rect 705829 872507 705897 872563
rect 705953 872507 706000 872563
rect 705512 872439 706000 872507
rect 705512 872383 705525 872439
rect 705581 872383 705649 872439
rect 705705 872383 705773 872439
rect 705829 872383 705897 872439
rect 705953 872383 706000 872439
rect 705512 872315 706000 872383
rect 705512 872259 705525 872315
rect 705581 872259 705649 872315
rect 705705 872259 705773 872315
rect 705829 872259 705897 872315
rect 705953 872259 706000 872315
rect 705512 872191 706000 872259
rect 705512 872135 705525 872191
rect 705581 872135 705649 872191
rect 705705 872135 705773 872191
rect 705829 872135 705897 872191
rect 705953 872135 706000 872191
rect 705512 872067 706000 872135
rect 705512 872011 705525 872067
rect 705581 872011 705649 872067
rect 705705 872011 705773 872067
rect 705829 872011 705897 872067
rect 705953 872011 706000 872067
rect 705512 871943 706000 872011
rect 705512 871887 705525 871943
rect 705581 871887 705649 871943
rect 705705 871887 705773 871943
rect 705829 871887 705897 871943
rect 705953 871887 706000 871943
rect 705512 871819 706000 871887
rect 705512 871763 705525 871819
rect 705581 871763 705649 871819
rect 705705 871763 705773 871819
rect 705829 871763 705897 871819
rect 705953 871763 706000 871819
rect 705512 871695 706000 871763
rect 705512 871639 705525 871695
rect 705581 871639 705649 871695
rect 705705 871639 705773 871695
rect 705829 871639 705897 871695
rect 705953 871639 706000 871695
rect 705512 871571 706000 871639
rect 705512 871515 705525 871571
rect 705581 871515 705649 871571
rect 705705 871515 705773 871571
rect 705829 871515 705897 871571
rect 705953 871515 706000 871571
rect 705512 871447 706000 871515
rect 705512 871391 705525 871447
rect 705581 871391 705649 871447
rect 705705 871391 705773 871447
rect 705829 871391 705897 871447
rect 705953 871391 706000 871447
rect 705512 871323 706000 871391
rect 705512 871267 705525 871323
rect 705581 871267 705649 871323
rect 705705 871267 705773 871323
rect 705829 871267 705897 871323
rect 705953 871267 706000 871323
rect 705512 871199 706000 871267
rect 70000 871105 70488 871172
rect 70000 871049 70047 871105
rect 70103 871049 70171 871105
rect 70227 871049 70295 871105
rect 70351 871049 70419 871105
rect 70475 871049 70488 871105
rect 70000 870981 70488 871049
rect 70000 870925 70047 870981
rect 70103 870925 70171 870981
rect 70227 870925 70295 870981
rect 70351 870925 70419 870981
rect 70475 870925 70488 870981
rect 70000 870857 70488 870925
rect 70000 870801 70047 870857
rect 70103 870801 70171 870857
rect 70227 870801 70295 870857
rect 70351 870801 70419 870857
rect 70475 870801 70488 870857
rect 705512 871143 705525 871199
rect 705581 871143 705649 871199
rect 705705 871143 705773 871199
rect 705829 871143 705897 871199
rect 705953 871143 706000 871199
rect 705512 871075 706000 871143
rect 705512 871019 705525 871075
rect 705581 871019 705649 871075
rect 705705 871019 705773 871075
rect 705829 871019 705897 871075
rect 705953 871019 706000 871075
rect 705512 870951 706000 871019
rect 705512 870895 705525 870951
rect 705581 870895 705649 870951
rect 705705 870895 705773 870951
rect 705829 870895 705897 870951
rect 705953 870895 706000 870951
rect 705512 870828 706000 870895
rect 70000 870733 70488 870801
rect 70000 870677 70047 870733
rect 70103 870677 70171 870733
rect 70227 870677 70295 870733
rect 70351 870677 70419 870733
rect 70475 870677 70488 870733
rect 70000 870609 70488 870677
rect 70000 870553 70047 870609
rect 70103 870553 70171 870609
rect 70227 870553 70295 870609
rect 70351 870553 70419 870609
rect 70475 870553 70488 870609
rect 70000 870485 70488 870553
rect 70000 870429 70047 870485
rect 70103 870429 70171 870485
rect 70227 870429 70295 870485
rect 70351 870429 70419 870485
rect 70475 870429 70488 870485
rect 70000 870361 70488 870429
rect 70000 870305 70047 870361
rect 70103 870305 70171 870361
rect 70227 870305 70295 870361
rect 70351 870305 70419 870361
rect 70475 870305 70488 870361
rect 70000 870237 70488 870305
rect 70000 870181 70047 870237
rect 70103 870181 70171 870237
rect 70227 870181 70295 870237
rect 70351 870181 70419 870237
rect 70475 870181 70488 870237
rect 70000 870113 70488 870181
rect 70000 870057 70047 870113
rect 70103 870057 70171 870113
rect 70227 870057 70295 870113
rect 70351 870057 70419 870113
rect 70475 870057 70488 870113
rect 70000 869989 70488 870057
rect 70000 869933 70047 869989
rect 70103 869933 70171 869989
rect 70227 869933 70295 869989
rect 70351 869933 70419 869989
rect 70475 869933 70488 869989
rect 70000 869865 70488 869933
rect 70000 869809 70047 869865
rect 70103 869809 70171 869865
rect 70227 869809 70295 869865
rect 70351 869809 70419 869865
rect 70475 869809 70488 869865
rect 70000 869741 70488 869809
rect 70000 869685 70047 869741
rect 70103 869685 70171 869741
rect 70227 869685 70295 869741
rect 70351 869685 70419 869741
rect 70475 869685 70488 869741
rect 70000 869617 70488 869685
rect 70000 869561 70047 869617
rect 70103 869561 70171 869617
rect 70227 869561 70295 869617
rect 70351 869561 70419 869617
rect 70475 869561 70488 869617
rect 70000 869493 70488 869561
rect 70000 869437 70047 869493
rect 70103 869437 70171 869493
rect 70227 869437 70295 869493
rect 70351 869437 70419 869493
rect 70475 869437 70488 869493
rect 70000 869369 70488 869437
rect 70000 869313 70047 869369
rect 70103 869313 70171 869369
rect 70227 869313 70295 869369
rect 70351 869313 70419 869369
rect 70475 869313 70488 869369
rect 70000 869245 70488 869313
rect 70000 869189 70047 869245
rect 70103 869189 70171 869245
rect 70227 869189 70295 869245
rect 70351 869189 70419 869245
rect 70475 869189 70488 869245
rect 70000 869122 70488 869189
rect 705512 870105 706000 870172
rect 705512 870049 705525 870105
rect 705581 870049 705649 870105
rect 705705 870049 705773 870105
rect 705829 870049 705897 870105
rect 705953 870049 706000 870105
rect 705512 869981 706000 870049
rect 705512 869925 705525 869981
rect 705581 869925 705649 869981
rect 705705 869925 705773 869981
rect 705829 869925 705897 869981
rect 705953 869925 706000 869981
rect 705512 869857 706000 869925
rect 705512 869801 705525 869857
rect 705581 869801 705649 869857
rect 705705 869801 705773 869857
rect 705829 869801 705897 869857
rect 705953 869801 706000 869857
rect 705512 869733 706000 869801
rect 705512 869677 705525 869733
rect 705581 869677 705649 869733
rect 705705 869677 705773 869733
rect 705829 869677 705897 869733
rect 705953 869677 706000 869733
rect 705512 869609 706000 869677
rect 705512 869553 705525 869609
rect 705581 869553 705649 869609
rect 705705 869553 705773 869609
rect 705829 869553 705897 869609
rect 705953 869553 706000 869609
rect 705512 869485 706000 869553
rect 705512 869429 705525 869485
rect 705581 869429 705649 869485
rect 705705 869429 705773 869485
rect 705829 869429 705897 869485
rect 705953 869429 706000 869485
rect 705512 869361 706000 869429
rect 705512 869305 705525 869361
rect 705581 869305 705649 869361
rect 705705 869305 705773 869361
rect 705829 869305 705897 869361
rect 705953 869305 706000 869361
rect 705512 869237 706000 869305
rect 705512 869181 705525 869237
rect 705581 869181 705649 869237
rect 705705 869181 705773 869237
rect 705829 869181 705897 869237
rect 705953 869181 706000 869237
rect 705512 869113 706000 869181
rect 705512 869057 705525 869113
rect 705581 869057 705649 869113
rect 705705 869057 705773 869113
rect 705829 869057 705897 869113
rect 705953 869057 706000 869113
rect 705512 868989 706000 869057
rect 705512 868933 705525 868989
rect 705581 868933 705649 868989
rect 705705 868933 705773 868989
rect 705829 868933 705897 868989
rect 705953 868933 706000 868989
rect 705512 868865 706000 868933
rect 705512 868809 705525 868865
rect 705581 868809 705649 868865
rect 705705 868809 705773 868865
rect 705829 868809 705897 868865
rect 705953 868809 706000 868865
rect 70000 868735 70488 868802
rect 70000 868679 70047 868735
rect 70103 868679 70171 868735
rect 70227 868679 70295 868735
rect 70351 868679 70419 868735
rect 70475 868679 70488 868735
rect 70000 868611 70488 868679
rect 70000 868555 70047 868611
rect 70103 868555 70171 868611
rect 70227 868555 70295 868611
rect 70351 868555 70419 868611
rect 70475 868555 70488 868611
rect 70000 868487 70488 868555
rect 70000 868431 70047 868487
rect 70103 868431 70171 868487
rect 70227 868431 70295 868487
rect 70351 868431 70419 868487
rect 70475 868431 70488 868487
rect 70000 868363 70488 868431
rect 70000 868307 70047 868363
rect 70103 868307 70171 868363
rect 70227 868307 70295 868363
rect 70351 868307 70419 868363
rect 70475 868307 70488 868363
rect 70000 868239 70488 868307
rect 70000 868183 70047 868239
rect 70103 868183 70171 868239
rect 70227 868183 70295 868239
rect 70351 868183 70419 868239
rect 70475 868183 70488 868239
rect 70000 868115 70488 868183
rect 705512 868741 706000 868809
rect 705512 868685 705525 868741
rect 705581 868685 705649 868741
rect 705705 868685 705773 868741
rect 705829 868685 705897 868741
rect 705953 868685 706000 868741
rect 705512 868617 706000 868685
rect 705512 868561 705525 868617
rect 705581 868561 705649 868617
rect 705705 868561 705773 868617
rect 705829 868561 705897 868617
rect 705953 868561 706000 868617
rect 705512 868493 706000 868561
rect 705512 868437 705525 868493
rect 705581 868437 705649 868493
rect 705705 868437 705773 868493
rect 705829 868437 705897 868493
rect 705953 868437 706000 868493
rect 705512 868369 706000 868437
rect 705512 868313 705525 868369
rect 705581 868313 705649 868369
rect 705705 868313 705773 868369
rect 705829 868313 705897 868369
rect 705953 868313 706000 868369
rect 705512 868245 706000 868313
rect 705512 868189 705525 868245
rect 705581 868189 705649 868245
rect 705705 868189 705773 868245
rect 705829 868189 705897 868245
rect 705953 868189 706000 868245
rect 705512 868122 706000 868189
rect 70000 868059 70047 868115
rect 70103 868059 70171 868115
rect 70227 868059 70295 868115
rect 70351 868059 70419 868115
rect 70475 868059 70488 868115
rect 70000 867991 70488 868059
rect 70000 867935 70047 867991
rect 70103 867935 70171 867991
rect 70227 867935 70295 867991
rect 70351 867935 70419 867991
rect 70475 867935 70488 867991
rect 70000 867867 70488 867935
rect 70000 867811 70047 867867
rect 70103 867811 70171 867867
rect 70227 867811 70295 867867
rect 70351 867811 70419 867867
rect 70475 867811 70488 867867
rect 70000 867743 70488 867811
rect 70000 867687 70047 867743
rect 70103 867687 70171 867743
rect 70227 867687 70295 867743
rect 70351 867687 70419 867743
rect 70475 867687 70488 867743
rect 70000 867619 70488 867687
rect 70000 867563 70047 867619
rect 70103 867563 70171 867619
rect 70227 867563 70295 867619
rect 70351 867563 70419 867619
rect 70475 867563 70488 867619
rect 70000 867495 70488 867563
rect 70000 867439 70047 867495
rect 70103 867439 70171 867495
rect 70227 867439 70295 867495
rect 70351 867439 70419 867495
rect 70475 867439 70488 867495
rect 70000 867371 70488 867439
rect 70000 867315 70047 867371
rect 70103 867315 70171 867371
rect 70227 867315 70295 867371
rect 70351 867315 70419 867371
rect 70475 867315 70488 867371
rect 70000 867247 70488 867315
rect 70000 867191 70047 867247
rect 70103 867191 70171 867247
rect 70227 867191 70295 867247
rect 70351 867191 70419 867247
rect 70475 867191 70488 867247
rect 70000 867123 70488 867191
rect 70000 867067 70047 867123
rect 70103 867067 70171 867123
rect 70227 867067 70295 867123
rect 70351 867067 70419 867123
rect 70475 867067 70488 867123
rect 70000 866999 70488 867067
rect 70000 866943 70047 866999
rect 70103 866943 70171 866999
rect 70227 866943 70295 866999
rect 70351 866943 70419 866999
rect 70475 866943 70488 866999
rect 70000 866875 70488 866943
rect 70000 866819 70047 866875
rect 70103 866819 70171 866875
rect 70227 866819 70295 866875
rect 70351 866819 70419 866875
rect 70475 866819 70488 866875
rect 70000 866752 70488 866819
rect 705512 867735 706000 867802
rect 705512 867679 705525 867735
rect 705581 867679 705649 867735
rect 705705 867679 705773 867735
rect 705829 867679 705897 867735
rect 705953 867679 706000 867735
rect 705512 867611 706000 867679
rect 705512 867555 705525 867611
rect 705581 867555 705649 867611
rect 705705 867555 705773 867611
rect 705829 867555 705897 867611
rect 705953 867555 706000 867611
rect 705512 867487 706000 867555
rect 705512 867431 705525 867487
rect 705581 867431 705649 867487
rect 705705 867431 705773 867487
rect 705829 867431 705897 867487
rect 705953 867431 706000 867487
rect 705512 867363 706000 867431
rect 705512 867307 705525 867363
rect 705581 867307 705649 867363
rect 705705 867307 705773 867363
rect 705829 867307 705897 867363
rect 705953 867307 706000 867363
rect 705512 867239 706000 867307
rect 705512 867183 705525 867239
rect 705581 867183 705649 867239
rect 705705 867183 705773 867239
rect 705829 867183 705897 867239
rect 705953 867183 706000 867239
rect 705512 867115 706000 867183
rect 705512 867059 705525 867115
rect 705581 867059 705649 867115
rect 705705 867059 705773 867115
rect 705829 867059 705897 867115
rect 705953 867059 706000 867115
rect 705512 866991 706000 867059
rect 705512 866935 705525 866991
rect 705581 866935 705649 866991
rect 705705 866935 705773 866991
rect 705829 866935 705897 866991
rect 705953 866935 706000 866991
rect 705512 866867 706000 866935
rect 705512 866811 705525 866867
rect 705581 866811 705649 866867
rect 705705 866811 705773 866867
rect 705829 866811 705897 866867
rect 705953 866811 706000 866867
rect 705512 866743 706000 866811
rect 705512 866687 705525 866743
rect 705581 866687 705649 866743
rect 705705 866687 705773 866743
rect 705829 866687 705897 866743
rect 705953 866687 706000 866743
rect 705512 866619 706000 866687
rect 705512 866563 705525 866619
rect 705581 866563 705649 866619
rect 705705 866563 705773 866619
rect 705829 866563 705897 866619
rect 705953 866563 706000 866619
rect 705512 866495 706000 866563
rect 705512 866439 705525 866495
rect 705581 866439 705649 866495
rect 705705 866439 705773 866495
rect 705829 866439 705897 866495
rect 705953 866439 706000 866495
rect 705512 866371 706000 866439
rect 705512 866315 705525 866371
rect 705581 866315 705649 866371
rect 705705 866315 705773 866371
rect 705829 866315 705897 866371
rect 705953 866315 706000 866371
rect 705512 866247 706000 866315
rect 705512 866191 705525 866247
rect 705581 866191 705649 866247
rect 705705 866191 705773 866247
rect 705829 866191 705897 866247
rect 705953 866191 706000 866247
rect 70000 866105 70488 866172
rect 70000 866049 70047 866105
rect 70103 866049 70171 866105
rect 70227 866049 70295 866105
rect 70351 866049 70419 866105
rect 70475 866049 70488 866105
rect 70000 865981 70488 866049
rect 70000 865925 70047 865981
rect 70103 865925 70171 865981
rect 70227 865925 70295 865981
rect 70351 865925 70419 865981
rect 70475 865925 70488 865981
rect 70000 865857 70488 865925
rect 70000 865801 70047 865857
rect 70103 865801 70171 865857
rect 70227 865801 70295 865857
rect 70351 865801 70419 865857
rect 70475 865801 70488 865857
rect 70000 865733 70488 865801
rect 705512 866123 706000 866191
rect 705512 866067 705525 866123
rect 705581 866067 705649 866123
rect 705705 866067 705773 866123
rect 705829 866067 705897 866123
rect 705953 866067 706000 866123
rect 705512 865999 706000 866067
rect 705512 865943 705525 865999
rect 705581 865943 705649 865999
rect 705705 865943 705773 865999
rect 705829 865943 705897 865999
rect 705953 865943 706000 865999
rect 705512 865875 706000 865943
rect 705512 865819 705525 865875
rect 705581 865819 705649 865875
rect 705705 865819 705773 865875
rect 705829 865819 705897 865875
rect 705953 865819 706000 865875
rect 705512 865752 706000 865819
rect 70000 865677 70047 865733
rect 70103 865677 70171 865733
rect 70227 865677 70295 865733
rect 70351 865677 70419 865733
rect 70475 865677 70488 865733
rect 70000 865609 70488 865677
rect 70000 865553 70047 865609
rect 70103 865553 70171 865609
rect 70227 865553 70295 865609
rect 70351 865553 70419 865609
rect 70475 865553 70488 865609
rect 70000 865485 70488 865553
rect 70000 865429 70047 865485
rect 70103 865429 70171 865485
rect 70227 865429 70295 865485
rect 70351 865429 70419 865485
rect 70475 865429 70488 865485
rect 70000 865361 70488 865429
rect 70000 865305 70047 865361
rect 70103 865305 70171 865361
rect 70227 865305 70295 865361
rect 70351 865305 70419 865361
rect 70475 865305 70488 865361
rect 70000 865237 70488 865305
rect 70000 865181 70047 865237
rect 70103 865181 70171 865237
rect 70227 865181 70295 865237
rect 70351 865181 70419 865237
rect 70475 865181 70488 865237
rect 70000 865113 70488 865181
rect 70000 865057 70047 865113
rect 70103 865057 70171 865113
rect 70227 865057 70295 865113
rect 70351 865057 70419 865113
rect 70475 865057 70488 865113
rect 70000 864989 70488 865057
rect 70000 864933 70047 864989
rect 70103 864933 70171 864989
rect 70227 864933 70295 864989
rect 70351 864933 70419 864989
rect 70475 864933 70488 864989
rect 70000 864865 70488 864933
rect 70000 864809 70047 864865
rect 70103 864809 70171 864865
rect 70227 864809 70295 864865
rect 70351 864809 70419 864865
rect 70475 864809 70488 864865
rect 70000 864741 70488 864809
rect 70000 864685 70047 864741
rect 70103 864685 70171 864741
rect 70227 864685 70295 864741
rect 70351 864685 70419 864741
rect 70475 864685 70488 864741
rect 70000 864617 70488 864685
rect 70000 864561 70047 864617
rect 70103 864561 70171 864617
rect 70227 864561 70295 864617
rect 70351 864561 70419 864617
rect 70475 864561 70488 864617
rect 70000 864493 70488 864561
rect 70000 864437 70047 864493
rect 70103 864437 70171 864493
rect 70227 864437 70295 864493
rect 70351 864437 70419 864493
rect 70475 864437 70488 864493
rect 70000 864369 70488 864437
rect 70000 864313 70047 864369
rect 70103 864313 70171 864369
rect 70227 864313 70295 864369
rect 70351 864313 70419 864369
rect 70475 864313 70488 864369
rect 70000 864272 70488 864313
rect 705512 865131 706000 865172
rect 705512 865075 705525 865131
rect 705581 865075 705649 865131
rect 705705 865075 705773 865131
rect 705829 865075 705897 865131
rect 705953 865075 706000 865131
rect 705512 865007 706000 865075
rect 705512 864951 705525 865007
rect 705581 864951 705649 865007
rect 705705 864951 705773 865007
rect 705829 864951 705897 865007
rect 705953 864951 706000 865007
rect 705512 864883 706000 864951
rect 705512 864827 705525 864883
rect 705581 864827 705649 864883
rect 705705 864827 705773 864883
rect 705829 864827 705897 864883
rect 705953 864827 706000 864883
rect 705512 864759 706000 864827
rect 705512 864703 705525 864759
rect 705581 864703 705649 864759
rect 705705 864703 705773 864759
rect 705829 864703 705897 864759
rect 705953 864703 706000 864759
rect 705512 864635 706000 864703
rect 705512 864579 705525 864635
rect 705581 864579 705649 864635
rect 705705 864579 705773 864635
rect 705829 864579 705897 864635
rect 705953 864579 706000 864635
rect 705512 864511 706000 864579
rect 705512 864455 705525 864511
rect 705581 864455 705649 864511
rect 705705 864455 705773 864511
rect 705829 864455 705897 864511
rect 705953 864455 706000 864511
rect 705512 864387 706000 864455
rect 705512 864331 705525 864387
rect 705581 864331 705649 864387
rect 705705 864331 705773 864387
rect 705829 864331 705897 864387
rect 705953 864331 706000 864387
rect 705512 864263 706000 864331
rect 705512 864207 705525 864263
rect 705581 864207 705649 864263
rect 705705 864207 705773 864263
rect 705829 864207 705897 864263
rect 705953 864207 706000 864263
rect 705512 864139 706000 864207
rect 705512 864083 705525 864139
rect 705581 864083 705649 864139
rect 705705 864083 705773 864139
rect 705829 864083 705897 864139
rect 705953 864083 706000 864139
rect 705512 864015 706000 864083
rect 705512 863959 705525 864015
rect 705581 863959 705649 864015
rect 705705 863959 705773 864015
rect 705829 863959 705897 864015
rect 705953 863959 706000 864015
rect 705512 863891 706000 863959
rect 705512 863835 705525 863891
rect 705581 863835 705649 863891
rect 705705 863835 705773 863891
rect 705829 863835 705897 863891
rect 705953 863835 706000 863891
rect 705512 863767 706000 863835
rect 705512 863711 705525 863767
rect 705581 863711 705649 863767
rect 705705 863711 705773 863767
rect 705829 863711 705897 863767
rect 705953 863711 706000 863767
rect 705512 863643 706000 863711
rect 705512 863587 705525 863643
rect 705581 863587 705649 863643
rect 705705 863587 705773 863643
rect 705829 863587 705897 863643
rect 705953 863587 706000 863643
rect 705512 863519 706000 863587
rect 705512 863463 705525 863519
rect 705581 863463 705649 863519
rect 705705 863463 705773 863519
rect 705829 863463 705897 863519
rect 705953 863463 706000 863519
rect 705512 863395 706000 863463
rect 705512 863339 705525 863395
rect 705581 863339 705649 863395
rect 705705 863339 705773 863395
rect 705829 863339 705897 863395
rect 705953 863339 706000 863395
rect 705512 863272 706000 863339
rect 70000 837661 70488 837728
rect 70000 837605 70047 837661
rect 70103 837605 70171 837661
rect 70227 837605 70295 837661
rect 70351 837605 70419 837661
rect 70475 837605 70488 837661
rect 70000 837537 70488 837605
rect 70000 837481 70047 837537
rect 70103 837481 70171 837537
rect 70227 837481 70295 837537
rect 70351 837481 70419 837537
rect 70475 837481 70488 837537
rect 70000 837413 70488 837481
rect 70000 837357 70047 837413
rect 70103 837357 70171 837413
rect 70227 837357 70295 837413
rect 70351 837357 70419 837413
rect 70475 837357 70488 837413
rect 70000 837289 70488 837357
rect 70000 837233 70047 837289
rect 70103 837233 70171 837289
rect 70227 837233 70295 837289
rect 70351 837233 70419 837289
rect 70475 837233 70488 837289
rect 70000 837165 70488 837233
rect 70000 837109 70047 837165
rect 70103 837109 70171 837165
rect 70227 837109 70295 837165
rect 70351 837109 70419 837165
rect 70475 837109 70488 837165
rect 70000 837041 70488 837109
rect 70000 836985 70047 837041
rect 70103 836985 70171 837041
rect 70227 836985 70295 837041
rect 70351 836985 70419 837041
rect 70475 836985 70488 837041
rect 70000 836917 70488 836985
rect 70000 836861 70047 836917
rect 70103 836861 70171 836917
rect 70227 836861 70295 836917
rect 70351 836861 70419 836917
rect 70475 836861 70488 836917
rect 70000 836793 70488 836861
rect 70000 836737 70047 836793
rect 70103 836737 70171 836793
rect 70227 836737 70295 836793
rect 70351 836737 70419 836793
rect 70475 836737 70488 836793
rect 70000 836669 70488 836737
rect 70000 836613 70047 836669
rect 70103 836613 70171 836669
rect 70227 836613 70295 836669
rect 70351 836613 70419 836669
rect 70475 836613 70488 836669
rect 70000 836545 70488 836613
rect 70000 836489 70047 836545
rect 70103 836489 70171 836545
rect 70227 836489 70295 836545
rect 70351 836489 70419 836545
rect 70475 836489 70488 836545
rect 70000 836421 70488 836489
rect 70000 836365 70047 836421
rect 70103 836365 70171 836421
rect 70227 836365 70295 836421
rect 70351 836365 70419 836421
rect 70475 836365 70488 836421
rect 70000 836297 70488 836365
rect 70000 836241 70047 836297
rect 70103 836241 70171 836297
rect 70227 836241 70295 836297
rect 70351 836241 70419 836297
rect 70475 836241 70488 836297
rect 70000 836173 70488 836241
rect 70000 836117 70047 836173
rect 70103 836117 70171 836173
rect 70227 836117 70295 836173
rect 70351 836117 70419 836173
rect 70475 836117 70488 836173
rect 70000 836049 70488 836117
rect 70000 835993 70047 836049
rect 70103 835993 70171 836049
rect 70227 835993 70295 836049
rect 70351 835993 70419 836049
rect 70475 835993 70488 836049
rect 70000 835925 70488 835993
rect 70000 835869 70047 835925
rect 70103 835869 70171 835925
rect 70227 835869 70295 835925
rect 70351 835869 70419 835925
rect 70475 835869 70488 835925
rect 70000 835828 70488 835869
rect 70000 835181 70488 835248
rect 70000 835125 70047 835181
rect 70103 835125 70171 835181
rect 70227 835125 70295 835181
rect 70351 835125 70419 835181
rect 70475 835125 70488 835181
rect 70000 835057 70488 835125
rect 70000 835001 70047 835057
rect 70103 835001 70171 835057
rect 70227 835001 70295 835057
rect 70351 835001 70419 835057
rect 70475 835001 70488 835057
rect 70000 834933 70488 835001
rect 70000 834877 70047 834933
rect 70103 834877 70171 834933
rect 70227 834877 70295 834933
rect 70351 834877 70419 834933
rect 70475 834877 70488 834933
rect 70000 834809 70488 834877
rect 70000 834753 70047 834809
rect 70103 834753 70171 834809
rect 70227 834753 70295 834809
rect 70351 834753 70419 834809
rect 70475 834753 70488 834809
rect 70000 834685 70488 834753
rect 70000 834629 70047 834685
rect 70103 834629 70171 834685
rect 70227 834629 70295 834685
rect 70351 834629 70419 834685
rect 70475 834629 70488 834685
rect 70000 834561 70488 834629
rect 70000 834505 70047 834561
rect 70103 834505 70171 834561
rect 70227 834505 70295 834561
rect 70351 834505 70419 834561
rect 70475 834505 70488 834561
rect 70000 834437 70488 834505
rect 70000 834381 70047 834437
rect 70103 834381 70171 834437
rect 70227 834381 70295 834437
rect 70351 834381 70419 834437
rect 70475 834381 70488 834437
rect 70000 834313 70488 834381
rect 70000 834257 70047 834313
rect 70103 834257 70171 834313
rect 70227 834257 70295 834313
rect 70351 834257 70419 834313
rect 70475 834257 70488 834313
rect 70000 834189 70488 834257
rect 70000 834133 70047 834189
rect 70103 834133 70171 834189
rect 70227 834133 70295 834189
rect 70351 834133 70419 834189
rect 70475 834133 70488 834189
rect 70000 834065 70488 834133
rect 70000 834009 70047 834065
rect 70103 834009 70171 834065
rect 70227 834009 70295 834065
rect 70351 834009 70419 834065
rect 70475 834009 70488 834065
rect 70000 833941 70488 834009
rect 70000 833885 70047 833941
rect 70103 833885 70171 833941
rect 70227 833885 70295 833941
rect 70351 833885 70419 833941
rect 70475 833885 70488 833941
rect 70000 833817 70488 833885
rect 70000 833761 70047 833817
rect 70103 833761 70171 833817
rect 70227 833761 70295 833817
rect 70351 833761 70419 833817
rect 70475 833761 70488 833817
rect 70000 833693 70488 833761
rect 70000 833637 70047 833693
rect 70103 833637 70171 833693
rect 70227 833637 70295 833693
rect 70351 833637 70419 833693
rect 70475 833637 70488 833693
rect 70000 833569 70488 833637
rect 70000 833513 70047 833569
rect 70103 833513 70171 833569
rect 70227 833513 70295 833569
rect 70351 833513 70419 833569
rect 70475 833513 70488 833569
rect 70000 833445 70488 833513
rect 70000 833389 70047 833445
rect 70103 833389 70171 833445
rect 70227 833389 70295 833445
rect 70351 833389 70419 833445
rect 70475 833389 70488 833445
rect 70000 833321 70488 833389
rect 70000 833265 70047 833321
rect 70103 833265 70171 833321
rect 70227 833265 70295 833321
rect 70351 833265 70419 833321
rect 70475 833265 70488 833321
rect 70000 833198 70488 833265
rect 70000 832811 70488 832878
rect 70000 832755 70047 832811
rect 70103 832755 70171 832811
rect 70227 832755 70295 832811
rect 70351 832755 70419 832811
rect 70475 832755 70488 832811
rect 70000 832687 70488 832755
rect 70000 832631 70047 832687
rect 70103 832631 70171 832687
rect 70227 832631 70295 832687
rect 70351 832631 70419 832687
rect 70475 832631 70488 832687
rect 70000 832563 70488 832631
rect 70000 832507 70047 832563
rect 70103 832507 70171 832563
rect 70227 832507 70295 832563
rect 70351 832507 70419 832563
rect 70475 832507 70488 832563
rect 70000 832439 70488 832507
rect 70000 832383 70047 832439
rect 70103 832383 70171 832439
rect 70227 832383 70295 832439
rect 70351 832383 70419 832439
rect 70475 832383 70488 832439
rect 70000 832315 70488 832383
rect 70000 832259 70047 832315
rect 70103 832259 70171 832315
rect 70227 832259 70295 832315
rect 70351 832259 70419 832315
rect 70475 832259 70488 832315
rect 70000 832191 70488 832259
rect 70000 832135 70047 832191
rect 70103 832135 70171 832191
rect 70227 832135 70295 832191
rect 70351 832135 70419 832191
rect 70475 832135 70488 832191
rect 70000 832067 70488 832135
rect 70000 832011 70047 832067
rect 70103 832011 70171 832067
rect 70227 832011 70295 832067
rect 70351 832011 70419 832067
rect 70475 832011 70488 832067
rect 70000 831943 70488 832011
rect 70000 831887 70047 831943
rect 70103 831887 70171 831943
rect 70227 831887 70295 831943
rect 70351 831887 70419 831943
rect 70475 831887 70488 831943
rect 70000 831819 70488 831887
rect 70000 831763 70047 831819
rect 70103 831763 70171 831819
rect 70227 831763 70295 831819
rect 70351 831763 70419 831819
rect 70475 831763 70488 831819
rect 70000 831695 70488 831763
rect 70000 831639 70047 831695
rect 70103 831639 70171 831695
rect 70227 831639 70295 831695
rect 70351 831639 70419 831695
rect 70475 831639 70488 831695
rect 70000 831571 70488 831639
rect 70000 831515 70047 831571
rect 70103 831515 70171 831571
rect 70227 831515 70295 831571
rect 70351 831515 70419 831571
rect 70475 831515 70488 831571
rect 70000 831447 70488 831515
rect 70000 831391 70047 831447
rect 70103 831391 70171 831447
rect 70227 831391 70295 831447
rect 70351 831391 70419 831447
rect 70475 831391 70488 831447
rect 70000 831323 70488 831391
rect 70000 831267 70047 831323
rect 70103 831267 70171 831323
rect 70227 831267 70295 831323
rect 70351 831267 70419 831323
rect 70475 831267 70488 831323
rect 70000 831199 70488 831267
rect 70000 831143 70047 831199
rect 70103 831143 70171 831199
rect 70227 831143 70295 831199
rect 70351 831143 70419 831199
rect 70475 831143 70488 831199
rect 70000 831075 70488 831143
rect 70000 831019 70047 831075
rect 70103 831019 70171 831075
rect 70227 831019 70295 831075
rect 70351 831019 70419 831075
rect 70475 831019 70488 831075
rect 70000 830951 70488 831019
rect 70000 830895 70047 830951
rect 70103 830895 70171 830951
rect 70227 830895 70295 830951
rect 70351 830895 70419 830951
rect 70475 830895 70488 830951
rect 70000 830828 70488 830895
rect 70000 830105 70488 830172
rect 70000 830049 70047 830105
rect 70103 830049 70171 830105
rect 70227 830049 70295 830105
rect 70351 830049 70419 830105
rect 70475 830049 70488 830105
rect 70000 829981 70488 830049
rect 70000 829925 70047 829981
rect 70103 829925 70171 829981
rect 70227 829925 70295 829981
rect 70351 829925 70419 829981
rect 70475 829925 70488 829981
rect 70000 829857 70488 829925
rect 70000 829801 70047 829857
rect 70103 829801 70171 829857
rect 70227 829801 70295 829857
rect 70351 829801 70419 829857
rect 70475 829801 70488 829857
rect 70000 829733 70488 829801
rect 70000 829677 70047 829733
rect 70103 829677 70171 829733
rect 70227 829677 70295 829733
rect 70351 829677 70419 829733
rect 70475 829677 70488 829733
rect 70000 829609 70488 829677
rect 70000 829553 70047 829609
rect 70103 829553 70171 829609
rect 70227 829553 70295 829609
rect 70351 829553 70419 829609
rect 70475 829553 70488 829609
rect 70000 829485 70488 829553
rect 70000 829429 70047 829485
rect 70103 829429 70171 829485
rect 70227 829429 70295 829485
rect 70351 829429 70419 829485
rect 70475 829429 70488 829485
rect 70000 829361 70488 829429
rect 70000 829305 70047 829361
rect 70103 829305 70171 829361
rect 70227 829305 70295 829361
rect 70351 829305 70419 829361
rect 70475 829305 70488 829361
rect 70000 829237 70488 829305
rect 70000 829181 70047 829237
rect 70103 829181 70171 829237
rect 70227 829181 70295 829237
rect 70351 829181 70419 829237
rect 70475 829181 70488 829237
rect 70000 829113 70488 829181
rect 70000 829057 70047 829113
rect 70103 829057 70171 829113
rect 70227 829057 70295 829113
rect 70351 829057 70419 829113
rect 70475 829057 70488 829113
rect 70000 828989 70488 829057
rect 70000 828933 70047 828989
rect 70103 828933 70171 828989
rect 70227 828933 70295 828989
rect 70351 828933 70419 828989
rect 70475 828933 70488 828989
rect 70000 828865 70488 828933
rect 70000 828809 70047 828865
rect 70103 828809 70171 828865
rect 70227 828809 70295 828865
rect 70351 828809 70419 828865
rect 70475 828809 70488 828865
rect 70000 828741 70488 828809
rect 70000 828685 70047 828741
rect 70103 828685 70171 828741
rect 70227 828685 70295 828741
rect 70351 828685 70419 828741
rect 70475 828685 70488 828741
rect 70000 828617 70488 828685
rect 70000 828561 70047 828617
rect 70103 828561 70171 828617
rect 70227 828561 70295 828617
rect 70351 828561 70419 828617
rect 70475 828561 70488 828617
rect 70000 828493 70488 828561
rect 70000 828437 70047 828493
rect 70103 828437 70171 828493
rect 70227 828437 70295 828493
rect 70351 828437 70419 828493
rect 70475 828437 70488 828493
rect 70000 828369 70488 828437
rect 70000 828313 70047 828369
rect 70103 828313 70171 828369
rect 70227 828313 70295 828369
rect 70351 828313 70419 828369
rect 70475 828313 70488 828369
rect 70000 828245 70488 828313
rect 70000 828189 70047 828245
rect 70103 828189 70171 828245
rect 70227 828189 70295 828245
rect 70351 828189 70419 828245
rect 70475 828189 70488 828245
rect 70000 828122 70488 828189
rect 70000 827735 70488 827802
rect 70000 827679 70047 827735
rect 70103 827679 70171 827735
rect 70227 827679 70295 827735
rect 70351 827679 70419 827735
rect 70475 827679 70488 827735
rect 70000 827611 70488 827679
rect 70000 827555 70047 827611
rect 70103 827555 70171 827611
rect 70227 827555 70295 827611
rect 70351 827555 70419 827611
rect 70475 827555 70488 827611
rect 70000 827487 70488 827555
rect 70000 827431 70047 827487
rect 70103 827431 70171 827487
rect 70227 827431 70295 827487
rect 70351 827431 70419 827487
rect 70475 827431 70488 827487
rect 70000 827363 70488 827431
rect 70000 827307 70047 827363
rect 70103 827307 70171 827363
rect 70227 827307 70295 827363
rect 70351 827307 70419 827363
rect 70475 827307 70488 827363
rect 70000 827239 70488 827307
rect 70000 827183 70047 827239
rect 70103 827183 70171 827239
rect 70227 827183 70295 827239
rect 70351 827183 70419 827239
rect 70475 827183 70488 827239
rect 70000 827115 70488 827183
rect 70000 827059 70047 827115
rect 70103 827059 70171 827115
rect 70227 827059 70295 827115
rect 70351 827059 70419 827115
rect 70475 827059 70488 827115
rect 70000 826991 70488 827059
rect 70000 826935 70047 826991
rect 70103 826935 70171 826991
rect 70227 826935 70295 826991
rect 70351 826935 70419 826991
rect 70475 826935 70488 826991
rect 70000 826867 70488 826935
rect 70000 826811 70047 826867
rect 70103 826811 70171 826867
rect 70227 826811 70295 826867
rect 70351 826811 70419 826867
rect 70475 826811 70488 826867
rect 70000 826743 70488 826811
rect 70000 826687 70047 826743
rect 70103 826687 70171 826743
rect 70227 826687 70295 826743
rect 70351 826687 70419 826743
rect 70475 826687 70488 826743
rect 70000 826619 70488 826687
rect 70000 826563 70047 826619
rect 70103 826563 70171 826619
rect 70227 826563 70295 826619
rect 70351 826563 70419 826619
rect 70475 826563 70488 826619
rect 70000 826495 70488 826563
rect 70000 826439 70047 826495
rect 70103 826439 70171 826495
rect 70227 826439 70295 826495
rect 70351 826439 70419 826495
rect 70475 826439 70488 826495
rect 70000 826371 70488 826439
rect 70000 826315 70047 826371
rect 70103 826315 70171 826371
rect 70227 826315 70295 826371
rect 70351 826315 70419 826371
rect 70475 826315 70488 826371
rect 70000 826247 70488 826315
rect 70000 826191 70047 826247
rect 70103 826191 70171 826247
rect 70227 826191 70295 826247
rect 70351 826191 70419 826247
rect 70475 826191 70488 826247
rect 70000 826123 70488 826191
rect 70000 826067 70047 826123
rect 70103 826067 70171 826123
rect 70227 826067 70295 826123
rect 70351 826067 70419 826123
rect 70475 826067 70488 826123
rect 70000 825999 70488 826067
rect 70000 825943 70047 825999
rect 70103 825943 70171 825999
rect 70227 825943 70295 825999
rect 70351 825943 70419 825999
rect 70475 825943 70488 825999
rect 70000 825875 70488 825943
rect 70000 825819 70047 825875
rect 70103 825819 70171 825875
rect 70227 825819 70295 825875
rect 70351 825819 70419 825875
rect 70475 825819 70488 825875
rect 70000 825752 70488 825819
rect 70000 825105 70488 825172
rect 70000 825049 70047 825105
rect 70103 825049 70171 825105
rect 70227 825049 70295 825105
rect 70351 825049 70419 825105
rect 70475 825049 70488 825105
rect 70000 824981 70488 825049
rect 70000 824925 70047 824981
rect 70103 824925 70171 824981
rect 70227 824925 70295 824981
rect 70351 824925 70419 824981
rect 70475 824925 70488 824981
rect 70000 824857 70488 824925
rect 70000 824801 70047 824857
rect 70103 824801 70171 824857
rect 70227 824801 70295 824857
rect 70351 824801 70419 824857
rect 70475 824801 70488 824857
rect 70000 824733 70488 824801
rect 70000 824677 70047 824733
rect 70103 824677 70171 824733
rect 70227 824677 70295 824733
rect 70351 824677 70419 824733
rect 70475 824677 70488 824733
rect 70000 824609 70488 824677
rect 70000 824553 70047 824609
rect 70103 824553 70171 824609
rect 70227 824553 70295 824609
rect 70351 824553 70419 824609
rect 70475 824553 70488 824609
rect 70000 824485 70488 824553
rect 70000 824429 70047 824485
rect 70103 824429 70171 824485
rect 70227 824429 70295 824485
rect 70351 824429 70419 824485
rect 70475 824429 70488 824485
rect 70000 824361 70488 824429
rect 70000 824305 70047 824361
rect 70103 824305 70171 824361
rect 70227 824305 70295 824361
rect 70351 824305 70419 824361
rect 70475 824305 70488 824361
rect 70000 824237 70488 824305
rect 70000 824181 70047 824237
rect 70103 824181 70171 824237
rect 70227 824181 70295 824237
rect 70351 824181 70419 824237
rect 70475 824181 70488 824237
rect 70000 824113 70488 824181
rect 70000 824057 70047 824113
rect 70103 824057 70171 824113
rect 70227 824057 70295 824113
rect 70351 824057 70419 824113
rect 70475 824057 70488 824113
rect 70000 823989 70488 824057
rect 70000 823933 70047 823989
rect 70103 823933 70171 823989
rect 70227 823933 70295 823989
rect 70351 823933 70419 823989
rect 70475 823933 70488 823989
rect 70000 823865 70488 823933
rect 70000 823809 70047 823865
rect 70103 823809 70171 823865
rect 70227 823809 70295 823865
rect 70351 823809 70419 823865
rect 70475 823809 70488 823865
rect 70000 823741 70488 823809
rect 70000 823685 70047 823741
rect 70103 823685 70171 823741
rect 70227 823685 70295 823741
rect 70351 823685 70419 823741
rect 70475 823685 70488 823741
rect 70000 823617 70488 823685
rect 70000 823561 70047 823617
rect 70103 823561 70171 823617
rect 70227 823561 70295 823617
rect 70351 823561 70419 823617
rect 70475 823561 70488 823617
rect 70000 823493 70488 823561
rect 70000 823437 70047 823493
rect 70103 823437 70171 823493
rect 70227 823437 70295 823493
rect 70351 823437 70419 823493
rect 70475 823437 70488 823493
rect 70000 823369 70488 823437
rect 70000 823313 70047 823369
rect 70103 823313 70171 823369
rect 70227 823313 70295 823369
rect 70351 823313 70419 823369
rect 70475 823313 70488 823369
rect 70000 823272 70488 823313
rect 70000 796661 70488 796728
rect 70000 796605 70047 796661
rect 70103 796605 70171 796661
rect 70227 796605 70295 796661
rect 70351 796605 70419 796661
rect 70475 796605 70488 796661
rect 70000 796537 70488 796605
rect 70000 796481 70047 796537
rect 70103 796481 70171 796537
rect 70227 796481 70295 796537
rect 70351 796481 70419 796537
rect 70475 796481 70488 796537
rect 70000 796413 70488 796481
rect 70000 796357 70047 796413
rect 70103 796357 70171 796413
rect 70227 796357 70295 796413
rect 70351 796357 70419 796413
rect 70475 796357 70488 796413
rect 70000 796289 70488 796357
rect 70000 796233 70047 796289
rect 70103 796233 70171 796289
rect 70227 796233 70295 796289
rect 70351 796233 70419 796289
rect 70475 796233 70488 796289
rect 70000 796165 70488 796233
rect 70000 796109 70047 796165
rect 70103 796109 70171 796165
rect 70227 796109 70295 796165
rect 70351 796109 70419 796165
rect 70475 796109 70488 796165
rect 70000 796041 70488 796109
rect 70000 795985 70047 796041
rect 70103 795985 70171 796041
rect 70227 795985 70295 796041
rect 70351 795985 70419 796041
rect 70475 795985 70488 796041
rect 70000 795917 70488 795985
rect 70000 795861 70047 795917
rect 70103 795861 70171 795917
rect 70227 795861 70295 795917
rect 70351 795861 70419 795917
rect 70475 795861 70488 795917
rect 70000 795793 70488 795861
rect 70000 795737 70047 795793
rect 70103 795737 70171 795793
rect 70227 795737 70295 795793
rect 70351 795737 70419 795793
rect 70475 795737 70488 795793
rect 70000 795669 70488 795737
rect 70000 795613 70047 795669
rect 70103 795613 70171 795669
rect 70227 795613 70295 795669
rect 70351 795613 70419 795669
rect 70475 795613 70488 795669
rect 70000 795545 70488 795613
rect 70000 795489 70047 795545
rect 70103 795489 70171 795545
rect 70227 795489 70295 795545
rect 70351 795489 70419 795545
rect 70475 795489 70488 795545
rect 70000 795421 70488 795489
rect 70000 795365 70047 795421
rect 70103 795365 70171 795421
rect 70227 795365 70295 795421
rect 70351 795365 70419 795421
rect 70475 795365 70488 795421
rect 70000 795297 70488 795365
rect 70000 795241 70047 795297
rect 70103 795241 70171 795297
rect 70227 795241 70295 795297
rect 70351 795241 70419 795297
rect 70475 795241 70488 795297
rect 70000 795173 70488 795241
rect 70000 795117 70047 795173
rect 70103 795117 70171 795173
rect 70227 795117 70295 795173
rect 70351 795117 70419 795173
rect 70475 795117 70488 795173
rect 70000 795049 70488 795117
rect 70000 794993 70047 795049
rect 70103 794993 70171 795049
rect 70227 794993 70295 795049
rect 70351 794993 70419 795049
rect 70475 794993 70488 795049
rect 70000 794925 70488 794993
rect 70000 794869 70047 794925
rect 70103 794869 70171 794925
rect 70227 794869 70295 794925
rect 70351 794869 70419 794925
rect 70475 794869 70488 794925
rect 70000 794828 70488 794869
rect 70000 794181 70488 794248
rect 70000 794125 70047 794181
rect 70103 794125 70171 794181
rect 70227 794125 70295 794181
rect 70351 794125 70419 794181
rect 70475 794125 70488 794181
rect 70000 794057 70488 794125
rect 70000 794001 70047 794057
rect 70103 794001 70171 794057
rect 70227 794001 70295 794057
rect 70351 794001 70419 794057
rect 70475 794001 70488 794057
rect 70000 793933 70488 794001
rect 70000 793877 70047 793933
rect 70103 793877 70171 793933
rect 70227 793877 70295 793933
rect 70351 793877 70419 793933
rect 70475 793877 70488 793933
rect 70000 793809 70488 793877
rect 70000 793753 70047 793809
rect 70103 793753 70171 793809
rect 70227 793753 70295 793809
rect 70351 793753 70419 793809
rect 70475 793753 70488 793809
rect 70000 793685 70488 793753
rect 70000 793629 70047 793685
rect 70103 793629 70171 793685
rect 70227 793629 70295 793685
rect 70351 793629 70419 793685
rect 70475 793629 70488 793685
rect 70000 793561 70488 793629
rect 70000 793505 70047 793561
rect 70103 793505 70171 793561
rect 70227 793505 70295 793561
rect 70351 793505 70419 793561
rect 70475 793505 70488 793561
rect 70000 793437 70488 793505
rect 70000 793381 70047 793437
rect 70103 793381 70171 793437
rect 70227 793381 70295 793437
rect 70351 793381 70419 793437
rect 70475 793381 70488 793437
rect 70000 793313 70488 793381
rect 70000 793257 70047 793313
rect 70103 793257 70171 793313
rect 70227 793257 70295 793313
rect 70351 793257 70419 793313
rect 70475 793257 70488 793313
rect 70000 793189 70488 793257
rect 70000 793133 70047 793189
rect 70103 793133 70171 793189
rect 70227 793133 70295 793189
rect 70351 793133 70419 793189
rect 70475 793133 70488 793189
rect 70000 793065 70488 793133
rect 70000 793009 70047 793065
rect 70103 793009 70171 793065
rect 70227 793009 70295 793065
rect 70351 793009 70419 793065
rect 70475 793009 70488 793065
rect 70000 792941 70488 793009
rect 70000 792885 70047 792941
rect 70103 792885 70171 792941
rect 70227 792885 70295 792941
rect 70351 792885 70419 792941
rect 70475 792885 70488 792941
rect 70000 792817 70488 792885
rect 70000 792761 70047 792817
rect 70103 792761 70171 792817
rect 70227 792761 70295 792817
rect 70351 792761 70419 792817
rect 70475 792761 70488 792817
rect 70000 792693 70488 792761
rect 70000 792637 70047 792693
rect 70103 792637 70171 792693
rect 70227 792637 70295 792693
rect 70351 792637 70419 792693
rect 70475 792637 70488 792693
rect 70000 792569 70488 792637
rect 70000 792513 70047 792569
rect 70103 792513 70171 792569
rect 70227 792513 70295 792569
rect 70351 792513 70419 792569
rect 70475 792513 70488 792569
rect 70000 792445 70488 792513
rect 70000 792389 70047 792445
rect 70103 792389 70171 792445
rect 70227 792389 70295 792445
rect 70351 792389 70419 792445
rect 70475 792389 70488 792445
rect 70000 792321 70488 792389
rect 70000 792265 70047 792321
rect 70103 792265 70171 792321
rect 70227 792265 70295 792321
rect 70351 792265 70419 792321
rect 70475 792265 70488 792321
rect 70000 792198 70488 792265
rect 70000 791811 70488 791878
rect 70000 791755 70047 791811
rect 70103 791755 70171 791811
rect 70227 791755 70295 791811
rect 70351 791755 70419 791811
rect 70475 791755 70488 791811
rect 70000 791687 70488 791755
rect 70000 791631 70047 791687
rect 70103 791631 70171 791687
rect 70227 791631 70295 791687
rect 70351 791631 70419 791687
rect 70475 791631 70488 791687
rect 70000 791563 70488 791631
rect 70000 791507 70047 791563
rect 70103 791507 70171 791563
rect 70227 791507 70295 791563
rect 70351 791507 70419 791563
rect 70475 791507 70488 791563
rect 70000 791439 70488 791507
rect 70000 791383 70047 791439
rect 70103 791383 70171 791439
rect 70227 791383 70295 791439
rect 70351 791383 70419 791439
rect 70475 791383 70488 791439
rect 70000 791315 70488 791383
rect 70000 791259 70047 791315
rect 70103 791259 70171 791315
rect 70227 791259 70295 791315
rect 70351 791259 70419 791315
rect 70475 791259 70488 791315
rect 70000 791191 70488 791259
rect 70000 791135 70047 791191
rect 70103 791135 70171 791191
rect 70227 791135 70295 791191
rect 70351 791135 70419 791191
rect 70475 791135 70488 791191
rect 70000 791067 70488 791135
rect 70000 791011 70047 791067
rect 70103 791011 70171 791067
rect 70227 791011 70295 791067
rect 70351 791011 70419 791067
rect 70475 791011 70488 791067
rect 70000 790943 70488 791011
rect 70000 790887 70047 790943
rect 70103 790887 70171 790943
rect 70227 790887 70295 790943
rect 70351 790887 70419 790943
rect 70475 790887 70488 790943
rect 70000 790819 70488 790887
rect 70000 790763 70047 790819
rect 70103 790763 70171 790819
rect 70227 790763 70295 790819
rect 70351 790763 70419 790819
rect 70475 790763 70488 790819
rect 70000 790695 70488 790763
rect 70000 790639 70047 790695
rect 70103 790639 70171 790695
rect 70227 790639 70295 790695
rect 70351 790639 70419 790695
rect 70475 790639 70488 790695
rect 70000 790571 70488 790639
rect 70000 790515 70047 790571
rect 70103 790515 70171 790571
rect 70227 790515 70295 790571
rect 70351 790515 70419 790571
rect 70475 790515 70488 790571
rect 70000 790447 70488 790515
rect 70000 790391 70047 790447
rect 70103 790391 70171 790447
rect 70227 790391 70295 790447
rect 70351 790391 70419 790447
rect 70475 790391 70488 790447
rect 70000 790323 70488 790391
rect 70000 790267 70047 790323
rect 70103 790267 70171 790323
rect 70227 790267 70295 790323
rect 70351 790267 70419 790323
rect 70475 790267 70488 790323
rect 70000 790199 70488 790267
rect 70000 790143 70047 790199
rect 70103 790143 70171 790199
rect 70227 790143 70295 790199
rect 70351 790143 70419 790199
rect 70475 790143 70488 790199
rect 70000 790075 70488 790143
rect 70000 790019 70047 790075
rect 70103 790019 70171 790075
rect 70227 790019 70295 790075
rect 70351 790019 70419 790075
rect 70475 790019 70488 790075
rect 70000 789951 70488 790019
rect 70000 789895 70047 789951
rect 70103 789895 70171 789951
rect 70227 789895 70295 789951
rect 70351 789895 70419 789951
rect 70475 789895 70488 789951
rect 70000 789828 70488 789895
rect 705512 791687 706000 791728
rect 705512 791631 705525 791687
rect 705581 791631 705649 791687
rect 705705 791631 705773 791687
rect 705829 791631 705897 791687
rect 705953 791631 706000 791687
rect 705512 791563 706000 791631
rect 705512 791507 705525 791563
rect 705581 791507 705649 791563
rect 705705 791507 705773 791563
rect 705829 791507 705897 791563
rect 705953 791507 706000 791563
rect 705512 791439 706000 791507
rect 705512 791383 705525 791439
rect 705581 791383 705649 791439
rect 705705 791383 705773 791439
rect 705829 791383 705897 791439
rect 705953 791383 706000 791439
rect 705512 791315 706000 791383
rect 705512 791259 705525 791315
rect 705581 791259 705649 791315
rect 705705 791259 705773 791315
rect 705829 791259 705897 791315
rect 705953 791259 706000 791315
rect 705512 791191 706000 791259
rect 705512 791135 705525 791191
rect 705581 791135 705649 791191
rect 705705 791135 705773 791191
rect 705829 791135 705897 791191
rect 705953 791135 706000 791191
rect 705512 791067 706000 791135
rect 705512 791011 705525 791067
rect 705581 791011 705649 791067
rect 705705 791011 705773 791067
rect 705829 791011 705897 791067
rect 705953 791011 706000 791067
rect 705512 790943 706000 791011
rect 705512 790887 705525 790943
rect 705581 790887 705649 790943
rect 705705 790887 705773 790943
rect 705829 790887 705897 790943
rect 705953 790887 706000 790943
rect 705512 790819 706000 790887
rect 705512 790763 705525 790819
rect 705581 790763 705649 790819
rect 705705 790763 705773 790819
rect 705829 790763 705897 790819
rect 705953 790763 706000 790819
rect 705512 790695 706000 790763
rect 705512 790639 705525 790695
rect 705581 790639 705649 790695
rect 705705 790639 705773 790695
rect 705829 790639 705897 790695
rect 705953 790639 706000 790695
rect 705512 790571 706000 790639
rect 705512 790515 705525 790571
rect 705581 790515 705649 790571
rect 705705 790515 705773 790571
rect 705829 790515 705897 790571
rect 705953 790515 706000 790571
rect 705512 790447 706000 790515
rect 705512 790391 705525 790447
rect 705581 790391 705649 790447
rect 705705 790391 705773 790447
rect 705829 790391 705897 790447
rect 705953 790391 706000 790447
rect 705512 790323 706000 790391
rect 705512 790267 705525 790323
rect 705581 790267 705649 790323
rect 705705 790267 705773 790323
rect 705829 790267 705897 790323
rect 705953 790267 706000 790323
rect 705512 790199 706000 790267
rect 705512 790143 705525 790199
rect 705581 790143 705649 790199
rect 705705 790143 705773 790199
rect 705829 790143 705897 790199
rect 705953 790143 706000 790199
rect 705512 790075 706000 790143
rect 705512 790019 705525 790075
rect 705581 790019 705649 790075
rect 705705 790019 705773 790075
rect 705829 790019 705897 790075
rect 705953 790019 706000 790075
rect 705512 789951 706000 790019
rect 705512 789895 705525 789951
rect 705581 789895 705649 789951
rect 705705 789895 705773 789951
rect 705829 789895 705897 789951
rect 705953 789895 706000 789951
rect 705512 789828 706000 789895
rect 705512 789181 706000 789248
rect 70000 789105 70488 789172
rect 70000 789049 70047 789105
rect 70103 789049 70171 789105
rect 70227 789049 70295 789105
rect 70351 789049 70419 789105
rect 70475 789049 70488 789105
rect 70000 788981 70488 789049
rect 70000 788925 70047 788981
rect 70103 788925 70171 788981
rect 70227 788925 70295 788981
rect 70351 788925 70419 788981
rect 70475 788925 70488 788981
rect 70000 788857 70488 788925
rect 70000 788801 70047 788857
rect 70103 788801 70171 788857
rect 70227 788801 70295 788857
rect 70351 788801 70419 788857
rect 70475 788801 70488 788857
rect 70000 788733 70488 788801
rect 70000 788677 70047 788733
rect 70103 788677 70171 788733
rect 70227 788677 70295 788733
rect 70351 788677 70419 788733
rect 70475 788677 70488 788733
rect 70000 788609 70488 788677
rect 70000 788553 70047 788609
rect 70103 788553 70171 788609
rect 70227 788553 70295 788609
rect 70351 788553 70419 788609
rect 70475 788553 70488 788609
rect 70000 788485 70488 788553
rect 70000 788429 70047 788485
rect 70103 788429 70171 788485
rect 70227 788429 70295 788485
rect 70351 788429 70419 788485
rect 70475 788429 70488 788485
rect 70000 788361 70488 788429
rect 70000 788305 70047 788361
rect 70103 788305 70171 788361
rect 70227 788305 70295 788361
rect 70351 788305 70419 788361
rect 70475 788305 70488 788361
rect 70000 788237 70488 788305
rect 70000 788181 70047 788237
rect 70103 788181 70171 788237
rect 70227 788181 70295 788237
rect 70351 788181 70419 788237
rect 70475 788181 70488 788237
rect 70000 788113 70488 788181
rect 70000 788057 70047 788113
rect 70103 788057 70171 788113
rect 70227 788057 70295 788113
rect 70351 788057 70419 788113
rect 70475 788057 70488 788113
rect 70000 787989 70488 788057
rect 70000 787933 70047 787989
rect 70103 787933 70171 787989
rect 70227 787933 70295 787989
rect 70351 787933 70419 787989
rect 70475 787933 70488 787989
rect 70000 787865 70488 787933
rect 70000 787809 70047 787865
rect 70103 787809 70171 787865
rect 70227 787809 70295 787865
rect 70351 787809 70419 787865
rect 70475 787809 70488 787865
rect 70000 787741 70488 787809
rect 70000 787685 70047 787741
rect 70103 787685 70171 787741
rect 70227 787685 70295 787741
rect 70351 787685 70419 787741
rect 70475 787685 70488 787741
rect 70000 787617 70488 787685
rect 70000 787561 70047 787617
rect 70103 787561 70171 787617
rect 70227 787561 70295 787617
rect 70351 787561 70419 787617
rect 70475 787561 70488 787617
rect 70000 787493 70488 787561
rect 70000 787437 70047 787493
rect 70103 787437 70171 787493
rect 70227 787437 70295 787493
rect 70351 787437 70419 787493
rect 70475 787437 70488 787493
rect 70000 787369 70488 787437
rect 70000 787313 70047 787369
rect 70103 787313 70171 787369
rect 70227 787313 70295 787369
rect 70351 787313 70419 787369
rect 70475 787313 70488 787369
rect 70000 787245 70488 787313
rect 70000 787189 70047 787245
rect 70103 787189 70171 787245
rect 70227 787189 70295 787245
rect 70351 787189 70419 787245
rect 70475 787189 70488 787245
rect 705512 789125 705525 789181
rect 705581 789125 705649 789181
rect 705705 789125 705773 789181
rect 705829 789125 705897 789181
rect 705953 789125 706000 789181
rect 705512 789057 706000 789125
rect 705512 789001 705525 789057
rect 705581 789001 705649 789057
rect 705705 789001 705773 789057
rect 705829 789001 705897 789057
rect 705953 789001 706000 789057
rect 705512 788933 706000 789001
rect 705512 788877 705525 788933
rect 705581 788877 705649 788933
rect 705705 788877 705773 788933
rect 705829 788877 705897 788933
rect 705953 788877 706000 788933
rect 705512 788809 706000 788877
rect 705512 788753 705525 788809
rect 705581 788753 705649 788809
rect 705705 788753 705773 788809
rect 705829 788753 705897 788809
rect 705953 788753 706000 788809
rect 705512 788685 706000 788753
rect 705512 788629 705525 788685
rect 705581 788629 705649 788685
rect 705705 788629 705773 788685
rect 705829 788629 705897 788685
rect 705953 788629 706000 788685
rect 705512 788561 706000 788629
rect 705512 788505 705525 788561
rect 705581 788505 705649 788561
rect 705705 788505 705773 788561
rect 705829 788505 705897 788561
rect 705953 788505 706000 788561
rect 705512 788437 706000 788505
rect 705512 788381 705525 788437
rect 705581 788381 705649 788437
rect 705705 788381 705773 788437
rect 705829 788381 705897 788437
rect 705953 788381 706000 788437
rect 705512 788313 706000 788381
rect 705512 788257 705525 788313
rect 705581 788257 705649 788313
rect 705705 788257 705773 788313
rect 705829 788257 705897 788313
rect 705953 788257 706000 788313
rect 705512 788189 706000 788257
rect 705512 788133 705525 788189
rect 705581 788133 705649 788189
rect 705705 788133 705773 788189
rect 705829 788133 705897 788189
rect 705953 788133 706000 788189
rect 705512 788065 706000 788133
rect 705512 788009 705525 788065
rect 705581 788009 705649 788065
rect 705705 788009 705773 788065
rect 705829 788009 705897 788065
rect 705953 788009 706000 788065
rect 705512 787941 706000 788009
rect 705512 787885 705525 787941
rect 705581 787885 705649 787941
rect 705705 787885 705773 787941
rect 705829 787885 705897 787941
rect 705953 787885 706000 787941
rect 705512 787817 706000 787885
rect 705512 787761 705525 787817
rect 705581 787761 705649 787817
rect 705705 787761 705773 787817
rect 705829 787761 705897 787817
rect 705953 787761 706000 787817
rect 705512 787693 706000 787761
rect 705512 787637 705525 787693
rect 705581 787637 705649 787693
rect 705705 787637 705773 787693
rect 705829 787637 705897 787693
rect 705953 787637 706000 787693
rect 705512 787569 706000 787637
rect 705512 787513 705525 787569
rect 705581 787513 705649 787569
rect 705705 787513 705773 787569
rect 705829 787513 705897 787569
rect 705953 787513 706000 787569
rect 705512 787445 706000 787513
rect 705512 787389 705525 787445
rect 705581 787389 705649 787445
rect 705705 787389 705773 787445
rect 705829 787389 705897 787445
rect 705953 787389 706000 787445
rect 705512 787321 706000 787389
rect 705512 787265 705525 787321
rect 705581 787265 705649 787321
rect 705705 787265 705773 787321
rect 705829 787265 705897 787321
rect 705953 787265 706000 787321
rect 705512 787198 706000 787265
rect 70000 787122 70488 787189
rect 705512 786811 706000 786878
rect 70000 786735 70488 786802
rect 70000 786679 70047 786735
rect 70103 786679 70171 786735
rect 70227 786679 70295 786735
rect 70351 786679 70419 786735
rect 70475 786679 70488 786735
rect 70000 786611 70488 786679
rect 70000 786555 70047 786611
rect 70103 786555 70171 786611
rect 70227 786555 70295 786611
rect 70351 786555 70419 786611
rect 70475 786555 70488 786611
rect 70000 786487 70488 786555
rect 70000 786431 70047 786487
rect 70103 786431 70171 786487
rect 70227 786431 70295 786487
rect 70351 786431 70419 786487
rect 70475 786431 70488 786487
rect 70000 786363 70488 786431
rect 70000 786307 70047 786363
rect 70103 786307 70171 786363
rect 70227 786307 70295 786363
rect 70351 786307 70419 786363
rect 70475 786307 70488 786363
rect 70000 786239 70488 786307
rect 70000 786183 70047 786239
rect 70103 786183 70171 786239
rect 70227 786183 70295 786239
rect 70351 786183 70419 786239
rect 70475 786183 70488 786239
rect 70000 786115 70488 786183
rect 70000 786059 70047 786115
rect 70103 786059 70171 786115
rect 70227 786059 70295 786115
rect 70351 786059 70419 786115
rect 70475 786059 70488 786115
rect 70000 785991 70488 786059
rect 70000 785935 70047 785991
rect 70103 785935 70171 785991
rect 70227 785935 70295 785991
rect 70351 785935 70419 785991
rect 70475 785935 70488 785991
rect 70000 785867 70488 785935
rect 70000 785811 70047 785867
rect 70103 785811 70171 785867
rect 70227 785811 70295 785867
rect 70351 785811 70419 785867
rect 70475 785811 70488 785867
rect 70000 785743 70488 785811
rect 70000 785687 70047 785743
rect 70103 785687 70171 785743
rect 70227 785687 70295 785743
rect 70351 785687 70419 785743
rect 70475 785687 70488 785743
rect 70000 785619 70488 785687
rect 70000 785563 70047 785619
rect 70103 785563 70171 785619
rect 70227 785563 70295 785619
rect 70351 785563 70419 785619
rect 70475 785563 70488 785619
rect 70000 785495 70488 785563
rect 70000 785439 70047 785495
rect 70103 785439 70171 785495
rect 70227 785439 70295 785495
rect 70351 785439 70419 785495
rect 70475 785439 70488 785495
rect 70000 785371 70488 785439
rect 70000 785315 70047 785371
rect 70103 785315 70171 785371
rect 70227 785315 70295 785371
rect 70351 785315 70419 785371
rect 70475 785315 70488 785371
rect 70000 785247 70488 785315
rect 70000 785191 70047 785247
rect 70103 785191 70171 785247
rect 70227 785191 70295 785247
rect 70351 785191 70419 785247
rect 70475 785191 70488 785247
rect 70000 785123 70488 785191
rect 70000 785067 70047 785123
rect 70103 785067 70171 785123
rect 70227 785067 70295 785123
rect 70351 785067 70419 785123
rect 70475 785067 70488 785123
rect 70000 784999 70488 785067
rect 70000 784943 70047 784999
rect 70103 784943 70171 784999
rect 70227 784943 70295 784999
rect 70351 784943 70419 784999
rect 70475 784943 70488 784999
rect 70000 784875 70488 784943
rect 70000 784819 70047 784875
rect 70103 784819 70171 784875
rect 70227 784819 70295 784875
rect 70351 784819 70419 784875
rect 70475 784819 70488 784875
rect 705512 786755 705525 786811
rect 705581 786755 705649 786811
rect 705705 786755 705773 786811
rect 705829 786755 705897 786811
rect 705953 786755 706000 786811
rect 705512 786687 706000 786755
rect 705512 786631 705525 786687
rect 705581 786631 705649 786687
rect 705705 786631 705773 786687
rect 705829 786631 705897 786687
rect 705953 786631 706000 786687
rect 705512 786563 706000 786631
rect 705512 786507 705525 786563
rect 705581 786507 705649 786563
rect 705705 786507 705773 786563
rect 705829 786507 705897 786563
rect 705953 786507 706000 786563
rect 705512 786439 706000 786507
rect 705512 786383 705525 786439
rect 705581 786383 705649 786439
rect 705705 786383 705773 786439
rect 705829 786383 705897 786439
rect 705953 786383 706000 786439
rect 705512 786315 706000 786383
rect 705512 786259 705525 786315
rect 705581 786259 705649 786315
rect 705705 786259 705773 786315
rect 705829 786259 705897 786315
rect 705953 786259 706000 786315
rect 705512 786191 706000 786259
rect 705512 786135 705525 786191
rect 705581 786135 705649 786191
rect 705705 786135 705773 786191
rect 705829 786135 705897 786191
rect 705953 786135 706000 786191
rect 705512 786067 706000 786135
rect 705512 786011 705525 786067
rect 705581 786011 705649 786067
rect 705705 786011 705773 786067
rect 705829 786011 705897 786067
rect 705953 786011 706000 786067
rect 705512 785943 706000 786011
rect 705512 785887 705525 785943
rect 705581 785887 705649 785943
rect 705705 785887 705773 785943
rect 705829 785887 705897 785943
rect 705953 785887 706000 785943
rect 705512 785819 706000 785887
rect 705512 785763 705525 785819
rect 705581 785763 705649 785819
rect 705705 785763 705773 785819
rect 705829 785763 705897 785819
rect 705953 785763 706000 785819
rect 705512 785695 706000 785763
rect 705512 785639 705525 785695
rect 705581 785639 705649 785695
rect 705705 785639 705773 785695
rect 705829 785639 705897 785695
rect 705953 785639 706000 785695
rect 705512 785571 706000 785639
rect 705512 785515 705525 785571
rect 705581 785515 705649 785571
rect 705705 785515 705773 785571
rect 705829 785515 705897 785571
rect 705953 785515 706000 785571
rect 705512 785447 706000 785515
rect 705512 785391 705525 785447
rect 705581 785391 705649 785447
rect 705705 785391 705773 785447
rect 705829 785391 705897 785447
rect 705953 785391 706000 785447
rect 705512 785323 706000 785391
rect 705512 785267 705525 785323
rect 705581 785267 705649 785323
rect 705705 785267 705773 785323
rect 705829 785267 705897 785323
rect 705953 785267 706000 785323
rect 705512 785199 706000 785267
rect 705512 785143 705525 785199
rect 705581 785143 705649 785199
rect 705705 785143 705773 785199
rect 705829 785143 705897 785199
rect 705953 785143 706000 785199
rect 705512 785075 706000 785143
rect 705512 785019 705525 785075
rect 705581 785019 705649 785075
rect 705705 785019 705773 785075
rect 705829 785019 705897 785075
rect 705953 785019 706000 785075
rect 705512 784951 706000 785019
rect 705512 784895 705525 784951
rect 705581 784895 705649 784951
rect 705705 784895 705773 784951
rect 705829 784895 705897 784951
rect 705953 784895 706000 784951
rect 705512 784828 706000 784895
rect 70000 784752 70488 784819
rect 70000 784105 70488 784172
rect 70000 784049 70047 784105
rect 70103 784049 70171 784105
rect 70227 784049 70295 784105
rect 70351 784049 70419 784105
rect 70475 784049 70488 784105
rect 70000 783981 70488 784049
rect 70000 783925 70047 783981
rect 70103 783925 70171 783981
rect 70227 783925 70295 783981
rect 70351 783925 70419 783981
rect 70475 783925 70488 783981
rect 70000 783857 70488 783925
rect 70000 783801 70047 783857
rect 70103 783801 70171 783857
rect 70227 783801 70295 783857
rect 70351 783801 70419 783857
rect 70475 783801 70488 783857
rect 70000 783733 70488 783801
rect 70000 783677 70047 783733
rect 70103 783677 70171 783733
rect 70227 783677 70295 783733
rect 70351 783677 70419 783733
rect 70475 783677 70488 783733
rect 70000 783609 70488 783677
rect 70000 783553 70047 783609
rect 70103 783553 70171 783609
rect 70227 783553 70295 783609
rect 70351 783553 70419 783609
rect 70475 783553 70488 783609
rect 70000 783485 70488 783553
rect 70000 783429 70047 783485
rect 70103 783429 70171 783485
rect 70227 783429 70295 783485
rect 70351 783429 70419 783485
rect 70475 783429 70488 783485
rect 70000 783361 70488 783429
rect 70000 783305 70047 783361
rect 70103 783305 70171 783361
rect 70227 783305 70295 783361
rect 70351 783305 70419 783361
rect 70475 783305 70488 783361
rect 70000 783237 70488 783305
rect 70000 783181 70047 783237
rect 70103 783181 70171 783237
rect 70227 783181 70295 783237
rect 70351 783181 70419 783237
rect 70475 783181 70488 783237
rect 70000 783113 70488 783181
rect 70000 783057 70047 783113
rect 70103 783057 70171 783113
rect 70227 783057 70295 783113
rect 70351 783057 70419 783113
rect 70475 783057 70488 783113
rect 70000 782989 70488 783057
rect 70000 782933 70047 782989
rect 70103 782933 70171 782989
rect 70227 782933 70295 782989
rect 70351 782933 70419 782989
rect 70475 782933 70488 782989
rect 70000 782865 70488 782933
rect 70000 782809 70047 782865
rect 70103 782809 70171 782865
rect 70227 782809 70295 782865
rect 70351 782809 70419 782865
rect 70475 782809 70488 782865
rect 70000 782741 70488 782809
rect 70000 782685 70047 782741
rect 70103 782685 70171 782741
rect 70227 782685 70295 782741
rect 70351 782685 70419 782741
rect 70475 782685 70488 782741
rect 70000 782617 70488 782685
rect 70000 782561 70047 782617
rect 70103 782561 70171 782617
rect 70227 782561 70295 782617
rect 70351 782561 70419 782617
rect 70475 782561 70488 782617
rect 70000 782493 70488 782561
rect 70000 782437 70047 782493
rect 70103 782437 70171 782493
rect 70227 782437 70295 782493
rect 70351 782437 70419 782493
rect 70475 782437 70488 782493
rect 70000 782369 70488 782437
rect 70000 782313 70047 782369
rect 70103 782313 70171 782369
rect 70227 782313 70295 782369
rect 70351 782313 70419 782369
rect 70475 782313 70488 782369
rect 70000 782272 70488 782313
rect 705512 784105 706000 784172
rect 705512 784049 705525 784105
rect 705581 784049 705649 784105
rect 705705 784049 705773 784105
rect 705829 784049 705897 784105
rect 705953 784049 706000 784105
rect 705512 783981 706000 784049
rect 705512 783925 705525 783981
rect 705581 783925 705649 783981
rect 705705 783925 705773 783981
rect 705829 783925 705897 783981
rect 705953 783925 706000 783981
rect 705512 783857 706000 783925
rect 705512 783801 705525 783857
rect 705581 783801 705649 783857
rect 705705 783801 705773 783857
rect 705829 783801 705897 783857
rect 705953 783801 706000 783857
rect 705512 783733 706000 783801
rect 705512 783677 705525 783733
rect 705581 783677 705649 783733
rect 705705 783677 705773 783733
rect 705829 783677 705897 783733
rect 705953 783677 706000 783733
rect 705512 783609 706000 783677
rect 705512 783553 705525 783609
rect 705581 783553 705649 783609
rect 705705 783553 705773 783609
rect 705829 783553 705897 783609
rect 705953 783553 706000 783609
rect 705512 783485 706000 783553
rect 705512 783429 705525 783485
rect 705581 783429 705649 783485
rect 705705 783429 705773 783485
rect 705829 783429 705897 783485
rect 705953 783429 706000 783485
rect 705512 783361 706000 783429
rect 705512 783305 705525 783361
rect 705581 783305 705649 783361
rect 705705 783305 705773 783361
rect 705829 783305 705897 783361
rect 705953 783305 706000 783361
rect 705512 783237 706000 783305
rect 705512 783181 705525 783237
rect 705581 783181 705649 783237
rect 705705 783181 705773 783237
rect 705829 783181 705897 783237
rect 705953 783181 706000 783237
rect 705512 783113 706000 783181
rect 705512 783057 705525 783113
rect 705581 783057 705649 783113
rect 705705 783057 705773 783113
rect 705829 783057 705897 783113
rect 705953 783057 706000 783113
rect 705512 782989 706000 783057
rect 705512 782933 705525 782989
rect 705581 782933 705649 782989
rect 705705 782933 705773 782989
rect 705829 782933 705897 782989
rect 705953 782933 706000 782989
rect 705512 782865 706000 782933
rect 705512 782809 705525 782865
rect 705581 782809 705649 782865
rect 705705 782809 705773 782865
rect 705829 782809 705897 782865
rect 705953 782809 706000 782865
rect 705512 782741 706000 782809
rect 705512 782685 705525 782741
rect 705581 782685 705649 782741
rect 705705 782685 705773 782741
rect 705829 782685 705897 782741
rect 705953 782685 706000 782741
rect 705512 782617 706000 782685
rect 705512 782561 705525 782617
rect 705581 782561 705649 782617
rect 705705 782561 705773 782617
rect 705829 782561 705897 782617
rect 705953 782561 706000 782617
rect 705512 782493 706000 782561
rect 705512 782437 705525 782493
rect 705581 782437 705649 782493
rect 705705 782437 705773 782493
rect 705829 782437 705897 782493
rect 705953 782437 706000 782493
rect 705512 782369 706000 782437
rect 705512 782313 705525 782369
rect 705581 782313 705649 782369
rect 705705 782313 705773 782369
rect 705829 782313 705897 782369
rect 705953 782313 706000 782369
rect 705512 782245 706000 782313
rect 705512 782189 705525 782245
rect 705581 782189 705649 782245
rect 705705 782189 705773 782245
rect 705829 782189 705897 782245
rect 705953 782189 706000 782245
rect 705512 782122 706000 782189
rect 705512 781735 706000 781802
rect 705512 781679 705525 781735
rect 705581 781679 705649 781735
rect 705705 781679 705773 781735
rect 705829 781679 705897 781735
rect 705953 781679 706000 781735
rect 705512 781611 706000 781679
rect 705512 781555 705525 781611
rect 705581 781555 705649 781611
rect 705705 781555 705773 781611
rect 705829 781555 705897 781611
rect 705953 781555 706000 781611
rect 705512 781487 706000 781555
rect 705512 781431 705525 781487
rect 705581 781431 705649 781487
rect 705705 781431 705773 781487
rect 705829 781431 705897 781487
rect 705953 781431 706000 781487
rect 705512 781363 706000 781431
rect 705512 781307 705525 781363
rect 705581 781307 705649 781363
rect 705705 781307 705773 781363
rect 705829 781307 705897 781363
rect 705953 781307 706000 781363
rect 705512 781239 706000 781307
rect 705512 781183 705525 781239
rect 705581 781183 705649 781239
rect 705705 781183 705773 781239
rect 705829 781183 705897 781239
rect 705953 781183 706000 781239
rect 705512 781115 706000 781183
rect 705512 781059 705525 781115
rect 705581 781059 705649 781115
rect 705705 781059 705773 781115
rect 705829 781059 705897 781115
rect 705953 781059 706000 781115
rect 705512 780991 706000 781059
rect 705512 780935 705525 780991
rect 705581 780935 705649 780991
rect 705705 780935 705773 780991
rect 705829 780935 705897 780991
rect 705953 780935 706000 780991
rect 705512 780867 706000 780935
rect 705512 780811 705525 780867
rect 705581 780811 705649 780867
rect 705705 780811 705773 780867
rect 705829 780811 705897 780867
rect 705953 780811 706000 780867
rect 705512 780743 706000 780811
rect 705512 780687 705525 780743
rect 705581 780687 705649 780743
rect 705705 780687 705773 780743
rect 705829 780687 705897 780743
rect 705953 780687 706000 780743
rect 705512 780619 706000 780687
rect 705512 780563 705525 780619
rect 705581 780563 705649 780619
rect 705705 780563 705773 780619
rect 705829 780563 705897 780619
rect 705953 780563 706000 780619
rect 705512 780495 706000 780563
rect 705512 780439 705525 780495
rect 705581 780439 705649 780495
rect 705705 780439 705773 780495
rect 705829 780439 705897 780495
rect 705953 780439 706000 780495
rect 705512 780371 706000 780439
rect 705512 780315 705525 780371
rect 705581 780315 705649 780371
rect 705705 780315 705773 780371
rect 705829 780315 705897 780371
rect 705953 780315 706000 780371
rect 705512 780247 706000 780315
rect 705512 780191 705525 780247
rect 705581 780191 705649 780247
rect 705705 780191 705773 780247
rect 705829 780191 705897 780247
rect 705953 780191 706000 780247
rect 705512 780123 706000 780191
rect 705512 780067 705525 780123
rect 705581 780067 705649 780123
rect 705705 780067 705773 780123
rect 705829 780067 705897 780123
rect 705953 780067 706000 780123
rect 705512 779999 706000 780067
rect 705512 779943 705525 779999
rect 705581 779943 705649 779999
rect 705705 779943 705773 779999
rect 705829 779943 705897 779999
rect 705953 779943 706000 779999
rect 705512 779875 706000 779943
rect 705512 779819 705525 779875
rect 705581 779819 705649 779875
rect 705705 779819 705773 779875
rect 705829 779819 705897 779875
rect 705953 779819 706000 779875
rect 705512 779752 706000 779819
rect 705512 779131 706000 779172
rect 705512 779075 705525 779131
rect 705581 779075 705649 779131
rect 705705 779075 705773 779131
rect 705829 779075 705897 779131
rect 705953 779075 706000 779131
rect 705512 779007 706000 779075
rect 705512 778951 705525 779007
rect 705581 778951 705649 779007
rect 705705 778951 705773 779007
rect 705829 778951 705897 779007
rect 705953 778951 706000 779007
rect 705512 778883 706000 778951
rect 705512 778827 705525 778883
rect 705581 778827 705649 778883
rect 705705 778827 705773 778883
rect 705829 778827 705897 778883
rect 705953 778827 706000 778883
rect 705512 778759 706000 778827
rect 705512 778703 705525 778759
rect 705581 778703 705649 778759
rect 705705 778703 705773 778759
rect 705829 778703 705897 778759
rect 705953 778703 706000 778759
rect 705512 778635 706000 778703
rect 705512 778579 705525 778635
rect 705581 778579 705649 778635
rect 705705 778579 705773 778635
rect 705829 778579 705897 778635
rect 705953 778579 706000 778635
rect 705512 778511 706000 778579
rect 705512 778455 705525 778511
rect 705581 778455 705649 778511
rect 705705 778455 705773 778511
rect 705829 778455 705897 778511
rect 705953 778455 706000 778511
rect 705512 778387 706000 778455
rect 705512 778331 705525 778387
rect 705581 778331 705649 778387
rect 705705 778331 705773 778387
rect 705829 778331 705897 778387
rect 705953 778331 706000 778387
rect 705512 778263 706000 778331
rect 705512 778207 705525 778263
rect 705581 778207 705649 778263
rect 705705 778207 705773 778263
rect 705829 778207 705897 778263
rect 705953 778207 706000 778263
rect 705512 778139 706000 778207
rect 705512 778083 705525 778139
rect 705581 778083 705649 778139
rect 705705 778083 705773 778139
rect 705829 778083 705897 778139
rect 705953 778083 706000 778139
rect 705512 778015 706000 778083
rect 705512 777959 705525 778015
rect 705581 777959 705649 778015
rect 705705 777959 705773 778015
rect 705829 777959 705897 778015
rect 705953 777959 706000 778015
rect 705512 777891 706000 777959
rect 705512 777835 705525 777891
rect 705581 777835 705649 777891
rect 705705 777835 705773 777891
rect 705829 777835 705897 777891
rect 705953 777835 706000 777891
rect 705512 777767 706000 777835
rect 705512 777711 705525 777767
rect 705581 777711 705649 777767
rect 705705 777711 705773 777767
rect 705829 777711 705897 777767
rect 705953 777711 706000 777767
rect 705512 777643 706000 777711
rect 705512 777587 705525 777643
rect 705581 777587 705649 777643
rect 705705 777587 705773 777643
rect 705829 777587 705897 777643
rect 705953 777587 706000 777643
rect 705512 777519 706000 777587
rect 705512 777463 705525 777519
rect 705581 777463 705649 777519
rect 705705 777463 705773 777519
rect 705829 777463 705897 777519
rect 705953 777463 706000 777519
rect 705512 777395 706000 777463
rect 705512 777339 705525 777395
rect 705581 777339 705649 777395
rect 705705 777339 705773 777395
rect 705829 777339 705897 777395
rect 705953 777339 706000 777395
rect 705512 777272 706000 777339
rect 705512 490687 706000 490728
rect 705512 490631 705525 490687
rect 705581 490631 705649 490687
rect 705705 490631 705773 490687
rect 705829 490631 705897 490687
rect 705953 490631 706000 490687
rect 705512 490563 706000 490631
rect 705512 490507 705525 490563
rect 705581 490507 705649 490563
rect 705705 490507 705773 490563
rect 705829 490507 705897 490563
rect 705953 490507 706000 490563
rect 705512 490439 706000 490507
rect 705512 490383 705525 490439
rect 705581 490383 705649 490439
rect 705705 490383 705773 490439
rect 705829 490383 705897 490439
rect 705953 490383 706000 490439
rect 705512 490315 706000 490383
rect 705512 490259 705525 490315
rect 705581 490259 705649 490315
rect 705705 490259 705773 490315
rect 705829 490259 705897 490315
rect 705953 490259 706000 490315
rect 705512 490191 706000 490259
rect 705512 490135 705525 490191
rect 705581 490135 705649 490191
rect 705705 490135 705773 490191
rect 705829 490135 705897 490191
rect 705953 490135 706000 490191
rect 705512 490067 706000 490135
rect 705512 490011 705525 490067
rect 705581 490011 705649 490067
rect 705705 490011 705773 490067
rect 705829 490011 705897 490067
rect 705953 490011 706000 490067
rect 705512 489943 706000 490011
rect 705512 489887 705525 489943
rect 705581 489887 705649 489943
rect 705705 489887 705773 489943
rect 705829 489887 705897 489943
rect 705953 489887 706000 489943
rect 705512 489819 706000 489887
rect 705512 489763 705525 489819
rect 705581 489763 705649 489819
rect 705705 489763 705773 489819
rect 705829 489763 705897 489819
rect 705953 489763 706000 489819
rect 705512 489695 706000 489763
rect 705512 489639 705525 489695
rect 705581 489639 705649 489695
rect 705705 489639 705773 489695
rect 705829 489639 705897 489695
rect 705953 489639 706000 489695
rect 705512 489571 706000 489639
rect 705512 489515 705525 489571
rect 705581 489515 705649 489571
rect 705705 489515 705773 489571
rect 705829 489515 705897 489571
rect 705953 489515 706000 489571
rect 705512 489447 706000 489515
rect 705512 489391 705525 489447
rect 705581 489391 705649 489447
rect 705705 489391 705773 489447
rect 705829 489391 705897 489447
rect 705953 489391 706000 489447
rect 705512 489323 706000 489391
rect 705512 489267 705525 489323
rect 705581 489267 705649 489323
rect 705705 489267 705773 489323
rect 705829 489267 705897 489323
rect 705953 489267 706000 489323
rect 705512 489199 706000 489267
rect 705512 489143 705525 489199
rect 705581 489143 705649 489199
rect 705705 489143 705773 489199
rect 705829 489143 705897 489199
rect 705953 489143 706000 489199
rect 705512 489075 706000 489143
rect 705512 489019 705525 489075
rect 705581 489019 705649 489075
rect 705705 489019 705773 489075
rect 705829 489019 705897 489075
rect 705953 489019 706000 489075
rect 705512 488951 706000 489019
rect 705512 488895 705525 488951
rect 705581 488895 705649 488951
rect 705705 488895 705773 488951
rect 705829 488895 705897 488951
rect 705953 488895 706000 488951
rect 705512 488828 706000 488895
rect 705512 488181 706000 488248
rect 705512 488125 705525 488181
rect 705581 488125 705649 488181
rect 705705 488125 705773 488181
rect 705829 488125 705897 488181
rect 705953 488125 706000 488181
rect 705512 488057 706000 488125
rect 705512 488001 705525 488057
rect 705581 488001 705649 488057
rect 705705 488001 705773 488057
rect 705829 488001 705897 488057
rect 705953 488001 706000 488057
rect 705512 487933 706000 488001
rect 705512 487877 705525 487933
rect 705581 487877 705649 487933
rect 705705 487877 705773 487933
rect 705829 487877 705897 487933
rect 705953 487877 706000 487933
rect 705512 487809 706000 487877
rect 705512 487753 705525 487809
rect 705581 487753 705649 487809
rect 705705 487753 705773 487809
rect 705829 487753 705897 487809
rect 705953 487753 706000 487809
rect 705512 487685 706000 487753
rect 705512 487629 705525 487685
rect 705581 487629 705649 487685
rect 705705 487629 705773 487685
rect 705829 487629 705897 487685
rect 705953 487629 706000 487685
rect 705512 487561 706000 487629
rect 705512 487505 705525 487561
rect 705581 487505 705649 487561
rect 705705 487505 705773 487561
rect 705829 487505 705897 487561
rect 705953 487505 706000 487561
rect 705512 487437 706000 487505
rect 705512 487381 705525 487437
rect 705581 487381 705649 487437
rect 705705 487381 705773 487437
rect 705829 487381 705897 487437
rect 705953 487381 706000 487437
rect 705512 487313 706000 487381
rect 705512 487257 705525 487313
rect 705581 487257 705649 487313
rect 705705 487257 705773 487313
rect 705829 487257 705897 487313
rect 705953 487257 706000 487313
rect 705512 487189 706000 487257
rect 705512 487133 705525 487189
rect 705581 487133 705649 487189
rect 705705 487133 705773 487189
rect 705829 487133 705897 487189
rect 705953 487133 706000 487189
rect 705512 487065 706000 487133
rect 705512 487009 705525 487065
rect 705581 487009 705649 487065
rect 705705 487009 705773 487065
rect 705829 487009 705897 487065
rect 705953 487009 706000 487065
rect 705512 486941 706000 487009
rect 705512 486885 705525 486941
rect 705581 486885 705649 486941
rect 705705 486885 705773 486941
rect 705829 486885 705897 486941
rect 705953 486885 706000 486941
rect 705512 486817 706000 486885
rect 705512 486761 705525 486817
rect 705581 486761 705649 486817
rect 705705 486761 705773 486817
rect 705829 486761 705897 486817
rect 705953 486761 706000 486817
rect 705512 486693 706000 486761
rect 705512 486637 705525 486693
rect 705581 486637 705649 486693
rect 705705 486637 705773 486693
rect 705829 486637 705897 486693
rect 705953 486637 706000 486693
rect 705512 486569 706000 486637
rect 705512 486513 705525 486569
rect 705581 486513 705649 486569
rect 705705 486513 705773 486569
rect 705829 486513 705897 486569
rect 705953 486513 706000 486569
rect 705512 486445 706000 486513
rect 705512 486389 705525 486445
rect 705581 486389 705649 486445
rect 705705 486389 705773 486445
rect 705829 486389 705897 486445
rect 705953 486389 706000 486445
rect 705512 486321 706000 486389
rect 705512 486265 705525 486321
rect 705581 486265 705649 486321
rect 705705 486265 705773 486321
rect 705829 486265 705897 486321
rect 705953 486265 706000 486321
rect 705512 486198 706000 486265
rect 705512 485811 706000 485878
rect 705512 485755 705525 485811
rect 705581 485755 705649 485811
rect 705705 485755 705773 485811
rect 705829 485755 705897 485811
rect 705953 485755 706000 485811
rect 705512 485687 706000 485755
rect 705512 485631 705525 485687
rect 705581 485631 705649 485687
rect 705705 485631 705773 485687
rect 705829 485631 705897 485687
rect 705953 485631 706000 485687
rect 705512 485563 706000 485631
rect 705512 485507 705525 485563
rect 705581 485507 705649 485563
rect 705705 485507 705773 485563
rect 705829 485507 705897 485563
rect 705953 485507 706000 485563
rect 705512 485439 706000 485507
rect 705512 485383 705525 485439
rect 705581 485383 705649 485439
rect 705705 485383 705773 485439
rect 705829 485383 705897 485439
rect 705953 485383 706000 485439
rect 705512 485315 706000 485383
rect 705512 485259 705525 485315
rect 705581 485259 705649 485315
rect 705705 485259 705773 485315
rect 705829 485259 705897 485315
rect 705953 485259 706000 485315
rect 705512 485191 706000 485259
rect 705512 485135 705525 485191
rect 705581 485135 705649 485191
rect 705705 485135 705773 485191
rect 705829 485135 705897 485191
rect 705953 485135 706000 485191
rect 705512 485067 706000 485135
rect 705512 485011 705525 485067
rect 705581 485011 705649 485067
rect 705705 485011 705773 485067
rect 705829 485011 705897 485067
rect 705953 485011 706000 485067
rect 705512 484943 706000 485011
rect 705512 484887 705525 484943
rect 705581 484887 705649 484943
rect 705705 484887 705773 484943
rect 705829 484887 705897 484943
rect 705953 484887 706000 484943
rect 705512 484819 706000 484887
rect 705512 484763 705525 484819
rect 705581 484763 705649 484819
rect 705705 484763 705773 484819
rect 705829 484763 705897 484819
rect 705953 484763 706000 484819
rect 705512 484695 706000 484763
rect 705512 484639 705525 484695
rect 705581 484639 705649 484695
rect 705705 484639 705773 484695
rect 705829 484639 705897 484695
rect 705953 484639 706000 484695
rect 705512 484571 706000 484639
rect 705512 484515 705525 484571
rect 705581 484515 705649 484571
rect 705705 484515 705773 484571
rect 705829 484515 705897 484571
rect 705953 484515 706000 484571
rect 705512 484447 706000 484515
rect 705512 484391 705525 484447
rect 705581 484391 705649 484447
rect 705705 484391 705773 484447
rect 705829 484391 705897 484447
rect 705953 484391 706000 484447
rect 705512 484323 706000 484391
rect 705512 484267 705525 484323
rect 705581 484267 705649 484323
rect 705705 484267 705773 484323
rect 705829 484267 705897 484323
rect 705953 484267 706000 484323
rect 705512 484199 706000 484267
rect 705512 484143 705525 484199
rect 705581 484143 705649 484199
rect 705705 484143 705773 484199
rect 705829 484143 705897 484199
rect 705953 484143 706000 484199
rect 705512 484075 706000 484143
rect 705512 484019 705525 484075
rect 705581 484019 705649 484075
rect 705705 484019 705773 484075
rect 705829 484019 705897 484075
rect 705953 484019 706000 484075
rect 705512 483951 706000 484019
rect 705512 483895 705525 483951
rect 705581 483895 705649 483951
rect 705705 483895 705773 483951
rect 705829 483895 705897 483951
rect 705953 483895 706000 483951
rect 705512 483828 706000 483895
rect 705512 483105 706000 483172
rect 705512 483049 705525 483105
rect 705581 483049 705649 483105
rect 705705 483049 705773 483105
rect 705829 483049 705897 483105
rect 705953 483049 706000 483105
rect 705512 482981 706000 483049
rect 705512 482925 705525 482981
rect 705581 482925 705649 482981
rect 705705 482925 705773 482981
rect 705829 482925 705897 482981
rect 705953 482925 706000 482981
rect 705512 482857 706000 482925
rect 705512 482801 705525 482857
rect 705581 482801 705649 482857
rect 705705 482801 705773 482857
rect 705829 482801 705897 482857
rect 705953 482801 706000 482857
rect 705512 482733 706000 482801
rect 705512 482677 705525 482733
rect 705581 482677 705649 482733
rect 705705 482677 705773 482733
rect 705829 482677 705897 482733
rect 705953 482677 706000 482733
rect 705512 482609 706000 482677
rect 705512 482553 705525 482609
rect 705581 482553 705649 482609
rect 705705 482553 705773 482609
rect 705829 482553 705897 482609
rect 705953 482553 706000 482609
rect 705512 482485 706000 482553
rect 705512 482429 705525 482485
rect 705581 482429 705649 482485
rect 705705 482429 705773 482485
rect 705829 482429 705897 482485
rect 705953 482429 706000 482485
rect 705512 482361 706000 482429
rect 705512 482305 705525 482361
rect 705581 482305 705649 482361
rect 705705 482305 705773 482361
rect 705829 482305 705897 482361
rect 705953 482305 706000 482361
rect 705512 482237 706000 482305
rect 705512 482181 705525 482237
rect 705581 482181 705649 482237
rect 705705 482181 705773 482237
rect 705829 482181 705897 482237
rect 705953 482181 706000 482237
rect 705512 482113 706000 482181
rect 705512 482057 705525 482113
rect 705581 482057 705649 482113
rect 705705 482057 705773 482113
rect 705829 482057 705897 482113
rect 705953 482057 706000 482113
rect 705512 481989 706000 482057
rect 705512 481933 705525 481989
rect 705581 481933 705649 481989
rect 705705 481933 705773 481989
rect 705829 481933 705897 481989
rect 705953 481933 706000 481989
rect 705512 481865 706000 481933
rect 705512 481809 705525 481865
rect 705581 481809 705649 481865
rect 705705 481809 705773 481865
rect 705829 481809 705897 481865
rect 705953 481809 706000 481865
rect 705512 481741 706000 481809
rect 705512 481685 705525 481741
rect 705581 481685 705649 481741
rect 705705 481685 705773 481741
rect 705829 481685 705897 481741
rect 705953 481685 706000 481741
rect 705512 481617 706000 481685
rect 705512 481561 705525 481617
rect 705581 481561 705649 481617
rect 705705 481561 705773 481617
rect 705829 481561 705897 481617
rect 705953 481561 706000 481617
rect 705512 481493 706000 481561
rect 705512 481437 705525 481493
rect 705581 481437 705649 481493
rect 705705 481437 705773 481493
rect 705829 481437 705897 481493
rect 705953 481437 706000 481493
rect 705512 481369 706000 481437
rect 705512 481313 705525 481369
rect 705581 481313 705649 481369
rect 705705 481313 705773 481369
rect 705829 481313 705897 481369
rect 705953 481313 706000 481369
rect 705512 481245 706000 481313
rect 705512 481189 705525 481245
rect 705581 481189 705649 481245
rect 705705 481189 705773 481245
rect 705829 481189 705897 481245
rect 705953 481189 706000 481245
rect 705512 481122 706000 481189
rect 705512 480735 706000 480802
rect 705512 480679 705525 480735
rect 705581 480679 705649 480735
rect 705705 480679 705773 480735
rect 705829 480679 705897 480735
rect 705953 480679 706000 480735
rect 705512 480611 706000 480679
rect 705512 480555 705525 480611
rect 705581 480555 705649 480611
rect 705705 480555 705773 480611
rect 705829 480555 705897 480611
rect 705953 480555 706000 480611
rect 705512 480487 706000 480555
rect 705512 480431 705525 480487
rect 705581 480431 705649 480487
rect 705705 480431 705773 480487
rect 705829 480431 705897 480487
rect 705953 480431 706000 480487
rect 705512 480363 706000 480431
rect 705512 480307 705525 480363
rect 705581 480307 705649 480363
rect 705705 480307 705773 480363
rect 705829 480307 705897 480363
rect 705953 480307 706000 480363
rect 705512 480239 706000 480307
rect 705512 480183 705525 480239
rect 705581 480183 705649 480239
rect 705705 480183 705773 480239
rect 705829 480183 705897 480239
rect 705953 480183 706000 480239
rect 705512 480115 706000 480183
rect 705512 480059 705525 480115
rect 705581 480059 705649 480115
rect 705705 480059 705773 480115
rect 705829 480059 705897 480115
rect 705953 480059 706000 480115
rect 705512 479991 706000 480059
rect 705512 479935 705525 479991
rect 705581 479935 705649 479991
rect 705705 479935 705773 479991
rect 705829 479935 705897 479991
rect 705953 479935 706000 479991
rect 705512 479867 706000 479935
rect 705512 479811 705525 479867
rect 705581 479811 705649 479867
rect 705705 479811 705773 479867
rect 705829 479811 705897 479867
rect 705953 479811 706000 479867
rect 705512 479743 706000 479811
rect 705512 479687 705525 479743
rect 705581 479687 705649 479743
rect 705705 479687 705773 479743
rect 705829 479687 705897 479743
rect 705953 479687 706000 479743
rect 705512 479619 706000 479687
rect 705512 479563 705525 479619
rect 705581 479563 705649 479619
rect 705705 479563 705773 479619
rect 705829 479563 705897 479619
rect 705953 479563 706000 479619
rect 705512 479495 706000 479563
rect 705512 479439 705525 479495
rect 705581 479439 705649 479495
rect 705705 479439 705773 479495
rect 705829 479439 705897 479495
rect 705953 479439 706000 479495
rect 705512 479371 706000 479439
rect 705512 479315 705525 479371
rect 705581 479315 705649 479371
rect 705705 479315 705773 479371
rect 705829 479315 705897 479371
rect 705953 479315 706000 479371
rect 705512 479247 706000 479315
rect 705512 479191 705525 479247
rect 705581 479191 705649 479247
rect 705705 479191 705773 479247
rect 705829 479191 705897 479247
rect 705953 479191 706000 479247
rect 705512 479123 706000 479191
rect 705512 479067 705525 479123
rect 705581 479067 705649 479123
rect 705705 479067 705773 479123
rect 705829 479067 705897 479123
rect 705953 479067 706000 479123
rect 705512 478999 706000 479067
rect 705512 478943 705525 478999
rect 705581 478943 705649 478999
rect 705705 478943 705773 478999
rect 705829 478943 705897 478999
rect 705953 478943 706000 478999
rect 705512 478875 706000 478943
rect 705512 478819 705525 478875
rect 705581 478819 705649 478875
rect 705705 478819 705773 478875
rect 705829 478819 705897 478875
rect 705953 478819 706000 478875
rect 705512 478752 706000 478819
rect 705512 478131 706000 478172
rect 705512 478075 705525 478131
rect 705581 478075 705649 478131
rect 705705 478075 705773 478131
rect 705829 478075 705897 478131
rect 705953 478075 706000 478131
rect 705512 478007 706000 478075
rect 705512 477951 705525 478007
rect 705581 477951 705649 478007
rect 705705 477951 705773 478007
rect 705829 477951 705897 478007
rect 705953 477951 706000 478007
rect 705512 477883 706000 477951
rect 705512 477827 705525 477883
rect 705581 477827 705649 477883
rect 705705 477827 705773 477883
rect 705829 477827 705897 477883
rect 705953 477827 706000 477883
rect 705512 477759 706000 477827
rect 705512 477703 705525 477759
rect 705581 477703 705649 477759
rect 705705 477703 705773 477759
rect 705829 477703 705897 477759
rect 705953 477703 706000 477759
rect 705512 477635 706000 477703
rect 705512 477579 705525 477635
rect 705581 477579 705649 477635
rect 705705 477579 705773 477635
rect 705829 477579 705897 477635
rect 705953 477579 706000 477635
rect 705512 477511 706000 477579
rect 705512 477455 705525 477511
rect 705581 477455 705649 477511
rect 705705 477455 705773 477511
rect 705829 477455 705897 477511
rect 705953 477455 706000 477511
rect 705512 477387 706000 477455
rect 705512 477331 705525 477387
rect 705581 477331 705649 477387
rect 705705 477331 705773 477387
rect 705829 477331 705897 477387
rect 705953 477331 706000 477387
rect 705512 477263 706000 477331
rect 705512 477207 705525 477263
rect 705581 477207 705649 477263
rect 705705 477207 705773 477263
rect 705829 477207 705897 477263
rect 705953 477207 706000 477263
rect 705512 477139 706000 477207
rect 705512 477083 705525 477139
rect 705581 477083 705649 477139
rect 705705 477083 705773 477139
rect 705829 477083 705897 477139
rect 705953 477083 706000 477139
rect 705512 477015 706000 477083
rect 705512 476959 705525 477015
rect 705581 476959 705649 477015
rect 705705 476959 705773 477015
rect 705829 476959 705897 477015
rect 705953 476959 706000 477015
rect 705512 476891 706000 476959
rect 705512 476835 705525 476891
rect 705581 476835 705649 476891
rect 705705 476835 705773 476891
rect 705829 476835 705897 476891
rect 705953 476835 706000 476891
rect 705512 476767 706000 476835
rect 705512 476711 705525 476767
rect 705581 476711 705649 476767
rect 705705 476711 705773 476767
rect 705829 476711 705897 476767
rect 705953 476711 706000 476767
rect 705512 476643 706000 476711
rect 705512 476587 705525 476643
rect 705581 476587 705649 476643
rect 705705 476587 705773 476643
rect 705829 476587 705897 476643
rect 705953 476587 706000 476643
rect 705512 476519 706000 476587
rect 705512 476463 705525 476519
rect 705581 476463 705649 476519
rect 705705 476463 705773 476519
rect 705829 476463 705897 476519
rect 705953 476463 706000 476519
rect 705512 476395 706000 476463
rect 705512 476339 705525 476395
rect 705581 476339 705649 476395
rect 705705 476339 705773 476395
rect 705829 476339 705897 476395
rect 705953 476339 706000 476395
rect 705512 476272 706000 476339
rect 70000 468661 70488 468728
rect 70000 468605 70047 468661
rect 70103 468605 70171 468661
rect 70227 468605 70295 468661
rect 70351 468605 70419 468661
rect 70475 468605 70488 468661
rect 70000 468537 70488 468605
rect 70000 468481 70047 468537
rect 70103 468481 70171 468537
rect 70227 468481 70295 468537
rect 70351 468481 70419 468537
rect 70475 468481 70488 468537
rect 70000 468413 70488 468481
rect 70000 468357 70047 468413
rect 70103 468357 70171 468413
rect 70227 468357 70295 468413
rect 70351 468357 70419 468413
rect 70475 468357 70488 468413
rect 70000 468289 70488 468357
rect 70000 468233 70047 468289
rect 70103 468233 70171 468289
rect 70227 468233 70295 468289
rect 70351 468233 70419 468289
rect 70475 468233 70488 468289
rect 70000 468165 70488 468233
rect 70000 468109 70047 468165
rect 70103 468109 70171 468165
rect 70227 468109 70295 468165
rect 70351 468109 70419 468165
rect 70475 468109 70488 468165
rect 70000 468041 70488 468109
rect 70000 467985 70047 468041
rect 70103 467985 70171 468041
rect 70227 467985 70295 468041
rect 70351 467985 70419 468041
rect 70475 467985 70488 468041
rect 70000 467917 70488 467985
rect 70000 467861 70047 467917
rect 70103 467861 70171 467917
rect 70227 467861 70295 467917
rect 70351 467861 70419 467917
rect 70475 467861 70488 467917
rect 70000 467793 70488 467861
rect 70000 467737 70047 467793
rect 70103 467737 70171 467793
rect 70227 467737 70295 467793
rect 70351 467737 70419 467793
rect 70475 467737 70488 467793
rect 70000 467669 70488 467737
rect 70000 467613 70047 467669
rect 70103 467613 70171 467669
rect 70227 467613 70295 467669
rect 70351 467613 70419 467669
rect 70475 467613 70488 467669
rect 70000 467545 70488 467613
rect 70000 467489 70047 467545
rect 70103 467489 70171 467545
rect 70227 467489 70295 467545
rect 70351 467489 70419 467545
rect 70475 467489 70488 467545
rect 70000 467421 70488 467489
rect 70000 467365 70047 467421
rect 70103 467365 70171 467421
rect 70227 467365 70295 467421
rect 70351 467365 70419 467421
rect 70475 467365 70488 467421
rect 70000 467297 70488 467365
rect 70000 467241 70047 467297
rect 70103 467241 70171 467297
rect 70227 467241 70295 467297
rect 70351 467241 70419 467297
rect 70475 467241 70488 467297
rect 70000 467173 70488 467241
rect 70000 467117 70047 467173
rect 70103 467117 70171 467173
rect 70227 467117 70295 467173
rect 70351 467117 70419 467173
rect 70475 467117 70488 467173
rect 70000 467049 70488 467117
rect 70000 466993 70047 467049
rect 70103 466993 70171 467049
rect 70227 466993 70295 467049
rect 70351 466993 70419 467049
rect 70475 466993 70488 467049
rect 70000 466925 70488 466993
rect 70000 466869 70047 466925
rect 70103 466869 70171 466925
rect 70227 466869 70295 466925
rect 70351 466869 70419 466925
rect 70475 466869 70488 466925
rect 70000 466828 70488 466869
rect 70000 466181 70488 466248
rect 70000 466125 70047 466181
rect 70103 466125 70171 466181
rect 70227 466125 70295 466181
rect 70351 466125 70419 466181
rect 70475 466125 70488 466181
rect 70000 466057 70488 466125
rect 70000 466001 70047 466057
rect 70103 466001 70171 466057
rect 70227 466001 70295 466057
rect 70351 466001 70419 466057
rect 70475 466001 70488 466057
rect 70000 465933 70488 466001
rect 70000 465877 70047 465933
rect 70103 465877 70171 465933
rect 70227 465877 70295 465933
rect 70351 465877 70419 465933
rect 70475 465877 70488 465933
rect 70000 465809 70488 465877
rect 70000 465753 70047 465809
rect 70103 465753 70171 465809
rect 70227 465753 70295 465809
rect 70351 465753 70419 465809
rect 70475 465753 70488 465809
rect 70000 465685 70488 465753
rect 70000 465629 70047 465685
rect 70103 465629 70171 465685
rect 70227 465629 70295 465685
rect 70351 465629 70419 465685
rect 70475 465629 70488 465685
rect 70000 465561 70488 465629
rect 70000 465505 70047 465561
rect 70103 465505 70171 465561
rect 70227 465505 70295 465561
rect 70351 465505 70419 465561
rect 70475 465505 70488 465561
rect 70000 465437 70488 465505
rect 70000 465381 70047 465437
rect 70103 465381 70171 465437
rect 70227 465381 70295 465437
rect 70351 465381 70419 465437
rect 70475 465381 70488 465437
rect 70000 465313 70488 465381
rect 70000 465257 70047 465313
rect 70103 465257 70171 465313
rect 70227 465257 70295 465313
rect 70351 465257 70419 465313
rect 70475 465257 70488 465313
rect 70000 465189 70488 465257
rect 70000 465133 70047 465189
rect 70103 465133 70171 465189
rect 70227 465133 70295 465189
rect 70351 465133 70419 465189
rect 70475 465133 70488 465189
rect 70000 465065 70488 465133
rect 70000 465009 70047 465065
rect 70103 465009 70171 465065
rect 70227 465009 70295 465065
rect 70351 465009 70419 465065
rect 70475 465009 70488 465065
rect 70000 464941 70488 465009
rect 70000 464885 70047 464941
rect 70103 464885 70171 464941
rect 70227 464885 70295 464941
rect 70351 464885 70419 464941
rect 70475 464885 70488 464941
rect 70000 464817 70488 464885
rect 70000 464761 70047 464817
rect 70103 464761 70171 464817
rect 70227 464761 70295 464817
rect 70351 464761 70419 464817
rect 70475 464761 70488 464817
rect 70000 464693 70488 464761
rect 70000 464637 70047 464693
rect 70103 464637 70171 464693
rect 70227 464637 70295 464693
rect 70351 464637 70419 464693
rect 70475 464637 70488 464693
rect 70000 464569 70488 464637
rect 70000 464513 70047 464569
rect 70103 464513 70171 464569
rect 70227 464513 70295 464569
rect 70351 464513 70419 464569
rect 70475 464513 70488 464569
rect 70000 464445 70488 464513
rect 70000 464389 70047 464445
rect 70103 464389 70171 464445
rect 70227 464389 70295 464445
rect 70351 464389 70419 464445
rect 70475 464389 70488 464445
rect 70000 464321 70488 464389
rect 70000 464265 70047 464321
rect 70103 464265 70171 464321
rect 70227 464265 70295 464321
rect 70351 464265 70419 464321
rect 70475 464265 70488 464321
rect 70000 464198 70488 464265
rect 70000 463811 70488 463878
rect 70000 463755 70047 463811
rect 70103 463755 70171 463811
rect 70227 463755 70295 463811
rect 70351 463755 70419 463811
rect 70475 463755 70488 463811
rect 70000 463687 70488 463755
rect 70000 463631 70047 463687
rect 70103 463631 70171 463687
rect 70227 463631 70295 463687
rect 70351 463631 70419 463687
rect 70475 463631 70488 463687
rect 70000 463563 70488 463631
rect 70000 463507 70047 463563
rect 70103 463507 70171 463563
rect 70227 463507 70295 463563
rect 70351 463507 70419 463563
rect 70475 463507 70488 463563
rect 70000 463439 70488 463507
rect 70000 463383 70047 463439
rect 70103 463383 70171 463439
rect 70227 463383 70295 463439
rect 70351 463383 70419 463439
rect 70475 463383 70488 463439
rect 70000 463315 70488 463383
rect 70000 463259 70047 463315
rect 70103 463259 70171 463315
rect 70227 463259 70295 463315
rect 70351 463259 70419 463315
rect 70475 463259 70488 463315
rect 70000 463191 70488 463259
rect 70000 463135 70047 463191
rect 70103 463135 70171 463191
rect 70227 463135 70295 463191
rect 70351 463135 70419 463191
rect 70475 463135 70488 463191
rect 70000 463067 70488 463135
rect 70000 463011 70047 463067
rect 70103 463011 70171 463067
rect 70227 463011 70295 463067
rect 70351 463011 70419 463067
rect 70475 463011 70488 463067
rect 70000 462943 70488 463011
rect 70000 462887 70047 462943
rect 70103 462887 70171 462943
rect 70227 462887 70295 462943
rect 70351 462887 70419 462943
rect 70475 462887 70488 462943
rect 70000 462819 70488 462887
rect 70000 462763 70047 462819
rect 70103 462763 70171 462819
rect 70227 462763 70295 462819
rect 70351 462763 70419 462819
rect 70475 462763 70488 462819
rect 70000 462695 70488 462763
rect 70000 462639 70047 462695
rect 70103 462639 70171 462695
rect 70227 462639 70295 462695
rect 70351 462639 70419 462695
rect 70475 462639 70488 462695
rect 70000 462571 70488 462639
rect 70000 462515 70047 462571
rect 70103 462515 70171 462571
rect 70227 462515 70295 462571
rect 70351 462515 70419 462571
rect 70475 462515 70488 462571
rect 70000 462447 70488 462515
rect 70000 462391 70047 462447
rect 70103 462391 70171 462447
rect 70227 462391 70295 462447
rect 70351 462391 70419 462447
rect 70475 462391 70488 462447
rect 70000 462323 70488 462391
rect 70000 462267 70047 462323
rect 70103 462267 70171 462323
rect 70227 462267 70295 462323
rect 70351 462267 70419 462323
rect 70475 462267 70488 462323
rect 70000 462199 70488 462267
rect 70000 462143 70047 462199
rect 70103 462143 70171 462199
rect 70227 462143 70295 462199
rect 70351 462143 70419 462199
rect 70475 462143 70488 462199
rect 70000 462075 70488 462143
rect 70000 462019 70047 462075
rect 70103 462019 70171 462075
rect 70227 462019 70295 462075
rect 70351 462019 70419 462075
rect 70475 462019 70488 462075
rect 70000 461951 70488 462019
rect 70000 461895 70047 461951
rect 70103 461895 70171 461951
rect 70227 461895 70295 461951
rect 70351 461895 70419 461951
rect 70475 461895 70488 461951
rect 70000 461828 70488 461895
rect 70000 461105 70488 461172
rect 70000 461049 70047 461105
rect 70103 461049 70171 461105
rect 70227 461049 70295 461105
rect 70351 461049 70419 461105
rect 70475 461049 70488 461105
rect 70000 460981 70488 461049
rect 70000 460925 70047 460981
rect 70103 460925 70171 460981
rect 70227 460925 70295 460981
rect 70351 460925 70419 460981
rect 70475 460925 70488 460981
rect 70000 460857 70488 460925
rect 70000 460801 70047 460857
rect 70103 460801 70171 460857
rect 70227 460801 70295 460857
rect 70351 460801 70419 460857
rect 70475 460801 70488 460857
rect 70000 460733 70488 460801
rect 70000 460677 70047 460733
rect 70103 460677 70171 460733
rect 70227 460677 70295 460733
rect 70351 460677 70419 460733
rect 70475 460677 70488 460733
rect 70000 460609 70488 460677
rect 70000 460553 70047 460609
rect 70103 460553 70171 460609
rect 70227 460553 70295 460609
rect 70351 460553 70419 460609
rect 70475 460553 70488 460609
rect 70000 460485 70488 460553
rect 70000 460429 70047 460485
rect 70103 460429 70171 460485
rect 70227 460429 70295 460485
rect 70351 460429 70419 460485
rect 70475 460429 70488 460485
rect 70000 460361 70488 460429
rect 70000 460305 70047 460361
rect 70103 460305 70171 460361
rect 70227 460305 70295 460361
rect 70351 460305 70419 460361
rect 70475 460305 70488 460361
rect 70000 460237 70488 460305
rect 70000 460181 70047 460237
rect 70103 460181 70171 460237
rect 70227 460181 70295 460237
rect 70351 460181 70419 460237
rect 70475 460181 70488 460237
rect 70000 460113 70488 460181
rect 70000 460057 70047 460113
rect 70103 460057 70171 460113
rect 70227 460057 70295 460113
rect 70351 460057 70419 460113
rect 70475 460057 70488 460113
rect 70000 459989 70488 460057
rect 70000 459933 70047 459989
rect 70103 459933 70171 459989
rect 70227 459933 70295 459989
rect 70351 459933 70419 459989
rect 70475 459933 70488 459989
rect 70000 459865 70488 459933
rect 70000 459809 70047 459865
rect 70103 459809 70171 459865
rect 70227 459809 70295 459865
rect 70351 459809 70419 459865
rect 70475 459809 70488 459865
rect 70000 459741 70488 459809
rect 70000 459685 70047 459741
rect 70103 459685 70171 459741
rect 70227 459685 70295 459741
rect 70351 459685 70419 459741
rect 70475 459685 70488 459741
rect 70000 459617 70488 459685
rect 70000 459561 70047 459617
rect 70103 459561 70171 459617
rect 70227 459561 70295 459617
rect 70351 459561 70419 459617
rect 70475 459561 70488 459617
rect 70000 459493 70488 459561
rect 70000 459437 70047 459493
rect 70103 459437 70171 459493
rect 70227 459437 70295 459493
rect 70351 459437 70419 459493
rect 70475 459437 70488 459493
rect 70000 459369 70488 459437
rect 70000 459313 70047 459369
rect 70103 459313 70171 459369
rect 70227 459313 70295 459369
rect 70351 459313 70419 459369
rect 70475 459313 70488 459369
rect 70000 459245 70488 459313
rect 70000 459189 70047 459245
rect 70103 459189 70171 459245
rect 70227 459189 70295 459245
rect 70351 459189 70419 459245
rect 70475 459189 70488 459245
rect 70000 459122 70488 459189
rect 70000 458735 70488 458802
rect 70000 458679 70047 458735
rect 70103 458679 70171 458735
rect 70227 458679 70295 458735
rect 70351 458679 70419 458735
rect 70475 458679 70488 458735
rect 70000 458611 70488 458679
rect 70000 458555 70047 458611
rect 70103 458555 70171 458611
rect 70227 458555 70295 458611
rect 70351 458555 70419 458611
rect 70475 458555 70488 458611
rect 70000 458487 70488 458555
rect 70000 458431 70047 458487
rect 70103 458431 70171 458487
rect 70227 458431 70295 458487
rect 70351 458431 70419 458487
rect 70475 458431 70488 458487
rect 70000 458363 70488 458431
rect 70000 458307 70047 458363
rect 70103 458307 70171 458363
rect 70227 458307 70295 458363
rect 70351 458307 70419 458363
rect 70475 458307 70488 458363
rect 70000 458239 70488 458307
rect 70000 458183 70047 458239
rect 70103 458183 70171 458239
rect 70227 458183 70295 458239
rect 70351 458183 70419 458239
rect 70475 458183 70488 458239
rect 70000 458115 70488 458183
rect 70000 458059 70047 458115
rect 70103 458059 70171 458115
rect 70227 458059 70295 458115
rect 70351 458059 70419 458115
rect 70475 458059 70488 458115
rect 70000 457991 70488 458059
rect 70000 457935 70047 457991
rect 70103 457935 70171 457991
rect 70227 457935 70295 457991
rect 70351 457935 70419 457991
rect 70475 457935 70488 457991
rect 70000 457867 70488 457935
rect 70000 457811 70047 457867
rect 70103 457811 70171 457867
rect 70227 457811 70295 457867
rect 70351 457811 70419 457867
rect 70475 457811 70488 457867
rect 70000 457743 70488 457811
rect 70000 457687 70047 457743
rect 70103 457687 70171 457743
rect 70227 457687 70295 457743
rect 70351 457687 70419 457743
rect 70475 457687 70488 457743
rect 70000 457619 70488 457687
rect 70000 457563 70047 457619
rect 70103 457563 70171 457619
rect 70227 457563 70295 457619
rect 70351 457563 70419 457619
rect 70475 457563 70488 457619
rect 70000 457495 70488 457563
rect 70000 457439 70047 457495
rect 70103 457439 70171 457495
rect 70227 457439 70295 457495
rect 70351 457439 70419 457495
rect 70475 457439 70488 457495
rect 70000 457371 70488 457439
rect 70000 457315 70047 457371
rect 70103 457315 70171 457371
rect 70227 457315 70295 457371
rect 70351 457315 70419 457371
rect 70475 457315 70488 457371
rect 70000 457247 70488 457315
rect 70000 457191 70047 457247
rect 70103 457191 70171 457247
rect 70227 457191 70295 457247
rect 70351 457191 70419 457247
rect 70475 457191 70488 457247
rect 70000 457123 70488 457191
rect 70000 457067 70047 457123
rect 70103 457067 70171 457123
rect 70227 457067 70295 457123
rect 70351 457067 70419 457123
rect 70475 457067 70488 457123
rect 70000 456999 70488 457067
rect 70000 456943 70047 456999
rect 70103 456943 70171 456999
rect 70227 456943 70295 456999
rect 70351 456943 70419 456999
rect 70475 456943 70488 456999
rect 70000 456875 70488 456943
rect 70000 456819 70047 456875
rect 70103 456819 70171 456875
rect 70227 456819 70295 456875
rect 70351 456819 70419 456875
rect 70475 456819 70488 456875
rect 70000 456752 70488 456819
rect 70000 456105 70488 456172
rect 70000 456049 70047 456105
rect 70103 456049 70171 456105
rect 70227 456049 70295 456105
rect 70351 456049 70419 456105
rect 70475 456049 70488 456105
rect 70000 455981 70488 456049
rect 70000 455925 70047 455981
rect 70103 455925 70171 455981
rect 70227 455925 70295 455981
rect 70351 455925 70419 455981
rect 70475 455925 70488 455981
rect 70000 455857 70488 455925
rect 70000 455801 70047 455857
rect 70103 455801 70171 455857
rect 70227 455801 70295 455857
rect 70351 455801 70419 455857
rect 70475 455801 70488 455857
rect 70000 455733 70488 455801
rect 70000 455677 70047 455733
rect 70103 455677 70171 455733
rect 70227 455677 70295 455733
rect 70351 455677 70419 455733
rect 70475 455677 70488 455733
rect 70000 455609 70488 455677
rect 70000 455553 70047 455609
rect 70103 455553 70171 455609
rect 70227 455553 70295 455609
rect 70351 455553 70419 455609
rect 70475 455553 70488 455609
rect 70000 455485 70488 455553
rect 70000 455429 70047 455485
rect 70103 455429 70171 455485
rect 70227 455429 70295 455485
rect 70351 455429 70419 455485
rect 70475 455429 70488 455485
rect 70000 455361 70488 455429
rect 70000 455305 70047 455361
rect 70103 455305 70171 455361
rect 70227 455305 70295 455361
rect 70351 455305 70419 455361
rect 70475 455305 70488 455361
rect 70000 455237 70488 455305
rect 70000 455181 70047 455237
rect 70103 455181 70171 455237
rect 70227 455181 70295 455237
rect 70351 455181 70419 455237
rect 70475 455181 70488 455237
rect 70000 455113 70488 455181
rect 70000 455057 70047 455113
rect 70103 455057 70171 455113
rect 70227 455057 70295 455113
rect 70351 455057 70419 455113
rect 70475 455057 70488 455113
rect 70000 454989 70488 455057
rect 70000 454933 70047 454989
rect 70103 454933 70171 454989
rect 70227 454933 70295 454989
rect 70351 454933 70419 454989
rect 70475 454933 70488 454989
rect 70000 454865 70488 454933
rect 70000 454809 70047 454865
rect 70103 454809 70171 454865
rect 70227 454809 70295 454865
rect 70351 454809 70419 454865
rect 70475 454809 70488 454865
rect 70000 454741 70488 454809
rect 70000 454685 70047 454741
rect 70103 454685 70171 454741
rect 70227 454685 70295 454741
rect 70351 454685 70419 454741
rect 70475 454685 70488 454741
rect 70000 454617 70488 454685
rect 70000 454561 70047 454617
rect 70103 454561 70171 454617
rect 70227 454561 70295 454617
rect 70351 454561 70419 454617
rect 70475 454561 70488 454617
rect 70000 454493 70488 454561
rect 70000 454437 70047 454493
rect 70103 454437 70171 454493
rect 70227 454437 70295 454493
rect 70351 454437 70419 454493
rect 70475 454437 70488 454493
rect 70000 454369 70488 454437
rect 70000 454313 70047 454369
rect 70103 454313 70171 454369
rect 70227 454313 70295 454369
rect 70351 454313 70419 454369
rect 70475 454313 70488 454369
rect 70000 454272 70488 454313
rect 705512 447687 706000 447728
rect 705512 447631 705525 447687
rect 705581 447631 705649 447687
rect 705705 447631 705773 447687
rect 705829 447631 705897 447687
rect 705953 447631 706000 447687
rect 705512 447563 706000 447631
rect 705512 447507 705525 447563
rect 705581 447507 705649 447563
rect 705705 447507 705773 447563
rect 705829 447507 705897 447563
rect 705953 447507 706000 447563
rect 705512 447439 706000 447507
rect 705512 447383 705525 447439
rect 705581 447383 705649 447439
rect 705705 447383 705773 447439
rect 705829 447383 705897 447439
rect 705953 447383 706000 447439
rect 705512 447315 706000 447383
rect 705512 447259 705525 447315
rect 705581 447259 705649 447315
rect 705705 447259 705773 447315
rect 705829 447259 705897 447315
rect 705953 447259 706000 447315
rect 705512 447191 706000 447259
rect 705512 447135 705525 447191
rect 705581 447135 705649 447191
rect 705705 447135 705773 447191
rect 705829 447135 705897 447191
rect 705953 447135 706000 447191
rect 705512 447067 706000 447135
rect 705512 447011 705525 447067
rect 705581 447011 705649 447067
rect 705705 447011 705773 447067
rect 705829 447011 705897 447067
rect 705953 447011 706000 447067
rect 705512 446943 706000 447011
rect 705512 446887 705525 446943
rect 705581 446887 705649 446943
rect 705705 446887 705773 446943
rect 705829 446887 705897 446943
rect 705953 446887 706000 446943
rect 705512 446819 706000 446887
rect 705512 446763 705525 446819
rect 705581 446763 705649 446819
rect 705705 446763 705773 446819
rect 705829 446763 705897 446819
rect 705953 446763 706000 446819
rect 705512 446695 706000 446763
rect 705512 446639 705525 446695
rect 705581 446639 705649 446695
rect 705705 446639 705773 446695
rect 705829 446639 705897 446695
rect 705953 446639 706000 446695
rect 705512 446571 706000 446639
rect 705512 446515 705525 446571
rect 705581 446515 705649 446571
rect 705705 446515 705773 446571
rect 705829 446515 705897 446571
rect 705953 446515 706000 446571
rect 705512 446447 706000 446515
rect 705512 446391 705525 446447
rect 705581 446391 705649 446447
rect 705705 446391 705773 446447
rect 705829 446391 705897 446447
rect 705953 446391 706000 446447
rect 705512 446323 706000 446391
rect 705512 446267 705525 446323
rect 705581 446267 705649 446323
rect 705705 446267 705773 446323
rect 705829 446267 705897 446323
rect 705953 446267 706000 446323
rect 705512 446199 706000 446267
rect 705512 446143 705525 446199
rect 705581 446143 705649 446199
rect 705705 446143 705773 446199
rect 705829 446143 705897 446199
rect 705953 446143 706000 446199
rect 705512 446075 706000 446143
rect 705512 446019 705525 446075
rect 705581 446019 705649 446075
rect 705705 446019 705773 446075
rect 705829 446019 705897 446075
rect 705953 446019 706000 446075
rect 705512 445951 706000 446019
rect 705512 445895 705525 445951
rect 705581 445895 705649 445951
rect 705705 445895 705773 445951
rect 705829 445895 705897 445951
rect 705953 445895 706000 445951
rect 705512 445828 706000 445895
rect 705512 445181 706000 445248
rect 705512 445125 705525 445181
rect 705581 445125 705649 445181
rect 705705 445125 705773 445181
rect 705829 445125 705897 445181
rect 705953 445125 706000 445181
rect 705512 445057 706000 445125
rect 705512 445001 705525 445057
rect 705581 445001 705649 445057
rect 705705 445001 705773 445057
rect 705829 445001 705897 445057
rect 705953 445001 706000 445057
rect 705512 444933 706000 445001
rect 705512 444877 705525 444933
rect 705581 444877 705649 444933
rect 705705 444877 705773 444933
rect 705829 444877 705897 444933
rect 705953 444877 706000 444933
rect 705512 444809 706000 444877
rect 705512 444753 705525 444809
rect 705581 444753 705649 444809
rect 705705 444753 705773 444809
rect 705829 444753 705897 444809
rect 705953 444753 706000 444809
rect 705512 444685 706000 444753
rect 705512 444629 705525 444685
rect 705581 444629 705649 444685
rect 705705 444629 705773 444685
rect 705829 444629 705897 444685
rect 705953 444629 706000 444685
rect 705512 444561 706000 444629
rect 705512 444505 705525 444561
rect 705581 444505 705649 444561
rect 705705 444505 705773 444561
rect 705829 444505 705897 444561
rect 705953 444505 706000 444561
rect 705512 444437 706000 444505
rect 705512 444381 705525 444437
rect 705581 444381 705649 444437
rect 705705 444381 705773 444437
rect 705829 444381 705897 444437
rect 705953 444381 706000 444437
rect 705512 444313 706000 444381
rect 705512 444257 705525 444313
rect 705581 444257 705649 444313
rect 705705 444257 705773 444313
rect 705829 444257 705897 444313
rect 705953 444257 706000 444313
rect 705512 444189 706000 444257
rect 705512 444133 705525 444189
rect 705581 444133 705649 444189
rect 705705 444133 705773 444189
rect 705829 444133 705897 444189
rect 705953 444133 706000 444189
rect 705512 444065 706000 444133
rect 705512 444009 705525 444065
rect 705581 444009 705649 444065
rect 705705 444009 705773 444065
rect 705829 444009 705897 444065
rect 705953 444009 706000 444065
rect 705512 443941 706000 444009
rect 705512 443885 705525 443941
rect 705581 443885 705649 443941
rect 705705 443885 705773 443941
rect 705829 443885 705897 443941
rect 705953 443885 706000 443941
rect 705512 443817 706000 443885
rect 705512 443761 705525 443817
rect 705581 443761 705649 443817
rect 705705 443761 705773 443817
rect 705829 443761 705897 443817
rect 705953 443761 706000 443817
rect 705512 443693 706000 443761
rect 705512 443637 705525 443693
rect 705581 443637 705649 443693
rect 705705 443637 705773 443693
rect 705829 443637 705897 443693
rect 705953 443637 706000 443693
rect 705512 443569 706000 443637
rect 705512 443513 705525 443569
rect 705581 443513 705649 443569
rect 705705 443513 705773 443569
rect 705829 443513 705897 443569
rect 705953 443513 706000 443569
rect 705512 443445 706000 443513
rect 705512 443389 705525 443445
rect 705581 443389 705649 443445
rect 705705 443389 705773 443445
rect 705829 443389 705897 443445
rect 705953 443389 706000 443445
rect 705512 443321 706000 443389
rect 705512 443265 705525 443321
rect 705581 443265 705649 443321
rect 705705 443265 705773 443321
rect 705829 443265 705897 443321
rect 705953 443265 706000 443321
rect 705512 443198 706000 443265
rect 705512 442811 706000 442878
rect 705512 442755 705525 442811
rect 705581 442755 705649 442811
rect 705705 442755 705773 442811
rect 705829 442755 705897 442811
rect 705953 442755 706000 442811
rect 705512 442687 706000 442755
rect 705512 442631 705525 442687
rect 705581 442631 705649 442687
rect 705705 442631 705773 442687
rect 705829 442631 705897 442687
rect 705953 442631 706000 442687
rect 705512 442563 706000 442631
rect 705512 442507 705525 442563
rect 705581 442507 705649 442563
rect 705705 442507 705773 442563
rect 705829 442507 705897 442563
rect 705953 442507 706000 442563
rect 705512 442439 706000 442507
rect 705512 442383 705525 442439
rect 705581 442383 705649 442439
rect 705705 442383 705773 442439
rect 705829 442383 705897 442439
rect 705953 442383 706000 442439
rect 705512 442315 706000 442383
rect 705512 442259 705525 442315
rect 705581 442259 705649 442315
rect 705705 442259 705773 442315
rect 705829 442259 705897 442315
rect 705953 442259 706000 442315
rect 705512 442191 706000 442259
rect 705512 442135 705525 442191
rect 705581 442135 705649 442191
rect 705705 442135 705773 442191
rect 705829 442135 705897 442191
rect 705953 442135 706000 442191
rect 705512 442067 706000 442135
rect 705512 442011 705525 442067
rect 705581 442011 705649 442067
rect 705705 442011 705773 442067
rect 705829 442011 705897 442067
rect 705953 442011 706000 442067
rect 705512 441943 706000 442011
rect 705512 441887 705525 441943
rect 705581 441887 705649 441943
rect 705705 441887 705773 441943
rect 705829 441887 705897 441943
rect 705953 441887 706000 441943
rect 705512 441819 706000 441887
rect 705512 441763 705525 441819
rect 705581 441763 705649 441819
rect 705705 441763 705773 441819
rect 705829 441763 705897 441819
rect 705953 441763 706000 441819
rect 705512 441695 706000 441763
rect 705512 441639 705525 441695
rect 705581 441639 705649 441695
rect 705705 441639 705773 441695
rect 705829 441639 705897 441695
rect 705953 441639 706000 441695
rect 705512 441571 706000 441639
rect 705512 441515 705525 441571
rect 705581 441515 705649 441571
rect 705705 441515 705773 441571
rect 705829 441515 705897 441571
rect 705953 441515 706000 441571
rect 705512 441447 706000 441515
rect 705512 441391 705525 441447
rect 705581 441391 705649 441447
rect 705705 441391 705773 441447
rect 705829 441391 705897 441447
rect 705953 441391 706000 441447
rect 705512 441323 706000 441391
rect 705512 441267 705525 441323
rect 705581 441267 705649 441323
rect 705705 441267 705773 441323
rect 705829 441267 705897 441323
rect 705953 441267 706000 441323
rect 705512 441199 706000 441267
rect 705512 441143 705525 441199
rect 705581 441143 705649 441199
rect 705705 441143 705773 441199
rect 705829 441143 705897 441199
rect 705953 441143 706000 441199
rect 705512 441075 706000 441143
rect 705512 441019 705525 441075
rect 705581 441019 705649 441075
rect 705705 441019 705773 441075
rect 705829 441019 705897 441075
rect 705953 441019 706000 441075
rect 705512 440951 706000 441019
rect 705512 440895 705525 440951
rect 705581 440895 705649 440951
rect 705705 440895 705773 440951
rect 705829 440895 705897 440951
rect 705953 440895 706000 440951
rect 705512 440828 706000 440895
rect 705512 440105 706000 440172
rect 705512 440049 705525 440105
rect 705581 440049 705649 440105
rect 705705 440049 705773 440105
rect 705829 440049 705897 440105
rect 705953 440049 706000 440105
rect 705512 439981 706000 440049
rect 705512 439925 705525 439981
rect 705581 439925 705649 439981
rect 705705 439925 705773 439981
rect 705829 439925 705897 439981
rect 705953 439925 706000 439981
rect 705512 439857 706000 439925
rect 705512 439801 705525 439857
rect 705581 439801 705649 439857
rect 705705 439801 705773 439857
rect 705829 439801 705897 439857
rect 705953 439801 706000 439857
rect 705512 439733 706000 439801
rect 705512 439677 705525 439733
rect 705581 439677 705649 439733
rect 705705 439677 705773 439733
rect 705829 439677 705897 439733
rect 705953 439677 706000 439733
rect 705512 439609 706000 439677
rect 705512 439553 705525 439609
rect 705581 439553 705649 439609
rect 705705 439553 705773 439609
rect 705829 439553 705897 439609
rect 705953 439553 706000 439609
rect 705512 439485 706000 439553
rect 705512 439429 705525 439485
rect 705581 439429 705649 439485
rect 705705 439429 705773 439485
rect 705829 439429 705897 439485
rect 705953 439429 706000 439485
rect 705512 439361 706000 439429
rect 705512 439305 705525 439361
rect 705581 439305 705649 439361
rect 705705 439305 705773 439361
rect 705829 439305 705897 439361
rect 705953 439305 706000 439361
rect 705512 439237 706000 439305
rect 705512 439181 705525 439237
rect 705581 439181 705649 439237
rect 705705 439181 705773 439237
rect 705829 439181 705897 439237
rect 705953 439181 706000 439237
rect 705512 439113 706000 439181
rect 705512 439057 705525 439113
rect 705581 439057 705649 439113
rect 705705 439057 705773 439113
rect 705829 439057 705897 439113
rect 705953 439057 706000 439113
rect 705512 438989 706000 439057
rect 705512 438933 705525 438989
rect 705581 438933 705649 438989
rect 705705 438933 705773 438989
rect 705829 438933 705897 438989
rect 705953 438933 706000 438989
rect 705512 438865 706000 438933
rect 705512 438809 705525 438865
rect 705581 438809 705649 438865
rect 705705 438809 705773 438865
rect 705829 438809 705897 438865
rect 705953 438809 706000 438865
rect 705512 438741 706000 438809
rect 705512 438685 705525 438741
rect 705581 438685 705649 438741
rect 705705 438685 705773 438741
rect 705829 438685 705897 438741
rect 705953 438685 706000 438741
rect 705512 438617 706000 438685
rect 705512 438561 705525 438617
rect 705581 438561 705649 438617
rect 705705 438561 705773 438617
rect 705829 438561 705897 438617
rect 705953 438561 706000 438617
rect 705512 438493 706000 438561
rect 705512 438437 705525 438493
rect 705581 438437 705649 438493
rect 705705 438437 705773 438493
rect 705829 438437 705897 438493
rect 705953 438437 706000 438493
rect 705512 438369 706000 438437
rect 705512 438313 705525 438369
rect 705581 438313 705649 438369
rect 705705 438313 705773 438369
rect 705829 438313 705897 438369
rect 705953 438313 706000 438369
rect 705512 438245 706000 438313
rect 705512 438189 705525 438245
rect 705581 438189 705649 438245
rect 705705 438189 705773 438245
rect 705829 438189 705897 438245
rect 705953 438189 706000 438245
rect 705512 438122 706000 438189
rect 705512 437735 706000 437802
rect 705512 437679 705525 437735
rect 705581 437679 705649 437735
rect 705705 437679 705773 437735
rect 705829 437679 705897 437735
rect 705953 437679 706000 437735
rect 705512 437611 706000 437679
rect 705512 437555 705525 437611
rect 705581 437555 705649 437611
rect 705705 437555 705773 437611
rect 705829 437555 705897 437611
rect 705953 437555 706000 437611
rect 705512 437487 706000 437555
rect 705512 437431 705525 437487
rect 705581 437431 705649 437487
rect 705705 437431 705773 437487
rect 705829 437431 705897 437487
rect 705953 437431 706000 437487
rect 705512 437363 706000 437431
rect 705512 437307 705525 437363
rect 705581 437307 705649 437363
rect 705705 437307 705773 437363
rect 705829 437307 705897 437363
rect 705953 437307 706000 437363
rect 705512 437239 706000 437307
rect 705512 437183 705525 437239
rect 705581 437183 705649 437239
rect 705705 437183 705773 437239
rect 705829 437183 705897 437239
rect 705953 437183 706000 437239
rect 705512 437115 706000 437183
rect 705512 437059 705525 437115
rect 705581 437059 705649 437115
rect 705705 437059 705773 437115
rect 705829 437059 705897 437115
rect 705953 437059 706000 437115
rect 705512 436991 706000 437059
rect 705512 436935 705525 436991
rect 705581 436935 705649 436991
rect 705705 436935 705773 436991
rect 705829 436935 705897 436991
rect 705953 436935 706000 436991
rect 705512 436867 706000 436935
rect 705512 436811 705525 436867
rect 705581 436811 705649 436867
rect 705705 436811 705773 436867
rect 705829 436811 705897 436867
rect 705953 436811 706000 436867
rect 705512 436743 706000 436811
rect 705512 436687 705525 436743
rect 705581 436687 705649 436743
rect 705705 436687 705773 436743
rect 705829 436687 705897 436743
rect 705953 436687 706000 436743
rect 705512 436619 706000 436687
rect 705512 436563 705525 436619
rect 705581 436563 705649 436619
rect 705705 436563 705773 436619
rect 705829 436563 705897 436619
rect 705953 436563 706000 436619
rect 705512 436495 706000 436563
rect 705512 436439 705525 436495
rect 705581 436439 705649 436495
rect 705705 436439 705773 436495
rect 705829 436439 705897 436495
rect 705953 436439 706000 436495
rect 705512 436371 706000 436439
rect 705512 436315 705525 436371
rect 705581 436315 705649 436371
rect 705705 436315 705773 436371
rect 705829 436315 705897 436371
rect 705953 436315 706000 436371
rect 705512 436247 706000 436315
rect 705512 436191 705525 436247
rect 705581 436191 705649 436247
rect 705705 436191 705773 436247
rect 705829 436191 705897 436247
rect 705953 436191 706000 436247
rect 705512 435752 706000 436191
rect 705512 435131 706000 435172
rect 705512 435075 705525 435131
rect 705581 435075 705649 435131
rect 705705 435075 705773 435131
rect 705829 435075 705897 435131
rect 705953 435075 706000 435131
rect 705512 435007 706000 435075
rect 705512 434951 705525 435007
rect 705581 434951 705649 435007
rect 705705 434951 705773 435007
rect 705829 434951 705897 435007
rect 705953 434951 706000 435007
rect 705512 434883 706000 434951
rect 705512 434827 705525 434883
rect 705581 434827 705649 434883
rect 705705 434827 705773 434883
rect 705829 434827 705897 434883
rect 705953 434827 706000 434883
rect 705512 434759 706000 434827
rect 705512 434703 705525 434759
rect 705581 434703 705649 434759
rect 705705 434703 705773 434759
rect 705829 434703 705897 434759
rect 705953 434703 706000 434759
rect 705512 434635 706000 434703
rect 705512 434579 705525 434635
rect 705581 434579 705649 434635
rect 705705 434579 705773 434635
rect 705829 434579 705897 434635
rect 705953 434579 706000 434635
rect 705512 434511 706000 434579
rect 705512 434455 705525 434511
rect 705581 434455 705649 434511
rect 705705 434455 705773 434511
rect 705829 434455 705897 434511
rect 705953 434455 706000 434511
rect 705512 434387 706000 434455
rect 705512 434331 705525 434387
rect 705581 434331 705649 434387
rect 705705 434331 705773 434387
rect 705829 434331 705897 434387
rect 705953 434331 706000 434387
rect 705512 434263 706000 434331
rect 705512 434207 705525 434263
rect 705581 434207 705649 434263
rect 705705 434207 705773 434263
rect 705829 434207 705897 434263
rect 705953 434207 706000 434263
rect 705512 434139 706000 434207
rect 705512 434083 705525 434139
rect 705581 434083 705649 434139
rect 705705 434083 705773 434139
rect 705829 434083 705897 434139
rect 705953 434083 706000 434139
rect 705512 434015 706000 434083
rect 705512 433959 705525 434015
rect 705581 433959 705649 434015
rect 705705 433959 705773 434015
rect 705829 433959 705897 434015
rect 705953 433959 706000 434015
rect 705512 433891 706000 433959
rect 705512 433835 705525 433891
rect 705581 433835 705649 433891
rect 705705 433835 705773 433891
rect 705829 433835 705897 433891
rect 705953 433835 706000 433891
rect 705512 433767 706000 433835
rect 705512 433711 705525 433767
rect 705581 433711 705649 433767
rect 705705 433711 705773 433767
rect 705829 433711 705897 433767
rect 705953 433711 706000 433767
rect 705512 433643 706000 433711
rect 705512 433587 705525 433643
rect 705581 433587 705649 433643
rect 705705 433587 705773 433643
rect 705829 433587 705897 433643
rect 705953 433587 706000 433643
rect 705512 433519 706000 433587
rect 705512 433463 705525 433519
rect 705581 433463 705649 433519
rect 705705 433463 705773 433519
rect 705829 433463 705897 433519
rect 705953 433463 706000 433519
rect 705512 433395 706000 433463
rect 705512 433339 705525 433395
rect 705581 433339 705649 433395
rect 705705 433339 705773 433395
rect 705829 433339 705897 433395
rect 705953 433339 706000 433395
rect 705512 433272 706000 433339
rect 70000 427661 70488 427728
rect 70000 427605 70047 427661
rect 70103 427605 70171 427661
rect 70227 427605 70295 427661
rect 70351 427605 70419 427661
rect 70475 427605 70488 427661
rect 70000 427537 70488 427605
rect 70000 427481 70047 427537
rect 70103 427481 70171 427537
rect 70227 427481 70295 427537
rect 70351 427481 70419 427537
rect 70475 427481 70488 427537
rect 70000 427413 70488 427481
rect 70000 427357 70047 427413
rect 70103 427357 70171 427413
rect 70227 427357 70295 427413
rect 70351 427357 70419 427413
rect 70475 427357 70488 427413
rect 70000 427289 70488 427357
rect 70000 427233 70047 427289
rect 70103 427233 70171 427289
rect 70227 427233 70295 427289
rect 70351 427233 70419 427289
rect 70475 427233 70488 427289
rect 70000 427165 70488 427233
rect 70000 427109 70047 427165
rect 70103 427109 70171 427165
rect 70227 427109 70295 427165
rect 70351 427109 70419 427165
rect 70475 427109 70488 427165
rect 70000 427041 70488 427109
rect 70000 426985 70047 427041
rect 70103 426985 70171 427041
rect 70227 426985 70295 427041
rect 70351 426985 70419 427041
rect 70475 426985 70488 427041
rect 70000 426917 70488 426985
rect 70000 426861 70047 426917
rect 70103 426861 70171 426917
rect 70227 426861 70295 426917
rect 70351 426861 70419 426917
rect 70475 426861 70488 426917
rect 70000 426793 70488 426861
rect 70000 426737 70047 426793
rect 70103 426737 70171 426793
rect 70227 426737 70295 426793
rect 70351 426737 70419 426793
rect 70475 426737 70488 426793
rect 70000 426669 70488 426737
rect 70000 426613 70047 426669
rect 70103 426613 70171 426669
rect 70227 426613 70295 426669
rect 70351 426613 70419 426669
rect 70475 426613 70488 426669
rect 70000 426545 70488 426613
rect 70000 426489 70047 426545
rect 70103 426489 70171 426545
rect 70227 426489 70295 426545
rect 70351 426489 70419 426545
rect 70475 426489 70488 426545
rect 70000 426421 70488 426489
rect 70000 426365 70047 426421
rect 70103 426365 70171 426421
rect 70227 426365 70295 426421
rect 70351 426365 70419 426421
rect 70475 426365 70488 426421
rect 70000 426297 70488 426365
rect 70000 426241 70047 426297
rect 70103 426241 70171 426297
rect 70227 426241 70295 426297
rect 70351 426241 70419 426297
rect 70475 426241 70488 426297
rect 70000 426173 70488 426241
rect 70000 426117 70047 426173
rect 70103 426117 70171 426173
rect 70227 426117 70295 426173
rect 70351 426117 70419 426173
rect 70475 426117 70488 426173
rect 70000 426049 70488 426117
rect 70000 425993 70047 426049
rect 70103 425993 70171 426049
rect 70227 425993 70295 426049
rect 70351 425993 70419 426049
rect 70475 425993 70488 426049
rect 70000 425925 70488 425993
rect 70000 425869 70047 425925
rect 70103 425869 70171 425925
rect 70227 425869 70295 425925
rect 70351 425869 70419 425925
rect 70475 425869 70488 425925
rect 70000 425828 70488 425869
rect 70000 425181 70488 425248
rect 70000 425125 70047 425181
rect 70103 425125 70171 425181
rect 70227 425125 70295 425181
rect 70351 425125 70419 425181
rect 70475 425125 70488 425181
rect 70000 425057 70488 425125
rect 70000 425001 70047 425057
rect 70103 425001 70171 425057
rect 70227 425001 70295 425057
rect 70351 425001 70419 425057
rect 70475 425001 70488 425057
rect 70000 424933 70488 425001
rect 70000 424877 70047 424933
rect 70103 424877 70171 424933
rect 70227 424877 70295 424933
rect 70351 424877 70419 424933
rect 70475 424877 70488 424933
rect 70000 424809 70488 424877
rect 70000 424753 70047 424809
rect 70103 424753 70171 424809
rect 70227 424753 70295 424809
rect 70351 424753 70419 424809
rect 70475 424753 70488 424809
rect 70000 424685 70488 424753
rect 70000 424629 70047 424685
rect 70103 424629 70171 424685
rect 70227 424629 70295 424685
rect 70351 424629 70419 424685
rect 70475 424629 70488 424685
rect 70000 424561 70488 424629
rect 70000 424505 70047 424561
rect 70103 424505 70171 424561
rect 70227 424505 70295 424561
rect 70351 424505 70419 424561
rect 70475 424505 70488 424561
rect 70000 424437 70488 424505
rect 70000 424381 70047 424437
rect 70103 424381 70171 424437
rect 70227 424381 70295 424437
rect 70351 424381 70419 424437
rect 70475 424381 70488 424437
rect 70000 424313 70488 424381
rect 70000 424257 70047 424313
rect 70103 424257 70171 424313
rect 70227 424257 70295 424313
rect 70351 424257 70419 424313
rect 70475 424257 70488 424313
rect 70000 424189 70488 424257
rect 70000 424133 70047 424189
rect 70103 424133 70171 424189
rect 70227 424133 70295 424189
rect 70351 424133 70419 424189
rect 70475 424133 70488 424189
rect 70000 424065 70488 424133
rect 70000 424009 70047 424065
rect 70103 424009 70171 424065
rect 70227 424009 70295 424065
rect 70351 424009 70419 424065
rect 70475 424009 70488 424065
rect 70000 423941 70488 424009
rect 70000 423885 70047 423941
rect 70103 423885 70171 423941
rect 70227 423885 70295 423941
rect 70351 423885 70419 423941
rect 70475 423885 70488 423941
rect 70000 423817 70488 423885
rect 70000 423761 70047 423817
rect 70103 423761 70171 423817
rect 70227 423761 70295 423817
rect 70351 423761 70419 423817
rect 70475 423761 70488 423817
rect 70000 423693 70488 423761
rect 70000 423637 70047 423693
rect 70103 423637 70171 423693
rect 70227 423637 70295 423693
rect 70351 423637 70419 423693
rect 70475 423637 70488 423693
rect 70000 423569 70488 423637
rect 70000 423513 70047 423569
rect 70103 423513 70171 423569
rect 70227 423513 70295 423569
rect 70351 423513 70419 423569
rect 70475 423513 70488 423569
rect 70000 423445 70488 423513
rect 70000 423389 70047 423445
rect 70103 423389 70171 423445
rect 70227 423389 70295 423445
rect 70351 423389 70419 423445
rect 70475 423389 70488 423445
rect 70000 423321 70488 423389
rect 70000 423265 70047 423321
rect 70103 423265 70171 423321
rect 70227 423265 70295 423321
rect 70351 423265 70419 423321
rect 70475 423265 70488 423321
rect 70000 423198 70488 423265
rect 70000 422811 70488 422878
rect 70000 422755 70047 422811
rect 70103 422755 70171 422811
rect 70227 422755 70295 422811
rect 70351 422755 70419 422811
rect 70475 422755 70488 422811
rect 70000 422687 70488 422755
rect 70000 422631 70047 422687
rect 70103 422631 70171 422687
rect 70227 422631 70295 422687
rect 70351 422631 70419 422687
rect 70475 422631 70488 422687
rect 70000 422563 70488 422631
rect 70000 422507 70047 422563
rect 70103 422507 70171 422563
rect 70227 422507 70295 422563
rect 70351 422507 70419 422563
rect 70475 422507 70488 422563
rect 70000 422439 70488 422507
rect 70000 422383 70047 422439
rect 70103 422383 70171 422439
rect 70227 422383 70295 422439
rect 70351 422383 70419 422439
rect 70475 422383 70488 422439
rect 70000 422315 70488 422383
rect 70000 422259 70047 422315
rect 70103 422259 70171 422315
rect 70227 422259 70295 422315
rect 70351 422259 70419 422315
rect 70475 422259 70488 422315
rect 70000 422191 70488 422259
rect 70000 422135 70047 422191
rect 70103 422135 70171 422191
rect 70227 422135 70295 422191
rect 70351 422135 70419 422191
rect 70475 422135 70488 422191
rect 70000 422067 70488 422135
rect 70000 422011 70047 422067
rect 70103 422011 70171 422067
rect 70227 422011 70295 422067
rect 70351 422011 70419 422067
rect 70475 422011 70488 422067
rect 70000 421943 70488 422011
rect 70000 421887 70047 421943
rect 70103 421887 70171 421943
rect 70227 421887 70295 421943
rect 70351 421887 70419 421943
rect 70475 421887 70488 421943
rect 70000 421819 70488 421887
rect 70000 421763 70047 421819
rect 70103 421763 70171 421819
rect 70227 421763 70295 421819
rect 70351 421763 70419 421819
rect 70475 421763 70488 421819
rect 70000 421695 70488 421763
rect 70000 421639 70047 421695
rect 70103 421639 70171 421695
rect 70227 421639 70295 421695
rect 70351 421639 70419 421695
rect 70475 421639 70488 421695
rect 70000 421571 70488 421639
rect 70000 421515 70047 421571
rect 70103 421515 70171 421571
rect 70227 421515 70295 421571
rect 70351 421515 70419 421571
rect 70475 421515 70488 421571
rect 70000 421447 70488 421515
rect 70000 421391 70047 421447
rect 70103 421391 70171 421447
rect 70227 421391 70295 421447
rect 70351 421391 70419 421447
rect 70475 421391 70488 421447
rect 70000 421323 70488 421391
rect 70000 421267 70047 421323
rect 70103 421267 70171 421323
rect 70227 421267 70295 421323
rect 70351 421267 70419 421323
rect 70475 421267 70488 421323
rect 70000 421199 70488 421267
rect 70000 421143 70047 421199
rect 70103 421143 70171 421199
rect 70227 421143 70295 421199
rect 70351 421143 70419 421199
rect 70475 421143 70488 421199
rect 70000 421075 70488 421143
rect 70000 421019 70047 421075
rect 70103 421019 70171 421075
rect 70227 421019 70295 421075
rect 70351 421019 70419 421075
rect 70475 421019 70488 421075
rect 70000 420951 70488 421019
rect 70000 420895 70047 420951
rect 70103 420895 70171 420951
rect 70227 420895 70295 420951
rect 70351 420895 70419 420951
rect 70475 420895 70488 420951
rect 70000 420828 70488 420895
rect 70000 420105 70488 420172
rect 70000 420049 70047 420105
rect 70103 420049 70171 420105
rect 70227 420049 70295 420105
rect 70351 420049 70419 420105
rect 70475 420049 70488 420105
rect 70000 419981 70488 420049
rect 70000 419925 70047 419981
rect 70103 419925 70171 419981
rect 70227 419925 70295 419981
rect 70351 419925 70419 419981
rect 70475 419925 70488 419981
rect 70000 419857 70488 419925
rect 70000 419801 70047 419857
rect 70103 419801 70171 419857
rect 70227 419801 70295 419857
rect 70351 419801 70419 419857
rect 70475 419801 70488 419857
rect 70000 419733 70488 419801
rect 70000 419677 70047 419733
rect 70103 419677 70171 419733
rect 70227 419677 70295 419733
rect 70351 419677 70419 419733
rect 70475 419677 70488 419733
rect 70000 419609 70488 419677
rect 70000 419553 70047 419609
rect 70103 419553 70171 419609
rect 70227 419553 70295 419609
rect 70351 419553 70419 419609
rect 70475 419553 70488 419609
rect 70000 419485 70488 419553
rect 70000 419429 70047 419485
rect 70103 419429 70171 419485
rect 70227 419429 70295 419485
rect 70351 419429 70419 419485
rect 70475 419429 70488 419485
rect 70000 419361 70488 419429
rect 70000 419305 70047 419361
rect 70103 419305 70171 419361
rect 70227 419305 70295 419361
rect 70351 419305 70419 419361
rect 70475 419305 70488 419361
rect 70000 419237 70488 419305
rect 70000 419181 70047 419237
rect 70103 419181 70171 419237
rect 70227 419181 70295 419237
rect 70351 419181 70419 419237
rect 70475 419181 70488 419237
rect 70000 419113 70488 419181
rect 70000 419057 70047 419113
rect 70103 419057 70171 419113
rect 70227 419057 70295 419113
rect 70351 419057 70419 419113
rect 70475 419057 70488 419113
rect 70000 418989 70488 419057
rect 70000 418933 70047 418989
rect 70103 418933 70171 418989
rect 70227 418933 70295 418989
rect 70351 418933 70419 418989
rect 70475 418933 70488 418989
rect 70000 418865 70488 418933
rect 70000 418809 70047 418865
rect 70103 418809 70171 418865
rect 70227 418809 70295 418865
rect 70351 418809 70419 418865
rect 70475 418809 70488 418865
rect 70000 418741 70488 418809
rect 70000 418685 70047 418741
rect 70103 418685 70171 418741
rect 70227 418685 70295 418741
rect 70351 418685 70419 418741
rect 70475 418685 70488 418741
rect 70000 418617 70488 418685
rect 70000 418561 70047 418617
rect 70103 418561 70171 418617
rect 70227 418561 70295 418617
rect 70351 418561 70419 418617
rect 70475 418561 70488 418617
rect 70000 418493 70488 418561
rect 70000 418437 70047 418493
rect 70103 418437 70171 418493
rect 70227 418437 70295 418493
rect 70351 418437 70419 418493
rect 70475 418437 70488 418493
rect 70000 418369 70488 418437
rect 70000 418313 70047 418369
rect 70103 418313 70171 418369
rect 70227 418313 70295 418369
rect 70351 418313 70419 418369
rect 70475 418313 70488 418369
rect 70000 418245 70488 418313
rect 70000 418189 70047 418245
rect 70103 418189 70171 418245
rect 70227 418189 70295 418245
rect 70351 418189 70419 418245
rect 70475 418189 70488 418245
rect 70000 418122 70488 418189
rect 70000 417735 70488 417802
rect 70000 417679 70047 417735
rect 70103 417679 70171 417735
rect 70227 417679 70295 417735
rect 70351 417679 70419 417735
rect 70475 417679 70488 417735
rect 70000 417611 70488 417679
rect 70000 417555 70047 417611
rect 70103 417555 70171 417611
rect 70227 417555 70295 417611
rect 70351 417555 70419 417611
rect 70475 417555 70488 417611
rect 70000 417487 70488 417555
rect 70000 417431 70047 417487
rect 70103 417431 70171 417487
rect 70227 417431 70295 417487
rect 70351 417431 70419 417487
rect 70475 417431 70488 417487
rect 70000 417363 70488 417431
rect 70000 417307 70047 417363
rect 70103 417307 70171 417363
rect 70227 417307 70295 417363
rect 70351 417307 70419 417363
rect 70475 417307 70488 417363
rect 70000 417239 70488 417307
rect 70000 417183 70047 417239
rect 70103 417183 70171 417239
rect 70227 417183 70295 417239
rect 70351 417183 70419 417239
rect 70475 417183 70488 417239
rect 70000 417115 70488 417183
rect 70000 417059 70047 417115
rect 70103 417059 70171 417115
rect 70227 417059 70295 417115
rect 70351 417059 70419 417115
rect 70475 417059 70488 417115
rect 70000 416991 70488 417059
rect 70000 416935 70047 416991
rect 70103 416935 70171 416991
rect 70227 416935 70295 416991
rect 70351 416935 70419 416991
rect 70475 416935 70488 416991
rect 70000 416867 70488 416935
rect 70000 416811 70047 416867
rect 70103 416811 70171 416867
rect 70227 416811 70295 416867
rect 70351 416811 70419 416867
rect 70475 416811 70488 416867
rect 70000 416743 70488 416811
rect 70000 416687 70047 416743
rect 70103 416687 70171 416743
rect 70227 416687 70295 416743
rect 70351 416687 70419 416743
rect 70475 416687 70488 416743
rect 70000 416619 70488 416687
rect 70000 416563 70047 416619
rect 70103 416563 70171 416619
rect 70227 416563 70295 416619
rect 70351 416563 70419 416619
rect 70475 416563 70488 416619
rect 70000 416495 70488 416563
rect 70000 416439 70047 416495
rect 70103 416439 70171 416495
rect 70227 416439 70295 416495
rect 70351 416439 70419 416495
rect 70475 416439 70488 416495
rect 70000 416371 70488 416439
rect 70000 416315 70047 416371
rect 70103 416315 70171 416371
rect 70227 416315 70295 416371
rect 70351 416315 70419 416371
rect 70475 416315 70488 416371
rect 70000 416247 70488 416315
rect 70000 416191 70047 416247
rect 70103 416191 70171 416247
rect 70227 416191 70295 416247
rect 70351 416191 70419 416247
rect 70475 416191 70488 416247
rect 70000 416123 70488 416191
rect 70000 416067 70047 416123
rect 70103 416067 70171 416123
rect 70227 416067 70295 416123
rect 70351 416067 70419 416123
rect 70475 416067 70488 416123
rect 70000 415999 70488 416067
rect 70000 415943 70047 415999
rect 70103 415943 70171 415999
rect 70227 415943 70295 415999
rect 70351 415943 70419 415999
rect 70475 415943 70488 415999
rect 70000 415875 70488 415943
rect 70000 415819 70047 415875
rect 70103 415819 70171 415875
rect 70227 415819 70295 415875
rect 70351 415819 70419 415875
rect 70475 415819 70488 415875
rect 70000 415752 70488 415819
rect 70000 415105 70488 415172
rect 70000 415049 70047 415105
rect 70103 415049 70171 415105
rect 70227 415049 70295 415105
rect 70351 415049 70419 415105
rect 70475 415049 70488 415105
rect 70000 414981 70488 415049
rect 70000 414925 70047 414981
rect 70103 414925 70171 414981
rect 70227 414925 70295 414981
rect 70351 414925 70419 414981
rect 70475 414925 70488 414981
rect 70000 414857 70488 414925
rect 70000 414801 70047 414857
rect 70103 414801 70171 414857
rect 70227 414801 70295 414857
rect 70351 414801 70419 414857
rect 70475 414801 70488 414857
rect 70000 414733 70488 414801
rect 70000 414677 70047 414733
rect 70103 414677 70171 414733
rect 70227 414677 70295 414733
rect 70351 414677 70419 414733
rect 70475 414677 70488 414733
rect 70000 414609 70488 414677
rect 70000 414553 70047 414609
rect 70103 414553 70171 414609
rect 70227 414553 70295 414609
rect 70351 414553 70419 414609
rect 70475 414553 70488 414609
rect 70000 414485 70488 414553
rect 70000 414429 70047 414485
rect 70103 414429 70171 414485
rect 70227 414429 70295 414485
rect 70351 414429 70419 414485
rect 70475 414429 70488 414485
rect 70000 414361 70488 414429
rect 70000 414305 70047 414361
rect 70103 414305 70171 414361
rect 70227 414305 70295 414361
rect 70351 414305 70419 414361
rect 70475 414305 70488 414361
rect 70000 414237 70488 414305
rect 70000 414181 70047 414237
rect 70103 414181 70171 414237
rect 70227 414181 70295 414237
rect 70351 414181 70419 414237
rect 70475 414181 70488 414237
rect 70000 414113 70488 414181
rect 70000 414057 70047 414113
rect 70103 414057 70171 414113
rect 70227 414057 70295 414113
rect 70351 414057 70419 414113
rect 70475 414057 70488 414113
rect 70000 413989 70488 414057
rect 70000 413933 70047 413989
rect 70103 413933 70171 413989
rect 70227 413933 70295 413989
rect 70351 413933 70419 413989
rect 70475 413933 70488 413989
rect 70000 413865 70488 413933
rect 70000 413809 70047 413865
rect 70103 413809 70171 413865
rect 70227 413809 70295 413865
rect 70351 413809 70419 413865
rect 70475 413809 70488 413865
rect 70000 413741 70488 413809
rect 70000 413685 70047 413741
rect 70103 413685 70171 413741
rect 70227 413685 70295 413741
rect 70351 413685 70419 413741
rect 70475 413685 70488 413741
rect 70000 413617 70488 413685
rect 70000 413561 70047 413617
rect 70103 413561 70171 413617
rect 70227 413561 70295 413617
rect 70351 413561 70419 413617
rect 70475 413561 70488 413617
rect 70000 413493 70488 413561
rect 70000 413437 70047 413493
rect 70103 413437 70171 413493
rect 70227 413437 70295 413493
rect 70351 413437 70419 413493
rect 70475 413437 70488 413493
rect 70000 413369 70488 413437
rect 70000 413313 70047 413369
rect 70103 413313 70171 413369
rect 70227 413313 70295 413369
rect 70351 413313 70419 413369
rect 70475 413313 70488 413369
rect 70000 413272 70488 413313
rect 705512 404687 706000 404728
rect 705512 404631 705525 404687
rect 705581 404631 705649 404687
rect 705705 404631 705773 404687
rect 705829 404631 705897 404687
rect 705953 404631 706000 404687
rect 705512 404563 706000 404631
rect 705512 404507 705525 404563
rect 705581 404507 705649 404563
rect 705705 404507 705773 404563
rect 705829 404507 705897 404563
rect 705953 404507 706000 404563
rect 705512 404439 706000 404507
rect 705512 404383 705525 404439
rect 705581 404383 705649 404439
rect 705705 404383 705773 404439
rect 705829 404383 705897 404439
rect 705953 404383 706000 404439
rect 705512 404315 706000 404383
rect 705512 404259 705525 404315
rect 705581 404259 705649 404315
rect 705705 404259 705773 404315
rect 705829 404259 705897 404315
rect 705953 404259 706000 404315
rect 705512 404191 706000 404259
rect 705512 404135 705525 404191
rect 705581 404135 705649 404191
rect 705705 404135 705773 404191
rect 705829 404135 705897 404191
rect 705953 404135 706000 404191
rect 705512 404067 706000 404135
rect 705512 404011 705525 404067
rect 705581 404011 705649 404067
rect 705705 404011 705773 404067
rect 705829 404011 705897 404067
rect 705953 404011 706000 404067
rect 705512 403943 706000 404011
rect 705512 403887 705525 403943
rect 705581 403887 705649 403943
rect 705705 403887 705773 403943
rect 705829 403887 705897 403943
rect 705953 403887 706000 403943
rect 705512 403819 706000 403887
rect 705512 403763 705525 403819
rect 705581 403763 705649 403819
rect 705705 403763 705773 403819
rect 705829 403763 705897 403819
rect 705953 403763 706000 403819
rect 705512 403695 706000 403763
rect 705512 403639 705525 403695
rect 705581 403639 705649 403695
rect 705705 403639 705773 403695
rect 705829 403639 705897 403695
rect 705953 403639 706000 403695
rect 705512 403571 706000 403639
rect 705512 403515 705525 403571
rect 705581 403515 705649 403571
rect 705705 403515 705773 403571
rect 705829 403515 705897 403571
rect 705953 403515 706000 403571
rect 705512 403447 706000 403515
rect 705512 403391 705525 403447
rect 705581 403391 705649 403447
rect 705705 403391 705773 403447
rect 705829 403391 705897 403447
rect 705953 403391 706000 403447
rect 705512 403323 706000 403391
rect 705512 403267 705525 403323
rect 705581 403267 705649 403323
rect 705705 403267 705773 403323
rect 705829 403267 705897 403323
rect 705953 403267 706000 403323
rect 705512 403199 706000 403267
rect 705512 403143 705525 403199
rect 705581 403143 705649 403199
rect 705705 403143 705773 403199
rect 705829 403143 705897 403199
rect 705953 403143 706000 403199
rect 705512 403075 706000 403143
rect 705512 403019 705525 403075
rect 705581 403019 705649 403075
rect 705705 403019 705773 403075
rect 705829 403019 705897 403075
rect 705953 403019 706000 403075
rect 705512 402951 706000 403019
rect 705512 402895 705525 402951
rect 705581 402895 705649 402951
rect 705705 402895 705773 402951
rect 705829 402895 705897 402951
rect 705953 402895 706000 402951
rect 705512 402828 706000 402895
rect 705512 402181 706000 402248
rect 705512 402125 705525 402181
rect 705581 402125 705649 402181
rect 705705 402125 705773 402181
rect 705829 402125 705897 402181
rect 705953 402125 706000 402181
rect 705512 402057 706000 402125
rect 705512 402001 705525 402057
rect 705581 402001 705649 402057
rect 705705 402001 705773 402057
rect 705829 402001 705897 402057
rect 705953 402001 706000 402057
rect 705512 401933 706000 402001
rect 705512 401877 705525 401933
rect 705581 401877 705649 401933
rect 705705 401877 705773 401933
rect 705829 401877 705897 401933
rect 705953 401877 706000 401933
rect 705512 401809 706000 401877
rect 705512 401753 705525 401809
rect 705581 401753 705649 401809
rect 705705 401753 705773 401809
rect 705829 401753 705897 401809
rect 705953 401753 706000 401809
rect 705512 401685 706000 401753
rect 705512 401629 705525 401685
rect 705581 401629 705649 401685
rect 705705 401629 705773 401685
rect 705829 401629 705897 401685
rect 705953 401629 706000 401685
rect 705512 401561 706000 401629
rect 705512 401505 705525 401561
rect 705581 401505 705649 401561
rect 705705 401505 705773 401561
rect 705829 401505 705897 401561
rect 705953 401505 706000 401561
rect 705512 401437 706000 401505
rect 705512 401381 705525 401437
rect 705581 401381 705649 401437
rect 705705 401381 705773 401437
rect 705829 401381 705897 401437
rect 705953 401381 706000 401437
rect 705512 401313 706000 401381
rect 705512 401257 705525 401313
rect 705581 401257 705649 401313
rect 705705 401257 705773 401313
rect 705829 401257 705897 401313
rect 705953 401257 706000 401313
rect 705512 401189 706000 401257
rect 705512 401133 705525 401189
rect 705581 401133 705649 401189
rect 705705 401133 705773 401189
rect 705829 401133 705897 401189
rect 705953 401133 706000 401189
rect 705512 401065 706000 401133
rect 705512 401009 705525 401065
rect 705581 401009 705649 401065
rect 705705 401009 705773 401065
rect 705829 401009 705897 401065
rect 705953 401009 706000 401065
rect 705512 400941 706000 401009
rect 705512 400885 705525 400941
rect 705581 400885 705649 400941
rect 705705 400885 705773 400941
rect 705829 400885 705897 400941
rect 705953 400885 706000 400941
rect 705512 400817 706000 400885
rect 705512 400761 705525 400817
rect 705581 400761 705649 400817
rect 705705 400761 705773 400817
rect 705829 400761 705897 400817
rect 705953 400761 706000 400817
rect 705512 400693 706000 400761
rect 705512 400637 705525 400693
rect 705581 400637 705649 400693
rect 705705 400637 705773 400693
rect 705829 400637 705897 400693
rect 705953 400637 706000 400693
rect 705512 400569 706000 400637
rect 705512 400513 705525 400569
rect 705581 400513 705649 400569
rect 705705 400513 705773 400569
rect 705829 400513 705897 400569
rect 705953 400513 706000 400569
rect 705512 400445 706000 400513
rect 705512 400389 705525 400445
rect 705581 400389 705649 400445
rect 705705 400389 705773 400445
rect 705829 400389 705897 400445
rect 705953 400389 706000 400445
rect 705512 400321 706000 400389
rect 705512 400265 705525 400321
rect 705581 400265 705649 400321
rect 705705 400265 705773 400321
rect 705829 400265 705897 400321
rect 705953 400265 706000 400321
rect 705512 400198 706000 400265
rect 705512 399811 706000 399878
rect 705512 399755 705525 399811
rect 705581 399755 705649 399811
rect 705705 399755 705773 399811
rect 705829 399755 705897 399811
rect 705953 399755 706000 399811
rect 705512 399687 706000 399755
rect 705512 399631 705525 399687
rect 705581 399631 705649 399687
rect 705705 399631 705773 399687
rect 705829 399631 705897 399687
rect 705953 399631 706000 399687
rect 705512 399563 706000 399631
rect 705512 399507 705525 399563
rect 705581 399507 705649 399563
rect 705705 399507 705773 399563
rect 705829 399507 705897 399563
rect 705953 399507 706000 399563
rect 705512 399439 706000 399507
rect 705512 399383 705525 399439
rect 705581 399383 705649 399439
rect 705705 399383 705773 399439
rect 705829 399383 705897 399439
rect 705953 399383 706000 399439
rect 705512 399315 706000 399383
rect 705512 399259 705525 399315
rect 705581 399259 705649 399315
rect 705705 399259 705773 399315
rect 705829 399259 705897 399315
rect 705953 399259 706000 399315
rect 705512 399191 706000 399259
rect 705512 399135 705525 399191
rect 705581 399135 705649 399191
rect 705705 399135 705773 399191
rect 705829 399135 705897 399191
rect 705953 399135 706000 399191
rect 705512 399067 706000 399135
rect 705512 399011 705525 399067
rect 705581 399011 705649 399067
rect 705705 399011 705773 399067
rect 705829 399011 705897 399067
rect 705953 399011 706000 399067
rect 705512 398943 706000 399011
rect 705512 398887 705525 398943
rect 705581 398887 705649 398943
rect 705705 398887 705773 398943
rect 705829 398887 705897 398943
rect 705953 398887 706000 398943
rect 705512 398819 706000 398887
rect 705512 398763 705525 398819
rect 705581 398763 705649 398819
rect 705705 398763 705773 398819
rect 705829 398763 705897 398819
rect 705953 398763 706000 398819
rect 705512 398695 706000 398763
rect 705512 398639 705525 398695
rect 705581 398639 705649 398695
rect 705705 398639 705773 398695
rect 705829 398639 705897 398695
rect 705953 398639 706000 398695
rect 705512 398571 706000 398639
rect 705512 398515 705525 398571
rect 705581 398515 705649 398571
rect 705705 398515 705773 398571
rect 705829 398515 705897 398571
rect 705953 398515 706000 398571
rect 705512 398447 706000 398515
rect 705512 398391 705525 398447
rect 705581 398391 705649 398447
rect 705705 398391 705773 398447
rect 705829 398391 705897 398447
rect 705953 398391 706000 398447
rect 705512 398323 706000 398391
rect 705512 398267 705525 398323
rect 705581 398267 705649 398323
rect 705705 398267 705773 398323
rect 705829 398267 705897 398323
rect 705953 398267 706000 398323
rect 705512 398199 706000 398267
rect 705512 398143 705525 398199
rect 705581 398143 705649 398199
rect 705705 398143 705773 398199
rect 705829 398143 705897 398199
rect 705953 398143 706000 398199
rect 705512 398075 706000 398143
rect 705512 398019 705525 398075
rect 705581 398019 705649 398075
rect 705705 398019 705773 398075
rect 705829 398019 705897 398075
rect 705953 398019 706000 398075
rect 705512 397951 706000 398019
rect 705512 397895 705525 397951
rect 705581 397895 705649 397951
rect 705705 397895 705773 397951
rect 705829 397895 705897 397951
rect 705953 397895 706000 397951
rect 705512 397828 706000 397895
rect 705512 397105 706000 397172
rect 705512 397049 705525 397105
rect 705581 397049 705649 397105
rect 705705 397049 705773 397105
rect 705829 397049 705897 397105
rect 705953 397049 706000 397105
rect 705512 396981 706000 397049
rect 705512 396925 705525 396981
rect 705581 396925 705649 396981
rect 705705 396925 705773 396981
rect 705829 396925 705897 396981
rect 705953 396925 706000 396981
rect 705512 396857 706000 396925
rect 705512 396801 705525 396857
rect 705581 396801 705649 396857
rect 705705 396801 705773 396857
rect 705829 396801 705897 396857
rect 705953 396801 706000 396857
rect 705512 396733 706000 396801
rect 705512 396677 705525 396733
rect 705581 396677 705649 396733
rect 705705 396677 705773 396733
rect 705829 396677 705897 396733
rect 705953 396677 706000 396733
rect 705512 396609 706000 396677
rect 705512 396553 705525 396609
rect 705581 396553 705649 396609
rect 705705 396553 705773 396609
rect 705829 396553 705897 396609
rect 705953 396553 706000 396609
rect 705512 396485 706000 396553
rect 705512 396429 705525 396485
rect 705581 396429 705649 396485
rect 705705 396429 705773 396485
rect 705829 396429 705897 396485
rect 705953 396429 706000 396485
rect 705512 396361 706000 396429
rect 705512 396305 705525 396361
rect 705581 396305 705649 396361
rect 705705 396305 705773 396361
rect 705829 396305 705897 396361
rect 705953 396305 706000 396361
rect 705512 396237 706000 396305
rect 705512 396181 705525 396237
rect 705581 396181 705649 396237
rect 705705 396181 705773 396237
rect 705829 396181 705897 396237
rect 705953 396181 706000 396237
rect 705512 396113 706000 396181
rect 705512 396057 705525 396113
rect 705581 396057 705649 396113
rect 705705 396057 705773 396113
rect 705829 396057 705897 396113
rect 705953 396057 706000 396113
rect 705512 395989 706000 396057
rect 705512 395933 705525 395989
rect 705581 395933 705649 395989
rect 705705 395933 705773 395989
rect 705829 395933 705897 395989
rect 705953 395933 706000 395989
rect 705512 395865 706000 395933
rect 705512 395809 705525 395865
rect 705581 395809 705649 395865
rect 705705 395809 705773 395865
rect 705829 395809 705897 395865
rect 705953 395809 706000 395865
rect 705512 395741 706000 395809
rect 705512 395685 705525 395741
rect 705581 395685 705649 395741
rect 705705 395685 705773 395741
rect 705829 395685 705897 395741
rect 705953 395685 706000 395741
rect 705512 395617 706000 395685
rect 705512 395561 705525 395617
rect 705581 395561 705649 395617
rect 705705 395561 705773 395617
rect 705829 395561 705897 395617
rect 705953 395561 706000 395617
rect 705512 395493 706000 395561
rect 705512 395437 705525 395493
rect 705581 395437 705649 395493
rect 705705 395437 705773 395493
rect 705829 395437 705897 395493
rect 705953 395437 706000 395493
rect 705512 395369 706000 395437
rect 705512 395313 705525 395369
rect 705581 395313 705649 395369
rect 705705 395313 705773 395369
rect 705829 395313 705897 395369
rect 705953 395313 706000 395369
rect 705512 395245 706000 395313
rect 705512 395189 705525 395245
rect 705581 395189 705649 395245
rect 705705 395189 705773 395245
rect 705829 395189 705897 395245
rect 705953 395189 706000 395245
rect 705512 395122 706000 395189
rect 705512 394735 706000 394802
rect 705512 394679 705525 394735
rect 705581 394679 705649 394735
rect 705705 394679 705773 394735
rect 705829 394679 705897 394735
rect 705953 394679 706000 394735
rect 705512 394611 706000 394679
rect 705512 394555 705525 394611
rect 705581 394555 705649 394611
rect 705705 394555 705773 394611
rect 705829 394555 705897 394611
rect 705953 394555 706000 394611
rect 705512 394487 706000 394555
rect 705512 394431 705525 394487
rect 705581 394431 705649 394487
rect 705705 394431 705773 394487
rect 705829 394431 705897 394487
rect 705953 394431 706000 394487
rect 705512 394363 706000 394431
rect 705512 394307 705525 394363
rect 705581 394307 705649 394363
rect 705705 394307 705773 394363
rect 705829 394307 705897 394363
rect 705953 394307 706000 394363
rect 705512 394239 706000 394307
rect 705512 394183 705525 394239
rect 705581 394183 705649 394239
rect 705705 394183 705773 394239
rect 705829 394183 705897 394239
rect 705953 394183 706000 394239
rect 705512 394115 706000 394183
rect 705512 394059 705525 394115
rect 705581 394059 705649 394115
rect 705705 394059 705773 394115
rect 705829 394059 705897 394115
rect 705953 394059 706000 394115
rect 705512 393991 706000 394059
rect 705512 393935 705525 393991
rect 705581 393935 705649 393991
rect 705705 393935 705773 393991
rect 705829 393935 705897 393991
rect 705953 393935 706000 393991
rect 705512 393867 706000 393935
rect 705512 393811 705525 393867
rect 705581 393811 705649 393867
rect 705705 393811 705773 393867
rect 705829 393811 705897 393867
rect 705953 393811 706000 393867
rect 705512 393743 706000 393811
rect 705512 393687 705525 393743
rect 705581 393687 705649 393743
rect 705705 393687 705773 393743
rect 705829 393687 705897 393743
rect 705953 393687 706000 393743
rect 705512 393619 706000 393687
rect 705512 393563 705525 393619
rect 705581 393563 705649 393619
rect 705705 393563 705773 393619
rect 705829 393563 705897 393619
rect 705953 393563 706000 393619
rect 705512 393495 706000 393563
rect 705512 393439 705525 393495
rect 705581 393439 705649 393495
rect 705705 393439 705773 393495
rect 705829 393439 705897 393495
rect 705953 393439 706000 393495
rect 705512 393371 706000 393439
rect 705512 393315 705525 393371
rect 705581 393315 705649 393371
rect 705705 393315 705773 393371
rect 705829 393315 705897 393371
rect 705953 393315 706000 393371
rect 705512 393247 706000 393315
rect 705512 393191 705525 393247
rect 705581 393191 705649 393247
rect 705705 393191 705773 393247
rect 705829 393191 705897 393247
rect 705953 393191 706000 393247
rect 705512 393123 706000 393191
rect 705512 393067 705525 393123
rect 705581 393067 705649 393123
rect 705705 393067 705773 393123
rect 705829 393067 705897 393123
rect 705953 393067 706000 393123
rect 705512 392999 706000 393067
rect 705512 392943 705525 392999
rect 705581 392943 705649 392999
rect 705705 392943 705773 392999
rect 705829 392943 705897 392999
rect 705953 392943 706000 392999
rect 705512 392875 706000 392943
rect 705512 392819 705525 392875
rect 705581 392819 705649 392875
rect 705705 392819 705773 392875
rect 705829 392819 705897 392875
rect 705953 392819 706000 392875
rect 705512 392752 706000 392819
rect 705512 392131 706000 392172
rect 705512 392075 705525 392131
rect 705581 392075 705649 392131
rect 705705 392075 705773 392131
rect 705829 392075 705897 392131
rect 705953 392075 706000 392131
rect 705512 392007 706000 392075
rect 705512 391951 705525 392007
rect 705581 391951 705649 392007
rect 705705 391951 705773 392007
rect 705829 391951 705897 392007
rect 705953 391951 706000 392007
rect 705512 391883 706000 391951
rect 705512 391827 705525 391883
rect 705581 391827 705649 391883
rect 705705 391827 705773 391883
rect 705829 391827 705897 391883
rect 705953 391827 706000 391883
rect 705512 391759 706000 391827
rect 705512 391703 705525 391759
rect 705581 391703 705649 391759
rect 705705 391703 705773 391759
rect 705829 391703 705897 391759
rect 705953 391703 706000 391759
rect 705512 391635 706000 391703
rect 705512 391579 705525 391635
rect 705581 391579 705649 391635
rect 705705 391579 705773 391635
rect 705829 391579 705897 391635
rect 705953 391579 706000 391635
rect 705512 391511 706000 391579
rect 705512 391455 705525 391511
rect 705581 391455 705649 391511
rect 705705 391455 705773 391511
rect 705829 391455 705897 391511
rect 705953 391455 706000 391511
rect 705512 391387 706000 391455
rect 705512 391331 705525 391387
rect 705581 391331 705649 391387
rect 705705 391331 705773 391387
rect 705829 391331 705897 391387
rect 705953 391331 706000 391387
rect 705512 391263 706000 391331
rect 705512 391207 705525 391263
rect 705581 391207 705649 391263
rect 705705 391207 705773 391263
rect 705829 391207 705897 391263
rect 705953 391207 706000 391263
rect 705512 391139 706000 391207
rect 705512 391083 705525 391139
rect 705581 391083 705649 391139
rect 705705 391083 705773 391139
rect 705829 391083 705897 391139
rect 705953 391083 706000 391139
rect 705512 391015 706000 391083
rect 705512 390959 705525 391015
rect 705581 390959 705649 391015
rect 705705 390959 705773 391015
rect 705829 390959 705897 391015
rect 705953 390959 706000 391015
rect 705512 390891 706000 390959
rect 705512 390835 705525 390891
rect 705581 390835 705649 390891
rect 705705 390835 705773 390891
rect 705829 390835 705897 390891
rect 705953 390835 706000 390891
rect 705512 390767 706000 390835
rect 705512 390711 705525 390767
rect 705581 390711 705649 390767
rect 705705 390711 705773 390767
rect 705829 390711 705897 390767
rect 705953 390711 706000 390767
rect 705512 390643 706000 390711
rect 705512 390587 705525 390643
rect 705581 390587 705649 390643
rect 705705 390587 705773 390643
rect 705829 390587 705897 390643
rect 705953 390587 706000 390643
rect 705512 390519 706000 390587
rect 705512 390463 705525 390519
rect 705581 390463 705649 390519
rect 705705 390463 705773 390519
rect 705829 390463 705897 390519
rect 705953 390463 706000 390519
rect 705512 390395 706000 390463
rect 705512 390339 705525 390395
rect 705581 390339 705649 390395
rect 705705 390339 705773 390395
rect 705829 390339 705897 390395
rect 705953 390339 706000 390395
rect 705512 390272 706000 390339
rect 70000 140661 70488 140728
rect 70000 140605 70047 140661
rect 70103 140605 70171 140661
rect 70227 140605 70295 140661
rect 70351 140605 70419 140661
rect 70475 140605 70488 140661
rect 70000 140537 70488 140605
rect 70000 140481 70047 140537
rect 70103 140481 70171 140537
rect 70227 140481 70295 140537
rect 70351 140481 70419 140537
rect 70475 140481 70488 140537
rect 70000 140413 70488 140481
rect 70000 140357 70047 140413
rect 70103 140357 70171 140413
rect 70227 140357 70295 140413
rect 70351 140357 70419 140413
rect 70475 140357 70488 140413
rect 70000 140289 70488 140357
rect 70000 140233 70047 140289
rect 70103 140233 70171 140289
rect 70227 140233 70295 140289
rect 70351 140233 70419 140289
rect 70475 140233 70488 140289
rect 70000 140165 70488 140233
rect 70000 140109 70047 140165
rect 70103 140109 70171 140165
rect 70227 140109 70295 140165
rect 70351 140109 70419 140165
rect 70475 140109 70488 140165
rect 70000 140041 70488 140109
rect 70000 139985 70047 140041
rect 70103 139985 70171 140041
rect 70227 139985 70295 140041
rect 70351 139985 70419 140041
rect 70475 139985 70488 140041
rect 70000 139917 70488 139985
rect 70000 139861 70047 139917
rect 70103 139861 70171 139917
rect 70227 139861 70295 139917
rect 70351 139861 70419 139917
rect 70475 139861 70488 139917
rect 70000 139793 70488 139861
rect 70000 139737 70047 139793
rect 70103 139737 70171 139793
rect 70227 139737 70295 139793
rect 70351 139737 70419 139793
rect 70475 139737 70488 139793
rect 70000 139669 70488 139737
rect 70000 139613 70047 139669
rect 70103 139613 70171 139669
rect 70227 139613 70295 139669
rect 70351 139613 70419 139669
rect 70475 139613 70488 139669
rect 70000 139545 70488 139613
rect 70000 139489 70047 139545
rect 70103 139489 70171 139545
rect 70227 139489 70295 139545
rect 70351 139489 70419 139545
rect 70475 139489 70488 139545
rect 70000 139421 70488 139489
rect 70000 139365 70047 139421
rect 70103 139365 70171 139421
rect 70227 139365 70295 139421
rect 70351 139365 70419 139421
rect 70475 139365 70488 139421
rect 70000 139297 70488 139365
rect 70000 139241 70047 139297
rect 70103 139241 70171 139297
rect 70227 139241 70295 139297
rect 70351 139241 70419 139297
rect 70475 139241 70488 139297
rect 70000 139173 70488 139241
rect 70000 139117 70047 139173
rect 70103 139117 70171 139173
rect 70227 139117 70295 139173
rect 70351 139117 70419 139173
rect 70475 139117 70488 139173
rect 70000 139049 70488 139117
rect 70000 138993 70047 139049
rect 70103 138993 70171 139049
rect 70227 138993 70295 139049
rect 70351 138993 70419 139049
rect 70475 138993 70488 139049
rect 70000 138925 70488 138993
rect 70000 138869 70047 138925
rect 70103 138869 70171 138925
rect 70227 138869 70295 138925
rect 70351 138869 70419 138925
rect 70475 138869 70488 138925
rect 70000 138828 70488 138869
rect 70000 138181 70488 138248
rect 70000 138125 70047 138181
rect 70103 138125 70171 138181
rect 70227 138125 70295 138181
rect 70351 138125 70419 138181
rect 70475 138125 70488 138181
rect 70000 138057 70488 138125
rect 70000 138001 70047 138057
rect 70103 138001 70171 138057
rect 70227 138001 70295 138057
rect 70351 138001 70419 138057
rect 70475 138001 70488 138057
rect 70000 137933 70488 138001
rect 70000 137877 70047 137933
rect 70103 137877 70171 137933
rect 70227 137877 70295 137933
rect 70351 137877 70419 137933
rect 70475 137877 70488 137933
rect 70000 137809 70488 137877
rect 70000 137753 70047 137809
rect 70103 137753 70171 137809
rect 70227 137753 70295 137809
rect 70351 137753 70419 137809
rect 70475 137753 70488 137809
rect 70000 137685 70488 137753
rect 70000 137629 70047 137685
rect 70103 137629 70171 137685
rect 70227 137629 70295 137685
rect 70351 137629 70419 137685
rect 70475 137629 70488 137685
rect 70000 137561 70488 137629
rect 70000 137505 70047 137561
rect 70103 137505 70171 137561
rect 70227 137505 70295 137561
rect 70351 137505 70419 137561
rect 70475 137505 70488 137561
rect 70000 137437 70488 137505
rect 70000 137381 70047 137437
rect 70103 137381 70171 137437
rect 70227 137381 70295 137437
rect 70351 137381 70419 137437
rect 70475 137381 70488 137437
rect 70000 137313 70488 137381
rect 70000 137257 70047 137313
rect 70103 137257 70171 137313
rect 70227 137257 70295 137313
rect 70351 137257 70419 137313
rect 70475 137257 70488 137313
rect 70000 137189 70488 137257
rect 70000 137133 70047 137189
rect 70103 137133 70171 137189
rect 70227 137133 70295 137189
rect 70351 137133 70419 137189
rect 70475 137133 70488 137189
rect 70000 137065 70488 137133
rect 70000 137009 70047 137065
rect 70103 137009 70171 137065
rect 70227 137009 70295 137065
rect 70351 137009 70419 137065
rect 70475 137009 70488 137065
rect 70000 136941 70488 137009
rect 70000 136885 70047 136941
rect 70103 136885 70171 136941
rect 70227 136885 70295 136941
rect 70351 136885 70419 136941
rect 70475 136885 70488 136941
rect 70000 136817 70488 136885
rect 70000 136761 70047 136817
rect 70103 136761 70171 136817
rect 70227 136761 70295 136817
rect 70351 136761 70419 136817
rect 70475 136761 70488 136817
rect 70000 136693 70488 136761
rect 70000 136637 70047 136693
rect 70103 136637 70171 136693
rect 70227 136637 70295 136693
rect 70351 136637 70419 136693
rect 70475 136637 70488 136693
rect 70000 136569 70488 136637
rect 70000 136513 70047 136569
rect 70103 136513 70171 136569
rect 70227 136513 70295 136569
rect 70351 136513 70419 136569
rect 70475 136513 70488 136569
rect 70000 136445 70488 136513
rect 70000 136389 70047 136445
rect 70103 136389 70171 136445
rect 70227 136389 70295 136445
rect 70351 136389 70419 136445
rect 70475 136389 70488 136445
rect 70000 136321 70488 136389
rect 70000 136265 70047 136321
rect 70103 136265 70171 136321
rect 70227 136265 70295 136321
rect 70351 136265 70419 136321
rect 70475 136265 70488 136321
rect 70000 136198 70488 136265
rect 70000 135811 70488 135878
rect 70000 135755 70047 135811
rect 70103 135755 70171 135811
rect 70227 135755 70295 135811
rect 70351 135755 70419 135811
rect 70475 135755 70488 135811
rect 70000 135687 70488 135755
rect 70000 135631 70047 135687
rect 70103 135631 70171 135687
rect 70227 135631 70295 135687
rect 70351 135631 70419 135687
rect 70475 135631 70488 135687
rect 70000 135563 70488 135631
rect 70000 135507 70047 135563
rect 70103 135507 70171 135563
rect 70227 135507 70295 135563
rect 70351 135507 70419 135563
rect 70475 135507 70488 135563
rect 70000 135439 70488 135507
rect 70000 135383 70047 135439
rect 70103 135383 70171 135439
rect 70227 135383 70295 135439
rect 70351 135383 70419 135439
rect 70475 135383 70488 135439
rect 70000 135315 70488 135383
rect 70000 135259 70047 135315
rect 70103 135259 70171 135315
rect 70227 135259 70295 135315
rect 70351 135259 70419 135315
rect 70475 135259 70488 135315
rect 70000 135191 70488 135259
rect 70000 135135 70047 135191
rect 70103 135135 70171 135191
rect 70227 135135 70295 135191
rect 70351 135135 70419 135191
rect 70475 135135 70488 135191
rect 70000 135067 70488 135135
rect 70000 135011 70047 135067
rect 70103 135011 70171 135067
rect 70227 135011 70295 135067
rect 70351 135011 70419 135067
rect 70475 135011 70488 135067
rect 70000 134943 70488 135011
rect 70000 134887 70047 134943
rect 70103 134887 70171 134943
rect 70227 134887 70295 134943
rect 70351 134887 70419 134943
rect 70475 134887 70488 134943
rect 70000 134819 70488 134887
rect 70000 134763 70047 134819
rect 70103 134763 70171 134819
rect 70227 134763 70295 134819
rect 70351 134763 70419 134819
rect 70475 134763 70488 134819
rect 70000 134695 70488 134763
rect 70000 134639 70047 134695
rect 70103 134639 70171 134695
rect 70227 134639 70295 134695
rect 70351 134639 70419 134695
rect 70475 134639 70488 134695
rect 70000 134571 70488 134639
rect 70000 134515 70047 134571
rect 70103 134515 70171 134571
rect 70227 134515 70295 134571
rect 70351 134515 70419 134571
rect 70475 134515 70488 134571
rect 70000 134447 70488 134515
rect 70000 134391 70047 134447
rect 70103 134391 70171 134447
rect 70227 134391 70295 134447
rect 70351 134391 70419 134447
rect 70475 134391 70488 134447
rect 70000 134323 70488 134391
rect 70000 134267 70047 134323
rect 70103 134267 70171 134323
rect 70227 134267 70295 134323
rect 70351 134267 70419 134323
rect 70475 134267 70488 134323
rect 70000 134199 70488 134267
rect 70000 134143 70047 134199
rect 70103 134143 70171 134199
rect 70227 134143 70295 134199
rect 70351 134143 70419 134199
rect 70475 134143 70488 134199
rect 70000 134075 70488 134143
rect 70000 134019 70047 134075
rect 70103 134019 70171 134075
rect 70227 134019 70295 134075
rect 70351 134019 70419 134075
rect 70475 134019 70488 134075
rect 70000 133951 70488 134019
rect 70000 133895 70047 133951
rect 70103 133895 70171 133951
rect 70227 133895 70295 133951
rect 70351 133895 70419 133951
rect 70475 133895 70488 133951
rect 70000 133828 70488 133895
rect 70000 133105 70488 133172
rect 70000 133049 70047 133105
rect 70103 133049 70171 133105
rect 70227 133049 70295 133105
rect 70351 133049 70419 133105
rect 70475 133049 70488 133105
rect 70000 132981 70488 133049
rect 70000 132925 70047 132981
rect 70103 132925 70171 132981
rect 70227 132925 70295 132981
rect 70351 132925 70419 132981
rect 70475 132925 70488 132981
rect 70000 132857 70488 132925
rect 70000 132801 70047 132857
rect 70103 132801 70171 132857
rect 70227 132801 70295 132857
rect 70351 132801 70419 132857
rect 70475 132801 70488 132857
rect 70000 132733 70488 132801
rect 70000 132677 70047 132733
rect 70103 132677 70171 132733
rect 70227 132677 70295 132733
rect 70351 132677 70419 132733
rect 70475 132677 70488 132733
rect 70000 132609 70488 132677
rect 70000 132553 70047 132609
rect 70103 132553 70171 132609
rect 70227 132553 70295 132609
rect 70351 132553 70419 132609
rect 70475 132553 70488 132609
rect 70000 132485 70488 132553
rect 70000 132429 70047 132485
rect 70103 132429 70171 132485
rect 70227 132429 70295 132485
rect 70351 132429 70419 132485
rect 70475 132429 70488 132485
rect 70000 132361 70488 132429
rect 70000 132305 70047 132361
rect 70103 132305 70171 132361
rect 70227 132305 70295 132361
rect 70351 132305 70419 132361
rect 70475 132305 70488 132361
rect 70000 132237 70488 132305
rect 70000 132181 70047 132237
rect 70103 132181 70171 132237
rect 70227 132181 70295 132237
rect 70351 132181 70419 132237
rect 70475 132181 70488 132237
rect 70000 132113 70488 132181
rect 70000 132057 70047 132113
rect 70103 132057 70171 132113
rect 70227 132057 70295 132113
rect 70351 132057 70419 132113
rect 70475 132057 70488 132113
rect 70000 131989 70488 132057
rect 70000 131933 70047 131989
rect 70103 131933 70171 131989
rect 70227 131933 70295 131989
rect 70351 131933 70419 131989
rect 70475 131933 70488 131989
rect 70000 131865 70488 131933
rect 70000 131809 70047 131865
rect 70103 131809 70171 131865
rect 70227 131809 70295 131865
rect 70351 131809 70419 131865
rect 70475 131809 70488 131865
rect 70000 131741 70488 131809
rect 70000 131685 70047 131741
rect 70103 131685 70171 131741
rect 70227 131685 70295 131741
rect 70351 131685 70419 131741
rect 70475 131685 70488 131741
rect 70000 131617 70488 131685
rect 70000 131561 70047 131617
rect 70103 131561 70171 131617
rect 70227 131561 70295 131617
rect 70351 131561 70419 131617
rect 70475 131561 70488 131617
rect 70000 131493 70488 131561
rect 70000 131437 70047 131493
rect 70103 131437 70171 131493
rect 70227 131437 70295 131493
rect 70351 131437 70419 131493
rect 70475 131437 70488 131493
rect 70000 131369 70488 131437
rect 70000 131313 70047 131369
rect 70103 131313 70171 131369
rect 70227 131313 70295 131369
rect 70351 131313 70419 131369
rect 70475 131313 70488 131369
rect 70000 131245 70488 131313
rect 70000 131189 70047 131245
rect 70103 131189 70171 131245
rect 70227 131189 70295 131245
rect 70351 131189 70419 131245
rect 70475 131189 70488 131245
rect 70000 131122 70488 131189
rect 70000 130735 70488 130802
rect 70000 130679 70047 130735
rect 70103 130679 70171 130735
rect 70227 130679 70295 130735
rect 70351 130679 70419 130735
rect 70475 130679 70488 130735
rect 70000 130611 70488 130679
rect 70000 130555 70047 130611
rect 70103 130555 70171 130611
rect 70227 130555 70295 130611
rect 70351 130555 70419 130611
rect 70475 130555 70488 130611
rect 70000 130487 70488 130555
rect 70000 130431 70047 130487
rect 70103 130431 70171 130487
rect 70227 130431 70295 130487
rect 70351 130431 70419 130487
rect 70475 130431 70488 130487
rect 70000 130363 70488 130431
rect 70000 130307 70047 130363
rect 70103 130307 70171 130363
rect 70227 130307 70295 130363
rect 70351 130307 70419 130363
rect 70475 130307 70488 130363
rect 70000 130239 70488 130307
rect 70000 130183 70047 130239
rect 70103 130183 70171 130239
rect 70227 130183 70295 130239
rect 70351 130183 70419 130239
rect 70475 130183 70488 130239
rect 70000 130115 70488 130183
rect 70000 130059 70047 130115
rect 70103 130059 70171 130115
rect 70227 130059 70295 130115
rect 70351 130059 70419 130115
rect 70475 130059 70488 130115
rect 70000 129991 70488 130059
rect 70000 129935 70047 129991
rect 70103 129935 70171 129991
rect 70227 129935 70295 129991
rect 70351 129935 70419 129991
rect 70475 129935 70488 129991
rect 70000 129867 70488 129935
rect 70000 129811 70047 129867
rect 70103 129811 70171 129867
rect 70227 129811 70295 129867
rect 70351 129811 70419 129867
rect 70475 129811 70488 129867
rect 70000 129743 70488 129811
rect 70000 129687 70047 129743
rect 70103 129687 70171 129743
rect 70227 129687 70295 129743
rect 70351 129687 70419 129743
rect 70475 129687 70488 129743
rect 70000 129619 70488 129687
rect 70000 129563 70047 129619
rect 70103 129563 70171 129619
rect 70227 129563 70295 129619
rect 70351 129563 70419 129619
rect 70475 129563 70488 129619
rect 70000 129495 70488 129563
rect 70000 129439 70047 129495
rect 70103 129439 70171 129495
rect 70227 129439 70295 129495
rect 70351 129439 70419 129495
rect 70475 129439 70488 129495
rect 70000 129371 70488 129439
rect 70000 129315 70047 129371
rect 70103 129315 70171 129371
rect 70227 129315 70295 129371
rect 70351 129315 70419 129371
rect 70475 129315 70488 129371
rect 70000 129247 70488 129315
rect 70000 129191 70047 129247
rect 70103 129191 70171 129247
rect 70227 129191 70295 129247
rect 70351 129191 70419 129247
rect 70475 129191 70488 129247
rect 70000 129123 70488 129191
rect 70000 129067 70047 129123
rect 70103 129067 70171 129123
rect 70227 129067 70295 129123
rect 70351 129067 70419 129123
rect 70475 129067 70488 129123
rect 70000 128999 70488 129067
rect 70000 128943 70047 128999
rect 70103 128943 70171 128999
rect 70227 128943 70295 128999
rect 70351 128943 70419 128999
rect 70475 128943 70488 128999
rect 70000 128875 70488 128943
rect 70000 128819 70047 128875
rect 70103 128819 70171 128875
rect 70227 128819 70295 128875
rect 70351 128819 70419 128875
rect 70475 128819 70488 128875
rect 70000 128752 70488 128819
rect 70000 128105 70488 128172
rect 70000 128049 70047 128105
rect 70103 128049 70171 128105
rect 70227 128049 70295 128105
rect 70351 128049 70419 128105
rect 70475 128049 70488 128105
rect 70000 127981 70488 128049
rect 70000 127925 70047 127981
rect 70103 127925 70171 127981
rect 70227 127925 70295 127981
rect 70351 127925 70419 127981
rect 70475 127925 70488 127981
rect 70000 127857 70488 127925
rect 70000 127801 70047 127857
rect 70103 127801 70171 127857
rect 70227 127801 70295 127857
rect 70351 127801 70419 127857
rect 70475 127801 70488 127857
rect 70000 127733 70488 127801
rect 70000 127677 70047 127733
rect 70103 127677 70171 127733
rect 70227 127677 70295 127733
rect 70351 127677 70419 127733
rect 70475 127677 70488 127733
rect 70000 127609 70488 127677
rect 70000 127553 70047 127609
rect 70103 127553 70171 127609
rect 70227 127553 70295 127609
rect 70351 127553 70419 127609
rect 70475 127553 70488 127609
rect 70000 127485 70488 127553
rect 70000 127429 70047 127485
rect 70103 127429 70171 127485
rect 70227 127429 70295 127485
rect 70351 127429 70419 127485
rect 70475 127429 70488 127485
rect 70000 127361 70488 127429
rect 70000 127305 70047 127361
rect 70103 127305 70171 127361
rect 70227 127305 70295 127361
rect 70351 127305 70419 127361
rect 70475 127305 70488 127361
rect 70000 127237 70488 127305
rect 70000 127181 70047 127237
rect 70103 127181 70171 127237
rect 70227 127181 70295 127237
rect 70351 127181 70419 127237
rect 70475 127181 70488 127237
rect 70000 127113 70488 127181
rect 70000 127057 70047 127113
rect 70103 127057 70171 127113
rect 70227 127057 70295 127113
rect 70351 127057 70419 127113
rect 70475 127057 70488 127113
rect 70000 126989 70488 127057
rect 70000 126933 70047 126989
rect 70103 126933 70171 126989
rect 70227 126933 70295 126989
rect 70351 126933 70419 126989
rect 70475 126933 70488 126989
rect 70000 126865 70488 126933
rect 70000 126809 70047 126865
rect 70103 126809 70171 126865
rect 70227 126809 70295 126865
rect 70351 126809 70419 126865
rect 70475 126809 70488 126865
rect 70000 126741 70488 126809
rect 70000 126685 70047 126741
rect 70103 126685 70171 126741
rect 70227 126685 70295 126741
rect 70351 126685 70419 126741
rect 70475 126685 70488 126741
rect 70000 126617 70488 126685
rect 70000 126561 70047 126617
rect 70103 126561 70171 126617
rect 70227 126561 70295 126617
rect 70351 126561 70419 126617
rect 70475 126561 70488 126617
rect 70000 126493 70488 126561
rect 70000 126437 70047 126493
rect 70103 126437 70171 126493
rect 70227 126437 70295 126493
rect 70351 126437 70419 126493
rect 70475 126437 70488 126493
rect 70000 126369 70488 126437
rect 70000 126313 70047 126369
rect 70103 126313 70171 126369
rect 70227 126313 70295 126369
rect 70351 126313 70419 126369
rect 70475 126313 70488 126369
rect 70000 126272 70488 126313
rect 70000 99661 70488 99728
rect 70000 99605 70047 99661
rect 70103 99605 70171 99661
rect 70227 99605 70295 99661
rect 70351 99605 70419 99661
rect 70475 99605 70488 99661
rect 70000 99537 70488 99605
rect 70000 99481 70047 99537
rect 70103 99481 70171 99537
rect 70227 99481 70295 99537
rect 70351 99481 70419 99537
rect 70475 99481 70488 99537
rect 70000 99413 70488 99481
rect 70000 99357 70047 99413
rect 70103 99357 70171 99413
rect 70227 99357 70295 99413
rect 70351 99357 70419 99413
rect 70475 99357 70488 99413
rect 70000 99289 70488 99357
rect 70000 99233 70047 99289
rect 70103 99233 70171 99289
rect 70227 99233 70295 99289
rect 70351 99233 70419 99289
rect 70475 99233 70488 99289
rect 70000 99165 70488 99233
rect 70000 99109 70047 99165
rect 70103 99109 70171 99165
rect 70227 99109 70295 99165
rect 70351 99109 70419 99165
rect 70475 99109 70488 99165
rect 70000 99041 70488 99109
rect 70000 98985 70047 99041
rect 70103 98985 70171 99041
rect 70227 98985 70295 99041
rect 70351 98985 70419 99041
rect 70475 98985 70488 99041
rect 70000 98917 70488 98985
rect 70000 98861 70047 98917
rect 70103 98861 70171 98917
rect 70227 98861 70295 98917
rect 70351 98861 70419 98917
rect 70475 98861 70488 98917
rect 70000 98793 70488 98861
rect 70000 98737 70047 98793
rect 70103 98737 70171 98793
rect 70227 98737 70295 98793
rect 70351 98737 70419 98793
rect 70475 98737 70488 98793
rect 70000 98669 70488 98737
rect 70000 98613 70047 98669
rect 70103 98613 70171 98669
rect 70227 98613 70295 98669
rect 70351 98613 70419 98669
rect 70475 98613 70488 98669
rect 70000 98545 70488 98613
rect 70000 98489 70047 98545
rect 70103 98489 70171 98545
rect 70227 98489 70295 98545
rect 70351 98489 70419 98545
rect 70475 98489 70488 98545
rect 70000 98421 70488 98489
rect 70000 98365 70047 98421
rect 70103 98365 70171 98421
rect 70227 98365 70295 98421
rect 70351 98365 70419 98421
rect 70475 98365 70488 98421
rect 70000 98297 70488 98365
rect 70000 98241 70047 98297
rect 70103 98241 70171 98297
rect 70227 98241 70295 98297
rect 70351 98241 70419 98297
rect 70475 98241 70488 98297
rect 70000 98173 70488 98241
rect 70000 98117 70047 98173
rect 70103 98117 70171 98173
rect 70227 98117 70295 98173
rect 70351 98117 70419 98173
rect 70475 98117 70488 98173
rect 70000 98049 70488 98117
rect 70000 97993 70047 98049
rect 70103 97993 70171 98049
rect 70227 97993 70295 98049
rect 70351 97993 70419 98049
rect 70475 97993 70488 98049
rect 70000 97925 70488 97993
rect 70000 97869 70047 97925
rect 70103 97869 70171 97925
rect 70227 97869 70295 97925
rect 70351 97869 70419 97925
rect 70475 97869 70488 97925
rect 70000 97828 70488 97869
rect 70000 97181 70488 97248
rect 70000 97125 70047 97181
rect 70103 97125 70171 97181
rect 70227 97125 70295 97181
rect 70351 97125 70419 97181
rect 70475 97125 70488 97181
rect 70000 97057 70488 97125
rect 70000 97001 70047 97057
rect 70103 97001 70171 97057
rect 70227 97001 70295 97057
rect 70351 97001 70419 97057
rect 70475 97001 70488 97057
rect 70000 96933 70488 97001
rect 70000 96877 70047 96933
rect 70103 96877 70171 96933
rect 70227 96877 70295 96933
rect 70351 96877 70419 96933
rect 70475 96877 70488 96933
rect 70000 96809 70488 96877
rect 70000 96753 70047 96809
rect 70103 96753 70171 96809
rect 70227 96753 70295 96809
rect 70351 96753 70419 96809
rect 70475 96753 70488 96809
rect 70000 96685 70488 96753
rect 70000 96629 70047 96685
rect 70103 96629 70171 96685
rect 70227 96629 70295 96685
rect 70351 96629 70419 96685
rect 70475 96629 70488 96685
rect 70000 96561 70488 96629
rect 70000 96505 70047 96561
rect 70103 96505 70171 96561
rect 70227 96505 70295 96561
rect 70351 96505 70419 96561
rect 70475 96505 70488 96561
rect 70000 96437 70488 96505
rect 70000 96381 70047 96437
rect 70103 96381 70171 96437
rect 70227 96381 70295 96437
rect 70351 96381 70419 96437
rect 70475 96381 70488 96437
rect 70000 96313 70488 96381
rect 70000 96257 70047 96313
rect 70103 96257 70171 96313
rect 70227 96257 70295 96313
rect 70351 96257 70419 96313
rect 70475 96257 70488 96313
rect 70000 96189 70488 96257
rect 70000 96133 70047 96189
rect 70103 96133 70171 96189
rect 70227 96133 70295 96189
rect 70351 96133 70419 96189
rect 70475 96133 70488 96189
rect 70000 96065 70488 96133
rect 70000 96009 70047 96065
rect 70103 96009 70171 96065
rect 70227 96009 70295 96065
rect 70351 96009 70419 96065
rect 70475 96009 70488 96065
rect 70000 95941 70488 96009
rect 70000 95885 70047 95941
rect 70103 95885 70171 95941
rect 70227 95885 70295 95941
rect 70351 95885 70419 95941
rect 70475 95885 70488 95941
rect 70000 95817 70488 95885
rect 70000 95761 70047 95817
rect 70103 95761 70171 95817
rect 70227 95761 70295 95817
rect 70351 95761 70419 95817
rect 70475 95761 70488 95817
rect 70000 95693 70488 95761
rect 70000 95637 70047 95693
rect 70103 95637 70171 95693
rect 70227 95637 70295 95693
rect 70351 95637 70419 95693
rect 70475 95637 70488 95693
rect 70000 95569 70488 95637
rect 70000 95513 70047 95569
rect 70103 95513 70171 95569
rect 70227 95513 70295 95569
rect 70351 95513 70419 95569
rect 70475 95513 70488 95569
rect 70000 95445 70488 95513
rect 70000 95389 70047 95445
rect 70103 95389 70171 95445
rect 70227 95389 70295 95445
rect 70351 95389 70419 95445
rect 70475 95389 70488 95445
rect 70000 95321 70488 95389
rect 70000 95265 70047 95321
rect 70103 95265 70171 95321
rect 70227 95265 70295 95321
rect 70351 95265 70419 95321
rect 70475 95265 70488 95321
rect 70000 95198 70488 95265
rect 70000 94811 70488 94878
rect 70000 94755 70047 94811
rect 70103 94755 70171 94811
rect 70227 94755 70295 94811
rect 70351 94755 70419 94811
rect 70475 94755 70488 94811
rect 70000 94687 70488 94755
rect 70000 94631 70047 94687
rect 70103 94631 70171 94687
rect 70227 94631 70295 94687
rect 70351 94631 70419 94687
rect 70475 94631 70488 94687
rect 70000 94563 70488 94631
rect 70000 94507 70047 94563
rect 70103 94507 70171 94563
rect 70227 94507 70295 94563
rect 70351 94507 70419 94563
rect 70475 94507 70488 94563
rect 70000 94439 70488 94507
rect 70000 94383 70047 94439
rect 70103 94383 70171 94439
rect 70227 94383 70295 94439
rect 70351 94383 70419 94439
rect 70475 94383 70488 94439
rect 70000 94315 70488 94383
rect 70000 94259 70047 94315
rect 70103 94259 70171 94315
rect 70227 94259 70295 94315
rect 70351 94259 70419 94315
rect 70475 94259 70488 94315
rect 70000 94191 70488 94259
rect 70000 94135 70047 94191
rect 70103 94135 70171 94191
rect 70227 94135 70295 94191
rect 70351 94135 70419 94191
rect 70475 94135 70488 94191
rect 70000 94067 70488 94135
rect 70000 94011 70047 94067
rect 70103 94011 70171 94067
rect 70227 94011 70295 94067
rect 70351 94011 70419 94067
rect 70475 94011 70488 94067
rect 70000 93943 70488 94011
rect 70000 93887 70047 93943
rect 70103 93887 70171 93943
rect 70227 93887 70295 93943
rect 70351 93887 70419 93943
rect 70475 93887 70488 93943
rect 70000 93819 70488 93887
rect 70000 93763 70047 93819
rect 70103 93763 70171 93819
rect 70227 93763 70295 93819
rect 70351 93763 70419 93819
rect 70475 93763 70488 93819
rect 70000 93695 70488 93763
rect 70000 93639 70047 93695
rect 70103 93639 70171 93695
rect 70227 93639 70295 93695
rect 70351 93639 70419 93695
rect 70475 93639 70488 93695
rect 70000 93571 70488 93639
rect 70000 93515 70047 93571
rect 70103 93515 70171 93571
rect 70227 93515 70295 93571
rect 70351 93515 70419 93571
rect 70475 93515 70488 93571
rect 70000 93447 70488 93515
rect 70000 93391 70047 93447
rect 70103 93391 70171 93447
rect 70227 93391 70295 93447
rect 70351 93391 70419 93447
rect 70475 93391 70488 93447
rect 70000 93323 70488 93391
rect 70000 93267 70047 93323
rect 70103 93267 70171 93323
rect 70227 93267 70295 93323
rect 70351 93267 70419 93323
rect 70475 93267 70488 93323
rect 70000 93199 70488 93267
rect 70000 93143 70047 93199
rect 70103 93143 70171 93199
rect 70227 93143 70295 93199
rect 70351 93143 70419 93199
rect 70475 93143 70488 93199
rect 70000 93075 70488 93143
rect 70000 93019 70047 93075
rect 70103 93019 70171 93075
rect 70227 93019 70295 93075
rect 70351 93019 70419 93075
rect 70475 93019 70488 93075
rect 70000 92951 70488 93019
rect 70000 92895 70047 92951
rect 70103 92895 70171 92951
rect 70227 92895 70295 92951
rect 70351 92895 70419 92951
rect 70475 92895 70488 92951
rect 70000 92828 70488 92895
rect 70000 92105 70488 92172
rect 70000 92049 70047 92105
rect 70103 92049 70171 92105
rect 70227 92049 70295 92105
rect 70351 92049 70419 92105
rect 70475 92049 70488 92105
rect 70000 91981 70488 92049
rect 70000 91925 70047 91981
rect 70103 91925 70171 91981
rect 70227 91925 70295 91981
rect 70351 91925 70419 91981
rect 70475 91925 70488 91981
rect 70000 91857 70488 91925
rect 70000 91801 70047 91857
rect 70103 91801 70171 91857
rect 70227 91801 70295 91857
rect 70351 91801 70419 91857
rect 70475 91801 70488 91857
rect 70000 91733 70488 91801
rect 70000 91677 70047 91733
rect 70103 91677 70171 91733
rect 70227 91677 70295 91733
rect 70351 91677 70419 91733
rect 70475 91677 70488 91733
rect 70000 91609 70488 91677
rect 70000 91553 70047 91609
rect 70103 91553 70171 91609
rect 70227 91553 70295 91609
rect 70351 91553 70419 91609
rect 70475 91553 70488 91609
rect 70000 91485 70488 91553
rect 70000 91429 70047 91485
rect 70103 91429 70171 91485
rect 70227 91429 70295 91485
rect 70351 91429 70419 91485
rect 70475 91429 70488 91485
rect 70000 91361 70488 91429
rect 70000 91305 70047 91361
rect 70103 91305 70171 91361
rect 70227 91305 70295 91361
rect 70351 91305 70419 91361
rect 70475 91305 70488 91361
rect 70000 91237 70488 91305
rect 70000 91181 70047 91237
rect 70103 91181 70171 91237
rect 70227 91181 70295 91237
rect 70351 91181 70419 91237
rect 70475 91181 70488 91237
rect 70000 91113 70488 91181
rect 70000 91057 70047 91113
rect 70103 91057 70171 91113
rect 70227 91057 70295 91113
rect 70351 91057 70419 91113
rect 70475 91057 70488 91113
rect 70000 90989 70488 91057
rect 70000 90933 70047 90989
rect 70103 90933 70171 90989
rect 70227 90933 70295 90989
rect 70351 90933 70419 90989
rect 70475 90933 70488 90989
rect 70000 90865 70488 90933
rect 70000 90809 70047 90865
rect 70103 90809 70171 90865
rect 70227 90809 70295 90865
rect 70351 90809 70419 90865
rect 70475 90809 70488 90865
rect 70000 90741 70488 90809
rect 70000 90685 70047 90741
rect 70103 90685 70171 90741
rect 70227 90685 70295 90741
rect 70351 90685 70419 90741
rect 70475 90685 70488 90741
rect 70000 90617 70488 90685
rect 70000 90561 70047 90617
rect 70103 90561 70171 90617
rect 70227 90561 70295 90617
rect 70351 90561 70419 90617
rect 70475 90561 70488 90617
rect 70000 90493 70488 90561
rect 70000 90437 70047 90493
rect 70103 90437 70171 90493
rect 70227 90437 70295 90493
rect 70351 90437 70419 90493
rect 70475 90437 70488 90493
rect 70000 90369 70488 90437
rect 70000 90313 70047 90369
rect 70103 90313 70171 90369
rect 70227 90313 70295 90369
rect 70351 90313 70419 90369
rect 70475 90313 70488 90369
rect 70000 90245 70488 90313
rect 70000 90189 70047 90245
rect 70103 90189 70171 90245
rect 70227 90189 70295 90245
rect 70351 90189 70419 90245
rect 70475 90189 70488 90245
rect 70000 90122 70488 90189
rect 70000 89735 70488 89802
rect 70000 89679 70047 89735
rect 70103 89679 70171 89735
rect 70227 89679 70295 89735
rect 70351 89679 70419 89735
rect 70475 89679 70488 89735
rect 70000 89611 70488 89679
rect 70000 89555 70047 89611
rect 70103 89555 70171 89611
rect 70227 89555 70295 89611
rect 70351 89555 70419 89611
rect 70475 89555 70488 89611
rect 70000 89487 70488 89555
rect 70000 89431 70047 89487
rect 70103 89431 70171 89487
rect 70227 89431 70295 89487
rect 70351 89431 70419 89487
rect 70475 89431 70488 89487
rect 70000 89363 70488 89431
rect 70000 89307 70047 89363
rect 70103 89307 70171 89363
rect 70227 89307 70295 89363
rect 70351 89307 70419 89363
rect 70475 89307 70488 89363
rect 70000 89239 70488 89307
rect 70000 89183 70047 89239
rect 70103 89183 70171 89239
rect 70227 89183 70295 89239
rect 70351 89183 70419 89239
rect 70475 89183 70488 89239
rect 70000 89115 70488 89183
rect 70000 89059 70047 89115
rect 70103 89059 70171 89115
rect 70227 89059 70295 89115
rect 70351 89059 70419 89115
rect 70475 89059 70488 89115
rect 70000 88991 70488 89059
rect 70000 88935 70047 88991
rect 70103 88935 70171 88991
rect 70227 88935 70295 88991
rect 70351 88935 70419 88991
rect 70475 88935 70488 88991
rect 70000 88867 70488 88935
rect 70000 88811 70047 88867
rect 70103 88811 70171 88867
rect 70227 88811 70295 88867
rect 70351 88811 70419 88867
rect 70475 88811 70488 88867
rect 70000 88743 70488 88811
rect 70000 88687 70047 88743
rect 70103 88687 70171 88743
rect 70227 88687 70295 88743
rect 70351 88687 70419 88743
rect 70475 88687 70488 88743
rect 70000 88619 70488 88687
rect 70000 88563 70047 88619
rect 70103 88563 70171 88619
rect 70227 88563 70295 88619
rect 70351 88563 70419 88619
rect 70475 88563 70488 88619
rect 70000 88495 70488 88563
rect 70000 88439 70047 88495
rect 70103 88439 70171 88495
rect 70227 88439 70295 88495
rect 70351 88439 70419 88495
rect 70475 88439 70488 88495
rect 70000 88371 70488 88439
rect 70000 88315 70047 88371
rect 70103 88315 70171 88371
rect 70227 88315 70295 88371
rect 70351 88315 70419 88371
rect 70475 88315 70488 88371
rect 70000 88247 70488 88315
rect 70000 88191 70047 88247
rect 70103 88191 70171 88247
rect 70227 88191 70295 88247
rect 70351 88191 70419 88247
rect 70475 88191 70488 88247
rect 70000 88123 70488 88191
rect 70000 88067 70047 88123
rect 70103 88067 70171 88123
rect 70227 88067 70295 88123
rect 70351 88067 70419 88123
rect 70475 88067 70488 88123
rect 70000 87999 70488 88067
rect 70000 87943 70047 87999
rect 70103 87943 70171 87999
rect 70227 87943 70295 87999
rect 70351 87943 70419 87999
rect 70475 87943 70488 87999
rect 70000 87875 70488 87943
rect 70000 87819 70047 87875
rect 70103 87819 70171 87875
rect 70227 87819 70295 87875
rect 70351 87819 70419 87875
rect 70475 87819 70488 87875
rect 70000 87752 70488 87819
rect 70000 87105 70488 87172
rect 70000 87049 70047 87105
rect 70103 87049 70171 87105
rect 70227 87049 70295 87105
rect 70351 87049 70419 87105
rect 70475 87049 70488 87105
rect 70000 86981 70488 87049
rect 70000 86925 70047 86981
rect 70103 86925 70171 86981
rect 70227 86925 70295 86981
rect 70351 86925 70419 86981
rect 70475 86925 70488 86981
rect 70000 86857 70488 86925
rect 70000 86801 70047 86857
rect 70103 86801 70171 86857
rect 70227 86801 70295 86857
rect 70351 86801 70419 86857
rect 70475 86801 70488 86857
rect 70000 86733 70488 86801
rect 70000 86677 70047 86733
rect 70103 86677 70171 86733
rect 70227 86677 70295 86733
rect 70351 86677 70419 86733
rect 70475 86677 70488 86733
rect 70000 86609 70488 86677
rect 70000 86553 70047 86609
rect 70103 86553 70171 86609
rect 70227 86553 70295 86609
rect 70351 86553 70419 86609
rect 70475 86553 70488 86609
rect 70000 86485 70488 86553
rect 70000 86429 70047 86485
rect 70103 86429 70171 86485
rect 70227 86429 70295 86485
rect 70351 86429 70419 86485
rect 70475 86429 70488 86485
rect 70000 86361 70488 86429
rect 70000 86305 70047 86361
rect 70103 86305 70171 86361
rect 70227 86305 70295 86361
rect 70351 86305 70419 86361
rect 70475 86305 70488 86361
rect 70000 86237 70488 86305
rect 70000 86181 70047 86237
rect 70103 86181 70171 86237
rect 70227 86181 70295 86237
rect 70351 86181 70419 86237
rect 70475 86181 70488 86237
rect 70000 86113 70488 86181
rect 70000 86057 70047 86113
rect 70103 86057 70171 86113
rect 70227 86057 70295 86113
rect 70351 86057 70419 86113
rect 70475 86057 70488 86113
rect 70000 85989 70488 86057
rect 70000 85933 70047 85989
rect 70103 85933 70171 85989
rect 70227 85933 70295 85989
rect 70351 85933 70419 85989
rect 70475 85933 70488 85989
rect 70000 85865 70488 85933
rect 70000 85809 70047 85865
rect 70103 85809 70171 85865
rect 70227 85809 70295 85865
rect 70351 85809 70419 85865
rect 70475 85809 70488 85865
rect 70000 85741 70488 85809
rect 70000 85685 70047 85741
rect 70103 85685 70171 85741
rect 70227 85685 70295 85741
rect 70351 85685 70419 85741
rect 70475 85685 70488 85741
rect 70000 85617 70488 85685
rect 70000 85561 70047 85617
rect 70103 85561 70171 85617
rect 70227 85561 70295 85617
rect 70351 85561 70419 85617
rect 70475 85561 70488 85617
rect 70000 85493 70488 85561
rect 70000 85437 70047 85493
rect 70103 85437 70171 85493
rect 70227 85437 70295 85493
rect 70351 85437 70419 85493
rect 70475 85437 70488 85493
rect 70000 85369 70488 85437
rect 70000 85313 70047 85369
rect 70103 85313 70171 85369
rect 70227 85313 70295 85369
rect 70351 85313 70419 85369
rect 70475 85313 70488 85369
rect 70000 85272 70488 85313
rect 655272 75945 657172 76088
rect 655272 75889 655326 75945
rect 655382 75889 655450 75945
rect 655506 75889 655574 75945
rect 655630 75889 655698 75945
rect 655754 75889 655822 75945
rect 655878 75889 655946 75945
rect 656002 75889 656070 75945
rect 656126 75889 656194 75945
rect 656250 75889 656318 75945
rect 656374 75889 657172 75945
rect 655272 75821 657172 75889
rect 655272 75765 655326 75821
rect 655382 75765 655450 75821
rect 655506 75765 655574 75821
rect 655630 75765 655698 75821
rect 655754 75765 655822 75821
rect 655878 75765 655946 75821
rect 656002 75765 656070 75821
rect 656126 75765 656194 75821
rect 656250 75765 656318 75821
rect 656374 75765 657172 75821
rect 655272 75697 657172 75765
rect 655272 75641 655326 75697
rect 655382 75641 655450 75697
rect 655506 75641 655574 75697
rect 655630 75641 655698 75697
rect 655754 75641 655822 75697
rect 655878 75641 655946 75697
rect 656002 75641 656070 75697
rect 656126 75641 656194 75697
rect 656250 75641 656318 75697
rect 656374 75641 657172 75697
rect 655272 75573 657172 75641
rect 655272 75517 655326 75573
rect 655382 75517 655450 75573
rect 655506 75517 655574 75573
rect 655630 75517 655698 75573
rect 655754 75517 655822 75573
rect 655878 75517 655946 75573
rect 656002 75517 656070 75573
rect 656126 75517 656194 75573
rect 656250 75517 656318 75573
rect 656374 75517 657172 75573
rect 655272 75449 657172 75517
rect 655272 75393 655326 75449
rect 655382 75393 655450 75449
rect 655506 75393 655574 75449
rect 655630 75393 655698 75449
rect 655754 75393 655822 75449
rect 655878 75393 655946 75449
rect 656002 75393 656070 75449
rect 656126 75393 656194 75449
rect 656250 75393 656318 75449
rect 656374 75393 657172 75449
rect 655272 75325 657172 75393
rect 655272 75269 655326 75325
rect 655382 75269 655450 75325
rect 655506 75269 655574 75325
rect 655630 75269 655698 75325
rect 655754 75269 655822 75325
rect 655878 75269 655946 75325
rect 656002 75269 656070 75325
rect 656126 75269 656194 75325
rect 656250 75269 656318 75325
rect 656374 75269 657172 75325
rect 655272 75201 657172 75269
rect 655272 75145 655326 75201
rect 655382 75145 655450 75201
rect 655506 75145 655574 75201
rect 655630 75145 655698 75201
rect 655754 75145 655822 75201
rect 655878 75145 655946 75201
rect 656002 75145 656070 75201
rect 656126 75145 656194 75201
rect 656250 75145 656318 75201
rect 656374 75145 657172 75201
rect 655272 75077 657172 75145
rect 655272 75021 655326 75077
rect 655382 75021 655450 75077
rect 655506 75021 655574 75077
rect 655630 75021 655698 75077
rect 655754 75021 655822 75077
rect 655878 75021 655946 75077
rect 656002 75021 656070 75077
rect 656126 75021 656194 75077
rect 656250 75021 656318 75077
rect 656374 75021 657172 75077
rect 655272 74953 657172 75021
rect 655272 74897 655326 74953
rect 655382 74897 655450 74953
rect 655506 74897 655574 74953
rect 655630 74897 655698 74953
rect 655754 74897 655822 74953
rect 655878 74897 655946 74953
rect 656002 74897 656070 74953
rect 656126 74897 656194 74953
rect 656250 74897 656318 74953
rect 656374 74897 657172 74953
rect 655272 74829 657172 74897
rect 655272 74773 655326 74829
rect 655382 74773 655450 74829
rect 655506 74773 655574 74829
rect 655630 74773 655698 74829
rect 655754 74773 655822 74829
rect 655878 74773 655946 74829
rect 656002 74773 656070 74829
rect 656126 74773 656194 74829
rect 656250 74773 656318 74829
rect 656374 74773 657172 74829
rect 655272 74705 657172 74773
rect 655272 74649 655326 74705
rect 655382 74649 655450 74705
rect 655506 74649 655574 74705
rect 655630 74649 655698 74705
rect 655754 74649 655822 74705
rect 655878 74649 655946 74705
rect 656002 74649 656070 74705
rect 656126 74649 656194 74705
rect 656250 74649 656318 74705
rect 656374 74649 657172 74705
rect 655272 74581 657172 74649
rect 655272 74525 655326 74581
rect 655382 74525 655450 74581
rect 655506 74525 655574 74581
rect 655630 74525 655698 74581
rect 655754 74525 655822 74581
rect 655878 74525 655946 74581
rect 656002 74525 656070 74581
rect 656126 74525 656194 74581
rect 656250 74525 656318 74581
rect 656374 74525 657172 74581
rect 105272 73945 107172 74088
rect 105272 73889 105326 73945
rect 105382 73889 105450 73945
rect 105506 73889 105574 73945
rect 105630 73889 105698 73945
rect 105754 73889 105822 73945
rect 105878 73889 105946 73945
rect 106002 73889 106070 73945
rect 106126 73889 106194 73945
rect 106250 73889 106318 73945
rect 106374 73889 106442 73945
rect 106498 73889 106566 73945
rect 106622 73889 106690 73945
rect 106746 73889 106814 73945
rect 106870 73889 106938 73945
rect 106994 73889 107062 73945
rect 107118 73889 107172 73945
rect 105272 73821 107172 73889
rect 105272 73765 105326 73821
rect 105382 73765 105450 73821
rect 105506 73765 105574 73821
rect 105630 73765 105698 73821
rect 105754 73765 105822 73821
rect 105878 73765 105946 73821
rect 106002 73765 106070 73821
rect 106126 73765 106194 73821
rect 106250 73765 106318 73821
rect 106374 73765 106442 73821
rect 106498 73765 106566 73821
rect 106622 73765 106690 73821
rect 106746 73765 106814 73821
rect 106870 73765 106938 73821
rect 106994 73765 107062 73821
rect 107118 73765 107172 73821
rect 105272 73697 107172 73765
rect 105272 73641 105326 73697
rect 105382 73641 105450 73697
rect 105506 73641 105574 73697
rect 105630 73641 105698 73697
rect 105754 73641 105822 73697
rect 105878 73641 105946 73697
rect 106002 73641 106070 73697
rect 106126 73641 106194 73697
rect 106250 73641 106318 73697
rect 106374 73641 106442 73697
rect 106498 73641 106566 73697
rect 106622 73641 106690 73697
rect 106746 73641 106814 73697
rect 106870 73641 106938 73697
rect 106994 73641 107062 73697
rect 107118 73641 107172 73697
rect 105272 73573 107172 73641
rect 105272 73517 105326 73573
rect 105382 73517 105450 73573
rect 105506 73517 105574 73573
rect 105630 73517 105698 73573
rect 105754 73517 105822 73573
rect 105878 73517 105946 73573
rect 106002 73517 106070 73573
rect 106126 73517 106194 73573
rect 106250 73517 106318 73573
rect 106374 73517 106442 73573
rect 106498 73517 106566 73573
rect 106622 73517 106690 73573
rect 106746 73517 106814 73573
rect 106870 73517 106938 73573
rect 106994 73517 107062 73573
rect 107118 73517 107172 73573
rect 105272 73449 107172 73517
rect 105272 73393 105326 73449
rect 105382 73393 105450 73449
rect 105506 73393 105574 73449
rect 105630 73393 105698 73449
rect 105754 73393 105822 73449
rect 105878 73393 105946 73449
rect 106002 73393 106070 73449
rect 106126 73393 106194 73449
rect 106250 73393 106318 73449
rect 106374 73393 106442 73449
rect 106498 73393 106566 73449
rect 106622 73393 106690 73449
rect 106746 73393 106814 73449
rect 106870 73393 106938 73449
rect 106994 73393 107062 73449
rect 107118 73393 107172 73449
rect 105272 73325 107172 73393
rect 105272 73269 105326 73325
rect 105382 73269 105450 73325
rect 105506 73269 105574 73325
rect 105630 73269 105698 73325
rect 105754 73269 105822 73325
rect 105878 73269 105946 73325
rect 106002 73269 106070 73325
rect 106126 73269 106194 73325
rect 106250 73269 106318 73325
rect 106374 73269 106442 73325
rect 106498 73269 106566 73325
rect 106622 73269 106690 73325
rect 106746 73269 106814 73325
rect 106870 73269 106938 73325
rect 106994 73269 107062 73325
rect 107118 73269 107172 73325
rect 105272 73201 107172 73269
rect 105272 73145 105326 73201
rect 105382 73145 105450 73201
rect 105506 73145 105574 73201
rect 105630 73145 105698 73201
rect 105754 73145 105822 73201
rect 105878 73145 105946 73201
rect 106002 73145 106070 73201
rect 106126 73145 106194 73201
rect 106250 73145 106318 73201
rect 106374 73145 106442 73201
rect 106498 73145 106566 73201
rect 106622 73145 106690 73201
rect 106746 73145 106814 73201
rect 106870 73145 106938 73201
rect 106994 73145 107062 73201
rect 107118 73145 107172 73201
rect 105272 73077 107172 73145
rect 105272 73021 105326 73077
rect 105382 73021 105450 73077
rect 105506 73021 105574 73077
rect 105630 73021 105698 73077
rect 105754 73021 105822 73077
rect 105878 73021 105946 73077
rect 106002 73021 106070 73077
rect 106126 73021 106194 73077
rect 106250 73021 106318 73077
rect 106374 73021 106442 73077
rect 106498 73021 106566 73077
rect 106622 73021 106690 73077
rect 106746 73021 106814 73077
rect 106870 73021 106938 73077
rect 106994 73021 107062 73077
rect 107118 73021 107172 73077
rect 105272 72953 107172 73021
rect 105272 72897 105326 72953
rect 105382 72897 105450 72953
rect 105506 72897 105574 72953
rect 105630 72897 105698 72953
rect 105754 72897 105822 72953
rect 105878 72897 105946 72953
rect 106002 72897 106070 72953
rect 106126 72897 106194 72953
rect 106250 72897 106318 72953
rect 106374 72897 106442 72953
rect 106498 72897 106566 72953
rect 106622 72897 106690 72953
rect 106746 72897 106814 72953
rect 106870 72897 106938 72953
rect 106994 72897 107062 72953
rect 107118 72897 107172 72953
rect 105272 72829 107172 72897
rect 105272 72773 105326 72829
rect 105382 72773 105450 72829
rect 105506 72773 105574 72829
rect 105630 72773 105698 72829
rect 105754 72773 105822 72829
rect 105878 72773 105946 72829
rect 106002 72773 106070 72829
rect 106126 72773 106194 72829
rect 106250 72773 106318 72829
rect 106374 72773 106442 72829
rect 106498 72773 106566 72829
rect 106622 72773 106690 72829
rect 106746 72773 106814 72829
rect 106870 72773 106938 72829
rect 106994 72773 107062 72829
rect 107118 72773 107172 72829
rect 105272 72705 107172 72773
rect 105272 72649 105326 72705
rect 105382 72649 105450 72705
rect 105506 72649 105574 72705
rect 105630 72649 105698 72705
rect 105754 72649 105822 72705
rect 105878 72649 105946 72705
rect 106002 72649 106070 72705
rect 106126 72649 106194 72705
rect 106250 72649 106318 72705
rect 106374 72649 106442 72705
rect 106498 72649 106566 72705
rect 106622 72649 106690 72705
rect 106746 72649 106814 72705
rect 106870 72649 106938 72705
rect 106994 72649 107062 72705
rect 107118 72649 107172 72705
rect 105272 72581 107172 72649
rect 105272 72525 105326 72581
rect 105382 72525 105450 72581
rect 105506 72525 105574 72581
rect 105630 72525 105698 72581
rect 105754 72525 105822 72581
rect 105878 72525 105946 72581
rect 106002 72525 106070 72581
rect 106126 72525 106194 72581
rect 106250 72525 106318 72581
rect 106374 72525 106442 72581
rect 106498 72525 106566 72581
rect 106622 72525 106690 72581
rect 106746 72525 106814 72581
rect 106870 72525 106938 72581
rect 106994 72525 107062 72581
rect 107118 72525 107172 72581
rect 105272 72457 107172 72525
rect 105272 72401 105326 72457
rect 105382 72401 105450 72457
rect 105506 72401 105574 72457
rect 105630 72401 105698 72457
rect 105754 72401 105822 72457
rect 105878 72401 105946 72457
rect 106002 72401 106070 72457
rect 106126 72401 106194 72457
rect 106250 72401 106318 72457
rect 106374 72401 106442 72457
rect 106498 72401 106566 72457
rect 106622 72401 106690 72457
rect 106746 72401 106814 72457
rect 106870 72401 106938 72457
rect 106994 72401 107062 72457
rect 107118 72401 107172 72457
rect 105272 72333 107172 72401
rect 105272 72277 105326 72333
rect 105382 72277 105450 72333
rect 105506 72277 105574 72333
rect 105630 72277 105698 72333
rect 105754 72277 105822 72333
rect 105878 72277 105946 72333
rect 106002 72277 106070 72333
rect 106126 72277 106194 72333
rect 106250 72277 106318 72333
rect 106374 72277 106442 72333
rect 106498 72277 106566 72333
rect 106622 72277 106690 72333
rect 106746 72277 106814 72333
rect 106870 72277 106938 72333
rect 106994 72277 107062 72333
rect 107118 72277 107172 72333
rect 105272 72209 107172 72277
rect 105272 72153 105326 72209
rect 105382 72153 105450 72209
rect 105506 72153 105574 72209
rect 105630 72153 105698 72209
rect 105754 72153 105822 72209
rect 105878 72153 105946 72209
rect 106002 72153 106070 72209
rect 106126 72153 106194 72209
rect 106250 72153 106318 72209
rect 106374 72153 106442 72209
rect 106498 72153 106566 72209
rect 106622 72153 106690 72209
rect 106746 72153 106814 72209
rect 106870 72153 106938 72209
rect 106994 72153 107062 72209
rect 107118 72153 107172 72209
rect 105272 70000 107172 72153
rect 107752 73945 109802 74088
rect 107752 73889 109046 73945
rect 109102 73889 109170 73945
rect 109226 73889 109294 73945
rect 109350 73889 109418 73945
rect 109474 73889 109542 73945
rect 109598 73889 109666 73945
rect 109722 73889 109802 73945
rect 107752 73821 109802 73889
rect 107752 73765 109046 73821
rect 109102 73765 109170 73821
rect 109226 73765 109294 73821
rect 109350 73765 109418 73821
rect 109474 73765 109542 73821
rect 109598 73765 109666 73821
rect 109722 73765 109802 73821
rect 107752 73697 109802 73765
rect 107752 73641 109046 73697
rect 109102 73641 109170 73697
rect 109226 73641 109294 73697
rect 109350 73641 109418 73697
rect 109474 73641 109542 73697
rect 109598 73641 109666 73697
rect 109722 73641 109802 73697
rect 107752 73573 109802 73641
rect 107752 73517 109046 73573
rect 109102 73517 109170 73573
rect 109226 73517 109294 73573
rect 109350 73517 109418 73573
rect 109474 73517 109542 73573
rect 109598 73517 109666 73573
rect 109722 73517 109802 73573
rect 107752 73449 109802 73517
rect 107752 73393 109046 73449
rect 109102 73393 109170 73449
rect 109226 73393 109294 73449
rect 109350 73393 109418 73449
rect 109474 73393 109542 73449
rect 109598 73393 109666 73449
rect 109722 73393 109802 73449
rect 107752 73325 109802 73393
rect 107752 73269 109046 73325
rect 109102 73269 109170 73325
rect 109226 73269 109294 73325
rect 109350 73269 109418 73325
rect 109474 73269 109542 73325
rect 109598 73269 109666 73325
rect 109722 73269 109802 73325
rect 107752 73201 109802 73269
rect 107752 73145 109046 73201
rect 109102 73145 109170 73201
rect 109226 73145 109294 73201
rect 109350 73145 109418 73201
rect 109474 73145 109542 73201
rect 109598 73145 109666 73201
rect 109722 73145 109802 73201
rect 107752 73077 109802 73145
rect 107752 73021 109046 73077
rect 109102 73021 109170 73077
rect 109226 73021 109294 73077
rect 109350 73021 109418 73077
rect 109474 73021 109542 73077
rect 109598 73021 109666 73077
rect 109722 73021 109802 73077
rect 107752 72953 109802 73021
rect 107752 72897 109046 72953
rect 109102 72897 109170 72953
rect 109226 72897 109294 72953
rect 109350 72897 109418 72953
rect 109474 72897 109542 72953
rect 109598 72897 109666 72953
rect 109722 72897 109802 72953
rect 107752 72829 109802 72897
rect 107752 72773 109046 72829
rect 109102 72773 109170 72829
rect 109226 72773 109294 72829
rect 109350 72773 109418 72829
rect 109474 72773 109542 72829
rect 109598 72773 109666 72829
rect 109722 72773 109802 72829
rect 107752 72705 109802 72773
rect 107752 72649 109046 72705
rect 109102 72649 109170 72705
rect 109226 72649 109294 72705
rect 109350 72649 109418 72705
rect 109474 72649 109542 72705
rect 109598 72649 109666 72705
rect 109722 72649 109802 72705
rect 107752 72581 109802 72649
rect 107752 72525 109046 72581
rect 109102 72525 109170 72581
rect 109226 72525 109294 72581
rect 109350 72525 109418 72581
rect 109474 72525 109542 72581
rect 109598 72525 109666 72581
rect 109722 72525 109802 72581
rect 107752 72457 109802 72525
rect 107752 72401 109046 72457
rect 109102 72401 109170 72457
rect 109226 72401 109294 72457
rect 109350 72401 109418 72457
rect 109474 72401 109542 72457
rect 109598 72401 109666 72457
rect 109722 72401 109802 72457
rect 107752 72333 109802 72401
rect 107752 72277 109046 72333
rect 109102 72277 109170 72333
rect 109226 72277 109294 72333
rect 109350 72277 109418 72333
rect 109474 72277 109542 72333
rect 109598 72277 109666 72333
rect 109722 72277 109802 72333
rect 107752 72209 109802 72277
rect 107752 72153 109046 72209
rect 109102 72153 109170 72209
rect 109226 72153 109294 72209
rect 109350 72153 109418 72209
rect 109474 72153 109542 72209
rect 109598 72153 109666 72209
rect 109722 72153 109802 72209
rect 107752 70000 109802 72153
rect 110122 73945 112172 74088
rect 110122 73889 110176 73945
rect 110232 73889 110300 73945
rect 110356 73889 110424 73945
rect 110480 73889 110548 73945
rect 110604 73889 110672 73945
rect 110728 73889 110796 73945
rect 110852 73889 110920 73945
rect 110976 73889 111044 73945
rect 111100 73889 111168 73945
rect 111224 73889 111292 73945
rect 111348 73889 111416 73945
rect 111472 73889 111540 73945
rect 111596 73889 111664 73945
rect 111720 73889 111788 73945
rect 111844 73889 111912 73945
rect 111968 73889 112036 73945
rect 112092 73889 112172 73945
rect 110122 73821 112172 73889
rect 110122 73765 110176 73821
rect 110232 73765 110300 73821
rect 110356 73765 110424 73821
rect 110480 73765 110548 73821
rect 110604 73765 110672 73821
rect 110728 73765 110796 73821
rect 110852 73765 110920 73821
rect 110976 73765 111044 73821
rect 111100 73765 111168 73821
rect 111224 73765 111292 73821
rect 111348 73765 111416 73821
rect 111472 73765 111540 73821
rect 111596 73765 111664 73821
rect 111720 73765 111788 73821
rect 111844 73765 111912 73821
rect 111968 73765 112036 73821
rect 112092 73765 112172 73821
rect 110122 73697 112172 73765
rect 110122 73641 110176 73697
rect 110232 73641 110300 73697
rect 110356 73641 110424 73697
rect 110480 73641 110548 73697
rect 110604 73641 110672 73697
rect 110728 73641 110796 73697
rect 110852 73641 110920 73697
rect 110976 73641 111044 73697
rect 111100 73641 111168 73697
rect 111224 73641 111292 73697
rect 111348 73641 111416 73697
rect 111472 73641 111540 73697
rect 111596 73641 111664 73697
rect 111720 73641 111788 73697
rect 111844 73641 111912 73697
rect 111968 73641 112036 73697
rect 112092 73641 112172 73697
rect 110122 73573 112172 73641
rect 110122 73517 110176 73573
rect 110232 73517 110300 73573
rect 110356 73517 110424 73573
rect 110480 73517 110548 73573
rect 110604 73517 110672 73573
rect 110728 73517 110796 73573
rect 110852 73517 110920 73573
rect 110976 73517 111044 73573
rect 111100 73517 111168 73573
rect 111224 73517 111292 73573
rect 111348 73517 111416 73573
rect 111472 73517 111540 73573
rect 111596 73517 111664 73573
rect 111720 73517 111788 73573
rect 111844 73517 111912 73573
rect 111968 73517 112036 73573
rect 112092 73517 112172 73573
rect 110122 73449 112172 73517
rect 110122 73393 110176 73449
rect 110232 73393 110300 73449
rect 110356 73393 110424 73449
rect 110480 73393 110548 73449
rect 110604 73393 110672 73449
rect 110728 73393 110796 73449
rect 110852 73393 110920 73449
rect 110976 73393 111044 73449
rect 111100 73393 111168 73449
rect 111224 73393 111292 73449
rect 111348 73393 111416 73449
rect 111472 73393 111540 73449
rect 111596 73393 111664 73449
rect 111720 73393 111788 73449
rect 111844 73393 111912 73449
rect 111968 73393 112036 73449
rect 112092 73393 112172 73449
rect 110122 73325 112172 73393
rect 110122 73269 110176 73325
rect 110232 73269 110300 73325
rect 110356 73269 110424 73325
rect 110480 73269 110548 73325
rect 110604 73269 110672 73325
rect 110728 73269 110796 73325
rect 110852 73269 110920 73325
rect 110976 73269 111044 73325
rect 111100 73269 111168 73325
rect 111224 73269 111292 73325
rect 111348 73269 111416 73325
rect 111472 73269 111540 73325
rect 111596 73269 111664 73325
rect 111720 73269 111788 73325
rect 111844 73269 111912 73325
rect 111968 73269 112036 73325
rect 112092 73269 112172 73325
rect 110122 73201 112172 73269
rect 110122 73145 110176 73201
rect 110232 73145 110300 73201
rect 110356 73145 110424 73201
rect 110480 73145 110548 73201
rect 110604 73145 110672 73201
rect 110728 73145 110796 73201
rect 110852 73145 110920 73201
rect 110976 73145 111044 73201
rect 111100 73145 111168 73201
rect 111224 73145 111292 73201
rect 111348 73145 111416 73201
rect 111472 73145 111540 73201
rect 111596 73145 111664 73201
rect 111720 73145 111788 73201
rect 111844 73145 111912 73201
rect 111968 73145 112036 73201
rect 112092 73145 112172 73201
rect 110122 73077 112172 73145
rect 110122 73021 110176 73077
rect 110232 73021 110300 73077
rect 110356 73021 110424 73077
rect 110480 73021 110548 73077
rect 110604 73021 110672 73077
rect 110728 73021 110796 73077
rect 110852 73021 110920 73077
rect 110976 73021 111044 73077
rect 111100 73021 111168 73077
rect 111224 73021 111292 73077
rect 111348 73021 111416 73077
rect 111472 73021 111540 73077
rect 111596 73021 111664 73077
rect 111720 73021 111788 73077
rect 111844 73021 111912 73077
rect 111968 73021 112036 73077
rect 112092 73021 112172 73077
rect 110122 72953 112172 73021
rect 110122 72897 110176 72953
rect 110232 72897 110300 72953
rect 110356 72897 110424 72953
rect 110480 72897 110548 72953
rect 110604 72897 110672 72953
rect 110728 72897 110796 72953
rect 110852 72897 110920 72953
rect 110976 72897 111044 72953
rect 111100 72897 111168 72953
rect 111224 72897 111292 72953
rect 111348 72897 111416 72953
rect 111472 72897 111540 72953
rect 111596 72897 111664 72953
rect 111720 72897 111788 72953
rect 111844 72897 111912 72953
rect 111968 72897 112036 72953
rect 112092 72897 112172 72953
rect 110122 72829 112172 72897
rect 110122 72773 110176 72829
rect 110232 72773 110300 72829
rect 110356 72773 110424 72829
rect 110480 72773 110548 72829
rect 110604 72773 110672 72829
rect 110728 72773 110796 72829
rect 110852 72773 110920 72829
rect 110976 72773 111044 72829
rect 111100 72773 111168 72829
rect 111224 72773 111292 72829
rect 111348 72773 111416 72829
rect 111472 72773 111540 72829
rect 111596 72773 111664 72829
rect 111720 72773 111788 72829
rect 111844 72773 111912 72829
rect 111968 72773 112036 72829
rect 112092 72773 112172 72829
rect 110122 72705 112172 72773
rect 110122 72649 110176 72705
rect 110232 72649 110300 72705
rect 110356 72649 110424 72705
rect 110480 72649 110548 72705
rect 110604 72649 110672 72705
rect 110728 72649 110796 72705
rect 110852 72649 110920 72705
rect 110976 72649 111044 72705
rect 111100 72649 111168 72705
rect 111224 72649 111292 72705
rect 111348 72649 111416 72705
rect 111472 72649 111540 72705
rect 111596 72649 111664 72705
rect 111720 72649 111788 72705
rect 111844 72649 111912 72705
rect 111968 72649 112036 72705
rect 112092 72649 112172 72705
rect 110122 72581 112172 72649
rect 110122 72525 110176 72581
rect 110232 72525 110300 72581
rect 110356 72525 110424 72581
rect 110480 72525 110548 72581
rect 110604 72525 110672 72581
rect 110728 72525 110796 72581
rect 110852 72525 110920 72581
rect 110976 72525 111044 72581
rect 111100 72525 111168 72581
rect 111224 72525 111292 72581
rect 111348 72525 111416 72581
rect 111472 72525 111540 72581
rect 111596 72525 111664 72581
rect 111720 72525 111788 72581
rect 111844 72525 111912 72581
rect 111968 72525 112036 72581
rect 112092 72525 112172 72581
rect 110122 72457 112172 72525
rect 110122 72401 110176 72457
rect 110232 72401 110300 72457
rect 110356 72401 110424 72457
rect 110480 72401 110548 72457
rect 110604 72401 110672 72457
rect 110728 72401 110796 72457
rect 110852 72401 110920 72457
rect 110976 72401 111044 72457
rect 111100 72401 111168 72457
rect 111224 72401 111292 72457
rect 111348 72401 111416 72457
rect 111472 72401 111540 72457
rect 111596 72401 111664 72457
rect 111720 72401 111788 72457
rect 111844 72401 111912 72457
rect 111968 72401 112036 72457
rect 112092 72401 112172 72457
rect 110122 72333 112172 72401
rect 110122 72277 110176 72333
rect 110232 72277 110300 72333
rect 110356 72277 110424 72333
rect 110480 72277 110548 72333
rect 110604 72277 110672 72333
rect 110728 72277 110796 72333
rect 110852 72277 110920 72333
rect 110976 72277 111044 72333
rect 111100 72277 111168 72333
rect 111224 72277 111292 72333
rect 111348 72277 111416 72333
rect 111472 72277 111540 72333
rect 111596 72277 111664 72333
rect 111720 72277 111788 72333
rect 111844 72277 111912 72333
rect 111968 72277 112036 72333
rect 112092 72277 112172 72333
rect 110122 72209 112172 72277
rect 110122 72153 110176 72209
rect 110232 72153 110300 72209
rect 110356 72153 110424 72209
rect 110480 72153 110548 72209
rect 110604 72153 110672 72209
rect 110728 72153 110796 72209
rect 110852 72153 110920 72209
rect 110976 72153 111044 72209
rect 111100 72153 111168 72209
rect 111224 72153 111292 72209
rect 111348 72153 111416 72209
rect 111472 72153 111540 72209
rect 111596 72153 111664 72209
rect 111720 72153 111788 72209
rect 111844 72153 111912 72209
rect 111968 72153 112036 72209
rect 112092 72153 112172 72209
rect 110122 70000 112172 72153
rect 112828 73945 114878 74088
rect 112828 73889 112882 73945
rect 112938 73889 113006 73945
rect 113062 73889 113130 73945
rect 113186 73889 113254 73945
rect 113310 73889 113378 73945
rect 113434 73889 113502 73945
rect 113558 73889 113626 73945
rect 113682 73889 113750 73945
rect 113806 73889 113874 73945
rect 113930 73889 113998 73945
rect 114054 73889 114122 73945
rect 114178 73889 114246 73945
rect 114302 73889 114370 73945
rect 114426 73889 114494 73945
rect 114550 73889 114618 73945
rect 114674 73889 114742 73945
rect 114798 73889 114878 73945
rect 112828 73821 114878 73889
rect 112828 73765 112882 73821
rect 112938 73765 113006 73821
rect 113062 73765 113130 73821
rect 113186 73765 113254 73821
rect 113310 73765 113378 73821
rect 113434 73765 113502 73821
rect 113558 73765 113626 73821
rect 113682 73765 113750 73821
rect 113806 73765 113874 73821
rect 113930 73765 113998 73821
rect 114054 73765 114122 73821
rect 114178 73765 114246 73821
rect 114302 73765 114370 73821
rect 114426 73765 114494 73821
rect 114550 73765 114618 73821
rect 114674 73765 114742 73821
rect 114798 73765 114878 73821
rect 112828 73697 114878 73765
rect 112828 73641 112882 73697
rect 112938 73641 113006 73697
rect 113062 73641 113130 73697
rect 113186 73641 113254 73697
rect 113310 73641 113378 73697
rect 113434 73641 113502 73697
rect 113558 73641 113626 73697
rect 113682 73641 113750 73697
rect 113806 73641 113874 73697
rect 113930 73641 113998 73697
rect 114054 73641 114122 73697
rect 114178 73641 114246 73697
rect 114302 73641 114370 73697
rect 114426 73641 114494 73697
rect 114550 73641 114618 73697
rect 114674 73641 114742 73697
rect 114798 73641 114878 73697
rect 112828 73573 114878 73641
rect 112828 73517 112882 73573
rect 112938 73517 113006 73573
rect 113062 73517 113130 73573
rect 113186 73517 113254 73573
rect 113310 73517 113378 73573
rect 113434 73517 113502 73573
rect 113558 73517 113626 73573
rect 113682 73517 113750 73573
rect 113806 73517 113874 73573
rect 113930 73517 113998 73573
rect 114054 73517 114122 73573
rect 114178 73517 114246 73573
rect 114302 73517 114370 73573
rect 114426 73517 114494 73573
rect 114550 73517 114618 73573
rect 114674 73517 114742 73573
rect 114798 73517 114878 73573
rect 112828 73449 114878 73517
rect 112828 73393 112882 73449
rect 112938 73393 113006 73449
rect 113062 73393 113130 73449
rect 113186 73393 113254 73449
rect 113310 73393 113378 73449
rect 113434 73393 113502 73449
rect 113558 73393 113626 73449
rect 113682 73393 113750 73449
rect 113806 73393 113874 73449
rect 113930 73393 113998 73449
rect 114054 73393 114122 73449
rect 114178 73393 114246 73449
rect 114302 73393 114370 73449
rect 114426 73393 114494 73449
rect 114550 73393 114618 73449
rect 114674 73393 114742 73449
rect 114798 73393 114878 73449
rect 112828 73325 114878 73393
rect 112828 73269 112882 73325
rect 112938 73269 113006 73325
rect 113062 73269 113130 73325
rect 113186 73269 113254 73325
rect 113310 73269 113378 73325
rect 113434 73269 113502 73325
rect 113558 73269 113626 73325
rect 113682 73269 113750 73325
rect 113806 73269 113874 73325
rect 113930 73269 113998 73325
rect 114054 73269 114122 73325
rect 114178 73269 114246 73325
rect 114302 73269 114370 73325
rect 114426 73269 114494 73325
rect 114550 73269 114618 73325
rect 114674 73269 114742 73325
rect 114798 73269 114878 73325
rect 112828 73201 114878 73269
rect 112828 73145 112882 73201
rect 112938 73145 113006 73201
rect 113062 73145 113130 73201
rect 113186 73145 113254 73201
rect 113310 73145 113378 73201
rect 113434 73145 113502 73201
rect 113558 73145 113626 73201
rect 113682 73145 113750 73201
rect 113806 73145 113874 73201
rect 113930 73145 113998 73201
rect 114054 73145 114122 73201
rect 114178 73145 114246 73201
rect 114302 73145 114370 73201
rect 114426 73145 114494 73201
rect 114550 73145 114618 73201
rect 114674 73145 114742 73201
rect 114798 73145 114878 73201
rect 112828 73077 114878 73145
rect 112828 73021 112882 73077
rect 112938 73021 113006 73077
rect 113062 73021 113130 73077
rect 113186 73021 113254 73077
rect 113310 73021 113378 73077
rect 113434 73021 113502 73077
rect 113558 73021 113626 73077
rect 113682 73021 113750 73077
rect 113806 73021 113874 73077
rect 113930 73021 113998 73077
rect 114054 73021 114122 73077
rect 114178 73021 114246 73077
rect 114302 73021 114370 73077
rect 114426 73021 114494 73077
rect 114550 73021 114618 73077
rect 114674 73021 114742 73077
rect 114798 73021 114878 73077
rect 112828 72953 114878 73021
rect 112828 72897 112882 72953
rect 112938 72897 113006 72953
rect 113062 72897 113130 72953
rect 113186 72897 113254 72953
rect 113310 72897 113378 72953
rect 113434 72897 113502 72953
rect 113558 72897 113626 72953
rect 113682 72897 113750 72953
rect 113806 72897 113874 72953
rect 113930 72897 113998 72953
rect 114054 72897 114122 72953
rect 114178 72897 114246 72953
rect 114302 72897 114370 72953
rect 114426 72897 114494 72953
rect 114550 72897 114618 72953
rect 114674 72897 114742 72953
rect 114798 72897 114878 72953
rect 112828 72829 114878 72897
rect 112828 72773 112882 72829
rect 112938 72773 113006 72829
rect 113062 72773 113130 72829
rect 113186 72773 113254 72829
rect 113310 72773 113378 72829
rect 113434 72773 113502 72829
rect 113558 72773 113626 72829
rect 113682 72773 113750 72829
rect 113806 72773 113874 72829
rect 113930 72773 113998 72829
rect 114054 72773 114122 72829
rect 114178 72773 114246 72829
rect 114302 72773 114370 72829
rect 114426 72773 114494 72829
rect 114550 72773 114618 72829
rect 114674 72773 114742 72829
rect 114798 72773 114878 72829
rect 112828 72705 114878 72773
rect 112828 72649 112882 72705
rect 112938 72649 113006 72705
rect 113062 72649 113130 72705
rect 113186 72649 113254 72705
rect 113310 72649 113378 72705
rect 113434 72649 113502 72705
rect 113558 72649 113626 72705
rect 113682 72649 113750 72705
rect 113806 72649 113874 72705
rect 113930 72649 113998 72705
rect 114054 72649 114122 72705
rect 114178 72649 114246 72705
rect 114302 72649 114370 72705
rect 114426 72649 114494 72705
rect 114550 72649 114618 72705
rect 114674 72649 114742 72705
rect 114798 72649 114878 72705
rect 112828 72581 114878 72649
rect 112828 72525 112882 72581
rect 112938 72525 113006 72581
rect 113062 72525 113130 72581
rect 113186 72525 113254 72581
rect 113310 72525 113378 72581
rect 113434 72525 113502 72581
rect 113558 72525 113626 72581
rect 113682 72525 113750 72581
rect 113806 72525 113874 72581
rect 113930 72525 113998 72581
rect 114054 72525 114122 72581
rect 114178 72525 114246 72581
rect 114302 72525 114370 72581
rect 114426 72525 114494 72581
rect 114550 72525 114618 72581
rect 114674 72525 114742 72581
rect 114798 72525 114878 72581
rect 112828 72457 114878 72525
rect 112828 72401 112882 72457
rect 112938 72401 113006 72457
rect 113062 72401 113130 72457
rect 113186 72401 113254 72457
rect 113310 72401 113378 72457
rect 113434 72401 113502 72457
rect 113558 72401 113626 72457
rect 113682 72401 113750 72457
rect 113806 72401 113874 72457
rect 113930 72401 113998 72457
rect 114054 72401 114122 72457
rect 114178 72401 114246 72457
rect 114302 72401 114370 72457
rect 114426 72401 114494 72457
rect 114550 72401 114618 72457
rect 114674 72401 114742 72457
rect 114798 72401 114878 72457
rect 112828 72333 114878 72401
rect 112828 72277 112882 72333
rect 112938 72277 113006 72333
rect 113062 72277 113130 72333
rect 113186 72277 113254 72333
rect 113310 72277 113378 72333
rect 113434 72277 113502 72333
rect 113558 72277 113626 72333
rect 113682 72277 113750 72333
rect 113806 72277 113874 72333
rect 113930 72277 113998 72333
rect 114054 72277 114122 72333
rect 114178 72277 114246 72333
rect 114302 72277 114370 72333
rect 114426 72277 114494 72333
rect 114550 72277 114618 72333
rect 114674 72277 114742 72333
rect 114798 72277 114878 72333
rect 112828 72209 114878 72277
rect 112828 72153 112882 72209
rect 112938 72153 113006 72209
rect 113062 72153 113130 72209
rect 113186 72153 113254 72209
rect 113310 72153 113378 72209
rect 113434 72153 113502 72209
rect 113558 72153 113626 72209
rect 113682 72153 113750 72209
rect 113806 72153 113874 72209
rect 113930 72153 113998 72209
rect 114054 72153 114122 72209
rect 114178 72153 114246 72209
rect 114302 72153 114370 72209
rect 114426 72153 114494 72209
rect 114550 72153 114618 72209
rect 114674 72153 114742 72209
rect 114798 72153 114878 72209
rect 112828 70000 114878 72153
rect 115198 73945 117248 74088
rect 115198 73889 115252 73945
rect 115308 73889 115376 73945
rect 115432 73889 115500 73945
rect 115556 73889 115624 73945
rect 115680 73889 115748 73945
rect 115804 73889 115872 73945
rect 115928 73889 115996 73945
rect 116052 73889 116120 73945
rect 116176 73889 116244 73945
rect 116300 73889 116368 73945
rect 116424 73889 116492 73945
rect 116548 73889 116616 73945
rect 116672 73889 116740 73945
rect 116796 73889 116864 73945
rect 116920 73889 116988 73945
rect 117044 73889 117112 73945
rect 117168 73889 117248 73945
rect 115198 73821 117248 73889
rect 115198 73765 115252 73821
rect 115308 73765 115376 73821
rect 115432 73765 115500 73821
rect 115556 73765 115624 73821
rect 115680 73765 115748 73821
rect 115804 73765 115872 73821
rect 115928 73765 115996 73821
rect 116052 73765 116120 73821
rect 116176 73765 116244 73821
rect 116300 73765 116368 73821
rect 116424 73765 116492 73821
rect 116548 73765 116616 73821
rect 116672 73765 116740 73821
rect 116796 73765 116864 73821
rect 116920 73765 116988 73821
rect 117044 73765 117112 73821
rect 117168 73765 117248 73821
rect 115198 73697 117248 73765
rect 115198 73641 115252 73697
rect 115308 73641 115376 73697
rect 115432 73641 115500 73697
rect 115556 73641 115624 73697
rect 115680 73641 115748 73697
rect 115804 73641 115872 73697
rect 115928 73641 115996 73697
rect 116052 73641 116120 73697
rect 116176 73641 116244 73697
rect 116300 73641 116368 73697
rect 116424 73641 116492 73697
rect 116548 73641 116616 73697
rect 116672 73641 116740 73697
rect 116796 73641 116864 73697
rect 116920 73641 116988 73697
rect 117044 73641 117112 73697
rect 117168 73641 117248 73697
rect 115198 73573 117248 73641
rect 115198 73517 115252 73573
rect 115308 73517 115376 73573
rect 115432 73517 115500 73573
rect 115556 73517 115624 73573
rect 115680 73517 115748 73573
rect 115804 73517 115872 73573
rect 115928 73517 115996 73573
rect 116052 73517 116120 73573
rect 116176 73517 116244 73573
rect 116300 73517 116368 73573
rect 116424 73517 116492 73573
rect 116548 73517 116616 73573
rect 116672 73517 116740 73573
rect 116796 73517 116864 73573
rect 116920 73517 116988 73573
rect 117044 73517 117112 73573
rect 117168 73517 117248 73573
rect 115198 73449 117248 73517
rect 115198 73393 115252 73449
rect 115308 73393 115376 73449
rect 115432 73393 115500 73449
rect 115556 73393 115624 73449
rect 115680 73393 115748 73449
rect 115804 73393 115872 73449
rect 115928 73393 115996 73449
rect 116052 73393 116120 73449
rect 116176 73393 116244 73449
rect 116300 73393 116368 73449
rect 116424 73393 116492 73449
rect 116548 73393 116616 73449
rect 116672 73393 116740 73449
rect 116796 73393 116864 73449
rect 116920 73393 116988 73449
rect 117044 73393 117112 73449
rect 117168 73393 117248 73449
rect 115198 73325 117248 73393
rect 115198 73269 115252 73325
rect 115308 73269 115376 73325
rect 115432 73269 115500 73325
rect 115556 73269 115624 73325
rect 115680 73269 115748 73325
rect 115804 73269 115872 73325
rect 115928 73269 115996 73325
rect 116052 73269 116120 73325
rect 116176 73269 116244 73325
rect 116300 73269 116368 73325
rect 116424 73269 116492 73325
rect 116548 73269 116616 73325
rect 116672 73269 116740 73325
rect 116796 73269 116864 73325
rect 116920 73269 116988 73325
rect 117044 73269 117112 73325
rect 117168 73269 117248 73325
rect 115198 73201 117248 73269
rect 115198 73145 115252 73201
rect 115308 73145 115376 73201
rect 115432 73145 115500 73201
rect 115556 73145 115624 73201
rect 115680 73145 115748 73201
rect 115804 73145 115872 73201
rect 115928 73145 115996 73201
rect 116052 73145 116120 73201
rect 116176 73145 116244 73201
rect 116300 73145 116368 73201
rect 116424 73145 116492 73201
rect 116548 73145 116616 73201
rect 116672 73145 116740 73201
rect 116796 73145 116864 73201
rect 116920 73145 116988 73201
rect 117044 73145 117112 73201
rect 117168 73145 117248 73201
rect 115198 73077 117248 73145
rect 115198 73021 115252 73077
rect 115308 73021 115376 73077
rect 115432 73021 115500 73077
rect 115556 73021 115624 73077
rect 115680 73021 115748 73077
rect 115804 73021 115872 73077
rect 115928 73021 115996 73077
rect 116052 73021 116120 73077
rect 116176 73021 116244 73077
rect 116300 73021 116368 73077
rect 116424 73021 116492 73077
rect 116548 73021 116616 73077
rect 116672 73021 116740 73077
rect 116796 73021 116864 73077
rect 116920 73021 116988 73077
rect 117044 73021 117112 73077
rect 117168 73021 117248 73077
rect 115198 72953 117248 73021
rect 115198 72897 115252 72953
rect 115308 72897 115376 72953
rect 115432 72897 115500 72953
rect 115556 72897 115624 72953
rect 115680 72897 115748 72953
rect 115804 72897 115872 72953
rect 115928 72897 115996 72953
rect 116052 72897 116120 72953
rect 116176 72897 116244 72953
rect 116300 72897 116368 72953
rect 116424 72897 116492 72953
rect 116548 72897 116616 72953
rect 116672 72897 116740 72953
rect 116796 72897 116864 72953
rect 116920 72897 116988 72953
rect 117044 72897 117112 72953
rect 117168 72897 117248 72953
rect 115198 72829 117248 72897
rect 115198 72773 115252 72829
rect 115308 72773 115376 72829
rect 115432 72773 115500 72829
rect 115556 72773 115624 72829
rect 115680 72773 115748 72829
rect 115804 72773 115872 72829
rect 115928 72773 115996 72829
rect 116052 72773 116120 72829
rect 116176 72773 116244 72829
rect 116300 72773 116368 72829
rect 116424 72773 116492 72829
rect 116548 72773 116616 72829
rect 116672 72773 116740 72829
rect 116796 72773 116864 72829
rect 116920 72773 116988 72829
rect 117044 72773 117112 72829
rect 117168 72773 117248 72829
rect 115198 72705 117248 72773
rect 115198 72649 115252 72705
rect 115308 72649 115376 72705
rect 115432 72649 115500 72705
rect 115556 72649 115624 72705
rect 115680 72649 115748 72705
rect 115804 72649 115872 72705
rect 115928 72649 115996 72705
rect 116052 72649 116120 72705
rect 116176 72649 116244 72705
rect 116300 72649 116368 72705
rect 116424 72649 116492 72705
rect 116548 72649 116616 72705
rect 116672 72649 116740 72705
rect 116796 72649 116864 72705
rect 116920 72649 116988 72705
rect 117044 72649 117112 72705
rect 117168 72649 117248 72705
rect 115198 72581 117248 72649
rect 115198 72525 115252 72581
rect 115308 72525 115376 72581
rect 115432 72525 115500 72581
rect 115556 72525 115624 72581
rect 115680 72525 115748 72581
rect 115804 72525 115872 72581
rect 115928 72525 115996 72581
rect 116052 72525 116120 72581
rect 116176 72525 116244 72581
rect 116300 72525 116368 72581
rect 116424 72525 116492 72581
rect 116548 72525 116616 72581
rect 116672 72525 116740 72581
rect 116796 72525 116864 72581
rect 116920 72525 116988 72581
rect 117044 72525 117112 72581
rect 117168 72525 117248 72581
rect 115198 72457 117248 72525
rect 115198 72401 115252 72457
rect 115308 72401 115376 72457
rect 115432 72401 115500 72457
rect 115556 72401 115624 72457
rect 115680 72401 115748 72457
rect 115804 72401 115872 72457
rect 115928 72401 115996 72457
rect 116052 72401 116120 72457
rect 116176 72401 116244 72457
rect 116300 72401 116368 72457
rect 116424 72401 116492 72457
rect 116548 72401 116616 72457
rect 116672 72401 116740 72457
rect 116796 72401 116864 72457
rect 116920 72401 116988 72457
rect 117044 72401 117112 72457
rect 117168 72401 117248 72457
rect 115198 72333 117248 72401
rect 115198 72277 115252 72333
rect 115308 72277 115376 72333
rect 115432 72277 115500 72333
rect 115556 72277 115624 72333
rect 115680 72277 115748 72333
rect 115804 72277 115872 72333
rect 115928 72277 115996 72333
rect 116052 72277 116120 72333
rect 116176 72277 116244 72333
rect 116300 72277 116368 72333
rect 116424 72277 116492 72333
rect 116548 72277 116616 72333
rect 116672 72277 116740 72333
rect 116796 72277 116864 72333
rect 116920 72277 116988 72333
rect 117044 72277 117112 72333
rect 117168 72277 117248 72333
rect 115198 72209 117248 72277
rect 115198 72153 115252 72209
rect 115308 72153 115376 72209
rect 115432 72153 115500 72209
rect 115556 72153 115624 72209
rect 115680 72153 115748 72209
rect 115804 72153 115872 72209
rect 115928 72153 115996 72209
rect 116052 72153 116120 72209
rect 116176 72153 116244 72209
rect 116300 72153 116368 72209
rect 116424 72153 116492 72209
rect 116548 72153 116616 72209
rect 116672 72153 116740 72209
rect 116796 72153 116864 72209
rect 116920 72153 116988 72209
rect 117044 72153 117112 72209
rect 117168 72153 117248 72209
rect 115198 70000 117248 72153
rect 117828 73945 119728 74088
rect 117828 73889 117882 73945
rect 117938 73889 118006 73945
rect 118062 73889 118130 73945
rect 118186 73889 118254 73945
rect 118310 73889 118378 73945
rect 118434 73889 118502 73945
rect 118558 73889 118626 73945
rect 118682 73889 118750 73945
rect 118806 73889 118874 73945
rect 118930 73889 118998 73945
rect 119054 73889 119122 73945
rect 119178 73889 119246 73945
rect 119302 73889 119370 73945
rect 119426 73889 119494 73945
rect 119550 73889 119618 73945
rect 119674 73889 119728 73945
rect 117828 73821 119728 73889
rect 117828 73765 117882 73821
rect 117938 73765 118006 73821
rect 118062 73765 118130 73821
rect 118186 73765 118254 73821
rect 118310 73765 118378 73821
rect 118434 73765 118502 73821
rect 118558 73765 118626 73821
rect 118682 73765 118750 73821
rect 118806 73765 118874 73821
rect 118930 73765 118998 73821
rect 119054 73765 119122 73821
rect 119178 73765 119246 73821
rect 119302 73765 119370 73821
rect 119426 73765 119494 73821
rect 119550 73765 119618 73821
rect 119674 73765 119728 73821
rect 117828 73697 119728 73765
rect 117828 73641 117882 73697
rect 117938 73641 118006 73697
rect 118062 73641 118130 73697
rect 118186 73641 118254 73697
rect 118310 73641 118378 73697
rect 118434 73641 118502 73697
rect 118558 73641 118626 73697
rect 118682 73641 118750 73697
rect 118806 73641 118874 73697
rect 118930 73641 118998 73697
rect 119054 73641 119122 73697
rect 119178 73641 119246 73697
rect 119302 73641 119370 73697
rect 119426 73641 119494 73697
rect 119550 73641 119618 73697
rect 119674 73641 119728 73697
rect 117828 73573 119728 73641
rect 117828 73517 117882 73573
rect 117938 73517 118006 73573
rect 118062 73517 118130 73573
rect 118186 73517 118254 73573
rect 118310 73517 118378 73573
rect 118434 73517 118502 73573
rect 118558 73517 118626 73573
rect 118682 73517 118750 73573
rect 118806 73517 118874 73573
rect 118930 73517 118998 73573
rect 119054 73517 119122 73573
rect 119178 73517 119246 73573
rect 119302 73517 119370 73573
rect 119426 73517 119494 73573
rect 119550 73517 119618 73573
rect 119674 73517 119728 73573
rect 117828 73449 119728 73517
rect 117828 73393 117882 73449
rect 117938 73393 118006 73449
rect 118062 73393 118130 73449
rect 118186 73393 118254 73449
rect 118310 73393 118378 73449
rect 118434 73393 118502 73449
rect 118558 73393 118626 73449
rect 118682 73393 118750 73449
rect 118806 73393 118874 73449
rect 118930 73393 118998 73449
rect 119054 73393 119122 73449
rect 119178 73393 119246 73449
rect 119302 73393 119370 73449
rect 119426 73393 119494 73449
rect 119550 73393 119618 73449
rect 119674 73393 119728 73449
rect 117828 73325 119728 73393
rect 117828 73269 117882 73325
rect 117938 73269 118006 73325
rect 118062 73269 118130 73325
rect 118186 73269 118254 73325
rect 118310 73269 118378 73325
rect 118434 73269 118502 73325
rect 118558 73269 118626 73325
rect 118682 73269 118750 73325
rect 118806 73269 118874 73325
rect 118930 73269 118998 73325
rect 119054 73269 119122 73325
rect 119178 73269 119246 73325
rect 119302 73269 119370 73325
rect 119426 73269 119494 73325
rect 119550 73269 119618 73325
rect 119674 73269 119728 73325
rect 117828 73201 119728 73269
rect 117828 73145 117882 73201
rect 117938 73145 118006 73201
rect 118062 73145 118130 73201
rect 118186 73145 118254 73201
rect 118310 73145 118378 73201
rect 118434 73145 118502 73201
rect 118558 73145 118626 73201
rect 118682 73145 118750 73201
rect 118806 73145 118874 73201
rect 118930 73145 118998 73201
rect 119054 73145 119122 73201
rect 119178 73145 119246 73201
rect 119302 73145 119370 73201
rect 119426 73145 119494 73201
rect 119550 73145 119618 73201
rect 119674 73145 119728 73201
rect 117828 73077 119728 73145
rect 117828 73021 117882 73077
rect 117938 73021 118006 73077
rect 118062 73021 118130 73077
rect 118186 73021 118254 73077
rect 118310 73021 118378 73077
rect 118434 73021 118502 73077
rect 118558 73021 118626 73077
rect 118682 73021 118750 73077
rect 118806 73021 118874 73077
rect 118930 73021 118998 73077
rect 119054 73021 119122 73077
rect 119178 73021 119246 73077
rect 119302 73021 119370 73077
rect 119426 73021 119494 73077
rect 119550 73021 119618 73077
rect 119674 73021 119728 73077
rect 117828 72953 119728 73021
rect 117828 72897 117882 72953
rect 117938 72897 118006 72953
rect 118062 72897 118130 72953
rect 118186 72897 118254 72953
rect 118310 72897 118378 72953
rect 118434 72897 118502 72953
rect 118558 72897 118626 72953
rect 118682 72897 118750 72953
rect 118806 72897 118874 72953
rect 118930 72897 118998 72953
rect 119054 72897 119122 72953
rect 119178 72897 119246 72953
rect 119302 72897 119370 72953
rect 119426 72897 119494 72953
rect 119550 72897 119618 72953
rect 119674 72897 119728 72953
rect 117828 72829 119728 72897
rect 117828 72773 117882 72829
rect 117938 72773 118006 72829
rect 118062 72773 118130 72829
rect 118186 72773 118254 72829
rect 118310 72773 118378 72829
rect 118434 72773 118502 72829
rect 118558 72773 118626 72829
rect 118682 72773 118750 72829
rect 118806 72773 118874 72829
rect 118930 72773 118998 72829
rect 119054 72773 119122 72829
rect 119178 72773 119246 72829
rect 119302 72773 119370 72829
rect 119426 72773 119494 72829
rect 119550 72773 119618 72829
rect 119674 72773 119728 72829
rect 117828 72705 119728 72773
rect 117828 72649 117882 72705
rect 117938 72649 118006 72705
rect 118062 72649 118130 72705
rect 118186 72649 118254 72705
rect 118310 72649 118378 72705
rect 118434 72649 118502 72705
rect 118558 72649 118626 72705
rect 118682 72649 118750 72705
rect 118806 72649 118874 72705
rect 118930 72649 118998 72705
rect 119054 72649 119122 72705
rect 119178 72649 119246 72705
rect 119302 72649 119370 72705
rect 119426 72649 119494 72705
rect 119550 72649 119618 72705
rect 119674 72649 119728 72705
rect 117828 72581 119728 72649
rect 117828 72525 117882 72581
rect 117938 72525 118006 72581
rect 118062 72525 118130 72581
rect 118186 72525 118254 72581
rect 118310 72525 118378 72581
rect 118434 72525 118502 72581
rect 118558 72525 118626 72581
rect 118682 72525 118750 72581
rect 118806 72525 118874 72581
rect 118930 72525 118998 72581
rect 119054 72525 119122 72581
rect 119178 72525 119246 72581
rect 119302 72525 119370 72581
rect 119426 72525 119494 72581
rect 119550 72525 119618 72581
rect 119674 72525 119728 72581
rect 117828 72457 119728 72525
rect 117828 72401 117882 72457
rect 117938 72401 118006 72457
rect 118062 72401 118130 72457
rect 118186 72401 118254 72457
rect 118310 72401 118378 72457
rect 118434 72401 118502 72457
rect 118558 72401 118626 72457
rect 118682 72401 118750 72457
rect 118806 72401 118874 72457
rect 118930 72401 118998 72457
rect 119054 72401 119122 72457
rect 119178 72401 119246 72457
rect 119302 72401 119370 72457
rect 119426 72401 119494 72457
rect 119550 72401 119618 72457
rect 119674 72401 119728 72457
rect 117828 72333 119728 72401
rect 117828 72277 117882 72333
rect 117938 72277 118006 72333
rect 118062 72277 118130 72333
rect 118186 72277 118254 72333
rect 118310 72277 118378 72333
rect 118434 72277 118502 72333
rect 118558 72277 118626 72333
rect 118682 72277 118750 72333
rect 118806 72277 118874 72333
rect 118930 72277 118998 72333
rect 119054 72277 119122 72333
rect 119178 72277 119246 72333
rect 119302 72277 119370 72333
rect 119426 72277 119494 72333
rect 119550 72277 119618 72333
rect 119674 72277 119728 72333
rect 117828 72209 119728 72277
rect 117828 72153 117882 72209
rect 117938 72153 118006 72209
rect 118062 72153 118130 72209
rect 118186 72153 118254 72209
rect 118310 72153 118378 72209
rect 118434 72153 118502 72209
rect 118558 72153 118626 72209
rect 118682 72153 118750 72209
rect 118806 72153 118874 72209
rect 118930 72153 118998 72209
rect 119054 72153 119122 72209
rect 119178 72153 119246 72209
rect 119302 72153 119370 72209
rect 119426 72153 119494 72209
rect 119550 72153 119618 72209
rect 119674 72153 119728 72209
rect 117828 70000 119728 72153
rect 270272 73945 272172 74088
rect 270272 73889 270326 73945
rect 270382 73889 270450 73945
rect 270506 73889 270574 73945
rect 270630 73889 270698 73945
rect 270754 73889 270822 73945
rect 270878 73889 270946 73945
rect 271002 73889 271070 73945
rect 271126 73889 271194 73945
rect 271250 73889 271318 73945
rect 271374 73889 271442 73945
rect 271498 73889 271566 73945
rect 271622 73889 271690 73945
rect 271746 73889 271814 73945
rect 271870 73889 271938 73945
rect 271994 73889 272062 73945
rect 272118 73889 272172 73945
rect 270272 73821 272172 73889
rect 270272 73765 270326 73821
rect 270382 73765 270450 73821
rect 270506 73765 270574 73821
rect 270630 73765 270698 73821
rect 270754 73765 270822 73821
rect 270878 73765 270946 73821
rect 271002 73765 271070 73821
rect 271126 73765 271194 73821
rect 271250 73765 271318 73821
rect 271374 73765 271442 73821
rect 271498 73765 271566 73821
rect 271622 73765 271690 73821
rect 271746 73765 271814 73821
rect 271870 73765 271938 73821
rect 271994 73765 272062 73821
rect 272118 73765 272172 73821
rect 270272 73697 272172 73765
rect 270272 73641 270326 73697
rect 270382 73641 270450 73697
rect 270506 73641 270574 73697
rect 270630 73641 270698 73697
rect 270754 73641 270822 73697
rect 270878 73641 270946 73697
rect 271002 73641 271070 73697
rect 271126 73641 271194 73697
rect 271250 73641 271318 73697
rect 271374 73641 271442 73697
rect 271498 73641 271566 73697
rect 271622 73641 271690 73697
rect 271746 73641 271814 73697
rect 271870 73641 271938 73697
rect 271994 73641 272062 73697
rect 272118 73641 272172 73697
rect 270272 73573 272172 73641
rect 270272 73517 270326 73573
rect 270382 73517 270450 73573
rect 270506 73517 270574 73573
rect 270630 73517 270698 73573
rect 270754 73517 270822 73573
rect 270878 73517 270946 73573
rect 271002 73517 271070 73573
rect 271126 73517 271194 73573
rect 271250 73517 271318 73573
rect 271374 73517 271442 73573
rect 271498 73517 271566 73573
rect 271622 73517 271690 73573
rect 271746 73517 271814 73573
rect 271870 73517 271938 73573
rect 271994 73517 272062 73573
rect 272118 73517 272172 73573
rect 270272 73449 272172 73517
rect 270272 73393 270326 73449
rect 270382 73393 270450 73449
rect 270506 73393 270574 73449
rect 270630 73393 270698 73449
rect 270754 73393 270822 73449
rect 270878 73393 270946 73449
rect 271002 73393 271070 73449
rect 271126 73393 271194 73449
rect 271250 73393 271318 73449
rect 271374 73393 271442 73449
rect 271498 73393 271566 73449
rect 271622 73393 271690 73449
rect 271746 73393 271814 73449
rect 271870 73393 271938 73449
rect 271994 73393 272062 73449
rect 272118 73393 272172 73449
rect 270272 73325 272172 73393
rect 270272 73269 270326 73325
rect 270382 73269 270450 73325
rect 270506 73269 270574 73325
rect 270630 73269 270698 73325
rect 270754 73269 270822 73325
rect 270878 73269 270946 73325
rect 271002 73269 271070 73325
rect 271126 73269 271194 73325
rect 271250 73269 271318 73325
rect 271374 73269 271442 73325
rect 271498 73269 271566 73325
rect 271622 73269 271690 73325
rect 271746 73269 271814 73325
rect 271870 73269 271938 73325
rect 271994 73269 272062 73325
rect 272118 73269 272172 73325
rect 270272 73201 272172 73269
rect 270272 73145 270326 73201
rect 270382 73145 270450 73201
rect 270506 73145 270574 73201
rect 270630 73145 270698 73201
rect 270754 73145 270822 73201
rect 270878 73145 270946 73201
rect 271002 73145 271070 73201
rect 271126 73145 271194 73201
rect 271250 73145 271318 73201
rect 271374 73145 271442 73201
rect 271498 73145 271566 73201
rect 271622 73145 271690 73201
rect 271746 73145 271814 73201
rect 271870 73145 271938 73201
rect 271994 73145 272062 73201
rect 272118 73145 272172 73201
rect 270272 73077 272172 73145
rect 270272 73021 270326 73077
rect 270382 73021 270450 73077
rect 270506 73021 270574 73077
rect 270630 73021 270698 73077
rect 270754 73021 270822 73077
rect 270878 73021 270946 73077
rect 271002 73021 271070 73077
rect 271126 73021 271194 73077
rect 271250 73021 271318 73077
rect 271374 73021 271442 73077
rect 271498 73021 271566 73077
rect 271622 73021 271690 73077
rect 271746 73021 271814 73077
rect 271870 73021 271938 73077
rect 271994 73021 272062 73077
rect 272118 73021 272172 73077
rect 270272 72953 272172 73021
rect 270272 72897 270326 72953
rect 270382 72897 270450 72953
rect 270506 72897 270574 72953
rect 270630 72897 270698 72953
rect 270754 72897 270822 72953
rect 270878 72897 270946 72953
rect 271002 72897 271070 72953
rect 271126 72897 271194 72953
rect 271250 72897 271318 72953
rect 271374 72897 271442 72953
rect 271498 72897 271566 72953
rect 271622 72897 271690 72953
rect 271746 72897 271814 72953
rect 271870 72897 271938 72953
rect 271994 72897 272062 72953
rect 272118 72897 272172 72953
rect 270272 72829 272172 72897
rect 270272 72773 270326 72829
rect 270382 72773 270450 72829
rect 270506 72773 270574 72829
rect 270630 72773 270698 72829
rect 270754 72773 270822 72829
rect 270878 72773 270946 72829
rect 271002 72773 271070 72829
rect 271126 72773 271194 72829
rect 271250 72773 271318 72829
rect 271374 72773 271442 72829
rect 271498 72773 271566 72829
rect 271622 72773 271690 72829
rect 271746 72773 271814 72829
rect 271870 72773 271938 72829
rect 271994 72773 272062 72829
rect 272118 72773 272172 72829
rect 270272 72705 272172 72773
rect 270272 72649 270326 72705
rect 270382 72649 270450 72705
rect 270506 72649 270574 72705
rect 270630 72649 270698 72705
rect 270754 72649 270822 72705
rect 270878 72649 270946 72705
rect 271002 72649 271070 72705
rect 271126 72649 271194 72705
rect 271250 72649 271318 72705
rect 271374 72649 271442 72705
rect 271498 72649 271566 72705
rect 271622 72649 271690 72705
rect 271746 72649 271814 72705
rect 271870 72649 271938 72705
rect 271994 72649 272062 72705
rect 272118 72649 272172 72705
rect 270272 72581 272172 72649
rect 270272 72525 270326 72581
rect 270382 72525 270450 72581
rect 270506 72525 270574 72581
rect 270630 72525 270698 72581
rect 270754 72525 270822 72581
rect 270878 72525 270946 72581
rect 271002 72525 271070 72581
rect 271126 72525 271194 72581
rect 271250 72525 271318 72581
rect 271374 72525 271442 72581
rect 271498 72525 271566 72581
rect 271622 72525 271690 72581
rect 271746 72525 271814 72581
rect 271870 72525 271938 72581
rect 271994 72525 272062 72581
rect 272118 72525 272172 72581
rect 270272 72457 272172 72525
rect 270272 72401 270326 72457
rect 270382 72401 270450 72457
rect 270506 72401 270574 72457
rect 270630 72401 270698 72457
rect 270754 72401 270822 72457
rect 270878 72401 270946 72457
rect 271002 72401 271070 72457
rect 271126 72401 271194 72457
rect 271250 72401 271318 72457
rect 271374 72401 271442 72457
rect 271498 72401 271566 72457
rect 271622 72401 271690 72457
rect 271746 72401 271814 72457
rect 271870 72401 271938 72457
rect 271994 72401 272062 72457
rect 272118 72401 272172 72457
rect 270272 72333 272172 72401
rect 270272 72277 270326 72333
rect 270382 72277 270450 72333
rect 270506 72277 270574 72333
rect 270630 72277 270698 72333
rect 270754 72277 270822 72333
rect 270878 72277 270946 72333
rect 271002 72277 271070 72333
rect 271126 72277 271194 72333
rect 271250 72277 271318 72333
rect 271374 72277 271442 72333
rect 271498 72277 271566 72333
rect 271622 72277 271690 72333
rect 271746 72277 271814 72333
rect 271870 72277 271938 72333
rect 271994 72277 272062 72333
rect 272118 72277 272172 72333
rect 270272 72209 272172 72277
rect 270272 72153 270326 72209
rect 270382 72153 270450 72209
rect 270506 72153 270574 72209
rect 270630 72153 270698 72209
rect 270754 72153 270822 72209
rect 270878 72153 270946 72209
rect 271002 72153 271070 72209
rect 271126 72153 271194 72209
rect 271250 72153 271318 72209
rect 271374 72153 271442 72209
rect 271498 72153 271566 72209
rect 271622 72153 271690 72209
rect 271746 72153 271814 72209
rect 271870 72153 271938 72209
rect 271994 72153 272062 72209
rect 272118 72153 272172 72209
rect 270272 70000 272172 72153
rect 272752 73945 274802 74088
rect 272752 73889 272806 73945
rect 272862 73889 272930 73945
rect 272986 73889 273054 73945
rect 273110 73889 273178 73945
rect 273234 73889 273302 73945
rect 273358 73889 273426 73945
rect 273482 73889 273550 73945
rect 273606 73889 273674 73945
rect 273730 73889 273798 73945
rect 273854 73889 273922 73945
rect 273978 73889 274046 73945
rect 274102 73889 274170 73945
rect 274226 73889 274294 73945
rect 274350 73889 274418 73945
rect 274474 73889 274542 73945
rect 274598 73889 274666 73945
rect 274722 73889 274802 73945
rect 272752 73821 274802 73889
rect 272752 73765 272806 73821
rect 272862 73765 272930 73821
rect 272986 73765 273054 73821
rect 273110 73765 273178 73821
rect 273234 73765 273302 73821
rect 273358 73765 273426 73821
rect 273482 73765 273550 73821
rect 273606 73765 273674 73821
rect 273730 73765 273798 73821
rect 273854 73765 273922 73821
rect 273978 73765 274046 73821
rect 274102 73765 274170 73821
rect 274226 73765 274294 73821
rect 274350 73765 274418 73821
rect 274474 73765 274542 73821
rect 274598 73765 274666 73821
rect 274722 73765 274802 73821
rect 272752 73697 274802 73765
rect 272752 73641 272806 73697
rect 272862 73641 272930 73697
rect 272986 73641 273054 73697
rect 273110 73641 273178 73697
rect 273234 73641 273302 73697
rect 273358 73641 273426 73697
rect 273482 73641 273550 73697
rect 273606 73641 273674 73697
rect 273730 73641 273798 73697
rect 273854 73641 273922 73697
rect 273978 73641 274046 73697
rect 274102 73641 274170 73697
rect 274226 73641 274294 73697
rect 274350 73641 274418 73697
rect 274474 73641 274542 73697
rect 274598 73641 274666 73697
rect 274722 73641 274802 73697
rect 272752 73573 274802 73641
rect 272752 73517 272806 73573
rect 272862 73517 272930 73573
rect 272986 73517 273054 73573
rect 273110 73517 273178 73573
rect 273234 73517 273302 73573
rect 273358 73517 273426 73573
rect 273482 73517 273550 73573
rect 273606 73517 273674 73573
rect 273730 73517 273798 73573
rect 273854 73517 273922 73573
rect 273978 73517 274046 73573
rect 274102 73517 274170 73573
rect 274226 73517 274294 73573
rect 274350 73517 274418 73573
rect 274474 73517 274542 73573
rect 274598 73517 274666 73573
rect 274722 73517 274802 73573
rect 272752 73449 274802 73517
rect 272752 73393 272806 73449
rect 272862 73393 272930 73449
rect 272986 73393 273054 73449
rect 273110 73393 273178 73449
rect 273234 73393 273302 73449
rect 273358 73393 273426 73449
rect 273482 73393 273550 73449
rect 273606 73393 273674 73449
rect 273730 73393 273798 73449
rect 273854 73393 273922 73449
rect 273978 73393 274046 73449
rect 274102 73393 274170 73449
rect 274226 73393 274294 73449
rect 274350 73393 274418 73449
rect 274474 73393 274542 73449
rect 274598 73393 274666 73449
rect 274722 73393 274802 73449
rect 272752 73325 274802 73393
rect 272752 73269 272806 73325
rect 272862 73269 272930 73325
rect 272986 73269 273054 73325
rect 273110 73269 273178 73325
rect 273234 73269 273302 73325
rect 273358 73269 273426 73325
rect 273482 73269 273550 73325
rect 273606 73269 273674 73325
rect 273730 73269 273798 73325
rect 273854 73269 273922 73325
rect 273978 73269 274046 73325
rect 274102 73269 274170 73325
rect 274226 73269 274294 73325
rect 274350 73269 274418 73325
rect 274474 73269 274542 73325
rect 274598 73269 274666 73325
rect 274722 73269 274802 73325
rect 272752 73201 274802 73269
rect 272752 73145 272806 73201
rect 272862 73145 272930 73201
rect 272986 73145 273054 73201
rect 273110 73145 273178 73201
rect 273234 73145 273302 73201
rect 273358 73145 273426 73201
rect 273482 73145 273550 73201
rect 273606 73145 273674 73201
rect 273730 73145 273798 73201
rect 273854 73145 273922 73201
rect 273978 73145 274046 73201
rect 274102 73145 274170 73201
rect 274226 73145 274294 73201
rect 274350 73145 274418 73201
rect 274474 73145 274542 73201
rect 274598 73145 274666 73201
rect 274722 73145 274802 73201
rect 272752 73077 274802 73145
rect 272752 73021 272806 73077
rect 272862 73021 272930 73077
rect 272986 73021 273054 73077
rect 273110 73021 273178 73077
rect 273234 73021 273302 73077
rect 273358 73021 273426 73077
rect 273482 73021 273550 73077
rect 273606 73021 273674 73077
rect 273730 73021 273798 73077
rect 273854 73021 273922 73077
rect 273978 73021 274046 73077
rect 274102 73021 274170 73077
rect 274226 73021 274294 73077
rect 274350 73021 274418 73077
rect 274474 73021 274542 73077
rect 274598 73021 274666 73077
rect 274722 73021 274802 73077
rect 272752 72953 274802 73021
rect 272752 72897 272806 72953
rect 272862 72897 272930 72953
rect 272986 72897 273054 72953
rect 273110 72897 273178 72953
rect 273234 72897 273302 72953
rect 273358 72897 273426 72953
rect 273482 72897 273550 72953
rect 273606 72897 273674 72953
rect 273730 72897 273798 72953
rect 273854 72897 273922 72953
rect 273978 72897 274046 72953
rect 274102 72897 274170 72953
rect 274226 72897 274294 72953
rect 274350 72897 274418 72953
rect 274474 72897 274542 72953
rect 274598 72897 274666 72953
rect 274722 72897 274802 72953
rect 272752 72829 274802 72897
rect 272752 72773 272806 72829
rect 272862 72773 272930 72829
rect 272986 72773 273054 72829
rect 273110 72773 273178 72829
rect 273234 72773 273302 72829
rect 273358 72773 273426 72829
rect 273482 72773 273550 72829
rect 273606 72773 273674 72829
rect 273730 72773 273798 72829
rect 273854 72773 273922 72829
rect 273978 72773 274046 72829
rect 274102 72773 274170 72829
rect 274226 72773 274294 72829
rect 274350 72773 274418 72829
rect 274474 72773 274542 72829
rect 274598 72773 274666 72829
rect 274722 72773 274802 72829
rect 272752 72705 274802 72773
rect 272752 72649 272806 72705
rect 272862 72649 272930 72705
rect 272986 72649 273054 72705
rect 273110 72649 273178 72705
rect 273234 72649 273302 72705
rect 273358 72649 273426 72705
rect 273482 72649 273550 72705
rect 273606 72649 273674 72705
rect 273730 72649 273798 72705
rect 273854 72649 273922 72705
rect 273978 72649 274046 72705
rect 274102 72649 274170 72705
rect 274226 72649 274294 72705
rect 274350 72649 274418 72705
rect 274474 72649 274542 72705
rect 274598 72649 274666 72705
rect 274722 72649 274802 72705
rect 272752 72581 274802 72649
rect 272752 72525 272806 72581
rect 272862 72525 272930 72581
rect 272986 72525 273054 72581
rect 273110 72525 273178 72581
rect 273234 72525 273302 72581
rect 273358 72525 273426 72581
rect 273482 72525 273550 72581
rect 273606 72525 273674 72581
rect 273730 72525 273798 72581
rect 273854 72525 273922 72581
rect 273978 72525 274046 72581
rect 274102 72525 274170 72581
rect 274226 72525 274294 72581
rect 274350 72525 274418 72581
rect 274474 72525 274542 72581
rect 274598 72525 274666 72581
rect 274722 72525 274802 72581
rect 272752 72457 274802 72525
rect 272752 72401 272806 72457
rect 272862 72401 272930 72457
rect 272986 72401 273054 72457
rect 273110 72401 273178 72457
rect 273234 72401 273302 72457
rect 273358 72401 273426 72457
rect 273482 72401 273550 72457
rect 273606 72401 273674 72457
rect 273730 72401 273798 72457
rect 273854 72401 273922 72457
rect 273978 72401 274046 72457
rect 274102 72401 274170 72457
rect 274226 72401 274294 72457
rect 274350 72401 274418 72457
rect 274474 72401 274542 72457
rect 274598 72401 274666 72457
rect 274722 72401 274802 72457
rect 272752 72333 274802 72401
rect 272752 72277 272806 72333
rect 272862 72277 272930 72333
rect 272986 72277 273054 72333
rect 273110 72277 273178 72333
rect 273234 72277 273302 72333
rect 273358 72277 273426 72333
rect 273482 72277 273550 72333
rect 273606 72277 273674 72333
rect 273730 72277 273798 72333
rect 273854 72277 273922 72333
rect 273978 72277 274046 72333
rect 274102 72277 274170 72333
rect 274226 72277 274294 72333
rect 274350 72277 274418 72333
rect 274474 72277 274542 72333
rect 274598 72277 274666 72333
rect 274722 72277 274802 72333
rect 272752 72209 274802 72277
rect 272752 72153 272806 72209
rect 272862 72153 272930 72209
rect 272986 72153 273054 72209
rect 273110 72153 273178 72209
rect 273234 72153 273302 72209
rect 273358 72153 273426 72209
rect 273482 72153 273550 72209
rect 273606 72153 273674 72209
rect 273730 72153 273798 72209
rect 273854 72153 273922 72209
rect 273978 72153 274046 72209
rect 274102 72153 274170 72209
rect 274226 72153 274294 72209
rect 274350 72153 274418 72209
rect 274474 72153 274542 72209
rect 274598 72153 274666 72209
rect 274722 72153 274802 72209
rect 272752 70000 274802 72153
rect 275122 73945 277172 74088
rect 275122 73889 275176 73945
rect 275232 73889 275300 73945
rect 275356 73889 275424 73945
rect 275480 73889 275548 73945
rect 275604 73889 275672 73945
rect 275728 73889 275796 73945
rect 275852 73889 275920 73945
rect 275976 73889 276044 73945
rect 276100 73889 276168 73945
rect 276224 73889 276292 73945
rect 276348 73889 276416 73945
rect 276472 73889 276540 73945
rect 276596 73889 276664 73945
rect 276720 73889 276788 73945
rect 276844 73889 276912 73945
rect 276968 73889 277036 73945
rect 277092 73889 277172 73945
rect 275122 73821 277172 73889
rect 275122 73765 275176 73821
rect 275232 73765 275300 73821
rect 275356 73765 275424 73821
rect 275480 73765 275548 73821
rect 275604 73765 275672 73821
rect 275728 73765 275796 73821
rect 275852 73765 275920 73821
rect 275976 73765 276044 73821
rect 276100 73765 276168 73821
rect 276224 73765 276292 73821
rect 276348 73765 276416 73821
rect 276472 73765 276540 73821
rect 276596 73765 276664 73821
rect 276720 73765 276788 73821
rect 276844 73765 276912 73821
rect 276968 73765 277036 73821
rect 277092 73765 277172 73821
rect 275122 73697 277172 73765
rect 275122 73641 275176 73697
rect 275232 73641 275300 73697
rect 275356 73641 275424 73697
rect 275480 73641 275548 73697
rect 275604 73641 275672 73697
rect 275728 73641 275796 73697
rect 275852 73641 275920 73697
rect 275976 73641 276044 73697
rect 276100 73641 276168 73697
rect 276224 73641 276292 73697
rect 276348 73641 276416 73697
rect 276472 73641 276540 73697
rect 276596 73641 276664 73697
rect 276720 73641 276788 73697
rect 276844 73641 276912 73697
rect 276968 73641 277036 73697
rect 277092 73641 277172 73697
rect 275122 73573 277172 73641
rect 275122 73517 275176 73573
rect 275232 73517 275300 73573
rect 275356 73517 275424 73573
rect 275480 73517 275548 73573
rect 275604 73517 275672 73573
rect 275728 73517 275796 73573
rect 275852 73517 275920 73573
rect 275976 73517 276044 73573
rect 276100 73517 276168 73573
rect 276224 73517 276292 73573
rect 276348 73517 276416 73573
rect 276472 73517 276540 73573
rect 276596 73517 276664 73573
rect 276720 73517 276788 73573
rect 276844 73517 276912 73573
rect 276968 73517 277036 73573
rect 277092 73517 277172 73573
rect 275122 73449 277172 73517
rect 275122 73393 275176 73449
rect 275232 73393 275300 73449
rect 275356 73393 275424 73449
rect 275480 73393 275548 73449
rect 275604 73393 275672 73449
rect 275728 73393 275796 73449
rect 275852 73393 275920 73449
rect 275976 73393 276044 73449
rect 276100 73393 276168 73449
rect 276224 73393 276292 73449
rect 276348 73393 276416 73449
rect 276472 73393 276540 73449
rect 276596 73393 276664 73449
rect 276720 73393 276788 73449
rect 276844 73393 276912 73449
rect 276968 73393 277036 73449
rect 277092 73393 277172 73449
rect 275122 73325 277172 73393
rect 275122 73269 275176 73325
rect 275232 73269 275300 73325
rect 275356 73269 275424 73325
rect 275480 73269 275548 73325
rect 275604 73269 275672 73325
rect 275728 73269 275796 73325
rect 275852 73269 275920 73325
rect 275976 73269 276044 73325
rect 276100 73269 276168 73325
rect 276224 73269 276292 73325
rect 276348 73269 276416 73325
rect 276472 73269 276540 73325
rect 276596 73269 276664 73325
rect 276720 73269 276788 73325
rect 276844 73269 276912 73325
rect 276968 73269 277036 73325
rect 277092 73269 277172 73325
rect 275122 73201 277172 73269
rect 275122 73145 275176 73201
rect 275232 73145 275300 73201
rect 275356 73145 275424 73201
rect 275480 73145 275548 73201
rect 275604 73145 275672 73201
rect 275728 73145 275796 73201
rect 275852 73145 275920 73201
rect 275976 73145 276044 73201
rect 276100 73145 276168 73201
rect 276224 73145 276292 73201
rect 276348 73145 276416 73201
rect 276472 73145 276540 73201
rect 276596 73145 276664 73201
rect 276720 73145 276788 73201
rect 276844 73145 276912 73201
rect 276968 73145 277036 73201
rect 277092 73145 277172 73201
rect 275122 73077 277172 73145
rect 275122 73021 275176 73077
rect 275232 73021 275300 73077
rect 275356 73021 275424 73077
rect 275480 73021 275548 73077
rect 275604 73021 275672 73077
rect 275728 73021 275796 73077
rect 275852 73021 275920 73077
rect 275976 73021 276044 73077
rect 276100 73021 276168 73077
rect 276224 73021 276292 73077
rect 276348 73021 276416 73077
rect 276472 73021 276540 73077
rect 276596 73021 276664 73077
rect 276720 73021 276788 73077
rect 276844 73021 276912 73077
rect 276968 73021 277036 73077
rect 277092 73021 277172 73077
rect 275122 72953 277172 73021
rect 275122 72897 275176 72953
rect 275232 72897 275300 72953
rect 275356 72897 275424 72953
rect 275480 72897 275548 72953
rect 275604 72897 275672 72953
rect 275728 72897 275796 72953
rect 275852 72897 275920 72953
rect 275976 72897 276044 72953
rect 276100 72897 276168 72953
rect 276224 72897 276292 72953
rect 276348 72897 276416 72953
rect 276472 72897 276540 72953
rect 276596 72897 276664 72953
rect 276720 72897 276788 72953
rect 276844 72897 276912 72953
rect 276968 72897 277036 72953
rect 277092 72897 277172 72953
rect 275122 72829 277172 72897
rect 275122 72773 275176 72829
rect 275232 72773 275300 72829
rect 275356 72773 275424 72829
rect 275480 72773 275548 72829
rect 275604 72773 275672 72829
rect 275728 72773 275796 72829
rect 275852 72773 275920 72829
rect 275976 72773 276044 72829
rect 276100 72773 276168 72829
rect 276224 72773 276292 72829
rect 276348 72773 276416 72829
rect 276472 72773 276540 72829
rect 276596 72773 276664 72829
rect 276720 72773 276788 72829
rect 276844 72773 276912 72829
rect 276968 72773 277036 72829
rect 277092 72773 277172 72829
rect 275122 72705 277172 72773
rect 275122 72649 275176 72705
rect 275232 72649 275300 72705
rect 275356 72649 275424 72705
rect 275480 72649 275548 72705
rect 275604 72649 275672 72705
rect 275728 72649 275796 72705
rect 275852 72649 275920 72705
rect 275976 72649 276044 72705
rect 276100 72649 276168 72705
rect 276224 72649 276292 72705
rect 276348 72649 276416 72705
rect 276472 72649 276540 72705
rect 276596 72649 276664 72705
rect 276720 72649 276788 72705
rect 276844 72649 276912 72705
rect 276968 72649 277036 72705
rect 277092 72649 277172 72705
rect 275122 72581 277172 72649
rect 275122 72525 275176 72581
rect 275232 72525 275300 72581
rect 275356 72525 275424 72581
rect 275480 72525 275548 72581
rect 275604 72525 275672 72581
rect 275728 72525 275796 72581
rect 275852 72525 275920 72581
rect 275976 72525 276044 72581
rect 276100 72525 276168 72581
rect 276224 72525 276292 72581
rect 276348 72525 276416 72581
rect 276472 72525 276540 72581
rect 276596 72525 276664 72581
rect 276720 72525 276788 72581
rect 276844 72525 276912 72581
rect 276968 72525 277036 72581
rect 277092 72525 277172 72581
rect 275122 72457 277172 72525
rect 275122 72401 275176 72457
rect 275232 72401 275300 72457
rect 275356 72401 275424 72457
rect 275480 72401 275548 72457
rect 275604 72401 275672 72457
rect 275728 72401 275796 72457
rect 275852 72401 275920 72457
rect 275976 72401 276044 72457
rect 276100 72401 276168 72457
rect 276224 72401 276292 72457
rect 276348 72401 276416 72457
rect 276472 72401 276540 72457
rect 276596 72401 276664 72457
rect 276720 72401 276788 72457
rect 276844 72401 276912 72457
rect 276968 72401 277036 72457
rect 277092 72401 277172 72457
rect 275122 72333 277172 72401
rect 275122 72277 275176 72333
rect 275232 72277 275300 72333
rect 275356 72277 275424 72333
rect 275480 72277 275548 72333
rect 275604 72277 275672 72333
rect 275728 72277 275796 72333
rect 275852 72277 275920 72333
rect 275976 72277 276044 72333
rect 276100 72277 276168 72333
rect 276224 72277 276292 72333
rect 276348 72277 276416 72333
rect 276472 72277 276540 72333
rect 276596 72277 276664 72333
rect 276720 72277 276788 72333
rect 276844 72277 276912 72333
rect 276968 72277 277036 72333
rect 277092 72277 277172 72333
rect 275122 72209 277172 72277
rect 275122 72153 275176 72209
rect 275232 72153 275300 72209
rect 275356 72153 275424 72209
rect 275480 72153 275548 72209
rect 275604 72153 275672 72209
rect 275728 72153 275796 72209
rect 275852 72153 275920 72209
rect 275976 72153 276044 72209
rect 276100 72153 276168 72209
rect 276224 72153 276292 72209
rect 276348 72153 276416 72209
rect 276472 72153 276540 72209
rect 276596 72153 276664 72209
rect 276720 72153 276788 72209
rect 276844 72153 276912 72209
rect 276968 72153 277036 72209
rect 277092 72153 277172 72209
rect 275122 70000 277172 72153
rect 277828 73945 279878 74088
rect 277828 73889 277882 73945
rect 277938 73889 278006 73945
rect 278062 73889 278130 73945
rect 278186 73889 278254 73945
rect 278310 73889 278378 73945
rect 278434 73889 278502 73945
rect 278558 73889 278626 73945
rect 278682 73889 278750 73945
rect 278806 73889 278874 73945
rect 278930 73889 278998 73945
rect 279054 73889 279122 73945
rect 279178 73889 279246 73945
rect 279302 73889 279370 73945
rect 279426 73889 279494 73945
rect 279550 73889 279618 73945
rect 279674 73889 279742 73945
rect 279798 73889 279878 73945
rect 277828 73821 279878 73889
rect 277828 73765 277882 73821
rect 277938 73765 278006 73821
rect 278062 73765 278130 73821
rect 278186 73765 278254 73821
rect 278310 73765 278378 73821
rect 278434 73765 278502 73821
rect 278558 73765 278626 73821
rect 278682 73765 278750 73821
rect 278806 73765 278874 73821
rect 278930 73765 278998 73821
rect 279054 73765 279122 73821
rect 279178 73765 279246 73821
rect 279302 73765 279370 73821
rect 279426 73765 279494 73821
rect 279550 73765 279618 73821
rect 279674 73765 279742 73821
rect 279798 73765 279878 73821
rect 277828 73697 279878 73765
rect 277828 73641 277882 73697
rect 277938 73641 278006 73697
rect 278062 73641 278130 73697
rect 278186 73641 278254 73697
rect 278310 73641 278378 73697
rect 278434 73641 278502 73697
rect 278558 73641 278626 73697
rect 278682 73641 278750 73697
rect 278806 73641 278874 73697
rect 278930 73641 278998 73697
rect 279054 73641 279122 73697
rect 279178 73641 279246 73697
rect 279302 73641 279370 73697
rect 279426 73641 279494 73697
rect 279550 73641 279618 73697
rect 279674 73641 279742 73697
rect 279798 73641 279878 73697
rect 277828 73573 279878 73641
rect 277828 73517 277882 73573
rect 277938 73517 278006 73573
rect 278062 73517 278130 73573
rect 278186 73517 278254 73573
rect 278310 73517 278378 73573
rect 278434 73517 278502 73573
rect 278558 73517 278626 73573
rect 278682 73517 278750 73573
rect 278806 73517 278874 73573
rect 278930 73517 278998 73573
rect 279054 73517 279122 73573
rect 279178 73517 279246 73573
rect 279302 73517 279370 73573
rect 279426 73517 279494 73573
rect 279550 73517 279618 73573
rect 279674 73517 279742 73573
rect 279798 73517 279878 73573
rect 277828 73449 279878 73517
rect 277828 73393 277882 73449
rect 277938 73393 278006 73449
rect 278062 73393 278130 73449
rect 278186 73393 278254 73449
rect 278310 73393 278378 73449
rect 278434 73393 278502 73449
rect 278558 73393 278626 73449
rect 278682 73393 278750 73449
rect 278806 73393 278874 73449
rect 278930 73393 278998 73449
rect 279054 73393 279122 73449
rect 279178 73393 279246 73449
rect 279302 73393 279370 73449
rect 279426 73393 279494 73449
rect 279550 73393 279618 73449
rect 279674 73393 279742 73449
rect 279798 73393 279878 73449
rect 277828 73325 279878 73393
rect 277828 73269 277882 73325
rect 277938 73269 278006 73325
rect 278062 73269 278130 73325
rect 278186 73269 278254 73325
rect 278310 73269 278378 73325
rect 278434 73269 278502 73325
rect 278558 73269 278626 73325
rect 278682 73269 278750 73325
rect 278806 73269 278874 73325
rect 278930 73269 278998 73325
rect 279054 73269 279122 73325
rect 279178 73269 279246 73325
rect 279302 73269 279370 73325
rect 279426 73269 279494 73325
rect 279550 73269 279618 73325
rect 279674 73269 279742 73325
rect 279798 73269 279878 73325
rect 277828 73201 279878 73269
rect 277828 73145 277882 73201
rect 277938 73145 278006 73201
rect 278062 73145 278130 73201
rect 278186 73145 278254 73201
rect 278310 73145 278378 73201
rect 278434 73145 278502 73201
rect 278558 73145 278626 73201
rect 278682 73145 278750 73201
rect 278806 73145 278874 73201
rect 278930 73145 278998 73201
rect 279054 73145 279122 73201
rect 279178 73145 279246 73201
rect 279302 73145 279370 73201
rect 279426 73145 279494 73201
rect 279550 73145 279618 73201
rect 279674 73145 279742 73201
rect 279798 73145 279878 73201
rect 277828 73077 279878 73145
rect 277828 73021 277882 73077
rect 277938 73021 278006 73077
rect 278062 73021 278130 73077
rect 278186 73021 278254 73077
rect 278310 73021 278378 73077
rect 278434 73021 278502 73077
rect 278558 73021 278626 73077
rect 278682 73021 278750 73077
rect 278806 73021 278874 73077
rect 278930 73021 278998 73077
rect 279054 73021 279122 73077
rect 279178 73021 279246 73077
rect 279302 73021 279370 73077
rect 279426 73021 279494 73077
rect 279550 73021 279618 73077
rect 279674 73021 279742 73077
rect 279798 73021 279878 73077
rect 277828 72953 279878 73021
rect 277828 72897 277882 72953
rect 277938 72897 278006 72953
rect 278062 72897 278130 72953
rect 278186 72897 278254 72953
rect 278310 72897 278378 72953
rect 278434 72897 278502 72953
rect 278558 72897 278626 72953
rect 278682 72897 278750 72953
rect 278806 72897 278874 72953
rect 278930 72897 278998 72953
rect 279054 72897 279122 72953
rect 279178 72897 279246 72953
rect 279302 72897 279370 72953
rect 279426 72897 279494 72953
rect 279550 72897 279618 72953
rect 279674 72897 279742 72953
rect 279798 72897 279878 72953
rect 277828 72829 279878 72897
rect 277828 72773 277882 72829
rect 277938 72773 278006 72829
rect 278062 72773 278130 72829
rect 278186 72773 278254 72829
rect 278310 72773 278378 72829
rect 278434 72773 278502 72829
rect 278558 72773 278626 72829
rect 278682 72773 278750 72829
rect 278806 72773 278874 72829
rect 278930 72773 278998 72829
rect 279054 72773 279122 72829
rect 279178 72773 279246 72829
rect 279302 72773 279370 72829
rect 279426 72773 279494 72829
rect 279550 72773 279618 72829
rect 279674 72773 279742 72829
rect 279798 72773 279878 72829
rect 277828 72705 279878 72773
rect 277828 72649 277882 72705
rect 277938 72649 278006 72705
rect 278062 72649 278130 72705
rect 278186 72649 278254 72705
rect 278310 72649 278378 72705
rect 278434 72649 278502 72705
rect 278558 72649 278626 72705
rect 278682 72649 278750 72705
rect 278806 72649 278874 72705
rect 278930 72649 278998 72705
rect 279054 72649 279122 72705
rect 279178 72649 279246 72705
rect 279302 72649 279370 72705
rect 279426 72649 279494 72705
rect 279550 72649 279618 72705
rect 279674 72649 279742 72705
rect 279798 72649 279878 72705
rect 277828 72581 279878 72649
rect 277828 72525 277882 72581
rect 277938 72525 278006 72581
rect 278062 72525 278130 72581
rect 278186 72525 278254 72581
rect 278310 72525 278378 72581
rect 278434 72525 278502 72581
rect 278558 72525 278626 72581
rect 278682 72525 278750 72581
rect 278806 72525 278874 72581
rect 278930 72525 278998 72581
rect 279054 72525 279122 72581
rect 279178 72525 279246 72581
rect 279302 72525 279370 72581
rect 279426 72525 279494 72581
rect 279550 72525 279618 72581
rect 279674 72525 279742 72581
rect 279798 72525 279878 72581
rect 277828 72457 279878 72525
rect 277828 72401 277882 72457
rect 277938 72401 278006 72457
rect 278062 72401 278130 72457
rect 278186 72401 278254 72457
rect 278310 72401 278378 72457
rect 278434 72401 278502 72457
rect 278558 72401 278626 72457
rect 278682 72401 278750 72457
rect 278806 72401 278874 72457
rect 278930 72401 278998 72457
rect 279054 72401 279122 72457
rect 279178 72401 279246 72457
rect 279302 72401 279370 72457
rect 279426 72401 279494 72457
rect 279550 72401 279618 72457
rect 279674 72401 279742 72457
rect 279798 72401 279878 72457
rect 277828 72333 279878 72401
rect 277828 72277 277882 72333
rect 277938 72277 278006 72333
rect 278062 72277 278130 72333
rect 278186 72277 278254 72333
rect 278310 72277 278378 72333
rect 278434 72277 278502 72333
rect 278558 72277 278626 72333
rect 278682 72277 278750 72333
rect 278806 72277 278874 72333
rect 278930 72277 278998 72333
rect 279054 72277 279122 72333
rect 279178 72277 279246 72333
rect 279302 72277 279370 72333
rect 279426 72277 279494 72333
rect 279550 72277 279618 72333
rect 279674 72277 279742 72333
rect 279798 72277 279878 72333
rect 277828 72209 279878 72277
rect 277828 72153 277882 72209
rect 277938 72153 278006 72209
rect 278062 72153 278130 72209
rect 278186 72153 278254 72209
rect 278310 72153 278378 72209
rect 278434 72153 278502 72209
rect 278558 72153 278626 72209
rect 278682 72153 278750 72209
rect 278806 72153 278874 72209
rect 278930 72153 278998 72209
rect 279054 72153 279122 72209
rect 279178 72153 279246 72209
rect 279302 72153 279370 72209
rect 279426 72153 279494 72209
rect 279550 72153 279618 72209
rect 279674 72153 279742 72209
rect 279798 72153 279878 72209
rect 277828 70000 279878 72153
rect 280198 73945 282248 74088
rect 280198 73889 280252 73945
rect 280308 73889 280376 73945
rect 280432 73889 280500 73945
rect 280556 73889 280624 73945
rect 280680 73889 280748 73945
rect 280804 73889 280872 73945
rect 280928 73889 280996 73945
rect 281052 73889 281120 73945
rect 281176 73889 281244 73945
rect 281300 73889 281368 73945
rect 281424 73889 281492 73945
rect 281548 73889 281616 73945
rect 281672 73889 281740 73945
rect 281796 73889 281864 73945
rect 281920 73889 281988 73945
rect 282044 73889 282112 73945
rect 282168 73889 282248 73945
rect 280198 73821 282248 73889
rect 280198 73765 280252 73821
rect 280308 73765 280376 73821
rect 280432 73765 280500 73821
rect 280556 73765 280624 73821
rect 280680 73765 280748 73821
rect 280804 73765 280872 73821
rect 280928 73765 280996 73821
rect 281052 73765 281120 73821
rect 281176 73765 281244 73821
rect 281300 73765 281368 73821
rect 281424 73765 281492 73821
rect 281548 73765 281616 73821
rect 281672 73765 281740 73821
rect 281796 73765 281864 73821
rect 281920 73765 281988 73821
rect 282044 73765 282112 73821
rect 282168 73765 282248 73821
rect 280198 73697 282248 73765
rect 280198 73641 280252 73697
rect 280308 73641 280376 73697
rect 280432 73641 280500 73697
rect 280556 73641 280624 73697
rect 280680 73641 280748 73697
rect 280804 73641 280872 73697
rect 280928 73641 280996 73697
rect 281052 73641 281120 73697
rect 281176 73641 281244 73697
rect 281300 73641 281368 73697
rect 281424 73641 281492 73697
rect 281548 73641 281616 73697
rect 281672 73641 281740 73697
rect 281796 73641 281864 73697
rect 281920 73641 281988 73697
rect 282044 73641 282112 73697
rect 282168 73641 282248 73697
rect 280198 73573 282248 73641
rect 280198 73517 280252 73573
rect 280308 73517 280376 73573
rect 280432 73517 280500 73573
rect 280556 73517 280624 73573
rect 280680 73517 280748 73573
rect 280804 73517 280872 73573
rect 280928 73517 280996 73573
rect 281052 73517 281120 73573
rect 281176 73517 281244 73573
rect 281300 73517 281368 73573
rect 281424 73517 281492 73573
rect 281548 73517 281616 73573
rect 281672 73517 281740 73573
rect 281796 73517 281864 73573
rect 281920 73517 281988 73573
rect 282044 73517 282112 73573
rect 282168 73517 282248 73573
rect 280198 73449 282248 73517
rect 280198 73393 280252 73449
rect 280308 73393 280376 73449
rect 280432 73393 280500 73449
rect 280556 73393 280624 73449
rect 280680 73393 280748 73449
rect 280804 73393 280872 73449
rect 280928 73393 280996 73449
rect 281052 73393 281120 73449
rect 281176 73393 281244 73449
rect 281300 73393 281368 73449
rect 281424 73393 281492 73449
rect 281548 73393 281616 73449
rect 281672 73393 281740 73449
rect 281796 73393 281864 73449
rect 281920 73393 281988 73449
rect 282044 73393 282112 73449
rect 282168 73393 282248 73449
rect 280198 73325 282248 73393
rect 280198 73269 280252 73325
rect 280308 73269 280376 73325
rect 280432 73269 280500 73325
rect 280556 73269 280624 73325
rect 280680 73269 280748 73325
rect 280804 73269 280872 73325
rect 280928 73269 280996 73325
rect 281052 73269 281120 73325
rect 281176 73269 281244 73325
rect 281300 73269 281368 73325
rect 281424 73269 281492 73325
rect 281548 73269 281616 73325
rect 281672 73269 281740 73325
rect 281796 73269 281864 73325
rect 281920 73269 281988 73325
rect 282044 73269 282112 73325
rect 282168 73269 282248 73325
rect 280198 73201 282248 73269
rect 280198 73145 280252 73201
rect 280308 73145 280376 73201
rect 280432 73145 280500 73201
rect 280556 73145 280624 73201
rect 280680 73145 280748 73201
rect 280804 73145 280872 73201
rect 280928 73145 280996 73201
rect 281052 73145 281120 73201
rect 281176 73145 281244 73201
rect 281300 73145 281368 73201
rect 281424 73145 281492 73201
rect 281548 73145 281616 73201
rect 281672 73145 281740 73201
rect 281796 73145 281864 73201
rect 281920 73145 281988 73201
rect 282044 73145 282112 73201
rect 282168 73145 282248 73201
rect 280198 73077 282248 73145
rect 280198 73021 280252 73077
rect 280308 73021 280376 73077
rect 280432 73021 280500 73077
rect 280556 73021 280624 73077
rect 280680 73021 280748 73077
rect 280804 73021 280872 73077
rect 280928 73021 280996 73077
rect 281052 73021 281120 73077
rect 281176 73021 281244 73077
rect 281300 73021 281368 73077
rect 281424 73021 281492 73077
rect 281548 73021 281616 73077
rect 281672 73021 281740 73077
rect 281796 73021 281864 73077
rect 281920 73021 281988 73077
rect 282044 73021 282112 73077
rect 282168 73021 282248 73077
rect 280198 72953 282248 73021
rect 280198 72897 280252 72953
rect 280308 72897 280376 72953
rect 280432 72897 280500 72953
rect 280556 72897 280624 72953
rect 280680 72897 280748 72953
rect 280804 72897 280872 72953
rect 280928 72897 280996 72953
rect 281052 72897 281120 72953
rect 281176 72897 281244 72953
rect 281300 72897 281368 72953
rect 281424 72897 281492 72953
rect 281548 72897 281616 72953
rect 281672 72897 281740 72953
rect 281796 72897 281864 72953
rect 281920 72897 281988 72953
rect 282044 72897 282112 72953
rect 282168 72897 282248 72953
rect 280198 72829 282248 72897
rect 280198 72773 280252 72829
rect 280308 72773 280376 72829
rect 280432 72773 280500 72829
rect 280556 72773 280624 72829
rect 280680 72773 280748 72829
rect 280804 72773 280872 72829
rect 280928 72773 280996 72829
rect 281052 72773 281120 72829
rect 281176 72773 281244 72829
rect 281300 72773 281368 72829
rect 281424 72773 281492 72829
rect 281548 72773 281616 72829
rect 281672 72773 281740 72829
rect 281796 72773 281864 72829
rect 281920 72773 281988 72829
rect 282044 72773 282112 72829
rect 282168 72773 282248 72829
rect 280198 72705 282248 72773
rect 280198 72649 280252 72705
rect 280308 72649 280376 72705
rect 280432 72649 280500 72705
rect 280556 72649 280624 72705
rect 280680 72649 280748 72705
rect 280804 72649 280872 72705
rect 280928 72649 280996 72705
rect 281052 72649 281120 72705
rect 281176 72649 281244 72705
rect 281300 72649 281368 72705
rect 281424 72649 281492 72705
rect 281548 72649 281616 72705
rect 281672 72649 281740 72705
rect 281796 72649 281864 72705
rect 281920 72649 281988 72705
rect 282044 72649 282112 72705
rect 282168 72649 282248 72705
rect 280198 72581 282248 72649
rect 280198 72525 280252 72581
rect 280308 72525 280376 72581
rect 280432 72525 280500 72581
rect 280556 72525 280624 72581
rect 280680 72525 280748 72581
rect 280804 72525 280872 72581
rect 280928 72525 280996 72581
rect 281052 72525 281120 72581
rect 281176 72525 281244 72581
rect 281300 72525 281368 72581
rect 281424 72525 281492 72581
rect 281548 72525 281616 72581
rect 281672 72525 281740 72581
rect 281796 72525 281864 72581
rect 281920 72525 281988 72581
rect 282044 72525 282112 72581
rect 282168 72525 282248 72581
rect 280198 72457 282248 72525
rect 280198 72401 280252 72457
rect 280308 72401 280376 72457
rect 280432 72401 280500 72457
rect 280556 72401 280624 72457
rect 280680 72401 280748 72457
rect 280804 72401 280872 72457
rect 280928 72401 280996 72457
rect 281052 72401 281120 72457
rect 281176 72401 281244 72457
rect 281300 72401 281368 72457
rect 281424 72401 281492 72457
rect 281548 72401 281616 72457
rect 281672 72401 281740 72457
rect 281796 72401 281864 72457
rect 281920 72401 281988 72457
rect 282044 72401 282112 72457
rect 282168 72401 282248 72457
rect 280198 72333 282248 72401
rect 280198 72277 280252 72333
rect 280308 72277 280376 72333
rect 280432 72277 280500 72333
rect 280556 72277 280624 72333
rect 280680 72277 280748 72333
rect 280804 72277 280872 72333
rect 280928 72277 280996 72333
rect 281052 72277 281120 72333
rect 281176 72277 281244 72333
rect 281300 72277 281368 72333
rect 281424 72277 281492 72333
rect 281548 72277 281616 72333
rect 281672 72277 281740 72333
rect 281796 72277 281864 72333
rect 281920 72277 281988 72333
rect 282044 72277 282112 72333
rect 282168 72277 282248 72333
rect 280198 72209 282248 72277
rect 280198 72153 280252 72209
rect 280308 72153 280376 72209
rect 280432 72153 280500 72209
rect 280556 72153 280624 72209
rect 280680 72153 280748 72209
rect 280804 72153 280872 72209
rect 280928 72153 280996 72209
rect 281052 72153 281120 72209
rect 281176 72153 281244 72209
rect 281300 72153 281368 72209
rect 281424 72153 281492 72209
rect 281548 72153 281616 72209
rect 281672 72153 281740 72209
rect 281796 72153 281864 72209
rect 281920 72153 281988 72209
rect 282044 72153 282112 72209
rect 282168 72153 282248 72209
rect 280198 70000 282248 72153
rect 282828 73945 284728 74088
rect 282828 73889 282882 73945
rect 282938 73889 283006 73945
rect 283062 73889 283130 73945
rect 283186 73889 283254 73945
rect 283310 73889 283378 73945
rect 283434 73889 283502 73945
rect 283558 73889 283626 73945
rect 283682 73889 283750 73945
rect 283806 73889 283874 73945
rect 283930 73889 284728 73945
rect 282828 73821 284728 73889
rect 282828 73765 282882 73821
rect 282938 73765 283006 73821
rect 283062 73765 283130 73821
rect 283186 73765 283254 73821
rect 283310 73765 283378 73821
rect 283434 73765 283502 73821
rect 283558 73765 283626 73821
rect 283682 73765 283750 73821
rect 283806 73765 283874 73821
rect 283930 73765 284728 73821
rect 282828 73697 284728 73765
rect 282828 73641 282882 73697
rect 282938 73641 283006 73697
rect 283062 73641 283130 73697
rect 283186 73641 283254 73697
rect 283310 73641 283378 73697
rect 283434 73641 283502 73697
rect 283558 73641 283626 73697
rect 283682 73641 283750 73697
rect 283806 73641 283874 73697
rect 283930 73641 284728 73697
rect 282828 73573 284728 73641
rect 282828 73517 282882 73573
rect 282938 73517 283006 73573
rect 283062 73517 283130 73573
rect 283186 73517 283254 73573
rect 283310 73517 283378 73573
rect 283434 73517 283502 73573
rect 283558 73517 283626 73573
rect 283682 73517 283750 73573
rect 283806 73517 283874 73573
rect 283930 73517 284728 73573
rect 282828 73449 284728 73517
rect 282828 73393 282882 73449
rect 282938 73393 283006 73449
rect 283062 73393 283130 73449
rect 283186 73393 283254 73449
rect 283310 73393 283378 73449
rect 283434 73393 283502 73449
rect 283558 73393 283626 73449
rect 283682 73393 283750 73449
rect 283806 73393 283874 73449
rect 283930 73393 284728 73449
rect 282828 73325 284728 73393
rect 282828 73269 282882 73325
rect 282938 73269 283006 73325
rect 283062 73269 283130 73325
rect 283186 73269 283254 73325
rect 283310 73269 283378 73325
rect 283434 73269 283502 73325
rect 283558 73269 283626 73325
rect 283682 73269 283750 73325
rect 283806 73269 283874 73325
rect 283930 73269 284728 73325
rect 282828 73201 284728 73269
rect 282828 73145 282882 73201
rect 282938 73145 283006 73201
rect 283062 73145 283130 73201
rect 283186 73145 283254 73201
rect 283310 73145 283378 73201
rect 283434 73145 283502 73201
rect 283558 73145 283626 73201
rect 283682 73145 283750 73201
rect 283806 73145 283874 73201
rect 283930 73145 284728 73201
rect 282828 73077 284728 73145
rect 282828 73021 282882 73077
rect 282938 73021 283006 73077
rect 283062 73021 283130 73077
rect 283186 73021 283254 73077
rect 283310 73021 283378 73077
rect 283434 73021 283502 73077
rect 283558 73021 283626 73077
rect 283682 73021 283750 73077
rect 283806 73021 283874 73077
rect 283930 73021 284728 73077
rect 282828 72953 284728 73021
rect 282828 72897 282882 72953
rect 282938 72897 283006 72953
rect 283062 72897 283130 72953
rect 283186 72897 283254 72953
rect 283310 72897 283378 72953
rect 283434 72897 283502 72953
rect 283558 72897 283626 72953
rect 283682 72897 283750 72953
rect 283806 72897 283874 72953
rect 283930 72897 284728 72953
rect 282828 72829 284728 72897
rect 282828 72773 282882 72829
rect 282938 72773 283006 72829
rect 283062 72773 283130 72829
rect 283186 72773 283254 72829
rect 283310 72773 283378 72829
rect 283434 72773 283502 72829
rect 283558 72773 283626 72829
rect 283682 72773 283750 72829
rect 283806 72773 283874 72829
rect 283930 72773 284728 72829
rect 282828 72705 284728 72773
rect 282828 72649 282882 72705
rect 282938 72649 283006 72705
rect 283062 72649 283130 72705
rect 283186 72649 283254 72705
rect 283310 72649 283378 72705
rect 283434 72649 283502 72705
rect 283558 72649 283626 72705
rect 283682 72649 283750 72705
rect 283806 72649 283874 72705
rect 283930 72649 284728 72705
rect 282828 72581 284728 72649
rect 282828 72525 282882 72581
rect 282938 72525 283006 72581
rect 283062 72525 283130 72581
rect 283186 72525 283254 72581
rect 283310 72525 283378 72581
rect 283434 72525 283502 72581
rect 283558 72525 283626 72581
rect 283682 72525 283750 72581
rect 283806 72525 283874 72581
rect 283930 72525 284728 72581
rect 282828 72457 284728 72525
rect 282828 72401 282882 72457
rect 282938 72401 283006 72457
rect 283062 72401 283130 72457
rect 283186 72401 283254 72457
rect 283310 72401 283378 72457
rect 283434 72401 283502 72457
rect 283558 72401 283626 72457
rect 283682 72401 283750 72457
rect 283806 72401 283874 72457
rect 283930 72401 284728 72457
rect 282828 72333 284728 72401
rect 282828 72277 282882 72333
rect 282938 72277 283006 72333
rect 283062 72277 283130 72333
rect 283186 72277 283254 72333
rect 283310 72277 283378 72333
rect 283434 72277 283502 72333
rect 283558 72277 283626 72333
rect 283682 72277 283750 72333
rect 283806 72277 283874 72333
rect 283930 72277 284728 72333
rect 282828 72209 284728 72277
rect 282828 72153 282882 72209
rect 282938 72153 283006 72209
rect 283062 72153 283130 72209
rect 283186 72153 283254 72209
rect 283310 72153 283378 72209
rect 283434 72153 283502 72209
rect 283558 72153 283626 72209
rect 283682 72153 283750 72209
rect 283806 72153 283874 72209
rect 283930 72153 284728 72209
rect 282828 70000 284728 72153
rect 600272 73945 602172 74088
rect 600272 73889 600326 73945
rect 600382 73889 600450 73945
rect 600506 73889 600574 73945
rect 600630 73889 600698 73945
rect 600754 73889 600822 73945
rect 600878 73889 600946 73945
rect 601002 73889 601070 73945
rect 601126 73889 601194 73945
rect 601250 73889 601318 73945
rect 601374 73889 601442 73945
rect 601498 73889 601566 73945
rect 601622 73889 601690 73945
rect 601746 73889 601814 73945
rect 601870 73889 601938 73945
rect 601994 73889 602062 73945
rect 602118 73889 602172 73945
rect 600272 73821 602172 73889
rect 600272 73765 600326 73821
rect 600382 73765 600450 73821
rect 600506 73765 600574 73821
rect 600630 73765 600698 73821
rect 600754 73765 600822 73821
rect 600878 73765 600946 73821
rect 601002 73765 601070 73821
rect 601126 73765 601194 73821
rect 601250 73765 601318 73821
rect 601374 73765 601442 73821
rect 601498 73765 601566 73821
rect 601622 73765 601690 73821
rect 601746 73765 601814 73821
rect 601870 73765 601938 73821
rect 601994 73765 602062 73821
rect 602118 73765 602172 73821
rect 600272 73697 602172 73765
rect 600272 73641 600326 73697
rect 600382 73641 600450 73697
rect 600506 73641 600574 73697
rect 600630 73641 600698 73697
rect 600754 73641 600822 73697
rect 600878 73641 600946 73697
rect 601002 73641 601070 73697
rect 601126 73641 601194 73697
rect 601250 73641 601318 73697
rect 601374 73641 601442 73697
rect 601498 73641 601566 73697
rect 601622 73641 601690 73697
rect 601746 73641 601814 73697
rect 601870 73641 601938 73697
rect 601994 73641 602062 73697
rect 602118 73641 602172 73697
rect 600272 73573 602172 73641
rect 600272 73517 600326 73573
rect 600382 73517 600450 73573
rect 600506 73517 600574 73573
rect 600630 73517 600698 73573
rect 600754 73517 600822 73573
rect 600878 73517 600946 73573
rect 601002 73517 601070 73573
rect 601126 73517 601194 73573
rect 601250 73517 601318 73573
rect 601374 73517 601442 73573
rect 601498 73517 601566 73573
rect 601622 73517 601690 73573
rect 601746 73517 601814 73573
rect 601870 73517 601938 73573
rect 601994 73517 602062 73573
rect 602118 73517 602172 73573
rect 600272 73449 602172 73517
rect 600272 73393 600326 73449
rect 600382 73393 600450 73449
rect 600506 73393 600574 73449
rect 600630 73393 600698 73449
rect 600754 73393 600822 73449
rect 600878 73393 600946 73449
rect 601002 73393 601070 73449
rect 601126 73393 601194 73449
rect 601250 73393 601318 73449
rect 601374 73393 601442 73449
rect 601498 73393 601566 73449
rect 601622 73393 601690 73449
rect 601746 73393 601814 73449
rect 601870 73393 601938 73449
rect 601994 73393 602062 73449
rect 602118 73393 602172 73449
rect 600272 73325 602172 73393
rect 600272 73269 600326 73325
rect 600382 73269 600450 73325
rect 600506 73269 600574 73325
rect 600630 73269 600698 73325
rect 600754 73269 600822 73325
rect 600878 73269 600946 73325
rect 601002 73269 601070 73325
rect 601126 73269 601194 73325
rect 601250 73269 601318 73325
rect 601374 73269 601442 73325
rect 601498 73269 601566 73325
rect 601622 73269 601690 73325
rect 601746 73269 601814 73325
rect 601870 73269 601938 73325
rect 601994 73269 602062 73325
rect 602118 73269 602172 73325
rect 600272 73201 602172 73269
rect 600272 73145 600326 73201
rect 600382 73145 600450 73201
rect 600506 73145 600574 73201
rect 600630 73145 600698 73201
rect 600754 73145 600822 73201
rect 600878 73145 600946 73201
rect 601002 73145 601070 73201
rect 601126 73145 601194 73201
rect 601250 73145 601318 73201
rect 601374 73145 601442 73201
rect 601498 73145 601566 73201
rect 601622 73145 601690 73201
rect 601746 73145 601814 73201
rect 601870 73145 601938 73201
rect 601994 73145 602062 73201
rect 602118 73145 602172 73201
rect 600272 73077 602172 73145
rect 600272 73021 600326 73077
rect 600382 73021 600450 73077
rect 600506 73021 600574 73077
rect 600630 73021 600698 73077
rect 600754 73021 600822 73077
rect 600878 73021 600946 73077
rect 601002 73021 601070 73077
rect 601126 73021 601194 73077
rect 601250 73021 601318 73077
rect 601374 73021 601442 73077
rect 601498 73021 601566 73077
rect 601622 73021 601690 73077
rect 601746 73021 601814 73077
rect 601870 73021 601938 73077
rect 601994 73021 602062 73077
rect 602118 73021 602172 73077
rect 600272 72953 602172 73021
rect 600272 72897 600326 72953
rect 600382 72897 600450 72953
rect 600506 72897 600574 72953
rect 600630 72897 600698 72953
rect 600754 72897 600822 72953
rect 600878 72897 600946 72953
rect 601002 72897 601070 72953
rect 601126 72897 601194 72953
rect 601250 72897 601318 72953
rect 601374 72897 601442 72953
rect 601498 72897 601566 72953
rect 601622 72897 601690 72953
rect 601746 72897 601814 72953
rect 601870 72897 601938 72953
rect 601994 72897 602062 72953
rect 602118 72897 602172 72953
rect 600272 72829 602172 72897
rect 600272 72773 600326 72829
rect 600382 72773 600450 72829
rect 600506 72773 600574 72829
rect 600630 72773 600698 72829
rect 600754 72773 600822 72829
rect 600878 72773 600946 72829
rect 601002 72773 601070 72829
rect 601126 72773 601194 72829
rect 601250 72773 601318 72829
rect 601374 72773 601442 72829
rect 601498 72773 601566 72829
rect 601622 72773 601690 72829
rect 601746 72773 601814 72829
rect 601870 72773 601938 72829
rect 601994 72773 602062 72829
rect 602118 72773 602172 72829
rect 600272 72705 602172 72773
rect 600272 72649 600326 72705
rect 600382 72649 600450 72705
rect 600506 72649 600574 72705
rect 600630 72649 600698 72705
rect 600754 72649 600822 72705
rect 600878 72649 600946 72705
rect 601002 72649 601070 72705
rect 601126 72649 601194 72705
rect 601250 72649 601318 72705
rect 601374 72649 601442 72705
rect 601498 72649 601566 72705
rect 601622 72649 601690 72705
rect 601746 72649 601814 72705
rect 601870 72649 601938 72705
rect 601994 72649 602062 72705
rect 602118 72649 602172 72705
rect 600272 72581 602172 72649
rect 600272 72525 600326 72581
rect 600382 72525 600450 72581
rect 600506 72525 600574 72581
rect 600630 72525 600698 72581
rect 600754 72525 600822 72581
rect 600878 72525 600946 72581
rect 601002 72525 601070 72581
rect 601126 72525 601194 72581
rect 601250 72525 601318 72581
rect 601374 72525 601442 72581
rect 601498 72525 601566 72581
rect 601622 72525 601690 72581
rect 601746 72525 601814 72581
rect 601870 72525 601938 72581
rect 601994 72525 602062 72581
rect 602118 72525 602172 72581
rect 600272 72457 602172 72525
rect 600272 72401 600326 72457
rect 600382 72401 600450 72457
rect 600506 72401 600574 72457
rect 600630 72401 600698 72457
rect 600754 72401 600822 72457
rect 600878 72401 600946 72457
rect 601002 72401 601070 72457
rect 601126 72401 601194 72457
rect 601250 72401 601318 72457
rect 601374 72401 601442 72457
rect 601498 72401 601566 72457
rect 601622 72401 601690 72457
rect 601746 72401 601814 72457
rect 601870 72401 601938 72457
rect 601994 72401 602062 72457
rect 602118 72401 602172 72457
rect 600272 72333 602172 72401
rect 600272 72277 600326 72333
rect 600382 72277 600450 72333
rect 600506 72277 600574 72333
rect 600630 72277 600698 72333
rect 600754 72277 600822 72333
rect 600878 72277 600946 72333
rect 601002 72277 601070 72333
rect 601126 72277 601194 72333
rect 601250 72277 601318 72333
rect 601374 72277 601442 72333
rect 601498 72277 601566 72333
rect 601622 72277 601690 72333
rect 601746 72277 601814 72333
rect 601870 72277 601938 72333
rect 601994 72277 602062 72333
rect 602118 72277 602172 72333
rect 600272 72209 602172 72277
rect 600272 72153 600326 72209
rect 600382 72153 600450 72209
rect 600506 72153 600574 72209
rect 600630 72153 600698 72209
rect 600754 72153 600822 72209
rect 600878 72153 600946 72209
rect 601002 72153 601070 72209
rect 601126 72153 601194 72209
rect 601250 72153 601318 72209
rect 601374 72153 601442 72209
rect 601498 72153 601566 72209
rect 601622 72153 601690 72209
rect 601746 72153 601814 72209
rect 601870 72153 601938 72209
rect 601994 72153 602062 72209
rect 602118 72153 602172 72209
rect 600272 70000 602172 72153
rect 602752 73945 604802 74088
rect 602752 73889 602806 73945
rect 602862 73889 602930 73945
rect 602986 73889 603054 73945
rect 603110 73889 603178 73945
rect 603234 73889 603302 73945
rect 603358 73889 603426 73945
rect 603482 73889 603550 73945
rect 603606 73889 603674 73945
rect 603730 73889 603798 73945
rect 603854 73889 603922 73945
rect 603978 73889 604802 73945
rect 602752 73821 604802 73889
rect 602752 73765 602806 73821
rect 602862 73765 602930 73821
rect 602986 73765 603054 73821
rect 603110 73765 603178 73821
rect 603234 73765 603302 73821
rect 603358 73765 603426 73821
rect 603482 73765 603550 73821
rect 603606 73765 603674 73821
rect 603730 73765 603798 73821
rect 603854 73765 603922 73821
rect 603978 73765 604802 73821
rect 602752 73697 604802 73765
rect 602752 73641 602806 73697
rect 602862 73641 602930 73697
rect 602986 73641 603054 73697
rect 603110 73641 603178 73697
rect 603234 73641 603302 73697
rect 603358 73641 603426 73697
rect 603482 73641 603550 73697
rect 603606 73641 603674 73697
rect 603730 73641 603798 73697
rect 603854 73641 603922 73697
rect 603978 73641 604802 73697
rect 602752 73573 604802 73641
rect 602752 73517 602806 73573
rect 602862 73517 602930 73573
rect 602986 73517 603054 73573
rect 603110 73517 603178 73573
rect 603234 73517 603302 73573
rect 603358 73517 603426 73573
rect 603482 73517 603550 73573
rect 603606 73517 603674 73573
rect 603730 73517 603798 73573
rect 603854 73517 603922 73573
rect 603978 73517 604802 73573
rect 602752 73449 604802 73517
rect 602752 73393 602806 73449
rect 602862 73393 602930 73449
rect 602986 73393 603054 73449
rect 603110 73393 603178 73449
rect 603234 73393 603302 73449
rect 603358 73393 603426 73449
rect 603482 73393 603550 73449
rect 603606 73393 603674 73449
rect 603730 73393 603798 73449
rect 603854 73393 603922 73449
rect 603978 73393 604802 73449
rect 602752 73325 604802 73393
rect 602752 73269 602806 73325
rect 602862 73269 602930 73325
rect 602986 73269 603054 73325
rect 603110 73269 603178 73325
rect 603234 73269 603302 73325
rect 603358 73269 603426 73325
rect 603482 73269 603550 73325
rect 603606 73269 603674 73325
rect 603730 73269 603798 73325
rect 603854 73269 603922 73325
rect 603978 73269 604802 73325
rect 602752 73201 604802 73269
rect 602752 73145 602806 73201
rect 602862 73145 602930 73201
rect 602986 73145 603054 73201
rect 603110 73145 603178 73201
rect 603234 73145 603302 73201
rect 603358 73145 603426 73201
rect 603482 73145 603550 73201
rect 603606 73145 603674 73201
rect 603730 73145 603798 73201
rect 603854 73145 603922 73201
rect 603978 73145 604802 73201
rect 602752 73077 604802 73145
rect 602752 73021 602806 73077
rect 602862 73021 602930 73077
rect 602986 73021 603054 73077
rect 603110 73021 603178 73077
rect 603234 73021 603302 73077
rect 603358 73021 603426 73077
rect 603482 73021 603550 73077
rect 603606 73021 603674 73077
rect 603730 73021 603798 73077
rect 603854 73021 603922 73077
rect 603978 73021 604802 73077
rect 602752 72953 604802 73021
rect 602752 72897 602806 72953
rect 602862 72897 602930 72953
rect 602986 72897 603054 72953
rect 603110 72897 603178 72953
rect 603234 72897 603302 72953
rect 603358 72897 603426 72953
rect 603482 72897 603550 72953
rect 603606 72897 603674 72953
rect 603730 72897 603798 72953
rect 603854 72897 603922 72953
rect 603978 72897 604802 72953
rect 602752 72829 604802 72897
rect 602752 72773 602806 72829
rect 602862 72773 602930 72829
rect 602986 72773 603054 72829
rect 603110 72773 603178 72829
rect 603234 72773 603302 72829
rect 603358 72773 603426 72829
rect 603482 72773 603550 72829
rect 603606 72773 603674 72829
rect 603730 72773 603798 72829
rect 603854 72773 603922 72829
rect 603978 72773 604802 72829
rect 602752 72705 604802 72773
rect 602752 72649 602806 72705
rect 602862 72649 602930 72705
rect 602986 72649 603054 72705
rect 603110 72649 603178 72705
rect 603234 72649 603302 72705
rect 603358 72649 603426 72705
rect 603482 72649 603550 72705
rect 603606 72649 603674 72705
rect 603730 72649 603798 72705
rect 603854 72649 603922 72705
rect 603978 72649 604802 72705
rect 602752 72581 604802 72649
rect 602752 72525 602806 72581
rect 602862 72525 602930 72581
rect 602986 72525 603054 72581
rect 603110 72525 603178 72581
rect 603234 72525 603302 72581
rect 603358 72525 603426 72581
rect 603482 72525 603550 72581
rect 603606 72525 603674 72581
rect 603730 72525 603798 72581
rect 603854 72525 603922 72581
rect 603978 72525 604802 72581
rect 602752 72457 604802 72525
rect 602752 72401 602806 72457
rect 602862 72401 602930 72457
rect 602986 72401 603054 72457
rect 603110 72401 603178 72457
rect 603234 72401 603302 72457
rect 603358 72401 603426 72457
rect 603482 72401 603550 72457
rect 603606 72401 603674 72457
rect 603730 72401 603798 72457
rect 603854 72401 603922 72457
rect 603978 72401 604802 72457
rect 602752 72333 604802 72401
rect 602752 72277 602806 72333
rect 602862 72277 602930 72333
rect 602986 72277 603054 72333
rect 603110 72277 603178 72333
rect 603234 72277 603302 72333
rect 603358 72277 603426 72333
rect 603482 72277 603550 72333
rect 603606 72277 603674 72333
rect 603730 72277 603798 72333
rect 603854 72277 603922 72333
rect 603978 72277 604802 72333
rect 602752 72209 604802 72277
rect 602752 72153 602806 72209
rect 602862 72153 602930 72209
rect 602986 72153 603054 72209
rect 603110 72153 603178 72209
rect 603234 72153 603302 72209
rect 603358 72153 603426 72209
rect 603482 72153 603550 72209
rect 603606 72153 603674 72209
rect 603730 72153 603798 72209
rect 603854 72153 603922 72209
rect 603978 72153 604802 72209
rect 602752 70000 604802 72153
rect 605122 73945 607172 74088
rect 605122 73889 605176 73945
rect 605232 73889 605300 73945
rect 605356 73889 605424 73945
rect 605480 73889 605548 73945
rect 605604 73889 605672 73945
rect 605728 73889 605796 73945
rect 605852 73889 605920 73945
rect 605976 73889 606044 73945
rect 606100 73889 606168 73945
rect 606224 73889 606292 73945
rect 606348 73889 606416 73945
rect 606472 73889 606540 73945
rect 606596 73889 606664 73945
rect 606720 73889 606788 73945
rect 606844 73889 606912 73945
rect 606968 73889 607036 73945
rect 607092 73889 607172 73945
rect 605122 73821 607172 73889
rect 605122 73765 605176 73821
rect 605232 73765 605300 73821
rect 605356 73765 605424 73821
rect 605480 73765 605548 73821
rect 605604 73765 605672 73821
rect 605728 73765 605796 73821
rect 605852 73765 605920 73821
rect 605976 73765 606044 73821
rect 606100 73765 606168 73821
rect 606224 73765 606292 73821
rect 606348 73765 606416 73821
rect 606472 73765 606540 73821
rect 606596 73765 606664 73821
rect 606720 73765 606788 73821
rect 606844 73765 606912 73821
rect 606968 73765 607036 73821
rect 607092 73765 607172 73821
rect 605122 73697 607172 73765
rect 605122 73641 605176 73697
rect 605232 73641 605300 73697
rect 605356 73641 605424 73697
rect 605480 73641 605548 73697
rect 605604 73641 605672 73697
rect 605728 73641 605796 73697
rect 605852 73641 605920 73697
rect 605976 73641 606044 73697
rect 606100 73641 606168 73697
rect 606224 73641 606292 73697
rect 606348 73641 606416 73697
rect 606472 73641 606540 73697
rect 606596 73641 606664 73697
rect 606720 73641 606788 73697
rect 606844 73641 606912 73697
rect 606968 73641 607036 73697
rect 607092 73641 607172 73697
rect 605122 73573 607172 73641
rect 605122 73517 605176 73573
rect 605232 73517 605300 73573
rect 605356 73517 605424 73573
rect 605480 73517 605548 73573
rect 605604 73517 605672 73573
rect 605728 73517 605796 73573
rect 605852 73517 605920 73573
rect 605976 73517 606044 73573
rect 606100 73517 606168 73573
rect 606224 73517 606292 73573
rect 606348 73517 606416 73573
rect 606472 73517 606540 73573
rect 606596 73517 606664 73573
rect 606720 73517 606788 73573
rect 606844 73517 606912 73573
rect 606968 73517 607036 73573
rect 607092 73517 607172 73573
rect 605122 73449 607172 73517
rect 605122 73393 605176 73449
rect 605232 73393 605300 73449
rect 605356 73393 605424 73449
rect 605480 73393 605548 73449
rect 605604 73393 605672 73449
rect 605728 73393 605796 73449
rect 605852 73393 605920 73449
rect 605976 73393 606044 73449
rect 606100 73393 606168 73449
rect 606224 73393 606292 73449
rect 606348 73393 606416 73449
rect 606472 73393 606540 73449
rect 606596 73393 606664 73449
rect 606720 73393 606788 73449
rect 606844 73393 606912 73449
rect 606968 73393 607036 73449
rect 607092 73393 607172 73449
rect 605122 73325 607172 73393
rect 605122 73269 605176 73325
rect 605232 73269 605300 73325
rect 605356 73269 605424 73325
rect 605480 73269 605548 73325
rect 605604 73269 605672 73325
rect 605728 73269 605796 73325
rect 605852 73269 605920 73325
rect 605976 73269 606044 73325
rect 606100 73269 606168 73325
rect 606224 73269 606292 73325
rect 606348 73269 606416 73325
rect 606472 73269 606540 73325
rect 606596 73269 606664 73325
rect 606720 73269 606788 73325
rect 606844 73269 606912 73325
rect 606968 73269 607036 73325
rect 607092 73269 607172 73325
rect 605122 73201 607172 73269
rect 605122 73145 605176 73201
rect 605232 73145 605300 73201
rect 605356 73145 605424 73201
rect 605480 73145 605548 73201
rect 605604 73145 605672 73201
rect 605728 73145 605796 73201
rect 605852 73145 605920 73201
rect 605976 73145 606044 73201
rect 606100 73145 606168 73201
rect 606224 73145 606292 73201
rect 606348 73145 606416 73201
rect 606472 73145 606540 73201
rect 606596 73145 606664 73201
rect 606720 73145 606788 73201
rect 606844 73145 606912 73201
rect 606968 73145 607036 73201
rect 607092 73145 607172 73201
rect 605122 73077 607172 73145
rect 605122 73021 605176 73077
rect 605232 73021 605300 73077
rect 605356 73021 605424 73077
rect 605480 73021 605548 73077
rect 605604 73021 605672 73077
rect 605728 73021 605796 73077
rect 605852 73021 605920 73077
rect 605976 73021 606044 73077
rect 606100 73021 606168 73077
rect 606224 73021 606292 73077
rect 606348 73021 606416 73077
rect 606472 73021 606540 73077
rect 606596 73021 606664 73077
rect 606720 73021 606788 73077
rect 606844 73021 606912 73077
rect 606968 73021 607036 73077
rect 607092 73021 607172 73077
rect 605122 72953 607172 73021
rect 605122 72897 605176 72953
rect 605232 72897 605300 72953
rect 605356 72897 605424 72953
rect 605480 72897 605548 72953
rect 605604 72897 605672 72953
rect 605728 72897 605796 72953
rect 605852 72897 605920 72953
rect 605976 72897 606044 72953
rect 606100 72897 606168 72953
rect 606224 72897 606292 72953
rect 606348 72897 606416 72953
rect 606472 72897 606540 72953
rect 606596 72897 606664 72953
rect 606720 72897 606788 72953
rect 606844 72897 606912 72953
rect 606968 72897 607036 72953
rect 607092 72897 607172 72953
rect 605122 72829 607172 72897
rect 605122 72773 605176 72829
rect 605232 72773 605300 72829
rect 605356 72773 605424 72829
rect 605480 72773 605548 72829
rect 605604 72773 605672 72829
rect 605728 72773 605796 72829
rect 605852 72773 605920 72829
rect 605976 72773 606044 72829
rect 606100 72773 606168 72829
rect 606224 72773 606292 72829
rect 606348 72773 606416 72829
rect 606472 72773 606540 72829
rect 606596 72773 606664 72829
rect 606720 72773 606788 72829
rect 606844 72773 606912 72829
rect 606968 72773 607036 72829
rect 607092 72773 607172 72829
rect 605122 72705 607172 72773
rect 605122 72649 605176 72705
rect 605232 72649 605300 72705
rect 605356 72649 605424 72705
rect 605480 72649 605548 72705
rect 605604 72649 605672 72705
rect 605728 72649 605796 72705
rect 605852 72649 605920 72705
rect 605976 72649 606044 72705
rect 606100 72649 606168 72705
rect 606224 72649 606292 72705
rect 606348 72649 606416 72705
rect 606472 72649 606540 72705
rect 606596 72649 606664 72705
rect 606720 72649 606788 72705
rect 606844 72649 606912 72705
rect 606968 72649 607036 72705
rect 607092 72649 607172 72705
rect 605122 72581 607172 72649
rect 605122 72525 605176 72581
rect 605232 72525 605300 72581
rect 605356 72525 605424 72581
rect 605480 72525 605548 72581
rect 605604 72525 605672 72581
rect 605728 72525 605796 72581
rect 605852 72525 605920 72581
rect 605976 72525 606044 72581
rect 606100 72525 606168 72581
rect 606224 72525 606292 72581
rect 606348 72525 606416 72581
rect 606472 72525 606540 72581
rect 606596 72525 606664 72581
rect 606720 72525 606788 72581
rect 606844 72525 606912 72581
rect 606968 72525 607036 72581
rect 607092 72525 607172 72581
rect 605122 72457 607172 72525
rect 605122 72401 605176 72457
rect 605232 72401 605300 72457
rect 605356 72401 605424 72457
rect 605480 72401 605548 72457
rect 605604 72401 605672 72457
rect 605728 72401 605796 72457
rect 605852 72401 605920 72457
rect 605976 72401 606044 72457
rect 606100 72401 606168 72457
rect 606224 72401 606292 72457
rect 606348 72401 606416 72457
rect 606472 72401 606540 72457
rect 606596 72401 606664 72457
rect 606720 72401 606788 72457
rect 606844 72401 606912 72457
rect 606968 72401 607036 72457
rect 607092 72401 607172 72457
rect 605122 72333 607172 72401
rect 605122 72277 605176 72333
rect 605232 72277 605300 72333
rect 605356 72277 605424 72333
rect 605480 72277 605548 72333
rect 605604 72277 605672 72333
rect 605728 72277 605796 72333
rect 605852 72277 605920 72333
rect 605976 72277 606044 72333
rect 606100 72277 606168 72333
rect 606224 72277 606292 72333
rect 606348 72277 606416 72333
rect 606472 72277 606540 72333
rect 606596 72277 606664 72333
rect 606720 72277 606788 72333
rect 606844 72277 606912 72333
rect 606968 72277 607036 72333
rect 607092 72277 607172 72333
rect 605122 72209 607172 72277
rect 605122 72153 605176 72209
rect 605232 72153 605300 72209
rect 605356 72153 605424 72209
rect 605480 72153 605548 72209
rect 605604 72153 605672 72209
rect 605728 72153 605796 72209
rect 605852 72153 605920 72209
rect 605976 72153 606044 72209
rect 606100 72153 606168 72209
rect 606224 72153 606292 72209
rect 606348 72153 606416 72209
rect 606472 72153 606540 72209
rect 606596 72153 606664 72209
rect 606720 72153 606788 72209
rect 606844 72153 606912 72209
rect 606968 72153 607036 72209
rect 607092 72153 607172 72209
rect 605122 70000 607172 72153
rect 607828 73945 609878 74088
rect 607828 73889 607882 73945
rect 607938 73889 608006 73945
rect 608062 73889 608130 73945
rect 608186 73889 608254 73945
rect 608310 73889 608378 73945
rect 608434 73889 608502 73945
rect 608558 73889 608626 73945
rect 608682 73889 608750 73945
rect 608806 73889 608874 73945
rect 608930 73889 608998 73945
rect 609054 73889 609122 73945
rect 609178 73889 609246 73945
rect 609302 73889 609370 73945
rect 609426 73889 609494 73945
rect 609550 73889 609618 73945
rect 609674 73889 609742 73945
rect 609798 73889 609878 73945
rect 607828 73821 609878 73889
rect 607828 73765 607882 73821
rect 607938 73765 608006 73821
rect 608062 73765 608130 73821
rect 608186 73765 608254 73821
rect 608310 73765 608378 73821
rect 608434 73765 608502 73821
rect 608558 73765 608626 73821
rect 608682 73765 608750 73821
rect 608806 73765 608874 73821
rect 608930 73765 608998 73821
rect 609054 73765 609122 73821
rect 609178 73765 609246 73821
rect 609302 73765 609370 73821
rect 609426 73765 609494 73821
rect 609550 73765 609618 73821
rect 609674 73765 609742 73821
rect 609798 73765 609878 73821
rect 607828 73697 609878 73765
rect 607828 73641 607882 73697
rect 607938 73641 608006 73697
rect 608062 73641 608130 73697
rect 608186 73641 608254 73697
rect 608310 73641 608378 73697
rect 608434 73641 608502 73697
rect 608558 73641 608626 73697
rect 608682 73641 608750 73697
rect 608806 73641 608874 73697
rect 608930 73641 608998 73697
rect 609054 73641 609122 73697
rect 609178 73641 609246 73697
rect 609302 73641 609370 73697
rect 609426 73641 609494 73697
rect 609550 73641 609618 73697
rect 609674 73641 609742 73697
rect 609798 73641 609878 73697
rect 607828 73573 609878 73641
rect 607828 73517 607882 73573
rect 607938 73517 608006 73573
rect 608062 73517 608130 73573
rect 608186 73517 608254 73573
rect 608310 73517 608378 73573
rect 608434 73517 608502 73573
rect 608558 73517 608626 73573
rect 608682 73517 608750 73573
rect 608806 73517 608874 73573
rect 608930 73517 608998 73573
rect 609054 73517 609122 73573
rect 609178 73517 609246 73573
rect 609302 73517 609370 73573
rect 609426 73517 609494 73573
rect 609550 73517 609618 73573
rect 609674 73517 609742 73573
rect 609798 73517 609878 73573
rect 607828 73449 609878 73517
rect 607828 73393 607882 73449
rect 607938 73393 608006 73449
rect 608062 73393 608130 73449
rect 608186 73393 608254 73449
rect 608310 73393 608378 73449
rect 608434 73393 608502 73449
rect 608558 73393 608626 73449
rect 608682 73393 608750 73449
rect 608806 73393 608874 73449
rect 608930 73393 608998 73449
rect 609054 73393 609122 73449
rect 609178 73393 609246 73449
rect 609302 73393 609370 73449
rect 609426 73393 609494 73449
rect 609550 73393 609618 73449
rect 609674 73393 609742 73449
rect 609798 73393 609878 73449
rect 607828 73325 609878 73393
rect 607828 73269 607882 73325
rect 607938 73269 608006 73325
rect 608062 73269 608130 73325
rect 608186 73269 608254 73325
rect 608310 73269 608378 73325
rect 608434 73269 608502 73325
rect 608558 73269 608626 73325
rect 608682 73269 608750 73325
rect 608806 73269 608874 73325
rect 608930 73269 608998 73325
rect 609054 73269 609122 73325
rect 609178 73269 609246 73325
rect 609302 73269 609370 73325
rect 609426 73269 609494 73325
rect 609550 73269 609618 73325
rect 609674 73269 609742 73325
rect 609798 73269 609878 73325
rect 607828 73201 609878 73269
rect 607828 73145 607882 73201
rect 607938 73145 608006 73201
rect 608062 73145 608130 73201
rect 608186 73145 608254 73201
rect 608310 73145 608378 73201
rect 608434 73145 608502 73201
rect 608558 73145 608626 73201
rect 608682 73145 608750 73201
rect 608806 73145 608874 73201
rect 608930 73145 608998 73201
rect 609054 73145 609122 73201
rect 609178 73145 609246 73201
rect 609302 73145 609370 73201
rect 609426 73145 609494 73201
rect 609550 73145 609618 73201
rect 609674 73145 609742 73201
rect 609798 73145 609878 73201
rect 607828 73077 609878 73145
rect 607828 73021 607882 73077
rect 607938 73021 608006 73077
rect 608062 73021 608130 73077
rect 608186 73021 608254 73077
rect 608310 73021 608378 73077
rect 608434 73021 608502 73077
rect 608558 73021 608626 73077
rect 608682 73021 608750 73077
rect 608806 73021 608874 73077
rect 608930 73021 608998 73077
rect 609054 73021 609122 73077
rect 609178 73021 609246 73077
rect 609302 73021 609370 73077
rect 609426 73021 609494 73077
rect 609550 73021 609618 73077
rect 609674 73021 609742 73077
rect 609798 73021 609878 73077
rect 607828 72953 609878 73021
rect 607828 72897 607882 72953
rect 607938 72897 608006 72953
rect 608062 72897 608130 72953
rect 608186 72897 608254 72953
rect 608310 72897 608378 72953
rect 608434 72897 608502 72953
rect 608558 72897 608626 72953
rect 608682 72897 608750 72953
rect 608806 72897 608874 72953
rect 608930 72897 608998 72953
rect 609054 72897 609122 72953
rect 609178 72897 609246 72953
rect 609302 72897 609370 72953
rect 609426 72897 609494 72953
rect 609550 72897 609618 72953
rect 609674 72897 609742 72953
rect 609798 72897 609878 72953
rect 607828 72829 609878 72897
rect 607828 72773 607882 72829
rect 607938 72773 608006 72829
rect 608062 72773 608130 72829
rect 608186 72773 608254 72829
rect 608310 72773 608378 72829
rect 608434 72773 608502 72829
rect 608558 72773 608626 72829
rect 608682 72773 608750 72829
rect 608806 72773 608874 72829
rect 608930 72773 608998 72829
rect 609054 72773 609122 72829
rect 609178 72773 609246 72829
rect 609302 72773 609370 72829
rect 609426 72773 609494 72829
rect 609550 72773 609618 72829
rect 609674 72773 609742 72829
rect 609798 72773 609878 72829
rect 607828 72705 609878 72773
rect 607828 72649 607882 72705
rect 607938 72649 608006 72705
rect 608062 72649 608130 72705
rect 608186 72649 608254 72705
rect 608310 72649 608378 72705
rect 608434 72649 608502 72705
rect 608558 72649 608626 72705
rect 608682 72649 608750 72705
rect 608806 72649 608874 72705
rect 608930 72649 608998 72705
rect 609054 72649 609122 72705
rect 609178 72649 609246 72705
rect 609302 72649 609370 72705
rect 609426 72649 609494 72705
rect 609550 72649 609618 72705
rect 609674 72649 609742 72705
rect 609798 72649 609878 72705
rect 607828 72581 609878 72649
rect 607828 72525 607882 72581
rect 607938 72525 608006 72581
rect 608062 72525 608130 72581
rect 608186 72525 608254 72581
rect 608310 72525 608378 72581
rect 608434 72525 608502 72581
rect 608558 72525 608626 72581
rect 608682 72525 608750 72581
rect 608806 72525 608874 72581
rect 608930 72525 608998 72581
rect 609054 72525 609122 72581
rect 609178 72525 609246 72581
rect 609302 72525 609370 72581
rect 609426 72525 609494 72581
rect 609550 72525 609618 72581
rect 609674 72525 609742 72581
rect 609798 72525 609878 72581
rect 607828 72457 609878 72525
rect 607828 72401 607882 72457
rect 607938 72401 608006 72457
rect 608062 72401 608130 72457
rect 608186 72401 608254 72457
rect 608310 72401 608378 72457
rect 608434 72401 608502 72457
rect 608558 72401 608626 72457
rect 608682 72401 608750 72457
rect 608806 72401 608874 72457
rect 608930 72401 608998 72457
rect 609054 72401 609122 72457
rect 609178 72401 609246 72457
rect 609302 72401 609370 72457
rect 609426 72401 609494 72457
rect 609550 72401 609618 72457
rect 609674 72401 609742 72457
rect 609798 72401 609878 72457
rect 607828 72333 609878 72401
rect 607828 72277 607882 72333
rect 607938 72277 608006 72333
rect 608062 72277 608130 72333
rect 608186 72277 608254 72333
rect 608310 72277 608378 72333
rect 608434 72277 608502 72333
rect 608558 72277 608626 72333
rect 608682 72277 608750 72333
rect 608806 72277 608874 72333
rect 608930 72277 608998 72333
rect 609054 72277 609122 72333
rect 609178 72277 609246 72333
rect 609302 72277 609370 72333
rect 609426 72277 609494 72333
rect 609550 72277 609618 72333
rect 609674 72277 609742 72333
rect 609798 72277 609878 72333
rect 607828 72209 609878 72277
rect 607828 72153 607882 72209
rect 607938 72153 608006 72209
rect 608062 72153 608130 72209
rect 608186 72153 608254 72209
rect 608310 72153 608378 72209
rect 608434 72153 608502 72209
rect 608558 72153 608626 72209
rect 608682 72153 608750 72209
rect 608806 72153 608874 72209
rect 608930 72153 608998 72209
rect 609054 72153 609122 72209
rect 609178 72153 609246 72209
rect 609302 72153 609370 72209
rect 609426 72153 609494 72209
rect 609550 72153 609618 72209
rect 609674 72153 609742 72209
rect 609798 72153 609878 72209
rect 607828 70000 609878 72153
rect 610198 73945 612248 74088
rect 610198 73889 610252 73945
rect 610308 73889 610376 73945
rect 610432 73889 610500 73945
rect 610556 73889 610624 73945
rect 610680 73889 610748 73945
rect 610804 73889 610872 73945
rect 610928 73889 610996 73945
rect 611052 73889 611120 73945
rect 611176 73889 611244 73945
rect 611300 73889 611368 73945
rect 611424 73889 611492 73945
rect 611548 73889 611616 73945
rect 611672 73889 611740 73945
rect 611796 73889 611864 73945
rect 611920 73889 611988 73945
rect 612044 73889 612112 73945
rect 612168 73889 612248 73945
rect 610198 73821 612248 73889
rect 610198 73765 610252 73821
rect 610308 73765 610376 73821
rect 610432 73765 610500 73821
rect 610556 73765 610624 73821
rect 610680 73765 610748 73821
rect 610804 73765 610872 73821
rect 610928 73765 610996 73821
rect 611052 73765 611120 73821
rect 611176 73765 611244 73821
rect 611300 73765 611368 73821
rect 611424 73765 611492 73821
rect 611548 73765 611616 73821
rect 611672 73765 611740 73821
rect 611796 73765 611864 73821
rect 611920 73765 611988 73821
rect 612044 73765 612112 73821
rect 612168 73765 612248 73821
rect 610198 73697 612248 73765
rect 610198 73641 610252 73697
rect 610308 73641 610376 73697
rect 610432 73641 610500 73697
rect 610556 73641 610624 73697
rect 610680 73641 610748 73697
rect 610804 73641 610872 73697
rect 610928 73641 610996 73697
rect 611052 73641 611120 73697
rect 611176 73641 611244 73697
rect 611300 73641 611368 73697
rect 611424 73641 611492 73697
rect 611548 73641 611616 73697
rect 611672 73641 611740 73697
rect 611796 73641 611864 73697
rect 611920 73641 611988 73697
rect 612044 73641 612112 73697
rect 612168 73641 612248 73697
rect 610198 73573 612248 73641
rect 610198 73517 610252 73573
rect 610308 73517 610376 73573
rect 610432 73517 610500 73573
rect 610556 73517 610624 73573
rect 610680 73517 610748 73573
rect 610804 73517 610872 73573
rect 610928 73517 610996 73573
rect 611052 73517 611120 73573
rect 611176 73517 611244 73573
rect 611300 73517 611368 73573
rect 611424 73517 611492 73573
rect 611548 73517 611616 73573
rect 611672 73517 611740 73573
rect 611796 73517 611864 73573
rect 611920 73517 611988 73573
rect 612044 73517 612112 73573
rect 612168 73517 612248 73573
rect 610198 73449 612248 73517
rect 610198 73393 610252 73449
rect 610308 73393 610376 73449
rect 610432 73393 610500 73449
rect 610556 73393 610624 73449
rect 610680 73393 610748 73449
rect 610804 73393 610872 73449
rect 610928 73393 610996 73449
rect 611052 73393 611120 73449
rect 611176 73393 611244 73449
rect 611300 73393 611368 73449
rect 611424 73393 611492 73449
rect 611548 73393 611616 73449
rect 611672 73393 611740 73449
rect 611796 73393 611864 73449
rect 611920 73393 611988 73449
rect 612044 73393 612112 73449
rect 612168 73393 612248 73449
rect 610198 73325 612248 73393
rect 610198 73269 610252 73325
rect 610308 73269 610376 73325
rect 610432 73269 610500 73325
rect 610556 73269 610624 73325
rect 610680 73269 610748 73325
rect 610804 73269 610872 73325
rect 610928 73269 610996 73325
rect 611052 73269 611120 73325
rect 611176 73269 611244 73325
rect 611300 73269 611368 73325
rect 611424 73269 611492 73325
rect 611548 73269 611616 73325
rect 611672 73269 611740 73325
rect 611796 73269 611864 73325
rect 611920 73269 611988 73325
rect 612044 73269 612112 73325
rect 612168 73269 612248 73325
rect 610198 73201 612248 73269
rect 610198 73145 610252 73201
rect 610308 73145 610376 73201
rect 610432 73145 610500 73201
rect 610556 73145 610624 73201
rect 610680 73145 610748 73201
rect 610804 73145 610872 73201
rect 610928 73145 610996 73201
rect 611052 73145 611120 73201
rect 611176 73145 611244 73201
rect 611300 73145 611368 73201
rect 611424 73145 611492 73201
rect 611548 73145 611616 73201
rect 611672 73145 611740 73201
rect 611796 73145 611864 73201
rect 611920 73145 611988 73201
rect 612044 73145 612112 73201
rect 612168 73145 612248 73201
rect 610198 73077 612248 73145
rect 610198 73021 610252 73077
rect 610308 73021 610376 73077
rect 610432 73021 610500 73077
rect 610556 73021 610624 73077
rect 610680 73021 610748 73077
rect 610804 73021 610872 73077
rect 610928 73021 610996 73077
rect 611052 73021 611120 73077
rect 611176 73021 611244 73077
rect 611300 73021 611368 73077
rect 611424 73021 611492 73077
rect 611548 73021 611616 73077
rect 611672 73021 611740 73077
rect 611796 73021 611864 73077
rect 611920 73021 611988 73077
rect 612044 73021 612112 73077
rect 612168 73021 612248 73077
rect 610198 72953 612248 73021
rect 610198 72897 610252 72953
rect 610308 72897 610376 72953
rect 610432 72897 610500 72953
rect 610556 72897 610624 72953
rect 610680 72897 610748 72953
rect 610804 72897 610872 72953
rect 610928 72897 610996 72953
rect 611052 72897 611120 72953
rect 611176 72897 611244 72953
rect 611300 72897 611368 72953
rect 611424 72897 611492 72953
rect 611548 72897 611616 72953
rect 611672 72897 611740 72953
rect 611796 72897 611864 72953
rect 611920 72897 611988 72953
rect 612044 72897 612112 72953
rect 612168 72897 612248 72953
rect 610198 72829 612248 72897
rect 610198 72773 610252 72829
rect 610308 72773 610376 72829
rect 610432 72773 610500 72829
rect 610556 72773 610624 72829
rect 610680 72773 610748 72829
rect 610804 72773 610872 72829
rect 610928 72773 610996 72829
rect 611052 72773 611120 72829
rect 611176 72773 611244 72829
rect 611300 72773 611368 72829
rect 611424 72773 611492 72829
rect 611548 72773 611616 72829
rect 611672 72773 611740 72829
rect 611796 72773 611864 72829
rect 611920 72773 611988 72829
rect 612044 72773 612112 72829
rect 612168 72773 612248 72829
rect 610198 72705 612248 72773
rect 610198 72649 610252 72705
rect 610308 72649 610376 72705
rect 610432 72649 610500 72705
rect 610556 72649 610624 72705
rect 610680 72649 610748 72705
rect 610804 72649 610872 72705
rect 610928 72649 610996 72705
rect 611052 72649 611120 72705
rect 611176 72649 611244 72705
rect 611300 72649 611368 72705
rect 611424 72649 611492 72705
rect 611548 72649 611616 72705
rect 611672 72649 611740 72705
rect 611796 72649 611864 72705
rect 611920 72649 611988 72705
rect 612044 72649 612112 72705
rect 612168 72649 612248 72705
rect 610198 72581 612248 72649
rect 610198 72525 610252 72581
rect 610308 72525 610376 72581
rect 610432 72525 610500 72581
rect 610556 72525 610624 72581
rect 610680 72525 610748 72581
rect 610804 72525 610872 72581
rect 610928 72525 610996 72581
rect 611052 72525 611120 72581
rect 611176 72525 611244 72581
rect 611300 72525 611368 72581
rect 611424 72525 611492 72581
rect 611548 72525 611616 72581
rect 611672 72525 611740 72581
rect 611796 72525 611864 72581
rect 611920 72525 611988 72581
rect 612044 72525 612112 72581
rect 612168 72525 612248 72581
rect 610198 72457 612248 72525
rect 610198 72401 610252 72457
rect 610308 72401 610376 72457
rect 610432 72401 610500 72457
rect 610556 72401 610624 72457
rect 610680 72401 610748 72457
rect 610804 72401 610872 72457
rect 610928 72401 610996 72457
rect 611052 72401 611120 72457
rect 611176 72401 611244 72457
rect 611300 72401 611368 72457
rect 611424 72401 611492 72457
rect 611548 72401 611616 72457
rect 611672 72401 611740 72457
rect 611796 72401 611864 72457
rect 611920 72401 611988 72457
rect 612044 72401 612112 72457
rect 612168 72401 612248 72457
rect 610198 72333 612248 72401
rect 610198 72277 610252 72333
rect 610308 72277 610376 72333
rect 610432 72277 610500 72333
rect 610556 72277 610624 72333
rect 610680 72277 610748 72333
rect 610804 72277 610872 72333
rect 610928 72277 610996 72333
rect 611052 72277 611120 72333
rect 611176 72277 611244 72333
rect 611300 72277 611368 72333
rect 611424 72277 611492 72333
rect 611548 72277 611616 72333
rect 611672 72277 611740 72333
rect 611796 72277 611864 72333
rect 611920 72277 611988 72333
rect 612044 72277 612112 72333
rect 612168 72277 612248 72333
rect 610198 72209 612248 72277
rect 610198 72153 610252 72209
rect 610308 72153 610376 72209
rect 610432 72153 610500 72209
rect 610556 72153 610624 72209
rect 610680 72153 610748 72209
rect 610804 72153 610872 72209
rect 610928 72153 610996 72209
rect 611052 72153 611120 72209
rect 611176 72153 611244 72209
rect 611300 72153 611368 72209
rect 611424 72153 611492 72209
rect 611548 72153 611616 72209
rect 611672 72153 611740 72209
rect 611796 72153 611864 72209
rect 611920 72153 611988 72209
rect 612044 72153 612112 72209
rect 612168 72153 612248 72209
rect 610198 70000 612248 72153
rect 612828 73945 614728 74088
rect 612828 73889 612882 73945
rect 612938 73889 613006 73945
rect 613062 73889 613130 73945
rect 613186 73889 613254 73945
rect 613310 73889 613378 73945
rect 613434 73889 613502 73945
rect 613558 73889 613626 73945
rect 613682 73889 613750 73945
rect 613806 73889 613874 73945
rect 613930 73889 613998 73945
rect 614054 73889 614122 73945
rect 614178 73889 614246 73945
rect 614302 73889 614370 73945
rect 614426 73889 614494 73945
rect 614550 73889 614618 73945
rect 614674 73889 614728 73945
rect 612828 73821 614728 73889
rect 612828 73765 612882 73821
rect 612938 73765 613006 73821
rect 613062 73765 613130 73821
rect 613186 73765 613254 73821
rect 613310 73765 613378 73821
rect 613434 73765 613502 73821
rect 613558 73765 613626 73821
rect 613682 73765 613750 73821
rect 613806 73765 613874 73821
rect 613930 73765 613998 73821
rect 614054 73765 614122 73821
rect 614178 73765 614246 73821
rect 614302 73765 614370 73821
rect 614426 73765 614494 73821
rect 614550 73765 614618 73821
rect 614674 73765 614728 73821
rect 612828 73697 614728 73765
rect 612828 73641 612882 73697
rect 612938 73641 613006 73697
rect 613062 73641 613130 73697
rect 613186 73641 613254 73697
rect 613310 73641 613378 73697
rect 613434 73641 613502 73697
rect 613558 73641 613626 73697
rect 613682 73641 613750 73697
rect 613806 73641 613874 73697
rect 613930 73641 613998 73697
rect 614054 73641 614122 73697
rect 614178 73641 614246 73697
rect 614302 73641 614370 73697
rect 614426 73641 614494 73697
rect 614550 73641 614618 73697
rect 614674 73641 614728 73697
rect 612828 73573 614728 73641
rect 612828 73517 612882 73573
rect 612938 73517 613006 73573
rect 613062 73517 613130 73573
rect 613186 73517 613254 73573
rect 613310 73517 613378 73573
rect 613434 73517 613502 73573
rect 613558 73517 613626 73573
rect 613682 73517 613750 73573
rect 613806 73517 613874 73573
rect 613930 73517 613998 73573
rect 614054 73517 614122 73573
rect 614178 73517 614246 73573
rect 614302 73517 614370 73573
rect 614426 73517 614494 73573
rect 614550 73517 614618 73573
rect 614674 73517 614728 73573
rect 612828 73449 614728 73517
rect 612828 73393 612882 73449
rect 612938 73393 613006 73449
rect 613062 73393 613130 73449
rect 613186 73393 613254 73449
rect 613310 73393 613378 73449
rect 613434 73393 613502 73449
rect 613558 73393 613626 73449
rect 613682 73393 613750 73449
rect 613806 73393 613874 73449
rect 613930 73393 613998 73449
rect 614054 73393 614122 73449
rect 614178 73393 614246 73449
rect 614302 73393 614370 73449
rect 614426 73393 614494 73449
rect 614550 73393 614618 73449
rect 614674 73393 614728 73449
rect 612828 73325 614728 73393
rect 612828 73269 612882 73325
rect 612938 73269 613006 73325
rect 613062 73269 613130 73325
rect 613186 73269 613254 73325
rect 613310 73269 613378 73325
rect 613434 73269 613502 73325
rect 613558 73269 613626 73325
rect 613682 73269 613750 73325
rect 613806 73269 613874 73325
rect 613930 73269 613998 73325
rect 614054 73269 614122 73325
rect 614178 73269 614246 73325
rect 614302 73269 614370 73325
rect 614426 73269 614494 73325
rect 614550 73269 614618 73325
rect 614674 73269 614728 73325
rect 612828 73201 614728 73269
rect 612828 73145 612882 73201
rect 612938 73145 613006 73201
rect 613062 73145 613130 73201
rect 613186 73145 613254 73201
rect 613310 73145 613378 73201
rect 613434 73145 613502 73201
rect 613558 73145 613626 73201
rect 613682 73145 613750 73201
rect 613806 73145 613874 73201
rect 613930 73145 613998 73201
rect 614054 73145 614122 73201
rect 614178 73145 614246 73201
rect 614302 73145 614370 73201
rect 614426 73145 614494 73201
rect 614550 73145 614618 73201
rect 614674 73145 614728 73201
rect 612828 73077 614728 73145
rect 612828 73021 612882 73077
rect 612938 73021 613006 73077
rect 613062 73021 613130 73077
rect 613186 73021 613254 73077
rect 613310 73021 613378 73077
rect 613434 73021 613502 73077
rect 613558 73021 613626 73077
rect 613682 73021 613750 73077
rect 613806 73021 613874 73077
rect 613930 73021 613998 73077
rect 614054 73021 614122 73077
rect 614178 73021 614246 73077
rect 614302 73021 614370 73077
rect 614426 73021 614494 73077
rect 614550 73021 614618 73077
rect 614674 73021 614728 73077
rect 612828 72953 614728 73021
rect 612828 72897 612882 72953
rect 612938 72897 613006 72953
rect 613062 72897 613130 72953
rect 613186 72897 613254 72953
rect 613310 72897 613378 72953
rect 613434 72897 613502 72953
rect 613558 72897 613626 72953
rect 613682 72897 613750 72953
rect 613806 72897 613874 72953
rect 613930 72897 613998 72953
rect 614054 72897 614122 72953
rect 614178 72897 614246 72953
rect 614302 72897 614370 72953
rect 614426 72897 614494 72953
rect 614550 72897 614618 72953
rect 614674 72897 614728 72953
rect 612828 72829 614728 72897
rect 612828 72773 612882 72829
rect 612938 72773 613006 72829
rect 613062 72773 613130 72829
rect 613186 72773 613254 72829
rect 613310 72773 613378 72829
rect 613434 72773 613502 72829
rect 613558 72773 613626 72829
rect 613682 72773 613750 72829
rect 613806 72773 613874 72829
rect 613930 72773 613998 72829
rect 614054 72773 614122 72829
rect 614178 72773 614246 72829
rect 614302 72773 614370 72829
rect 614426 72773 614494 72829
rect 614550 72773 614618 72829
rect 614674 72773 614728 72829
rect 612828 72705 614728 72773
rect 612828 72649 612882 72705
rect 612938 72649 613006 72705
rect 613062 72649 613130 72705
rect 613186 72649 613254 72705
rect 613310 72649 613378 72705
rect 613434 72649 613502 72705
rect 613558 72649 613626 72705
rect 613682 72649 613750 72705
rect 613806 72649 613874 72705
rect 613930 72649 613998 72705
rect 614054 72649 614122 72705
rect 614178 72649 614246 72705
rect 614302 72649 614370 72705
rect 614426 72649 614494 72705
rect 614550 72649 614618 72705
rect 614674 72649 614728 72705
rect 612828 72581 614728 72649
rect 612828 72525 612882 72581
rect 612938 72525 613006 72581
rect 613062 72525 613130 72581
rect 613186 72525 613254 72581
rect 613310 72525 613378 72581
rect 613434 72525 613502 72581
rect 613558 72525 613626 72581
rect 613682 72525 613750 72581
rect 613806 72525 613874 72581
rect 613930 72525 613998 72581
rect 614054 72525 614122 72581
rect 614178 72525 614246 72581
rect 614302 72525 614370 72581
rect 614426 72525 614494 72581
rect 614550 72525 614618 72581
rect 614674 72525 614728 72581
rect 612828 72457 614728 72525
rect 612828 72401 612882 72457
rect 612938 72401 613006 72457
rect 613062 72401 613130 72457
rect 613186 72401 613254 72457
rect 613310 72401 613378 72457
rect 613434 72401 613502 72457
rect 613558 72401 613626 72457
rect 613682 72401 613750 72457
rect 613806 72401 613874 72457
rect 613930 72401 613998 72457
rect 614054 72401 614122 72457
rect 614178 72401 614246 72457
rect 614302 72401 614370 72457
rect 614426 72401 614494 72457
rect 614550 72401 614618 72457
rect 614674 72401 614728 72457
rect 612828 72333 614728 72401
rect 612828 72277 612882 72333
rect 612938 72277 613006 72333
rect 613062 72277 613130 72333
rect 613186 72277 613254 72333
rect 613310 72277 613378 72333
rect 613434 72277 613502 72333
rect 613558 72277 613626 72333
rect 613682 72277 613750 72333
rect 613806 72277 613874 72333
rect 613930 72277 613998 72333
rect 614054 72277 614122 72333
rect 614178 72277 614246 72333
rect 614302 72277 614370 72333
rect 614426 72277 614494 72333
rect 614550 72277 614618 72333
rect 614674 72277 614728 72333
rect 612828 72209 614728 72277
rect 612828 72153 612882 72209
rect 612938 72153 613006 72209
rect 613062 72153 613130 72209
rect 613186 72153 613254 72209
rect 613310 72153 613378 72209
rect 613434 72153 613502 72209
rect 613558 72153 613626 72209
rect 613682 72153 613750 72209
rect 613806 72153 613874 72209
rect 613930 72153 613998 72209
rect 614054 72153 614122 72209
rect 614178 72153 614246 72209
rect 614302 72153 614370 72209
rect 614426 72153 614494 72209
rect 614550 72153 614618 72209
rect 614674 72153 614728 72209
rect 612828 70000 614728 72153
rect 655272 70000 657172 74525
rect 657752 75945 659802 76088
rect 657752 75889 657806 75945
rect 657862 75889 657930 75945
rect 657986 75889 658054 75945
rect 658110 75889 658178 75945
rect 658234 75889 658302 75945
rect 658358 75889 658426 75945
rect 658482 75889 658550 75945
rect 658606 75889 658674 75945
rect 658730 75889 658798 75945
rect 658854 75889 658922 75945
rect 658978 75889 659046 75945
rect 659102 75889 659170 75945
rect 659226 75889 659294 75945
rect 659350 75889 659418 75945
rect 659474 75889 659542 75945
rect 659598 75889 659666 75945
rect 659722 75889 659802 75945
rect 657752 75821 659802 75889
rect 657752 75765 657806 75821
rect 657862 75765 657930 75821
rect 657986 75765 658054 75821
rect 658110 75765 658178 75821
rect 658234 75765 658302 75821
rect 658358 75765 658426 75821
rect 658482 75765 658550 75821
rect 658606 75765 658674 75821
rect 658730 75765 658798 75821
rect 658854 75765 658922 75821
rect 658978 75765 659046 75821
rect 659102 75765 659170 75821
rect 659226 75765 659294 75821
rect 659350 75765 659418 75821
rect 659474 75765 659542 75821
rect 659598 75765 659666 75821
rect 659722 75765 659802 75821
rect 657752 75697 659802 75765
rect 657752 75641 657806 75697
rect 657862 75641 657930 75697
rect 657986 75641 658054 75697
rect 658110 75641 658178 75697
rect 658234 75641 658302 75697
rect 658358 75641 658426 75697
rect 658482 75641 658550 75697
rect 658606 75641 658674 75697
rect 658730 75641 658798 75697
rect 658854 75641 658922 75697
rect 658978 75641 659046 75697
rect 659102 75641 659170 75697
rect 659226 75641 659294 75697
rect 659350 75641 659418 75697
rect 659474 75641 659542 75697
rect 659598 75641 659666 75697
rect 659722 75641 659802 75697
rect 657752 75573 659802 75641
rect 657752 75517 657806 75573
rect 657862 75517 657930 75573
rect 657986 75517 658054 75573
rect 658110 75517 658178 75573
rect 658234 75517 658302 75573
rect 658358 75517 658426 75573
rect 658482 75517 658550 75573
rect 658606 75517 658674 75573
rect 658730 75517 658798 75573
rect 658854 75517 658922 75573
rect 658978 75517 659046 75573
rect 659102 75517 659170 75573
rect 659226 75517 659294 75573
rect 659350 75517 659418 75573
rect 659474 75517 659542 75573
rect 659598 75517 659666 75573
rect 659722 75517 659802 75573
rect 657752 75449 659802 75517
rect 657752 75393 657806 75449
rect 657862 75393 657930 75449
rect 657986 75393 658054 75449
rect 658110 75393 658178 75449
rect 658234 75393 658302 75449
rect 658358 75393 658426 75449
rect 658482 75393 658550 75449
rect 658606 75393 658674 75449
rect 658730 75393 658798 75449
rect 658854 75393 658922 75449
rect 658978 75393 659046 75449
rect 659102 75393 659170 75449
rect 659226 75393 659294 75449
rect 659350 75393 659418 75449
rect 659474 75393 659542 75449
rect 659598 75393 659666 75449
rect 659722 75393 659802 75449
rect 657752 75325 659802 75393
rect 657752 75269 657806 75325
rect 657862 75269 657930 75325
rect 657986 75269 658054 75325
rect 658110 75269 658178 75325
rect 658234 75269 658302 75325
rect 658358 75269 658426 75325
rect 658482 75269 658550 75325
rect 658606 75269 658674 75325
rect 658730 75269 658798 75325
rect 658854 75269 658922 75325
rect 658978 75269 659046 75325
rect 659102 75269 659170 75325
rect 659226 75269 659294 75325
rect 659350 75269 659418 75325
rect 659474 75269 659542 75325
rect 659598 75269 659666 75325
rect 659722 75269 659802 75325
rect 657752 75201 659802 75269
rect 657752 75145 657806 75201
rect 657862 75145 657930 75201
rect 657986 75145 658054 75201
rect 658110 75145 658178 75201
rect 658234 75145 658302 75201
rect 658358 75145 658426 75201
rect 658482 75145 658550 75201
rect 658606 75145 658674 75201
rect 658730 75145 658798 75201
rect 658854 75145 658922 75201
rect 658978 75145 659046 75201
rect 659102 75145 659170 75201
rect 659226 75145 659294 75201
rect 659350 75145 659418 75201
rect 659474 75145 659542 75201
rect 659598 75145 659666 75201
rect 659722 75145 659802 75201
rect 657752 75077 659802 75145
rect 657752 75021 657806 75077
rect 657862 75021 657930 75077
rect 657986 75021 658054 75077
rect 658110 75021 658178 75077
rect 658234 75021 658302 75077
rect 658358 75021 658426 75077
rect 658482 75021 658550 75077
rect 658606 75021 658674 75077
rect 658730 75021 658798 75077
rect 658854 75021 658922 75077
rect 658978 75021 659046 75077
rect 659102 75021 659170 75077
rect 659226 75021 659294 75077
rect 659350 75021 659418 75077
rect 659474 75021 659542 75077
rect 659598 75021 659666 75077
rect 659722 75021 659802 75077
rect 657752 74953 659802 75021
rect 657752 74897 657806 74953
rect 657862 74897 657930 74953
rect 657986 74897 658054 74953
rect 658110 74897 658178 74953
rect 658234 74897 658302 74953
rect 658358 74897 658426 74953
rect 658482 74897 658550 74953
rect 658606 74897 658674 74953
rect 658730 74897 658798 74953
rect 658854 74897 658922 74953
rect 658978 74897 659046 74953
rect 659102 74897 659170 74953
rect 659226 74897 659294 74953
rect 659350 74897 659418 74953
rect 659474 74897 659542 74953
rect 659598 74897 659666 74953
rect 659722 74897 659802 74953
rect 657752 74829 659802 74897
rect 657752 74773 657806 74829
rect 657862 74773 657930 74829
rect 657986 74773 658054 74829
rect 658110 74773 658178 74829
rect 658234 74773 658302 74829
rect 658358 74773 658426 74829
rect 658482 74773 658550 74829
rect 658606 74773 658674 74829
rect 658730 74773 658798 74829
rect 658854 74773 658922 74829
rect 658978 74773 659046 74829
rect 659102 74773 659170 74829
rect 659226 74773 659294 74829
rect 659350 74773 659418 74829
rect 659474 74773 659542 74829
rect 659598 74773 659666 74829
rect 659722 74773 659802 74829
rect 657752 74705 659802 74773
rect 657752 74649 657806 74705
rect 657862 74649 657930 74705
rect 657986 74649 658054 74705
rect 658110 74649 658178 74705
rect 658234 74649 658302 74705
rect 658358 74649 658426 74705
rect 658482 74649 658550 74705
rect 658606 74649 658674 74705
rect 658730 74649 658798 74705
rect 658854 74649 658922 74705
rect 658978 74649 659046 74705
rect 659102 74649 659170 74705
rect 659226 74649 659294 74705
rect 659350 74649 659418 74705
rect 659474 74649 659542 74705
rect 659598 74649 659666 74705
rect 659722 74649 659802 74705
rect 657752 74581 659802 74649
rect 657752 74525 657806 74581
rect 657862 74525 657930 74581
rect 657986 74525 658054 74581
rect 658110 74525 658178 74581
rect 658234 74525 658302 74581
rect 658358 74525 658426 74581
rect 658482 74525 658550 74581
rect 658606 74525 658674 74581
rect 658730 74525 658798 74581
rect 658854 74525 658922 74581
rect 658978 74525 659046 74581
rect 659102 74525 659170 74581
rect 659226 74525 659294 74581
rect 659350 74525 659418 74581
rect 659474 74525 659542 74581
rect 659598 74525 659666 74581
rect 659722 74525 659802 74581
rect 657752 70000 659802 74525
rect 660122 75945 662172 76088
rect 660122 75889 660176 75945
rect 660232 75889 660300 75945
rect 660356 75889 660424 75945
rect 660480 75889 660548 75945
rect 660604 75889 660672 75945
rect 660728 75889 660796 75945
rect 660852 75889 660920 75945
rect 660976 75889 661044 75945
rect 661100 75889 661168 75945
rect 661224 75889 661292 75945
rect 661348 75889 661416 75945
rect 661472 75889 661540 75945
rect 661596 75889 661664 75945
rect 661720 75889 661788 75945
rect 661844 75889 661912 75945
rect 661968 75889 662036 75945
rect 662092 75889 662172 75945
rect 660122 75821 662172 75889
rect 660122 75765 660176 75821
rect 660232 75765 660300 75821
rect 660356 75765 660424 75821
rect 660480 75765 660548 75821
rect 660604 75765 660672 75821
rect 660728 75765 660796 75821
rect 660852 75765 660920 75821
rect 660976 75765 661044 75821
rect 661100 75765 661168 75821
rect 661224 75765 661292 75821
rect 661348 75765 661416 75821
rect 661472 75765 661540 75821
rect 661596 75765 661664 75821
rect 661720 75765 661788 75821
rect 661844 75765 661912 75821
rect 661968 75765 662036 75821
rect 662092 75765 662172 75821
rect 660122 75697 662172 75765
rect 660122 75641 660176 75697
rect 660232 75641 660300 75697
rect 660356 75641 660424 75697
rect 660480 75641 660548 75697
rect 660604 75641 660672 75697
rect 660728 75641 660796 75697
rect 660852 75641 660920 75697
rect 660976 75641 661044 75697
rect 661100 75641 661168 75697
rect 661224 75641 661292 75697
rect 661348 75641 661416 75697
rect 661472 75641 661540 75697
rect 661596 75641 661664 75697
rect 661720 75641 661788 75697
rect 661844 75641 661912 75697
rect 661968 75641 662036 75697
rect 662092 75641 662172 75697
rect 660122 75573 662172 75641
rect 660122 75517 660176 75573
rect 660232 75517 660300 75573
rect 660356 75517 660424 75573
rect 660480 75517 660548 75573
rect 660604 75517 660672 75573
rect 660728 75517 660796 75573
rect 660852 75517 660920 75573
rect 660976 75517 661044 75573
rect 661100 75517 661168 75573
rect 661224 75517 661292 75573
rect 661348 75517 661416 75573
rect 661472 75517 661540 75573
rect 661596 75517 661664 75573
rect 661720 75517 661788 75573
rect 661844 75517 661912 75573
rect 661968 75517 662036 75573
rect 662092 75517 662172 75573
rect 660122 75449 662172 75517
rect 660122 75393 660176 75449
rect 660232 75393 660300 75449
rect 660356 75393 660424 75449
rect 660480 75393 660548 75449
rect 660604 75393 660672 75449
rect 660728 75393 660796 75449
rect 660852 75393 660920 75449
rect 660976 75393 661044 75449
rect 661100 75393 661168 75449
rect 661224 75393 661292 75449
rect 661348 75393 661416 75449
rect 661472 75393 661540 75449
rect 661596 75393 661664 75449
rect 661720 75393 661788 75449
rect 661844 75393 661912 75449
rect 661968 75393 662036 75449
rect 662092 75393 662172 75449
rect 660122 75325 662172 75393
rect 660122 75269 660176 75325
rect 660232 75269 660300 75325
rect 660356 75269 660424 75325
rect 660480 75269 660548 75325
rect 660604 75269 660672 75325
rect 660728 75269 660796 75325
rect 660852 75269 660920 75325
rect 660976 75269 661044 75325
rect 661100 75269 661168 75325
rect 661224 75269 661292 75325
rect 661348 75269 661416 75325
rect 661472 75269 661540 75325
rect 661596 75269 661664 75325
rect 661720 75269 661788 75325
rect 661844 75269 661912 75325
rect 661968 75269 662036 75325
rect 662092 75269 662172 75325
rect 660122 75201 662172 75269
rect 660122 75145 660176 75201
rect 660232 75145 660300 75201
rect 660356 75145 660424 75201
rect 660480 75145 660548 75201
rect 660604 75145 660672 75201
rect 660728 75145 660796 75201
rect 660852 75145 660920 75201
rect 660976 75145 661044 75201
rect 661100 75145 661168 75201
rect 661224 75145 661292 75201
rect 661348 75145 661416 75201
rect 661472 75145 661540 75201
rect 661596 75145 661664 75201
rect 661720 75145 661788 75201
rect 661844 75145 661912 75201
rect 661968 75145 662036 75201
rect 662092 75145 662172 75201
rect 660122 75077 662172 75145
rect 660122 75021 660176 75077
rect 660232 75021 660300 75077
rect 660356 75021 660424 75077
rect 660480 75021 660548 75077
rect 660604 75021 660672 75077
rect 660728 75021 660796 75077
rect 660852 75021 660920 75077
rect 660976 75021 661044 75077
rect 661100 75021 661168 75077
rect 661224 75021 661292 75077
rect 661348 75021 661416 75077
rect 661472 75021 661540 75077
rect 661596 75021 661664 75077
rect 661720 75021 661788 75077
rect 661844 75021 661912 75077
rect 661968 75021 662036 75077
rect 662092 75021 662172 75077
rect 660122 74953 662172 75021
rect 660122 74897 660176 74953
rect 660232 74897 660300 74953
rect 660356 74897 660424 74953
rect 660480 74897 660548 74953
rect 660604 74897 660672 74953
rect 660728 74897 660796 74953
rect 660852 74897 660920 74953
rect 660976 74897 661044 74953
rect 661100 74897 661168 74953
rect 661224 74897 661292 74953
rect 661348 74897 661416 74953
rect 661472 74897 661540 74953
rect 661596 74897 661664 74953
rect 661720 74897 661788 74953
rect 661844 74897 661912 74953
rect 661968 74897 662036 74953
rect 662092 74897 662172 74953
rect 660122 74829 662172 74897
rect 660122 74773 660176 74829
rect 660232 74773 660300 74829
rect 660356 74773 660424 74829
rect 660480 74773 660548 74829
rect 660604 74773 660672 74829
rect 660728 74773 660796 74829
rect 660852 74773 660920 74829
rect 660976 74773 661044 74829
rect 661100 74773 661168 74829
rect 661224 74773 661292 74829
rect 661348 74773 661416 74829
rect 661472 74773 661540 74829
rect 661596 74773 661664 74829
rect 661720 74773 661788 74829
rect 661844 74773 661912 74829
rect 661968 74773 662036 74829
rect 662092 74773 662172 74829
rect 660122 74705 662172 74773
rect 660122 74649 660176 74705
rect 660232 74649 660300 74705
rect 660356 74649 660424 74705
rect 660480 74649 660548 74705
rect 660604 74649 660672 74705
rect 660728 74649 660796 74705
rect 660852 74649 660920 74705
rect 660976 74649 661044 74705
rect 661100 74649 661168 74705
rect 661224 74649 661292 74705
rect 661348 74649 661416 74705
rect 661472 74649 661540 74705
rect 661596 74649 661664 74705
rect 661720 74649 661788 74705
rect 661844 74649 661912 74705
rect 661968 74649 662036 74705
rect 662092 74649 662172 74705
rect 660122 74581 662172 74649
rect 660122 74525 660176 74581
rect 660232 74525 660300 74581
rect 660356 74525 660424 74581
rect 660480 74525 660548 74581
rect 660604 74525 660672 74581
rect 660728 74525 660796 74581
rect 660852 74525 660920 74581
rect 660976 74525 661044 74581
rect 661100 74525 661168 74581
rect 661224 74525 661292 74581
rect 661348 74525 661416 74581
rect 661472 74525 661540 74581
rect 661596 74525 661664 74581
rect 661720 74525 661788 74581
rect 661844 74525 661912 74581
rect 661968 74525 662036 74581
rect 662092 74525 662172 74581
rect 660122 70000 662172 74525
rect 662828 75945 664878 76088
rect 662828 75889 662882 75945
rect 662938 75889 663006 75945
rect 663062 75889 663130 75945
rect 663186 75889 663254 75945
rect 663310 75889 663378 75945
rect 663434 75889 663502 75945
rect 663558 75889 663626 75945
rect 663682 75889 663750 75945
rect 663806 75889 663874 75945
rect 663930 75889 663998 75945
rect 664054 75889 664122 75945
rect 664178 75889 664246 75945
rect 664302 75889 664370 75945
rect 664426 75889 664494 75945
rect 664550 75889 664618 75945
rect 664674 75889 664742 75945
rect 664798 75889 664878 75945
rect 662828 75821 664878 75889
rect 662828 75765 662882 75821
rect 662938 75765 663006 75821
rect 663062 75765 663130 75821
rect 663186 75765 663254 75821
rect 663310 75765 663378 75821
rect 663434 75765 663502 75821
rect 663558 75765 663626 75821
rect 663682 75765 663750 75821
rect 663806 75765 663874 75821
rect 663930 75765 663998 75821
rect 664054 75765 664122 75821
rect 664178 75765 664246 75821
rect 664302 75765 664370 75821
rect 664426 75765 664494 75821
rect 664550 75765 664618 75821
rect 664674 75765 664742 75821
rect 664798 75765 664878 75821
rect 662828 75697 664878 75765
rect 662828 75641 662882 75697
rect 662938 75641 663006 75697
rect 663062 75641 663130 75697
rect 663186 75641 663254 75697
rect 663310 75641 663378 75697
rect 663434 75641 663502 75697
rect 663558 75641 663626 75697
rect 663682 75641 663750 75697
rect 663806 75641 663874 75697
rect 663930 75641 663998 75697
rect 664054 75641 664122 75697
rect 664178 75641 664246 75697
rect 664302 75641 664370 75697
rect 664426 75641 664494 75697
rect 664550 75641 664618 75697
rect 664674 75641 664742 75697
rect 664798 75641 664878 75697
rect 662828 75573 664878 75641
rect 662828 75517 662882 75573
rect 662938 75517 663006 75573
rect 663062 75517 663130 75573
rect 663186 75517 663254 75573
rect 663310 75517 663378 75573
rect 663434 75517 663502 75573
rect 663558 75517 663626 75573
rect 663682 75517 663750 75573
rect 663806 75517 663874 75573
rect 663930 75517 663998 75573
rect 664054 75517 664122 75573
rect 664178 75517 664246 75573
rect 664302 75517 664370 75573
rect 664426 75517 664494 75573
rect 664550 75517 664618 75573
rect 664674 75517 664742 75573
rect 664798 75517 664878 75573
rect 662828 75449 664878 75517
rect 662828 75393 662882 75449
rect 662938 75393 663006 75449
rect 663062 75393 663130 75449
rect 663186 75393 663254 75449
rect 663310 75393 663378 75449
rect 663434 75393 663502 75449
rect 663558 75393 663626 75449
rect 663682 75393 663750 75449
rect 663806 75393 663874 75449
rect 663930 75393 663998 75449
rect 664054 75393 664122 75449
rect 664178 75393 664246 75449
rect 664302 75393 664370 75449
rect 664426 75393 664494 75449
rect 664550 75393 664618 75449
rect 664674 75393 664742 75449
rect 664798 75393 664878 75449
rect 662828 75325 664878 75393
rect 662828 75269 662882 75325
rect 662938 75269 663006 75325
rect 663062 75269 663130 75325
rect 663186 75269 663254 75325
rect 663310 75269 663378 75325
rect 663434 75269 663502 75325
rect 663558 75269 663626 75325
rect 663682 75269 663750 75325
rect 663806 75269 663874 75325
rect 663930 75269 663998 75325
rect 664054 75269 664122 75325
rect 664178 75269 664246 75325
rect 664302 75269 664370 75325
rect 664426 75269 664494 75325
rect 664550 75269 664618 75325
rect 664674 75269 664742 75325
rect 664798 75269 664878 75325
rect 662828 75201 664878 75269
rect 662828 75145 662882 75201
rect 662938 75145 663006 75201
rect 663062 75145 663130 75201
rect 663186 75145 663254 75201
rect 663310 75145 663378 75201
rect 663434 75145 663502 75201
rect 663558 75145 663626 75201
rect 663682 75145 663750 75201
rect 663806 75145 663874 75201
rect 663930 75145 663998 75201
rect 664054 75145 664122 75201
rect 664178 75145 664246 75201
rect 664302 75145 664370 75201
rect 664426 75145 664494 75201
rect 664550 75145 664618 75201
rect 664674 75145 664742 75201
rect 664798 75145 664878 75201
rect 662828 75077 664878 75145
rect 662828 75021 662882 75077
rect 662938 75021 663006 75077
rect 663062 75021 663130 75077
rect 663186 75021 663254 75077
rect 663310 75021 663378 75077
rect 663434 75021 663502 75077
rect 663558 75021 663626 75077
rect 663682 75021 663750 75077
rect 663806 75021 663874 75077
rect 663930 75021 663998 75077
rect 664054 75021 664122 75077
rect 664178 75021 664246 75077
rect 664302 75021 664370 75077
rect 664426 75021 664494 75077
rect 664550 75021 664618 75077
rect 664674 75021 664742 75077
rect 664798 75021 664878 75077
rect 662828 74953 664878 75021
rect 662828 74897 662882 74953
rect 662938 74897 663006 74953
rect 663062 74897 663130 74953
rect 663186 74897 663254 74953
rect 663310 74897 663378 74953
rect 663434 74897 663502 74953
rect 663558 74897 663626 74953
rect 663682 74897 663750 74953
rect 663806 74897 663874 74953
rect 663930 74897 663998 74953
rect 664054 74897 664122 74953
rect 664178 74897 664246 74953
rect 664302 74897 664370 74953
rect 664426 74897 664494 74953
rect 664550 74897 664618 74953
rect 664674 74897 664742 74953
rect 664798 74897 664878 74953
rect 662828 74829 664878 74897
rect 662828 74773 662882 74829
rect 662938 74773 663006 74829
rect 663062 74773 663130 74829
rect 663186 74773 663254 74829
rect 663310 74773 663378 74829
rect 663434 74773 663502 74829
rect 663558 74773 663626 74829
rect 663682 74773 663750 74829
rect 663806 74773 663874 74829
rect 663930 74773 663998 74829
rect 664054 74773 664122 74829
rect 664178 74773 664246 74829
rect 664302 74773 664370 74829
rect 664426 74773 664494 74829
rect 664550 74773 664618 74829
rect 664674 74773 664742 74829
rect 664798 74773 664878 74829
rect 662828 74705 664878 74773
rect 662828 74649 662882 74705
rect 662938 74649 663006 74705
rect 663062 74649 663130 74705
rect 663186 74649 663254 74705
rect 663310 74649 663378 74705
rect 663434 74649 663502 74705
rect 663558 74649 663626 74705
rect 663682 74649 663750 74705
rect 663806 74649 663874 74705
rect 663930 74649 663998 74705
rect 664054 74649 664122 74705
rect 664178 74649 664246 74705
rect 664302 74649 664370 74705
rect 664426 74649 664494 74705
rect 664550 74649 664618 74705
rect 664674 74649 664742 74705
rect 664798 74649 664878 74705
rect 662828 74581 664878 74649
rect 662828 74525 662882 74581
rect 662938 74525 663006 74581
rect 663062 74525 663130 74581
rect 663186 74525 663254 74581
rect 663310 74525 663378 74581
rect 663434 74525 663502 74581
rect 663558 74525 663626 74581
rect 663682 74525 663750 74581
rect 663806 74525 663874 74581
rect 663930 74525 663998 74581
rect 664054 74525 664122 74581
rect 664178 74525 664246 74581
rect 664302 74525 664370 74581
rect 664426 74525 664494 74581
rect 664550 74525 664618 74581
rect 664674 74525 664742 74581
rect 664798 74525 664878 74581
rect 662828 70000 664878 74525
rect 665198 75945 667248 76088
rect 665198 75889 665252 75945
rect 665308 75889 665376 75945
rect 665432 75889 665500 75945
rect 665556 75889 665624 75945
rect 665680 75889 665748 75945
rect 665804 75889 665872 75945
rect 665928 75889 665996 75945
rect 666052 75889 666120 75945
rect 666176 75889 666244 75945
rect 666300 75889 666368 75945
rect 666424 75889 666492 75945
rect 666548 75889 666616 75945
rect 666672 75889 666740 75945
rect 666796 75889 666864 75945
rect 666920 75889 666988 75945
rect 667044 75889 667112 75945
rect 667168 75889 667248 75945
rect 665198 75821 667248 75889
rect 665198 75765 665252 75821
rect 665308 75765 665376 75821
rect 665432 75765 665500 75821
rect 665556 75765 665624 75821
rect 665680 75765 665748 75821
rect 665804 75765 665872 75821
rect 665928 75765 665996 75821
rect 666052 75765 666120 75821
rect 666176 75765 666244 75821
rect 666300 75765 666368 75821
rect 666424 75765 666492 75821
rect 666548 75765 666616 75821
rect 666672 75765 666740 75821
rect 666796 75765 666864 75821
rect 666920 75765 666988 75821
rect 667044 75765 667112 75821
rect 667168 75765 667248 75821
rect 665198 75697 667248 75765
rect 665198 75641 665252 75697
rect 665308 75641 665376 75697
rect 665432 75641 665500 75697
rect 665556 75641 665624 75697
rect 665680 75641 665748 75697
rect 665804 75641 665872 75697
rect 665928 75641 665996 75697
rect 666052 75641 666120 75697
rect 666176 75641 666244 75697
rect 666300 75641 666368 75697
rect 666424 75641 666492 75697
rect 666548 75641 666616 75697
rect 666672 75641 666740 75697
rect 666796 75641 666864 75697
rect 666920 75641 666988 75697
rect 667044 75641 667112 75697
rect 667168 75641 667248 75697
rect 665198 75573 667248 75641
rect 665198 75517 665252 75573
rect 665308 75517 665376 75573
rect 665432 75517 665500 75573
rect 665556 75517 665624 75573
rect 665680 75517 665748 75573
rect 665804 75517 665872 75573
rect 665928 75517 665996 75573
rect 666052 75517 666120 75573
rect 666176 75517 666244 75573
rect 666300 75517 666368 75573
rect 666424 75517 666492 75573
rect 666548 75517 666616 75573
rect 666672 75517 666740 75573
rect 666796 75517 666864 75573
rect 666920 75517 666988 75573
rect 667044 75517 667112 75573
rect 667168 75517 667248 75573
rect 665198 75449 667248 75517
rect 665198 75393 665252 75449
rect 665308 75393 665376 75449
rect 665432 75393 665500 75449
rect 665556 75393 665624 75449
rect 665680 75393 665748 75449
rect 665804 75393 665872 75449
rect 665928 75393 665996 75449
rect 666052 75393 666120 75449
rect 666176 75393 666244 75449
rect 666300 75393 666368 75449
rect 666424 75393 666492 75449
rect 666548 75393 666616 75449
rect 666672 75393 666740 75449
rect 666796 75393 666864 75449
rect 666920 75393 666988 75449
rect 667044 75393 667112 75449
rect 667168 75393 667248 75449
rect 665198 75325 667248 75393
rect 665198 75269 665252 75325
rect 665308 75269 665376 75325
rect 665432 75269 665500 75325
rect 665556 75269 665624 75325
rect 665680 75269 665748 75325
rect 665804 75269 665872 75325
rect 665928 75269 665996 75325
rect 666052 75269 666120 75325
rect 666176 75269 666244 75325
rect 666300 75269 666368 75325
rect 666424 75269 666492 75325
rect 666548 75269 666616 75325
rect 666672 75269 666740 75325
rect 666796 75269 666864 75325
rect 666920 75269 666988 75325
rect 667044 75269 667112 75325
rect 667168 75269 667248 75325
rect 665198 75201 667248 75269
rect 665198 75145 665252 75201
rect 665308 75145 665376 75201
rect 665432 75145 665500 75201
rect 665556 75145 665624 75201
rect 665680 75145 665748 75201
rect 665804 75145 665872 75201
rect 665928 75145 665996 75201
rect 666052 75145 666120 75201
rect 666176 75145 666244 75201
rect 666300 75145 666368 75201
rect 666424 75145 666492 75201
rect 666548 75145 666616 75201
rect 666672 75145 666740 75201
rect 666796 75145 666864 75201
rect 666920 75145 666988 75201
rect 667044 75145 667112 75201
rect 667168 75145 667248 75201
rect 665198 75077 667248 75145
rect 665198 75021 665252 75077
rect 665308 75021 665376 75077
rect 665432 75021 665500 75077
rect 665556 75021 665624 75077
rect 665680 75021 665748 75077
rect 665804 75021 665872 75077
rect 665928 75021 665996 75077
rect 666052 75021 666120 75077
rect 666176 75021 666244 75077
rect 666300 75021 666368 75077
rect 666424 75021 666492 75077
rect 666548 75021 666616 75077
rect 666672 75021 666740 75077
rect 666796 75021 666864 75077
rect 666920 75021 666988 75077
rect 667044 75021 667112 75077
rect 667168 75021 667248 75077
rect 665198 74953 667248 75021
rect 665198 74897 665252 74953
rect 665308 74897 665376 74953
rect 665432 74897 665500 74953
rect 665556 74897 665624 74953
rect 665680 74897 665748 74953
rect 665804 74897 665872 74953
rect 665928 74897 665996 74953
rect 666052 74897 666120 74953
rect 666176 74897 666244 74953
rect 666300 74897 666368 74953
rect 666424 74897 666492 74953
rect 666548 74897 666616 74953
rect 666672 74897 666740 74953
rect 666796 74897 666864 74953
rect 666920 74897 666988 74953
rect 667044 74897 667112 74953
rect 667168 74897 667248 74953
rect 665198 74829 667248 74897
rect 665198 74773 665252 74829
rect 665308 74773 665376 74829
rect 665432 74773 665500 74829
rect 665556 74773 665624 74829
rect 665680 74773 665748 74829
rect 665804 74773 665872 74829
rect 665928 74773 665996 74829
rect 666052 74773 666120 74829
rect 666176 74773 666244 74829
rect 666300 74773 666368 74829
rect 666424 74773 666492 74829
rect 666548 74773 666616 74829
rect 666672 74773 666740 74829
rect 666796 74773 666864 74829
rect 666920 74773 666988 74829
rect 667044 74773 667112 74829
rect 667168 74773 667248 74829
rect 665198 74705 667248 74773
rect 665198 74649 665252 74705
rect 665308 74649 665376 74705
rect 665432 74649 665500 74705
rect 665556 74649 665624 74705
rect 665680 74649 665748 74705
rect 665804 74649 665872 74705
rect 665928 74649 665996 74705
rect 666052 74649 666120 74705
rect 666176 74649 666244 74705
rect 666300 74649 666368 74705
rect 666424 74649 666492 74705
rect 666548 74649 666616 74705
rect 666672 74649 666740 74705
rect 666796 74649 666864 74705
rect 666920 74649 666988 74705
rect 667044 74649 667112 74705
rect 667168 74649 667248 74705
rect 665198 74581 667248 74649
rect 665198 74525 665252 74581
rect 665308 74525 665376 74581
rect 665432 74525 665500 74581
rect 665556 74525 665624 74581
rect 665680 74525 665748 74581
rect 665804 74525 665872 74581
rect 665928 74525 665996 74581
rect 666052 74525 666120 74581
rect 666176 74525 666244 74581
rect 666300 74525 666368 74581
rect 666424 74525 666492 74581
rect 666548 74525 666616 74581
rect 666672 74525 666740 74581
rect 666796 74525 666864 74581
rect 666920 74525 666988 74581
rect 667044 74525 667112 74581
rect 667168 74525 667248 74581
rect 665198 70000 667248 74525
rect 667828 75945 669728 76088
rect 667828 75889 667882 75945
rect 667938 75889 668006 75945
rect 668062 75889 668130 75945
rect 668186 75889 668254 75945
rect 668310 75889 668378 75945
rect 668434 75889 668502 75945
rect 668558 75889 668626 75945
rect 668682 75889 668750 75945
rect 668806 75889 668874 75945
rect 668930 75889 668998 75945
rect 669054 75889 669122 75945
rect 669178 75889 669246 75945
rect 669302 75889 669370 75945
rect 669426 75889 669494 75945
rect 669550 75889 669618 75945
rect 669674 75889 669728 75945
rect 667828 75821 669728 75889
rect 667828 75765 667882 75821
rect 667938 75765 668006 75821
rect 668062 75765 668130 75821
rect 668186 75765 668254 75821
rect 668310 75765 668378 75821
rect 668434 75765 668502 75821
rect 668558 75765 668626 75821
rect 668682 75765 668750 75821
rect 668806 75765 668874 75821
rect 668930 75765 668998 75821
rect 669054 75765 669122 75821
rect 669178 75765 669246 75821
rect 669302 75765 669370 75821
rect 669426 75765 669494 75821
rect 669550 75765 669618 75821
rect 669674 75765 669728 75821
rect 667828 75697 669728 75765
rect 667828 75641 667882 75697
rect 667938 75641 668006 75697
rect 668062 75641 668130 75697
rect 668186 75641 668254 75697
rect 668310 75641 668378 75697
rect 668434 75641 668502 75697
rect 668558 75641 668626 75697
rect 668682 75641 668750 75697
rect 668806 75641 668874 75697
rect 668930 75641 668998 75697
rect 669054 75641 669122 75697
rect 669178 75641 669246 75697
rect 669302 75641 669370 75697
rect 669426 75641 669494 75697
rect 669550 75641 669618 75697
rect 669674 75641 669728 75697
rect 667828 75573 669728 75641
rect 667828 75517 667882 75573
rect 667938 75517 668006 75573
rect 668062 75517 668130 75573
rect 668186 75517 668254 75573
rect 668310 75517 668378 75573
rect 668434 75517 668502 75573
rect 668558 75517 668626 75573
rect 668682 75517 668750 75573
rect 668806 75517 668874 75573
rect 668930 75517 668998 75573
rect 669054 75517 669122 75573
rect 669178 75517 669246 75573
rect 669302 75517 669370 75573
rect 669426 75517 669494 75573
rect 669550 75517 669618 75573
rect 669674 75517 669728 75573
rect 667828 75449 669728 75517
rect 667828 75393 667882 75449
rect 667938 75393 668006 75449
rect 668062 75393 668130 75449
rect 668186 75393 668254 75449
rect 668310 75393 668378 75449
rect 668434 75393 668502 75449
rect 668558 75393 668626 75449
rect 668682 75393 668750 75449
rect 668806 75393 668874 75449
rect 668930 75393 668998 75449
rect 669054 75393 669122 75449
rect 669178 75393 669246 75449
rect 669302 75393 669370 75449
rect 669426 75393 669494 75449
rect 669550 75393 669618 75449
rect 669674 75393 669728 75449
rect 667828 75325 669728 75393
rect 667828 75269 667882 75325
rect 667938 75269 668006 75325
rect 668062 75269 668130 75325
rect 668186 75269 668254 75325
rect 668310 75269 668378 75325
rect 668434 75269 668502 75325
rect 668558 75269 668626 75325
rect 668682 75269 668750 75325
rect 668806 75269 668874 75325
rect 668930 75269 668998 75325
rect 669054 75269 669122 75325
rect 669178 75269 669246 75325
rect 669302 75269 669370 75325
rect 669426 75269 669494 75325
rect 669550 75269 669618 75325
rect 669674 75269 669728 75325
rect 667828 75201 669728 75269
rect 667828 75145 667882 75201
rect 667938 75145 668006 75201
rect 668062 75145 668130 75201
rect 668186 75145 668254 75201
rect 668310 75145 668378 75201
rect 668434 75145 668502 75201
rect 668558 75145 668626 75201
rect 668682 75145 668750 75201
rect 668806 75145 668874 75201
rect 668930 75145 668998 75201
rect 669054 75145 669122 75201
rect 669178 75145 669246 75201
rect 669302 75145 669370 75201
rect 669426 75145 669494 75201
rect 669550 75145 669618 75201
rect 669674 75145 669728 75201
rect 667828 75077 669728 75145
rect 667828 75021 667882 75077
rect 667938 75021 668006 75077
rect 668062 75021 668130 75077
rect 668186 75021 668254 75077
rect 668310 75021 668378 75077
rect 668434 75021 668502 75077
rect 668558 75021 668626 75077
rect 668682 75021 668750 75077
rect 668806 75021 668874 75077
rect 668930 75021 668998 75077
rect 669054 75021 669122 75077
rect 669178 75021 669246 75077
rect 669302 75021 669370 75077
rect 669426 75021 669494 75077
rect 669550 75021 669618 75077
rect 669674 75021 669728 75077
rect 667828 74953 669728 75021
rect 667828 74897 667882 74953
rect 667938 74897 668006 74953
rect 668062 74897 668130 74953
rect 668186 74897 668254 74953
rect 668310 74897 668378 74953
rect 668434 74897 668502 74953
rect 668558 74897 668626 74953
rect 668682 74897 668750 74953
rect 668806 74897 668874 74953
rect 668930 74897 668998 74953
rect 669054 74897 669122 74953
rect 669178 74897 669246 74953
rect 669302 74897 669370 74953
rect 669426 74897 669494 74953
rect 669550 74897 669618 74953
rect 669674 74897 669728 74953
rect 667828 74829 669728 74897
rect 667828 74773 667882 74829
rect 667938 74773 668006 74829
rect 668062 74773 668130 74829
rect 668186 74773 668254 74829
rect 668310 74773 668378 74829
rect 668434 74773 668502 74829
rect 668558 74773 668626 74829
rect 668682 74773 668750 74829
rect 668806 74773 668874 74829
rect 668930 74773 668998 74829
rect 669054 74773 669122 74829
rect 669178 74773 669246 74829
rect 669302 74773 669370 74829
rect 669426 74773 669494 74829
rect 669550 74773 669618 74829
rect 669674 74773 669728 74829
rect 667828 74705 669728 74773
rect 667828 74649 667882 74705
rect 667938 74649 668006 74705
rect 668062 74649 668130 74705
rect 668186 74649 668254 74705
rect 668310 74649 668378 74705
rect 668434 74649 668502 74705
rect 668558 74649 668626 74705
rect 668682 74649 668750 74705
rect 668806 74649 668874 74705
rect 668930 74649 668998 74705
rect 669054 74649 669122 74705
rect 669178 74649 669246 74705
rect 669302 74649 669370 74705
rect 669426 74649 669494 74705
rect 669550 74649 669618 74705
rect 669674 74649 669728 74705
rect 667828 74581 669728 74649
rect 667828 74525 667882 74581
rect 667938 74525 668006 74581
rect 668062 74525 668130 74581
rect 668186 74525 668254 74581
rect 668310 74525 668378 74581
rect 668434 74525 668502 74581
rect 668558 74525 668626 74581
rect 668682 74525 668750 74581
rect 668806 74525 668874 74581
rect 668930 74525 668998 74581
rect 669054 74525 669122 74581
rect 669178 74525 669246 74581
rect 669302 74525 669370 74581
rect 669426 74525 669494 74581
rect 669550 74525 669618 74581
rect 669674 74525 669728 74581
rect 667828 70000 669728 74525
<< via2 >>
rect 379326 941599 379382 941655
rect 379450 941599 379506 941655
rect 379574 941599 379630 941655
rect 379698 941599 379754 941655
rect 379822 941599 379878 941655
rect 379946 941599 380002 941655
rect 379326 941475 379382 941531
rect 379450 941475 379506 941531
rect 379574 941475 379630 941531
rect 379698 941475 379754 941531
rect 379822 941475 379878 941531
rect 379946 941475 380002 941531
rect 379326 941351 379382 941407
rect 379450 941351 379506 941407
rect 379574 941351 379630 941407
rect 379698 941351 379754 941407
rect 379822 941351 379878 941407
rect 379946 941351 380002 941407
rect 379326 941227 379382 941283
rect 379450 941227 379506 941283
rect 379574 941227 379630 941283
rect 379698 941227 379754 941283
rect 379822 941227 379878 941283
rect 379946 941227 380002 941283
rect 379326 941103 379382 941159
rect 379450 941103 379506 941159
rect 379574 941103 379630 941159
rect 379698 941103 379754 941159
rect 379822 941103 379878 941159
rect 379946 941103 380002 941159
rect 379326 940979 379382 941035
rect 379450 940979 379506 941035
rect 379574 940979 379630 941035
rect 379698 940979 379754 941035
rect 379822 940979 379878 941035
rect 379946 940979 380002 941035
rect 379326 940855 379382 940911
rect 379450 940855 379506 940911
rect 379574 940855 379630 940911
rect 379698 940855 379754 940911
rect 379822 940855 379878 940911
rect 379946 940855 380002 940911
rect 379326 940731 379382 940787
rect 379450 940731 379506 940787
rect 379574 940731 379630 940787
rect 379698 940731 379754 940787
rect 379822 940731 379878 940787
rect 379946 940731 380002 940787
rect 379326 940607 379382 940663
rect 379450 940607 379506 940663
rect 379574 940607 379630 940663
rect 379698 940607 379754 940663
rect 379822 940607 379878 940663
rect 379946 940607 380002 940663
rect 379326 940483 379382 940539
rect 379450 940483 379506 940539
rect 379574 940483 379630 940539
rect 379698 940483 379754 940539
rect 379822 940483 379878 940539
rect 379946 940483 380002 940539
rect 379326 940359 379382 940415
rect 379450 940359 379506 940415
rect 379574 940359 379630 940415
rect 379698 940359 379754 940415
rect 379822 940359 379878 940415
rect 379946 940359 380002 940415
rect 379326 940235 379382 940291
rect 379450 940235 379506 940291
rect 379574 940235 379630 940291
rect 379698 940235 379754 940291
rect 379822 940235 379878 940291
rect 379946 940235 380002 940291
rect 379326 940111 379382 940167
rect 379450 940111 379506 940167
rect 379574 940111 379630 940167
rect 379698 940111 379754 940167
rect 379822 940111 379878 940167
rect 379946 940111 380002 940167
rect 379326 939987 379382 940043
rect 379450 939987 379506 940043
rect 379574 939987 379630 940043
rect 379698 939987 379754 940043
rect 379822 939987 379878 940043
rect 379946 939987 380002 940043
rect 379326 939863 379382 939919
rect 379450 939863 379506 939919
rect 379574 939863 379630 939919
rect 379698 939863 379754 939919
rect 379822 939863 379878 939919
rect 379946 939863 380002 939919
rect 381832 941599 381888 941655
rect 381956 941599 382012 941655
rect 382080 941599 382136 941655
rect 382204 941599 382260 941655
rect 382328 941599 382384 941655
rect 382452 941599 382508 941655
rect 382576 941599 382632 941655
rect 382700 941599 382756 941655
rect 382824 941599 382880 941655
rect 382948 941599 383004 941655
rect 383072 941599 383128 941655
rect 383196 941599 383252 941655
rect 383320 941599 383376 941655
rect 383444 941599 383500 941655
rect 383568 941599 383624 941655
rect 383692 941599 383748 941655
rect 381832 941475 381888 941531
rect 381956 941475 382012 941531
rect 382080 941475 382136 941531
rect 382204 941475 382260 941531
rect 382328 941475 382384 941531
rect 382452 941475 382508 941531
rect 382576 941475 382632 941531
rect 382700 941475 382756 941531
rect 382824 941475 382880 941531
rect 382948 941475 383004 941531
rect 383072 941475 383128 941531
rect 383196 941475 383252 941531
rect 383320 941475 383376 941531
rect 383444 941475 383500 941531
rect 383568 941475 383624 941531
rect 383692 941475 383748 941531
rect 381832 941351 381888 941407
rect 381956 941351 382012 941407
rect 382080 941351 382136 941407
rect 382204 941351 382260 941407
rect 382328 941351 382384 941407
rect 382452 941351 382508 941407
rect 382576 941351 382632 941407
rect 382700 941351 382756 941407
rect 382824 941351 382880 941407
rect 382948 941351 383004 941407
rect 383072 941351 383128 941407
rect 383196 941351 383252 941407
rect 383320 941351 383376 941407
rect 383444 941351 383500 941407
rect 383568 941351 383624 941407
rect 383692 941351 383748 941407
rect 381832 941227 381888 941283
rect 381956 941227 382012 941283
rect 382080 941227 382136 941283
rect 382204 941227 382260 941283
rect 382328 941227 382384 941283
rect 382452 941227 382508 941283
rect 382576 941227 382632 941283
rect 382700 941227 382756 941283
rect 382824 941227 382880 941283
rect 382948 941227 383004 941283
rect 383072 941227 383128 941283
rect 383196 941227 383252 941283
rect 383320 941227 383376 941283
rect 383444 941227 383500 941283
rect 383568 941227 383624 941283
rect 383692 941227 383748 941283
rect 381832 941103 381888 941159
rect 381956 941103 382012 941159
rect 382080 941103 382136 941159
rect 382204 941103 382260 941159
rect 382328 941103 382384 941159
rect 382452 941103 382508 941159
rect 382576 941103 382632 941159
rect 382700 941103 382756 941159
rect 382824 941103 382880 941159
rect 382948 941103 383004 941159
rect 383072 941103 383128 941159
rect 383196 941103 383252 941159
rect 383320 941103 383376 941159
rect 383444 941103 383500 941159
rect 383568 941103 383624 941159
rect 383692 941103 383748 941159
rect 381832 940979 381888 941035
rect 381956 940979 382012 941035
rect 382080 940979 382136 941035
rect 382204 940979 382260 941035
rect 382328 940979 382384 941035
rect 382452 940979 382508 941035
rect 382576 940979 382632 941035
rect 382700 940979 382756 941035
rect 382824 940979 382880 941035
rect 382948 940979 383004 941035
rect 383072 940979 383128 941035
rect 383196 940979 383252 941035
rect 383320 940979 383376 941035
rect 383444 940979 383500 941035
rect 383568 940979 383624 941035
rect 383692 940979 383748 941035
rect 381832 940855 381888 940911
rect 381956 940855 382012 940911
rect 382080 940855 382136 940911
rect 382204 940855 382260 940911
rect 382328 940855 382384 940911
rect 382452 940855 382508 940911
rect 382576 940855 382632 940911
rect 382700 940855 382756 940911
rect 382824 940855 382880 940911
rect 382948 940855 383004 940911
rect 383072 940855 383128 940911
rect 383196 940855 383252 940911
rect 383320 940855 383376 940911
rect 383444 940855 383500 940911
rect 383568 940855 383624 940911
rect 383692 940855 383748 940911
rect 381832 940731 381888 940787
rect 381956 940731 382012 940787
rect 382080 940731 382136 940787
rect 382204 940731 382260 940787
rect 382328 940731 382384 940787
rect 382452 940731 382508 940787
rect 382576 940731 382632 940787
rect 382700 940731 382756 940787
rect 382824 940731 382880 940787
rect 382948 940731 383004 940787
rect 383072 940731 383128 940787
rect 383196 940731 383252 940787
rect 383320 940731 383376 940787
rect 383444 940731 383500 940787
rect 383568 940731 383624 940787
rect 383692 940731 383748 940787
rect 381832 940607 381888 940663
rect 381956 940607 382012 940663
rect 382080 940607 382136 940663
rect 382204 940607 382260 940663
rect 382328 940607 382384 940663
rect 382452 940607 382508 940663
rect 382576 940607 382632 940663
rect 382700 940607 382756 940663
rect 382824 940607 382880 940663
rect 382948 940607 383004 940663
rect 383072 940607 383128 940663
rect 383196 940607 383252 940663
rect 383320 940607 383376 940663
rect 383444 940607 383500 940663
rect 383568 940607 383624 940663
rect 383692 940607 383748 940663
rect 381832 940483 381888 940539
rect 381956 940483 382012 940539
rect 382080 940483 382136 940539
rect 382204 940483 382260 940539
rect 382328 940483 382384 940539
rect 382452 940483 382508 940539
rect 382576 940483 382632 940539
rect 382700 940483 382756 940539
rect 382824 940483 382880 940539
rect 382948 940483 383004 940539
rect 383072 940483 383128 940539
rect 383196 940483 383252 940539
rect 383320 940483 383376 940539
rect 383444 940483 383500 940539
rect 383568 940483 383624 940539
rect 383692 940483 383748 940539
rect 381832 940359 381888 940415
rect 381956 940359 382012 940415
rect 382080 940359 382136 940415
rect 382204 940359 382260 940415
rect 382328 940359 382384 940415
rect 382452 940359 382508 940415
rect 382576 940359 382632 940415
rect 382700 940359 382756 940415
rect 382824 940359 382880 940415
rect 382948 940359 383004 940415
rect 383072 940359 383128 940415
rect 383196 940359 383252 940415
rect 383320 940359 383376 940415
rect 383444 940359 383500 940415
rect 383568 940359 383624 940415
rect 383692 940359 383748 940415
rect 381832 940235 381888 940291
rect 381956 940235 382012 940291
rect 382080 940235 382136 940291
rect 382204 940235 382260 940291
rect 382328 940235 382384 940291
rect 382452 940235 382508 940291
rect 382576 940235 382632 940291
rect 382700 940235 382756 940291
rect 382824 940235 382880 940291
rect 382948 940235 383004 940291
rect 383072 940235 383128 940291
rect 383196 940235 383252 940291
rect 383320 940235 383376 940291
rect 383444 940235 383500 940291
rect 383568 940235 383624 940291
rect 383692 940235 383748 940291
rect 381832 940111 381888 940167
rect 381956 940111 382012 940167
rect 382080 940111 382136 940167
rect 382204 940111 382260 940167
rect 382328 940111 382384 940167
rect 382452 940111 382508 940167
rect 382576 940111 382632 940167
rect 382700 940111 382756 940167
rect 382824 940111 382880 940167
rect 382948 940111 383004 940167
rect 383072 940111 383128 940167
rect 383196 940111 383252 940167
rect 383320 940111 383376 940167
rect 383444 940111 383500 940167
rect 383568 940111 383624 940167
rect 383692 940111 383748 940167
rect 381832 939987 381888 940043
rect 381956 939987 382012 940043
rect 382080 939987 382136 940043
rect 382204 939987 382260 940043
rect 382328 939987 382384 940043
rect 382452 939987 382508 940043
rect 382576 939987 382632 940043
rect 382700 939987 382756 940043
rect 382824 939987 382880 940043
rect 382948 939987 383004 940043
rect 383072 939987 383128 940043
rect 383196 939987 383252 940043
rect 383320 939987 383376 940043
rect 383444 939987 383500 940043
rect 383568 939987 383624 940043
rect 383692 939987 383748 940043
rect 381832 939863 381888 939919
rect 381956 939863 382012 939919
rect 382080 939863 382136 939919
rect 382204 939863 382260 939919
rect 382328 939863 382384 939919
rect 382452 939863 382508 939919
rect 382576 939863 382632 939919
rect 382700 939863 382756 939919
rect 382824 939863 382880 939919
rect 382948 939863 383004 939919
rect 383072 939863 383128 939919
rect 383196 939863 383252 939919
rect 383320 939863 383376 939919
rect 383444 939863 383500 939919
rect 383568 939863 383624 939919
rect 383692 939863 383748 939919
rect 384202 941599 384258 941655
rect 384326 941599 384382 941655
rect 384450 941599 384506 941655
rect 384574 941599 384630 941655
rect 384698 941599 384754 941655
rect 384822 941599 384878 941655
rect 384946 941599 385002 941655
rect 385070 941599 385126 941655
rect 385194 941599 385250 941655
rect 385318 941599 385374 941655
rect 385442 941599 385498 941655
rect 385566 941599 385622 941655
rect 385690 941599 385746 941655
rect 385814 941599 385870 941655
rect 385938 941599 385994 941655
rect 386062 941599 386118 941655
rect 384202 941475 384258 941531
rect 384326 941475 384382 941531
rect 384450 941475 384506 941531
rect 384574 941475 384630 941531
rect 384698 941475 384754 941531
rect 384822 941475 384878 941531
rect 384946 941475 385002 941531
rect 385070 941475 385126 941531
rect 385194 941475 385250 941531
rect 385318 941475 385374 941531
rect 385442 941475 385498 941531
rect 385566 941475 385622 941531
rect 385690 941475 385746 941531
rect 385814 941475 385870 941531
rect 385938 941475 385994 941531
rect 386062 941475 386118 941531
rect 384202 941351 384258 941407
rect 384326 941351 384382 941407
rect 384450 941351 384506 941407
rect 384574 941351 384630 941407
rect 384698 941351 384754 941407
rect 384822 941351 384878 941407
rect 384946 941351 385002 941407
rect 385070 941351 385126 941407
rect 385194 941351 385250 941407
rect 385318 941351 385374 941407
rect 385442 941351 385498 941407
rect 385566 941351 385622 941407
rect 385690 941351 385746 941407
rect 385814 941351 385870 941407
rect 385938 941351 385994 941407
rect 386062 941351 386118 941407
rect 384202 941227 384258 941283
rect 384326 941227 384382 941283
rect 384450 941227 384506 941283
rect 384574 941227 384630 941283
rect 384698 941227 384754 941283
rect 384822 941227 384878 941283
rect 384946 941227 385002 941283
rect 385070 941227 385126 941283
rect 385194 941227 385250 941283
rect 385318 941227 385374 941283
rect 385442 941227 385498 941283
rect 385566 941227 385622 941283
rect 385690 941227 385746 941283
rect 385814 941227 385870 941283
rect 385938 941227 385994 941283
rect 386062 941227 386118 941283
rect 384202 941103 384258 941159
rect 384326 941103 384382 941159
rect 384450 941103 384506 941159
rect 384574 941103 384630 941159
rect 384698 941103 384754 941159
rect 384822 941103 384878 941159
rect 384946 941103 385002 941159
rect 385070 941103 385126 941159
rect 385194 941103 385250 941159
rect 385318 941103 385374 941159
rect 385442 941103 385498 941159
rect 385566 941103 385622 941159
rect 385690 941103 385746 941159
rect 385814 941103 385870 941159
rect 385938 941103 385994 941159
rect 386062 941103 386118 941159
rect 384202 940979 384258 941035
rect 384326 940979 384382 941035
rect 384450 940979 384506 941035
rect 384574 940979 384630 941035
rect 384698 940979 384754 941035
rect 384822 940979 384878 941035
rect 384946 940979 385002 941035
rect 385070 940979 385126 941035
rect 385194 940979 385250 941035
rect 385318 940979 385374 941035
rect 385442 940979 385498 941035
rect 385566 940979 385622 941035
rect 385690 940979 385746 941035
rect 385814 940979 385870 941035
rect 385938 940979 385994 941035
rect 386062 940979 386118 941035
rect 384202 940855 384258 940911
rect 384326 940855 384382 940911
rect 384450 940855 384506 940911
rect 384574 940855 384630 940911
rect 384698 940855 384754 940911
rect 384822 940855 384878 940911
rect 384946 940855 385002 940911
rect 385070 940855 385126 940911
rect 385194 940855 385250 940911
rect 385318 940855 385374 940911
rect 385442 940855 385498 940911
rect 385566 940855 385622 940911
rect 385690 940855 385746 940911
rect 385814 940855 385870 940911
rect 385938 940855 385994 940911
rect 386062 940855 386118 940911
rect 384202 940731 384258 940787
rect 384326 940731 384382 940787
rect 384450 940731 384506 940787
rect 384574 940731 384630 940787
rect 384698 940731 384754 940787
rect 384822 940731 384878 940787
rect 384946 940731 385002 940787
rect 385070 940731 385126 940787
rect 385194 940731 385250 940787
rect 385318 940731 385374 940787
rect 385442 940731 385498 940787
rect 385566 940731 385622 940787
rect 385690 940731 385746 940787
rect 385814 940731 385870 940787
rect 385938 940731 385994 940787
rect 386062 940731 386118 940787
rect 384202 940607 384258 940663
rect 384326 940607 384382 940663
rect 384450 940607 384506 940663
rect 384574 940607 384630 940663
rect 384698 940607 384754 940663
rect 384822 940607 384878 940663
rect 384946 940607 385002 940663
rect 385070 940607 385126 940663
rect 385194 940607 385250 940663
rect 385318 940607 385374 940663
rect 385442 940607 385498 940663
rect 385566 940607 385622 940663
rect 385690 940607 385746 940663
rect 385814 940607 385870 940663
rect 385938 940607 385994 940663
rect 386062 940607 386118 940663
rect 384202 940483 384258 940539
rect 384326 940483 384382 940539
rect 384450 940483 384506 940539
rect 384574 940483 384630 940539
rect 384698 940483 384754 940539
rect 384822 940483 384878 940539
rect 384946 940483 385002 940539
rect 385070 940483 385126 940539
rect 385194 940483 385250 940539
rect 385318 940483 385374 940539
rect 385442 940483 385498 940539
rect 385566 940483 385622 940539
rect 385690 940483 385746 940539
rect 385814 940483 385870 940539
rect 385938 940483 385994 940539
rect 386062 940483 386118 940539
rect 384202 940359 384258 940415
rect 384326 940359 384382 940415
rect 384450 940359 384506 940415
rect 384574 940359 384630 940415
rect 384698 940359 384754 940415
rect 384822 940359 384878 940415
rect 384946 940359 385002 940415
rect 385070 940359 385126 940415
rect 385194 940359 385250 940415
rect 385318 940359 385374 940415
rect 385442 940359 385498 940415
rect 385566 940359 385622 940415
rect 385690 940359 385746 940415
rect 385814 940359 385870 940415
rect 385938 940359 385994 940415
rect 386062 940359 386118 940415
rect 384202 940235 384258 940291
rect 384326 940235 384382 940291
rect 384450 940235 384506 940291
rect 384574 940235 384630 940291
rect 384698 940235 384754 940291
rect 384822 940235 384878 940291
rect 384946 940235 385002 940291
rect 385070 940235 385126 940291
rect 385194 940235 385250 940291
rect 385318 940235 385374 940291
rect 385442 940235 385498 940291
rect 385566 940235 385622 940291
rect 385690 940235 385746 940291
rect 385814 940235 385870 940291
rect 385938 940235 385994 940291
rect 386062 940235 386118 940291
rect 384202 940111 384258 940167
rect 384326 940111 384382 940167
rect 384450 940111 384506 940167
rect 384574 940111 384630 940167
rect 384698 940111 384754 940167
rect 384822 940111 384878 940167
rect 384946 940111 385002 940167
rect 385070 940111 385126 940167
rect 385194 940111 385250 940167
rect 385318 940111 385374 940167
rect 385442 940111 385498 940167
rect 385566 940111 385622 940167
rect 385690 940111 385746 940167
rect 385814 940111 385870 940167
rect 385938 940111 385994 940167
rect 386062 940111 386118 940167
rect 384202 939987 384258 940043
rect 384326 939987 384382 940043
rect 384450 939987 384506 940043
rect 384574 939987 384630 940043
rect 384698 939987 384754 940043
rect 384822 939987 384878 940043
rect 384946 939987 385002 940043
rect 385070 939987 385126 940043
rect 385194 939987 385250 940043
rect 385318 939987 385374 940043
rect 385442 939987 385498 940043
rect 385566 939987 385622 940043
rect 385690 939987 385746 940043
rect 385814 939987 385870 940043
rect 385938 939987 385994 940043
rect 386062 939987 386118 940043
rect 384202 939863 384258 939919
rect 384326 939863 384382 939919
rect 384450 939863 384506 939919
rect 384574 939863 384630 939919
rect 384698 939863 384754 939919
rect 384822 939863 384878 939919
rect 384946 939863 385002 939919
rect 385070 939863 385126 939919
rect 385194 939863 385250 939919
rect 385318 939863 385374 939919
rect 385442 939863 385498 939919
rect 385566 939863 385622 939919
rect 385690 939863 385746 939919
rect 385814 939863 385870 939919
rect 385938 939863 385994 939919
rect 386062 939863 386118 939919
rect 386908 941599 386964 941655
rect 387032 941599 387088 941655
rect 387156 941599 387212 941655
rect 387280 941599 387336 941655
rect 387404 941599 387460 941655
rect 387528 941599 387584 941655
rect 387652 941599 387708 941655
rect 387776 941599 387832 941655
rect 387900 941599 387956 941655
rect 388024 941599 388080 941655
rect 388148 941599 388204 941655
rect 388272 941599 388328 941655
rect 388396 941599 388452 941655
rect 388520 941599 388576 941655
rect 388644 941599 388700 941655
rect 388768 941599 388824 941655
rect 386908 941475 386964 941531
rect 387032 941475 387088 941531
rect 387156 941475 387212 941531
rect 387280 941475 387336 941531
rect 387404 941475 387460 941531
rect 387528 941475 387584 941531
rect 387652 941475 387708 941531
rect 387776 941475 387832 941531
rect 387900 941475 387956 941531
rect 388024 941475 388080 941531
rect 388148 941475 388204 941531
rect 388272 941475 388328 941531
rect 388396 941475 388452 941531
rect 388520 941475 388576 941531
rect 388644 941475 388700 941531
rect 388768 941475 388824 941531
rect 386908 941351 386964 941407
rect 387032 941351 387088 941407
rect 387156 941351 387212 941407
rect 387280 941351 387336 941407
rect 387404 941351 387460 941407
rect 387528 941351 387584 941407
rect 387652 941351 387708 941407
rect 387776 941351 387832 941407
rect 387900 941351 387956 941407
rect 388024 941351 388080 941407
rect 388148 941351 388204 941407
rect 388272 941351 388328 941407
rect 388396 941351 388452 941407
rect 388520 941351 388576 941407
rect 388644 941351 388700 941407
rect 388768 941351 388824 941407
rect 386908 941227 386964 941283
rect 387032 941227 387088 941283
rect 387156 941227 387212 941283
rect 387280 941227 387336 941283
rect 387404 941227 387460 941283
rect 387528 941227 387584 941283
rect 387652 941227 387708 941283
rect 387776 941227 387832 941283
rect 387900 941227 387956 941283
rect 388024 941227 388080 941283
rect 388148 941227 388204 941283
rect 388272 941227 388328 941283
rect 388396 941227 388452 941283
rect 388520 941227 388576 941283
rect 388644 941227 388700 941283
rect 388768 941227 388824 941283
rect 386908 941103 386964 941159
rect 387032 941103 387088 941159
rect 387156 941103 387212 941159
rect 387280 941103 387336 941159
rect 387404 941103 387460 941159
rect 387528 941103 387584 941159
rect 387652 941103 387708 941159
rect 387776 941103 387832 941159
rect 387900 941103 387956 941159
rect 388024 941103 388080 941159
rect 388148 941103 388204 941159
rect 388272 941103 388328 941159
rect 388396 941103 388452 941159
rect 388520 941103 388576 941159
rect 388644 941103 388700 941159
rect 388768 941103 388824 941159
rect 386908 940979 386964 941035
rect 387032 940979 387088 941035
rect 387156 940979 387212 941035
rect 387280 940979 387336 941035
rect 387404 940979 387460 941035
rect 387528 940979 387584 941035
rect 387652 940979 387708 941035
rect 387776 940979 387832 941035
rect 387900 940979 387956 941035
rect 388024 940979 388080 941035
rect 388148 940979 388204 941035
rect 388272 940979 388328 941035
rect 388396 940979 388452 941035
rect 388520 940979 388576 941035
rect 388644 940979 388700 941035
rect 388768 940979 388824 941035
rect 386908 940855 386964 940911
rect 387032 940855 387088 940911
rect 387156 940855 387212 940911
rect 387280 940855 387336 940911
rect 387404 940855 387460 940911
rect 387528 940855 387584 940911
rect 387652 940855 387708 940911
rect 387776 940855 387832 940911
rect 387900 940855 387956 940911
rect 388024 940855 388080 940911
rect 388148 940855 388204 940911
rect 388272 940855 388328 940911
rect 388396 940855 388452 940911
rect 388520 940855 388576 940911
rect 388644 940855 388700 940911
rect 388768 940855 388824 940911
rect 386908 940731 386964 940787
rect 387032 940731 387088 940787
rect 387156 940731 387212 940787
rect 387280 940731 387336 940787
rect 387404 940731 387460 940787
rect 387528 940731 387584 940787
rect 387652 940731 387708 940787
rect 387776 940731 387832 940787
rect 387900 940731 387956 940787
rect 388024 940731 388080 940787
rect 388148 940731 388204 940787
rect 388272 940731 388328 940787
rect 388396 940731 388452 940787
rect 388520 940731 388576 940787
rect 388644 940731 388700 940787
rect 388768 940731 388824 940787
rect 386908 940607 386964 940663
rect 387032 940607 387088 940663
rect 387156 940607 387212 940663
rect 387280 940607 387336 940663
rect 387404 940607 387460 940663
rect 387528 940607 387584 940663
rect 387652 940607 387708 940663
rect 387776 940607 387832 940663
rect 387900 940607 387956 940663
rect 388024 940607 388080 940663
rect 388148 940607 388204 940663
rect 388272 940607 388328 940663
rect 388396 940607 388452 940663
rect 388520 940607 388576 940663
rect 388644 940607 388700 940663
rect 388768 940607 388824 940663
rect 386908 940483 386964 940539
rect 387032 940483 387088 940539
rect 387156 940483 387212 940539
rect 387280 940483 387336 940539
rect 387404 940483 387460 940539
rect 387528 940483 387584 940539
rect 387652 940483 387708 940539
rect 387776 940483 387832 940539
rect 387900 940483 387956 940539
rect 388024 940483 388080 940539
rect 388148 940483 388204 940539
rect 388272 940483 388328 940539
rect 388396 940483 388452 940539
rect 388520 940483 388576 940539
rect 388644 940483 388700 940539
rect 388768 940483 388824 940539
rect 386908 940359 386964 940415
rect 387032 940359 387088 940415
rect 387156 940359 387212 940415
rect 387280 940359 387336 940415
rect 387404 940359 387460 940415
rect 387528 940359 387584 940415
rect 387652 940359 387708 940415
rect 387776 940359 387832 940415
rect 387900 940359 387956 940415
rect 388024 940359 388080 940415
rect 388148 940359 388204 940415
rect 388272 940359 388328 940415
rect 388396 940359 388452 940415
rect 388520 940359 388576 940415
rect 388644 940359 388700 940415
rect 388768 940359 388824 940415
rect 386908 940235 386964 940291
rect 387032 940235 387088 940291
rect 387156 940235 387212 940291
rect 387280 940235 387336 940291
rect 387404 940235 387460 940291
rect 387528 940235 387584 940291
rect 387652 940235 387708 940291
rect 387776 940235 387832 940291
rect 387900 940235 387956 940291
rect 388024 940235 388080 940291
rect 388148 940235 388204 940291
rect 388272 940235 388328 940291
rect 388396 940235 388452 940291
rect 388520 940235 388576 940291
rect 388644 940235 388700 940291
rect 388768 940235 388824 940291
rect 386908 940111 386964 940167
rect 387032 940111 387088 940167
rect 387156 940111 387212 940167
rect 387280 940111 387336 940167
rect 387404 940111 387460 940167
rect 387528 940111 387584 940167
rect 387652 940111 387708 940167
rect 387776 940111 387832 940167
rect 387900 940111 387956 940167
rect 388024 940111 388080 940167
rect 388148 940111 388204 940167
rect 388272 940111 388328 940167
rect 388396 940111 388452 940167
rect 388520 940111 388576 940167
rect 388644 940111 388700 940167
rect 388768 940111 388824 940167
rect 386908 939987 386964 940043
rect 387032 939987 387088 940043
rect 387156 939987 387212 940043
rect 387280 939987 387336 940043
rect 387404 939987 387460 940043
rect 387528 939987 387584 940043
rect 387652 939987 387708 940043
rect 387776 939987 387832 940043
rect 387900 939987 387956 940043
rect 388024 939987 388080 940043
rect 388148 939987 388204 940043
rect 388272 939987 388328 940043
rect 388396 939987 388452 940043
rect 388520 939987 388576 940043
rect 388644 939987 388700 940043
rect 388768 939987 388824 940043
rect 386908 939863 386964 939919
rect 387032 939863 387088 939919
rect 387156 939863 387212 939919
rect 387280 939863 387336 939919
rect 387404 939863 387460 939919
rect 387528 939863 387584 939919
rect 387652 939863 387708 939919
rect 387776 939863 387832 939919
rect 387900 939863 387956 939919
rect 388024 939863 388080 939919
rect 388148 939863 388204 939919
rect 388272 939863 388328 939919
rect 388396 939863 388452 939919
rect 388520 939863 388576 939919
rect 388644 939863 388700 939919
rect 388768 939863 388824 939919
rect 389278 941599 389334 941655
rect 389402 941599 389458 941655
rect 389526 941599 389582 941655
rect 389650 941599 389706 941655
rect 389774 941599 389830 941655
rect 389898 941599 389954 941655
rect 390022 941599 390078 941655
rect 390146 941599 390202 941655
rect 390270 941599 390326 941655
rect 390394 941599 390450 941655
rect 390518 941599 390574 941655
rect 390642 941599 390698 941655
rect 390766 941599 390822 941655
rect 390890 941599 390946 941655
rect 391014 941599 391070 941655
rect 391138 941599 391194 941655
rect 389278 941475 389334 941531
rect 389402 941475 389458 941531
rect 389526 941475 389582 941531
rect 389650 941475 389706 941531
rect 389774 941475 389830 941531
rect 389898 941475 389954 941531
rect 390022 941475 390078 941531
rect 390146 941475 390202 941531
rect 390270 941475 390326 941531
rect 390394 941475 390450 941531
rect 390518 941475 390574 941531
rect 390642 941475 390698 941531
rect 390766 941475 390822 941531
rect 390890 941475 390946 941531
rect 391014 941475 391070 941531
rect 391138 941475 391194 941531
rect 389278 941351 389334 941407
rect 389402 941351 389458 941407
rect 389526 941351 389582 941407
rect 389650 941351 389706 941407
rect 389774 941351 389830 941407
rect 389898 941351 389954 941407
rect 390022 941351 390078 941407
rect 390146 941351 390202 941407
rect 390270 941351 390326 941407
rect 390394 941351 390450 941407
rect 390518 941351 390574 941407
rect 390642 941351 390698 941407
rect 390766 941351 390822 941407
rect 390890 941351 390946 941407
rect 391014 941351 391070 941407
rect 391138 941351 391194 941407
rect 389278 941227 389334 941283
rect 389402 941227 389458 941283
rect 389526 941227 389582 941283
rect 389650 941227 389706 941283
rect 389774 941227 389830 941283
rect 389898 941227 389954 941283
rect 390022 941227 390078 941283
rect 390146 941227 390202 941283
rect 390270 941227 390326 941283
rect 390394 941227 390450 941283
rect 390518 941227 390574 941283
rect 390642 941227 390698 941283
rect 390766 941227 390822 941283
rect 390890 941227 390946 941283
rect 391014 941227 391070 941283
rect 391138 941227 391194 941283
rect 389278 941103 389334 941159
rect 389402 941103 389458 941159
rect 389526 941103 389582 941159
rect 389650 941103 389706 941159
rect 389774 941103 389830 941159
rect 389898 941103 389954 941159
rect 390022 941103 390078 941159
rect 390146 941103 390202 941159
rect 390270 941103 390326 941159
rect 390394 941103 390450 941159
rect 390518 941103 390574 941159
rect 390642 941103 390698 941159
rect 390766 941103 390822 941159
rect 390890 941103 390946 941159
rect 391014 941103 391070 941159
rect 391138 941103 391194 941159
rect 389278 940979 389334 941035
rect 389402 940979 389458 941035
rect 389526 940979 389582 941035
rect 389650 940979 389706 941035
rect 389774 940979 389830 941035
rect 389898 940979 389954 941035
rect 390022 940979 390078 941035
rect 390146 940979 390202 941035
rect 390270 940979 390326 941035
rect 390394 940979 390450 941035
rect 390518 940979 390574 941035
rect 390642 940979 390698 941035
rect 390766 940979 390822 941035
rect 390890 940979 390946 941035
rect 391014 940979 391070 941035
rect 391138 940979 391194 941035
rect 389278 940855 389334 940911
rect 389402 940855 389458 940911
rect 389526 940855 389582 940911
rect 389650 940855 389706 940911
rect 389774 940855 389830 940911
rect 389898 940855 389954 940911
rect 390022 940855 390078 940911
rect 390146 940855 390202 940911
rect 390270 940855 390326 940911
rect 390394 940855 390450 940911
rect 390518 940855 390574 940911
rect 390642 940855 390698 940911
rect 390766 940855 390822 940911
rect 390890 940855 390946 940911
rect 391014 940855 391070 940911
rect 391138 940855 391194 940911
rect 389278 940731 389334 940787
rect 389402 940731 389458 940787
rect 389526 940731 389582 940787
rect 389650 940731 389706 940787
rect 389774 940731 389830 940787
rect 389898 940731 389954 940787
rect 390022 940731 390078 940787
rect 390146 940731 390202 940787
rect 390270 940731 390326 940787
rect 390394 940731 390450 940787
rect 390518 940731 390574 940787
rect 390642 940731 390698 940787
rect 390766 940731 390822 940787
rect 390890 940731 390946 940787
rect 391014 940731 391070 940787
rect 391138 940731 391194 940787
rect 389278 940607 389334 940663
rect 389402 940607 389458 940663
rect 389526 940607 389582 940663
rect 389650 940607 389706 940663
rect 389774 940607 389830 940663
rect 389898 940607 389954 940663
rect 390022 940607 390078 940663
rect 390146 940607 390202 940663
rect 390270 940607 390326 940663
rect 390394 940607 390450 940663
rect 390518 940607 390574 940663
rect 390642 940607 390698 940663
rect 390766 940607 390822 940663
rect 390890 940607 390946 940663
rect 391014 940607 391070 940663
rect 391138 940607 391194 940663
rect 389278 940483 389334 940539
rect 389402 940483 389458 940539
rect 389526 940483 389582 940539
rect 389650 940483 389706 940539
rect 389774 940483 389830 940539
rect 389898 940483 389954 940539
rect 390022 940483 390078 940539
rect 390146 940483 390202 940539
rect 390270 940483 390326 940539
rect 390394 940483 390450 940539
rect 390518 940483 390574 940539
rect 390642 940483 390698 940539
rect 390766 940483 390822 940539
rect 390890 940483 390946 940539
rect 391014 940483 391070 940539
rect 391138 940483 391194 940539
rect 389278 940359 389334 940415
rect 389402 940359 389458 940415
rect 389526 940359 389582 940415
rect 389650 940359 389706 940415
rect 389774 940359 389830 940415
rect 389898 940359 389954 940415
rect 390022 940359 390078 940415
rect 390146 940359 390202 940415
rect 390270 940359 390326 940415
rect 390394 940359 390450 940415
rect 390518 940359 390574 940415
rect 390642 940359 390698 940415
rect 390766 940359 390822 940415
rect 390890 940359 390946 940415
rect 391014 940359 391070 940415
rect 391138 940359 391194 940415
rect 389278 940235 389334 940291
rect 389402 940235 389458 940291
rect 389526 940235 389582 940291
rect 389650 940235 389706 940291
rect 389774 940235 389830 940291
rect 389898 940235 389954 940291
rect 390022 940235 390078 940291
rect 390146 940235 390202 940291
rect 390270 940235 390326 940291
rect 390394 940235 390450 940291
rect 390518 940235 390574 940291
rect 390642 940235 390698 940291
rect 390766 940235 390822 940291
rect 390890 940235 390946 940291
rect 391014 940235 391070 940291
rect 391138 940235 391194 940291
rect 389278 940111 389334 940167
rect 389402 940111 389458 940167
rect 389526 940111 389582 940167
rect 389650 940111 389706 940167
rect 389774 940111 389830 940167
rect 389898 940111 389954 940167
rect 390022 940111 390078 940167
rect 390146 940111 390202 940167
rect 390270 940111 390326 940167
rect 390394 940111 390450 940167
rect 390518 940111 390574 940167
rect 390642 940111 390698 940167
rect 390766 940111 390822 940167
rect 390890 940111 390946 940167
rect 391014 940111 391070 940167
rect 391138 940111 391194 940167
rect 389278 939987 389334 940043
rect 389402 939987 389458 940043
rect 389526 939987 389582 940043
rect 389650 939987 389706 940043
rect 389774 939987 389830 940043
rect 389898 939987 389954 940043
rect 390022 939987 390078 940043
rect 390146 939987 390202 940043
rect 390270 939987 390326 940043
rect 390394 939987 390450 940043
rect 390518 939987 390574 940043
rect 390642 939987 390698 940043
rect 390766 939987 390822 940043
rect 390890 939987 390946 940043
rect 391014 939987 391070 940043
rect 391138 939987 391194 940043
rect 389278 939863 389334 939919
rect 389402 939863 389458 939919
rect 389526 939863 389582 939919
rect 389650 939863 389706 939919
rect 389774 939863 389830 939919
rect 389898 939863 389954 939919
rect 390022 939863 390078 939919
rect 390146 939863 390202 939919
rect 390270 939863 390326 939919
rect 390394 939863 390450 939919
rect 390518 939863 390574 939919
rect 390642 939863 390698 939919
rect 390766 939863 390822 939919
rect 390890 939863 390946 939919
rect 391014 939863 391070 939919
rect 391138 939863 391194 939919
rect 391882 941599 391938 941655
rect 392006 941599 392062 941655
rect 392130 941599 392186 941655
rect 392254 941599 392310 941655
rect 392378 941599 392434 941655
rect 392502 941599 392558 941655
rect 392626 941599 392682 941655
rect 392750 941599 392806 941655
rect 392874 941599 392930 941655
rect 392998 941599 393054 941655
rect 393122 941599 393178 941655
rect 393246 941599 393302 941655
rect 393370 941599 393426 941655
rect 393494 941599 393550 941655
rect 393618 941599 393674 941655
rect 391882 941475 391938 941531
rect 392006 941475 392062 941531
rect 392130 941475 392186 941531
rect 392254 941475 392310 941531
rect 392378 941475 392434 941531
rect 392502 941475 392558 941531
rect 392626 941475 392682 941531
rect 392750 941475 392806 941531
rect 392874 941475 392930 941531
rect 392998 941475 393054 941531
rect 393122 941475 393178 941531
rect 393246 941475 393302 941531
rect 393370 941475 393426 941531
rect 393494 941475 393550 941531
rect 393618 941475 393674 941531
rect 391882 941351 391938 941407
rect 392006 941351 392062 941407
rect 392130 941351 392186 941407
rect 392254 941351 392310 941407
rect 392378 941351 392434 941407
rect 392502 941351 392558 941407
rect 392626 941351 392682 941407
rect 392750 941351 392806 941407
rect 392874 941351 392930 941407
rect 392998 941351 393054 941407
rect 393122 941351 393178 941407
rect 393246 941351 393302 941407
rect 393370 941351 393426 941407
rect 393494 941351 393550 941407
rect 393618 941351 393674 941407
rect 391882 941227 391938 941283
rect 392006 941227 392062 941283
rect 392130 941227 392186 941283
rect 392254 941227 392310 941283
rect 392378 941227 392434 941283
rect 392502 941227 392558 941283
rect 392626 941227 392682 941283
rect 392750 941227 392806 941283
rect 392874 941227 392930 941283
rect 392998 941227 393054 941283
rect 393122 941227 393178 941283
rect 393246 941227 393302 941283
rect 393370 941227 393426 941283
rect 393494 941227 393550 941283
rect 393618 941227 393674 941283
rect 391882 941103 391938 941159
rect 392006 941103 392062 941159
rect 392130 941103 392186 941159
rect 392254 941103 392310 941159
rect 392378 941103 392434 941159
rect 392502 941103 392558 941159
rect 392626 941103 392682 941159
rect 392750 941103 392806 941159
rect 392874 941103 392930 941159
rect 392998 941103 393054 941159
rect 393122 941103 393178 941159
rect 393246 941103 393302 941159
rect 393370 941103 393426 941159
rect 393494 941103 393550 941159
rect 393618 941103 393674 941159
rect 391882 940979 391938 941035
rect 392006 940979 392062 941035
rect 392130 940979 392186 941035
rect 392254 940979 392310 941035
rect 392378 940979 392434 941035
rect 392502 940979 392558 941035
rect 392626 940979 392682 941035
rect 392750 940979 392806 941035
rect 392874 940979 392930 941035
rect 392998 940979 393054 941035
rect 393122 940979 393178 941035
rect 393246 940979 393302 941035
rect 393370 940979 393426 941035
rect 393494 940979 393550 941035
rect 393618 940979 393674 941035
rect 391882 940855 391938 940911
rect 392006 940855 392062 940911
rect 392130 940855 392186 940911
rect 392254 940855 392310 940911
rect 392378 940855 392434 940911
rect 392502 940855 392558 940911
rect 392626 940855 392682 940911
rect 392750 940855 392806 940911
rect 392874 940855 392930 940911
rect 392998 940855 393054 940911
rect 393122 940855 393178 940911
rect 393246 940855 393302 940911
rect 393370 940855 393426 940911
rect 393494 940855 393550 940911
rect 393618 940855 393674 940911
rect 391882 940731 391938 940787
rect 392006 940731 392062 940787
rect 392130 940731 392186 940787
rect 392254 940731 392310 940787
rect 392378 940731 392434 940787
rect 392502 940731 392558 940787
rect 392626 940731 392682 940787
rect 392750 940731 392806 940787
rect 392874 940731 392930 940787
rect 392998 940731 393054 940787
rect 393122 940731 393178 940787
rect 393246 940731 393302 940787
rect 393370 940731 393426 940787
rect 393494 940731 393550 940787
rect 393618 940731 393674 940787
rect 391882 940607 391938 940663
rect 392006 940607 392062 940663
rect 392130 940607 392186 940663
rect 392254 940607 392310 940663
rect 392378 940607 392434 940663
rect 392502 940607 392558 940663
rect 392626 940607 392682 940663
rect 392750 940607 392806 940663
rect 392874 940607 392930 940663
rect 392998 940607 393054 940663
rect 393122 940607 393178 940663
rect 393246 940607 393302 940663
rect 393370 940607 393426 940663
rect 393494 940607 393550 940663
rect 393618 940607 393674 940663
rect 391882 940483 391938 940539
rect 392006 940483 392062 940539
rect 392130 940483 392186 940539
rect 392254 940483 392310 940539
rect 392378 940483 392434 940539
rect 392502 940483 392558 940539
rect 392626 940483 392682 940539
rect 392750 940483 392806 940539
rect 392874 940483 392930 940539
rect 392998 940483 393054 940539
rect 393122 940483 393178 940539
rect 393246 940483 393302 940539
rect 393370 940483 393426 940539
rect 393494 940483 393550 940539
rect 393618 940483 393674 940539
rect 391882 940359 391938 940415
rect 392006 940359 392062 940415
rect 392130 940359 392186 940415
rect 392254 940359 392310 940415
rect 392378 940359 392434 940415
rect 392502 940359 392558 940415
rect 392626 940359 392682 940415
rect 392750 940359 392806 940415
rect 392874 940359 392930 940415
rect 392998 940359 393054 940415
rect 393122 940359 393178 940415
rect 393246 940359 393302 940415
rect 393370 940359 393426 940415
rect 393494 940359 393550 940415
rect 393618 940359 393674 940415
rect 391882 940235 391938 940291
rect 392006 940235 392062 940291
rect 392130 940235 392186 940291
rect 392254 940235 392310 940291
rect 392378 940235 392434 940291
rect 392502 940235 392558 940291
rect 392626 940235 392682 940291
rect 392750 940235 392806 940291
rect 392874 940235 392930 940291
rect 392998 940235 393054 940291
rect 393122 940235 393178 940291
rect 393246 940235 393302 940291
rect 393370 940235 393426 940291
rect 393494 940235 393550 940291
rect 393618 940235 393674 940291
rect 391882 940111 391938 940167
rect 392006 940111 392062 940167
rect 392130 940111 392186 940167
rect 392254 940111 392310 940167
rect 392378 940111 392434 940167
rect 392502 940111 392558 940167
rect 392626 940111 392682 940167
rect 392750 940111 392806 940167
rect 392874 940111 392930 940167
rect 392998 940111 393054 940167
rect 393122 940111 393178 940167
rect 393246 940111 393302 940167
rect 393370 940111 393426 940167
rect 393494 940111 393550 940167
rect 393618 940111 393674 940167
rect 391882 939987 391938 940043
rect 392006 939987 392062 940043
rect 392130 939987 392186 940043
rect 392254 939987 392310 940043
rect 392378 939987 392434 940043
rect 392502 939987 392558 940043
rect 392626 939987 392682 940043
rect 392750 939987 392806 940043
rect 392874 939987 392930 940043
rect 392998 939987 393054 940043
rect 393122 939987 393178 940043
rect 393246 939987 393302 940043
rect 393370 939987 393426 940043
rect 393494 939987 393550 940043
rect 393618 939987 393674 940043
rect 391882 939863 391938 939919
rect 392006 939863 392062 939919
rect 392130 939863 392186 939919
rect 392254 939863 392310 939919
rect 392378 939863 392434 939919
rect 392502 939863 392558 939919
rect 392626 939863 392682 939919
rect 392750 939863 392806 939919
rect 392874 939863 392930 939919
rect 392998 939863 393054 939919
rect 393122 939863 393178 939919
rect 393246 939863 393302 939919
rect 393370 939863 393426 939919
rect 393494 939863 393550 939919
rect 393618 939863 393674 939919
rect 599326 941599 599382 941655
rect 599450 941599 599506 941655
rect 599574 941599 599630 941655
rect 599698 941599 599754 941655
rect 599822 941599 599878 941655
rect 599946 941599 600002 941655
rect 600070 941599 600126 941655
rect 600194 941599 600250 941655
rect 600318 941599 600374 941655
rect 600442 941599 600498 941655
rect 600566 941599 600622 941655
rect 600690 941599 600746 941655
rect 600814 941599 600870 941655
rect 600938 941599 600994 941655
rect 601062 941599 601118 941655
rect 599326 941475 599382 941531
rect 599450 941475 599506 941531
rect 599574 941475 599630 941531
rect 599698 941475 599754 941531
rect 599822 941475 599878 941531
rect 599946 941475 600002 941531
rect 600070 941475 600126 941531
rect 600194 941475 600250 941531
rect 600318 941475 600374 941531
rect 600442 941475 600498 941531
rect 600566 941475 600622 941531
rect 600690 941475 600746 941531
rect 600814 941475 600870 941531
rect 600938 941475 600994 941531
rect 601062 941475 601118 941531
rect 599326 941351 599382 941407
rect 599450 941351 599506 941407
rect 599574 941351 599630 941407
rect 599698 941351 599754 941407
rect 599822 941351 599878 941407
rect 599946 941351 600002 941407
rect 600070 941351 600126 941407
rect 600194 941351 600250 941407
rect 600318 941351 600374 941407
rect 600442 941351 600498 941407
rect 600566 941351 600622 941407
rect 600690 941351 600746 941407
rect 600814 941351 600870 941407
rect 600938 941351 600994 941407
rect 601062 941351 601118 941407
rect 599326 941227 599382 941283
rect 599450 941227 599506 941283
rect 599574 941227 599630 941283
rect 599698 941227 599754 941283
rect 599822 941227 599878 941283
rect 599946 941227 600002 941283
rect 600070 941227 600126 941283
rect 600194 941227 600250 941283
rect 600318 941227 600374 941283
rect 600442 941227 600498 941283
rect 600566 941227 600622 941283
rect 600690 941227 600746 941283
rect 600814 941227 600870 941283
rect 600938 941227 600994 941283
rect 601062 941227 601118 941283
rect 599326 941103 599382 941159
rect 599450 941103 599506 941159
rect 599574 941103 599630 941159
rect 599698 941103 599754 941159
rect 599822 941103 599878 941159
rect 599946 941103 600002 941159
rect 600070 941103 600126 941159
rect 600194 941103 600250 941159
rect 600318 941103 600374 941159
rect 600442 941103 600498 941159
rect 600566 941103 600622 941159
rect 600690 941103 600746 941159
rect 600814 941103 600870 941159
rect 600938 941103 600994 941159
rect 601062 941103 601118 941159
rect 599326 940979 599382 941035
rect 599450 940979 599506 941035
rect 599574 940979 599630 941035
rect 599698 940979 599754 941035
rect 599822 940979 599878 941035
rect 599946 940979 600002 941035
rect 600070 940979 600126 941035
rect 600194 940979 600250 941035
rect 600318 940979 600374 941035
rect 600442 940979 600498 941035
rect 600566 940979 600622 941035
rect 600690 940979 600746 941035
rect 600814 940979 600870 941035
rect 600938 940979 600994 941035
rect 601062 940979 601118 941035
rect 599326 940855 599382 940911
rect 599450 940855 599506 940911
rect 599574 940855 599630 940911
rect 599698 940855 599754 940911
rect 599822 940855 599878 940911
rect 599946 940855 600002 940911
rect 600070 940855 600126 940911
rect 600194 940855 600250 940911
rect 600318 940855 600374 940911
rect 600442 940855 600498 940911
rect 600566 940855 600622 940911
rect 600690 940855 600746 940911
rect 600814 940855 600870 940911
rect 600938 940855 600994 940911
rect 601062 940855 601118 940911
rect 599326 940731 599382 940787
rect 599450 940731 599506 940787
rect 599574 940731 599630 940787
rect 599698 940731 599754 940787
rect 599822 940731 599878 940787
rect 599946 940731 600002 940787
rect 600070 940731 600126 940787
rect 600194 940731 600250 940787
rect 600318 940731 600374 940787
rect 600442 940731 600498 940787
rect 600566 940731 600622 940787
rect 600690 940731 600746 940787
rect 600814 940731 600870 940787
rect 600938 940731 600994 940787
rect 601062 940731 601118 940787
rect 599326 940607 599382 940663
rect 599450 940607 599506 940663
rect 599574 940607 599630 940663
rect 599698 940607 599754 940663
rect 599822 940607 599878 940663
rect 599946 940607 600002 940663
rect 600070 940607 600126 940663
rect 600194 940607 600250 940663
rect 600318 940607 600374 940663
rect 600442 940607 600498 940663
rect 600566 940607 600622 940663
rect 600690 940607 600746 940663
rect 600814 940607 600870 940663
rect 600938 940607 600994 940663
rect 601062 940607 601118 940663
rect 599326 940483 599382 940539
rect 599450 940483 599506 940539
rect 599574 940483 599630 940539
rect 599698 940483 599754 940539
rect 599822 940483 599878 940539
rect 599946 940483 600002 940539
rect 600070 940483 600126 940539
rect 600194 940483 600250 940539
rect 600318 940483 600374 940539
rect 600442 940483 600498 940539
rect 600566 940483 600622 940539
rect 600690 940483 600746 940539
rect 600814 940483 600870 940539
rect 600938 940483 600994 940539
rect 601062 940483 601118 940539
rect 599326 940359 599382 940415
rect 599450 940359 599506 940415
rect 599574 940359 599630 940415
rect 599698 940359 599754 940415
rect 599822 940359 599878 940415
rect 599946 940359 600002 940415
rect 600070 940359 600126 940415
rect 600194 940359 600250 940415
rect 600318 940359 600374 940415
rect 600442 940359 600498 940415
rect 600566 940359 600622 940415
rect 600690 940359 600746 940415
rect 600814 940359 600870 940415
rect 600938 940359 600994 940415
rect 601062 940359 601118 940415
rect 599326 940235 599382 940291
rect 599450 940235 599506 940291
rect 599574 940235 599630 940291
rect 599698 940235 599754 940291
rect 599822 940235 599878 940291
rect 599946 940235 600002 940291
rect 600070 940235 600126 940291
rect 600194 940235 600250 940291
rect 600318 940235 600374 940291
rect 600442 940235 600498 940291
rect 600566 940235 600622 940291
rect 600690 940235 600746 940291
rect 600814 940235 600870 940291
rect 600938 940235 600994 940291
rect 601062 940235 601118 940291
rect 599326 940111 599382 940167
rect 599450 940111 599506 940167
rect 599574 940111 599630 940167
rect 599698 940111 599754 940167
rect 599822 940111 599878 940167
rect 599946 940111 600002 940167
rect 600070 940111 600126 940167
rect 600194 940111 600250 940167
rect 600318 940111 600374 940167
rect 600442 940111 600498 940167
rect 600566 940111 600622 940167
rect 600690 940111 600746 940167
rect 600814 940111 600870 940167
rect 600938 940111 600994 940167
rect 601062 940111 601118 940167
rect 599326 939987 599382 940043
rect 599450 939987 599506 940043
rect 599574 939987 599630 940043
rect 599698 939987 599754 940043
rect 599822 939987 599878 940043
rect 599946 939987 600002 940043
rect 600070 939987 600126 940043
rect 600194 939987 600250 940043
rect 600318 939987 600374 940043
rect 600442 939987 600498 940043
rect 600566 939987 600622 940043
rect 600690 939987 600746 940043
rect 600814 939987 600870 940043
rect 600938 939987 600994 940043
rect 601062 939987 601118 940043
rect 599326 939863 599382 939919
rect 599450 939863 599506 939919
rect 599574 939863 599630 939919
rect 599698 939863 599754 939919
rect 599822 939863 599878 939919
rect 599946 939863 600002 939919
rect 600070 939863 600126 939919
rect 600194 939863 600250 939919
rect 600318 939863 600374 939919
rect 600442 939863 600498 939919
rect 600566 939863 600622 939919
rect 600690 939863 600746 939919
rect 600814 939863 600870 939919
rect 600938 939863 600994 939919
rect 601062 939863 601118 939919
rect 601832 941599 601888 941655
rect 601956 941599 602012 941655
rect 602080 941599 602136 941655
rect 602204 941599 602260 941655
rect 602328 941599 602384 941655
rect 602452 941599 602508 941655
rect 602576 941599 602632 941655
rect 602700 941599 602756 941655
rect 602824 941599 602880 941655
rect 602948 941599 603004 941655
rect 603072 941599 603128 941655
rect 603196 941599 603252 941655
rect 603320 941599 603376 941655
rect 603444 941599 603500 941655
rect 603568 941599 603624 941655
rect 603692 941599 603748 941655
rect 601832 941475 601888 941531
rect 601956 941475 602012 941531
rect 602080 941475 602136 941531
rect 602204 941475 602260 941531
rect 602328 941475 602384 941531
rect 602452 941475 602508 941531
rect 602576 941475 602632 941531
rect 602700 941475 602756 941531
rect 602824 941475 602880 941531
rect 602948 941475 603004 941531
rect 603072 941475 603128 941531
rect 603196 941475 603252 941531
rect 603320 941475 603376 941531
rect 603444 941475 603500 941531
rect 603568 941475 603624 941531
rect 603692 941475 603748 941531
rect 601832 941351 601888 941407
rect 601956 941351 602012 941407
rect 602080 941351 602136 941407
rect 602204 941351 602260 941407
rect 602328 941351 602384 941407
rect 602452 941351 602508 941407
rect 602576 941351 602632 941407
rect 602700 941351 602756 941407
rect 602824 941351 602880 941407
rect 602948 941351 603004 941407
rect 603072 941351 603128 941407
rect 603196 941351 603252 941407
rect 603320 941351 603376 941407
rect 603444 941351 603500 941407
rect 603568 941351 603624 941407
rect 603692 941351 603748 941407
rect 601832 941227 601888 941283
rect 601956 941227 602012 941283
rect 602080 941227 602136 941283
rect 602204 941227 602260 941283
rect 602328 941227 602384 941283
rect 602452 941227 602508 941283
rect 602576 941227 602632 941283
rect 602700 941227 602756 941283
rect 602824 941227 602880 941283
rect 602948 941227 603004 941283
rect 603072 941227 603128 941283
rect 603196 941227 603252 941283
rect 603320 941227 603376 941283
rect 603444 941227 603500 941283
rect 603568 941227 603624 941283
rect 603692 941227 603748 941283
rect 601832 941103 601888 941159
rect 601956 941103 602012 941159
rect 602080 941103 602136 941159
rect 602204 941103 602260 941159
rect 602328 941103 602384 941159
rect 602452 941103 602508 941159
rect 602576 941103 602632 941159
rect 602700 941103 602756 941159
rect 602824 941103 602880 941159
rect 602948 941103 603004 941159
rect 603072 941103 603128 941159
rect 603196 941103 603252 941159
rect 603320 941103 603376 941159
rect 603444 941103 603500 941159
rect 603568 941103 603624 941159
rect 603692 941103 603748 941159
rect 601832 940979 601888 941035
rect 601956 940979 602012 941035
rect 602080 940979 602136 941035
rect 602204 940979 602260 941035
rect 602328 940979 602384 941035
rect 602452 940979 602508 941035
rect 602576 940979 602632 941035
rect 602700 940979 602756 941035
rect 602824 940979 602880 941035
rect 602948 940979 603004 941035
rect 603072 940979 603128 941035
rect 603196 940979 603252 941035
rect 603320 940979 603376 941035
rect 603444 940979 603500 941035
rect 603568 940979 603624 941035
rect 603692 940979 603748 941035
rect 601832 940855 601888 940911
rect 601956 940855 602012 940911
rect 602080 940855 602136 940911
rect 602204 940855 602260 940911
rect 602328 940855 602384 940911
rect 602452 940855 602508 940911
rect 602576 940855 602632 940911
rect 602700 940855 602756 940911
rect 602824 940855 602880 940911
rect 602948 940855 603004 940911
rect 603072 940855 603128 940911
rect 603196 940855 603252 940911
rect 603320 940855 603376 940911
rect 603444 940855 603500 940911
rect 603568 940855 603624 940911
rect 603692 940855 603748 940911
rect 601832 940731 601888 940787
rect 601956 940731 602012 940787
rect 602080 940731 602136 940787
rect 602204 940731 602260 940787
rect 602328 940731 602384 940787
rect 602452 940731 602508 940787
rect 602576 940731 602632 940787
rect 602700 940731 602756 940787
rect 602824 940731 602880 940787
rect 602948 940731 603004 940787
rect 603072 940731 603128 940787
rect 603196 940731 603252 940787
rect 603320 940731 603376 940787
rect 603444 940731 603500 940787
rect 603568 940731 603624 940787
rect 603692 940731 603748 940787
rect 601832 940607 601888 940663
rect 601956 940607 602012 940663
rect 602080 940607 602136 940663
rect 602204 940607 602260 940663
rect 602328 940607 602384 940663
rect 602452 940607 602508 940663
rect 602576 940607 602632 940663
rect 602700 940607 602756 940663
rect 602824 940607 602880 940663
rect 602948 940607 603004 940663
rect 603072 940607 603128 940663
rect 603196 940607 603252 940663
rect 603320 940607 603376 940663
rect 603444 940607 603500 940663
rect 603568 940607 603624 940663
rect 603692 940607 603748 940663
rect 601832 940483 601888 940539
rect 601956 940483 602012 940539
rect 602080 940483 602136 940539
rect 602204 940483 602260 940539
rect 602328 940483 602384 940539
rect 602452 940483 602508 940539
rect 602576 940483 602632 940539
rect 602700 940483 602756 940539
rect 602824 940483 602880 940539
rect 602948 940483 603004 940539
rect 603072 940483 603128 940539
rect 603196 940483 603252 940539
rect 603320 940483 603376 940539
rect 603444 940483 603500 940539
rect 603568 940483 603624 940539
rect 603692 940483 603748 940539
rect 601832 940359 601888 940415
rect 601956 940359 602012 940415
rect 602080 940359 602136 940415
rect 602204 940359 602260 940415
rect 602328 940359 602384 940415
rect 602452 940359 602508 940415
rect 602576 940359 602632 940415
rect 602700 940359 602756 940415
rect 602824 940359 602880 940415
rect 602948 940359 603004 940415
rect 603072 940359 603128 940415
rect 603196 940359 603252 940415
rect 603320 940359 603376 940415
rect 603444 940359 603500 940415
rect 603568 940359 603624 940415
rect 603692 940359 603748 940415
rect 601832 940235 601888 940291
rect 601956 940235 602012 940291
rect 602080 940235 602136 940291
rect 602204 940235 602260 940291
rect 602328 940235 602384 940291
rect 602452 940235 602508 940291
rect 602576 940235 602632 940291
rect 602700 940235 602756 940291
rect 602824 940235 602880 940291
rect 602948 940235 603004 940291
rect 603072 940235 603128 940291
rect 603196 940235 603252 940291
rect 603320 940235 603376 940291
rect 603444 940235 603500 940291
rect 603568 940235 603624 940291
rect 603692 940235 603748 940291
rect 601832 940111 601888 940167
rect 601956 940111 602012 940167
rect 602080 940111 602136 940167
rect 602204 940111 602260 940167
rect 602328 940111 602384 940167
rect 602452 940111 602508 940167
rect 602576 940111 602632 940167
rect 602700 940111 602756 940167
rect 602824 940111 602880 940167
rect 602948 940111 603004 940167
rect 603072 940111 603128 940167
rect 603196 940111 603252 940167
rect 603320 940111 603376 940167
rect 603444 940111 603500 940167
rect 603568 940111 603624 940167
rect 603692 940111 603748 940167
rect 601832 939987 601888 940043
rect 601956 939987 602012 940043
rect 602080 939987 602136 940043
rect 602204 939987 602260 940043
rect 602328 939987 602384 940043
rect 602452 939987 602508 940043
rect 602576 939987 602632 940043
rect 602700 939987 602756 940043
rect 602824 939987 602880 940043
rect 602948 939987 603004 940043
rect 603072 939987 603128 940043
rect 603196 939987 603252 940043
rect 603320 939987 603376 940043
rect 603444 939987 603500 940043
rect 603568 939987 603624 940043
rect 603692 939987 603748 940043
rect 601832 939863 601888 939919
rect 601956 939863 602012 939919
rect 602080 939863 602136 939919
rect 602204 939863 602260 939919
rect 602328 939863 602384 939919
rect 602452 939863 602508 939919
rect 602576 939863 602632 939919
rect 602700 939863 602756 939919
rect 602824 939863 602880 939919
rect 602948 939863 603004 939919
rect 603072 939863 603128 939919
rect 603196 939863 603252 939919
rect 603320 939863 603376 939919
rect 603444 939863 603500 939919
rect 603568 939863 603624 939919
rect 603692 939863 603748 939919
rect 605070 941599 605126 941655
rect 605194 941599 605250 941655
rect 605318 941599 605374 941655
rect 605442 941599 605498 941655
rect 605566 941599 605622 941655
rect 605690 941599 605746 941655
rect 605814 941599 605870 941655
rect 605938 941599 605994 941655
rect 606062 941599 606118 941655
rect 605070 941475 605126 941531
rect 605194 941475 605250 941531
rect 605318 941475 605374 941531
rect 605442 941475 605498 941531
rect 605566 941475 605622 941531
rect 605690 941475 605746 941531
rect 605814 941475 605870 941531
rect 605938 941475 605994 941531
rect 606062 941475 606118 941531
rect 605070 941351 605126 941407
rect 605194 941351 605250 941407
rect 605318 941351 605374 941407
rect 605442 941351 605498 941407
rect 605566 941351 605622 941407
rect 605690 941351 605746 941407
rect 605814 941351 605870 941407
rect 605938 941351 605994 941407
rect 606062 941351 606118 941407
rect 605070 941227 605126 941283
rect 605194 941227 605250 941283
rect 605318 941227 605374 941283
rect 605442 941227 605498 941283
rect 605566 941227 605622 941283
rect 605690 941227 605746 941283
rect 605814 941227 605870 941283
rect 605938 941227 605994 941283
rect 606062 941227 606118 941283
rect 605070 941103 605126 941159
rect 605194 941103 605250 941159
rect 605318 941103 605374 941159
rect 605442 941103 605498 941159
rect 605566 941103 605622 941159
rect 605690 941103 605746 941159
rect 605814 941103 605870 941159
rect 605938 941103 605994 941159
rect 606062 941103 606118 941159
rect 605070 940979 605126 941035
rect 605194 940979 605250 941035
rect 605318 940979 605374 941035
rect 605442 940979 605498 941035
rect 605566 940979 605622 941035
rect 605690 940979 605746 941035
rect 605814 940979 605870 941035
rect 605938 940979 605994 941035
rect 606062 940979 606118 941035
rect 605070 940855 605126 940911
rect 605194 940855 605250 940911
rect 605318 940855 605374 940911
rect 605442 940855 605498 940911
rect 605566 940855 605622 940911
rect 605690 940855 605746 940911
rect 605814 940855 605870 940911
rect 605938 940855 605994 940911
rect 606062 940855 606118 940911
rect 605070 940731 605126 940787
rect 605194 940731 605250 940787
rect 605318 940731 605374 940787
rect 605442 940731 605498 940787
rect 605566 940731 605622 940787
rect 605690 940731 605746 940787
rect 605814 940731 605870 940787
rect 605938 940731 605994 940787
rect 606062 940731 606118 940787
rect 605070 940607 605126 940663
rect 605194 940607 605250 940663
rect 605318 940607 605374 940663
rect 605442 940607 605498 940663
rect 605566 940607 605622 940663
rect 605690 940607 605746 940663
rect 605814 940607 605870 940663
rect 605938 940607 605994 940663
rect 606062 940607 606118 940663
rect 605070 940483 605126 940539
rect 605194 940483 605250 940539
rect 605318 940483 605374 940539
rect 605442 940483 605498 940539
rect 605566 940483 605622 940539
rect 605690 940483 605746 940539
rect 605814 940483 605870 940539
rect 605938 940483 605994 940539
rect 606062 940483 606118 940539
rect 605070 940359 605126 940415
rect 605194 940359 605250 940415
rect 605318 940359 605374 940415
rect 605442 940359 605498 940415
rect 605566 940359 605622 940415
rect 605690 940359 605746 940415
rect 605814 940359 605870 940415
rect 605938 940359 605994 940415
rect 606062 940359 606118 940415
rect 605070 940235 605126 940291
rect 605194 940235 605250 940291
rect 605318 940235 605374 940291
rect 605442 940235 605498 940291
rect 605566 940235 605622 940291
rect 605690 940235 605746 940291
rect 605814 940235 605870 940291
rect 605938 940235 605994 940291
rect 606062 940235 606118 940291
rect 605070 940111 605126 940167
rect 605194 940111 605250 940167
rect 605318 940111 605374 940167
rect 605442 940111 605498 940167
rect 605566 940111 605622 940167
rect 605690 940111 605746 940167
rect 605814 940111 605870 940167
rect 605938 940111 605994 940167
rect 606062 940111 606118 940167
rect 605070 939987 605126 940043
rect 605194 939987 605250 940043
rect 605318 939987 605374 940043
rect 605442 939987 605498 940043
rect 605566 939987 605622 940043
rect 605690 939987 605746 940043
rect 605814 939987 605870 940043
rect 605938 939987 605994 940043
rect 606062 939987 606118 940043
rect 605070 939863 605126 939919
rect 605194 939863 605250 939919
rect 605318 939863 605374 939919
rect 605442 939863 605498 939919
rect 605566 939863 605622 939919
rect 605690 939863 605746 939919
rect 605814 939863 605870 939919
rect 605938 939863 605994 939919
rect 606062 939863 606118 939919
rect 606908 941599 606964 941655
rect 607032 941599 607088 941655
rect 607156 941599 607212 941655
rect 607280 941599 607336 941655
rect 607404 941599 607460 941655
rect 607528 941599 607584 941655
rect 607652 941599 607708 941655
rect 607776 941599 607832 941655
rect 607900 941599 607956 941655
rect 608024 941599 608080 941655
rect 608148 941599 608204 941655
rect 608272 941599 608328 941655
rect 608396 941599 608452 941655
rect 608520 941599 608576 941655
rect 608644 941599 608700 941655
rect 608768 941599 608824 941655
rect 606908 941475 606964 941531
rect 607032 941475 607088 941531
rect 607156 941475 607212 941531
rect 607280 941475 607336 941531
rect 607404 941475 607460 941531
rect 607528 941475 607584 941531
rect 607652 941475 607708 941531
rect 607776 941475 607832 941531
rect 607900 941475 607956 941531
rect 608024 941475 608080 941531
rect 608148 941475 608204 941531
rect 608272 941475 608328 941531
rect 608396 941475 608452 941531
rect 608520 941475 608576 941531
rect 608644 941475 608700 941531
rect 608768 941475 608824 941531
rect 606908 941351 606964 941407
rect 607032 941351 607088 941407
rect 607156 941351 607212 941407
rect 607280 941351 607336 941407
rect 607404 941351 607460 941407
rect 607528 941351 607584 941407
rect 607652 941351 607708 941407
rect 607776 941351 607832 941407
rect 607900 941351 607956 941407
rect 608024 941351 608080 941407
rect 608148 941351 608204 941407
rect 608272 941351 608328 941407
rect 608396 941351 608452 941407
rect 608520 941351 608576 941407
rect 608644 941351 608700 941407
rect 608768 941351 608824 941407
rect 606908 941227 606964 941283
rect 607032 941227 607088 941283
rect 607156 941227 607212 941283
rect 607280 941227 607336 941283
rect 607404 941227 607460 941283
rect 607528 941227 607584 941283
rect 607652 941227 607708 941283
rect 607776 941227 607832 941283
rect 607900 941227 607956 941283
rect 608024 941227 608080 941283
rect 608148 941227 608204 941283
rect 608272 941227 608328 941283
rect 608396 941227 608452 941283
rect 608520 941227 608576 941283
rect 608644 941227 608700 941283
rect 608768 941227 608824 941283
rect 606908 941103 606964 941159
rect 607032 941103 607088 941159
rect 607156 941103 607212 941159
rect 607280 941103 607336 941159
rect 607404 941103 607460 941159
rect 607528 941103 607584 941159
rect 607652 941103 607708 941159
rect 607776 941103 607832 941159
rect 607900 941103 607956 941159
rect 608024 941103 608080 941159
rect 608148 941103 608204 941159
rect 608272 941103 608328 941159
rect 608396 941103 608452 941159
rect 608520 941103 608576 941159
rect 608644 941103 608700 941159
rect 608768 941103 608824 941159
rect 606908 940979 606964 941035
rect 607032 940979 607088 941035
rect 607156 940979 607212 941035
rect 607280 940979 607336 941035
rect 607404 940979 607460 941035
rect 607528 940979 607584 941035
rect 607652 940979 607708 941035
rect 607776 940979 607832 941035
rect 607900 940979 607956 941035
rect 608024 940979 608080 941035
rect 608148 940979 608204 941035
rect 608272 940979 608328 941035
rect 608396 940979 608452 941035
rect 608520 940979 608576 941035
rect 608644 940979 608700 941035
rect 608768 940979 608824 941035
rect 606908 940855 606964 940911
rect 607032 940855 607088 940911
rect 607156 940855 607212 940911
rect 607280 940855 607336 940911
rect 607404 940855 607460 940911
rect 607528 940855 607584 940911
rect 607652 940855 607708 940911
rect 607776 940855 607832 940911
rect 607900 940855 607956 940911
rect 608024 940855 608080 940911
rect 608148 940855 608204 940911
rect 608272 940855 608328 940911
rect 608396 940855 608452 940911
rect 608520 940855 608576 940911
rect 608644 940855 608700 940911
rect 608768 940855 608824 940911
rect 606908 940731 606964 940787
rect 607032 940731 607088 940787
rect 607156 940731 607212 940787
rect 607280 940731 607336 940787
rect 607404 940731 607460 940787
rect 607528 940731 607584 940787
rect 607652 940731 607708 940787
rect 607776 940731 607832 940787
rect 607900 940731 607956 940787
rect 608024 940731 608080 940787
rect 608148 940731 608204 940787
rect 608272 940731 608328 940787
rect 608396 940731 608452 940787
rect 608520 940731 608576 940787
rect 608644 940731 608700 940787
rect 608768 940731 608824 940787
rect 606908 940607 606964 940663
rect 607032 940607 607088 940663
rect 607156 940607 607212 940663
rect 607280 940607 607336 940663
rect 607404 940607 607460 940663
rect 607528 940607 607584 940663
rect 607652 940607 607708 940663
rect 607776 940607 607832 940663
rect 607900 940607 607956 940663
rect 608024 940607 608080 940663
rect 608148 940607 608204 940663
rect 608272 940607 608328 940663
rect 608396 940607 608452 940663
rect 608520 940607 608576 940663
rect 608644 940607 608700 940663
rect 608768 940607 608824 940663
rect 606908 940483 606964 940539
rect 607032 940483 607088 940539
rect 607156 940483 607212 940539
rect 607280 940483 607336 940539
rect 607404 940483 607460 940539
rect 607528 940483 607584 940539
rect 607652 940483 607708 940539
rect 607776 940483 607832 940539
rect 607900 940483 607956 940539
rect 608024 940483 608080 940539
rect 608148 940483 608204 940539
rect 608272 940483 608328 940539
rect 608396 940483 608452 940539
rect 608520 940483 608576 940539
rect 608644 940483 608700 940539
rect 608768 940483 608824 940539
rect 606908 940359 606964 940415
rect 607032 940359 607088 940415
rect 607156 940359 607212 940415
rect 607280 940359 607336 940415
rect 607404 940359 607460 940415
rect 607528 940359 607584 940415
rect 607652 940359 607708 940415
rect 607776 940359 607832 940415
rect 607900 940359 607956 940415
rect 608024 940359 608080 940415
rect 608148 940359 608204 940415
rect 608272 940359 608328 940415
rect 608396 940359 608452 940415
rect 608520 940359 608576 940415
rect 608644 940359 608700 940415
rect 608768 940359 608824 940415
rect 606908 940235 606964 940291
rect 607032 940235 607088 940291
rect 607156 940235 607212 940291
rect 607280 940235 607336 940291
rect 607404 940235 607460 940291
rect 607528 940235 607584 940291
rect 607652 940235 607708 940291
rect 607776 940235 607832 940291
rect 607900 940235 607956 940291
rect 608024 940235 608080 940291
rect 608148 940235 608204 940291
rect 608272 940235 608328 940291
rect 608396 940235 608452 940291
rect 608520 940235 608576 940291
rect 608644 940235 608700 940291
rect 608768 940235 608824 940291
rect 606908 940111 606964 940167
rect 607032 940111 607088 940167
rect 607156 940111 607212 940167
rect 607280 940111 607336 940167
rect 607404 940111 607460 940167
rect 607528 940111 607584 940167
rect 607652 940111 607708 940167
rect 607776 940111 607832 940167
rect 607900 940111 607956 940167
rect 608024 940111 608080 940167
rect 608148 940111 608204 940167
rect 608272 940111 608328 940167
rect 608396 940111 608452 940167
rect 608520 940111 608576 940167
rect 608644 940111 608700 940167
rect 608768 940111 608824 940167
rect 606908 939987 606964 940043
rect 607032 939987 607088 940043
rect 607156 939987 607212 940043
rect 607280 939987 607336 940043
rect 607404 939987 607460 940043
rect 607528 939987 607584 940043
rect 607652 939987 607708 940043
rect 607776 939987 607832 940043
rect 607900 939987 607956 940043
rect 608024 939987 608080 940043
rect 608148 939987 608204 940043
rect 608272 939987 608328 940043
rect 608396 939987 608452 940043
rect 608520 939987 608576 940043
rect 608644 939987 608700 940043
rect 608768 939987 608824 940043
rect 606908 939863 606964 939919
rect 607032 939863 607088 939919
rect 607156 939863 607212 939919
rect 607280 939863 607336 939919
rect 607404 939863 607460 939919
rect 607528 939863 607584 939919
rect 607652 939863 607708 939919
rect 607776 939863 607832 939919
rect 607900 939863 607956 939919
rect 608024 939863 608080 939919
rect 608148 939863 608204 939919
rect 608272 939863 608328 939919
rect 608396 939863 608452 939919
rect 608520 939863 608576 939919
rect 608644 939863 608700 939919
rect 608768 939863 608824 939919
rect 609278 941599 609334 941655
rect 609402 941599 609458 941655
rect 609526 941599 609582 941655
rect 609650 941599 609706 941655
rect 609774 941599 609830 941655
rect 609898 941599 609954 941655
rect 610022 941599 610078 941655
rect 610146 941599 610202 941655
rect 610270 941599 610326 941655
rect 610394 941599 610450 941655
rect 610518 941599 610574 941655
rect 610642 941599 610698 941655
rect 610766 941599 610822 941655
rect 610890 941599 610946 941655
rect 611014 941599 611070 941655
rect 611138 941599 611194 941655
rect 609278 941475 609334 941531
rect 609402 941475 609458 941531
rect 609526 941475 609582 941531
rect 609650 941475 609706 941531
rect 609774 941475 609830 941531
rect 609898 941475 609954 941531
rect 610022 941475 610078 941531
rect 610146 941475 610202 941531
rect 610270 941475 610326 941531
rect 610394 941475 610450 941531
rect 610518 941475 610574 941531
rect 610642 941475 610698 941531
rect 610766 941475 610822 941531
rect 610890 941475 610946 941531
rect 611014 941475 611070 941531
rect 611138 941475 611194 941531
rect 609278 941351 609334 941407
rect 609402 941351 609458 941407
rect 609526 941351 609582 941407
rect 609650 941351 609706 941407
rect 609774 941351 609830 941407
rect 609898 941351 609954 941407
rect 610022 941351 610078 941407
rect 610146 941351 610202 941407
rect 610270 941351 610326 941407
rect 610394 941351 610450 941407
rect 610518 941351 610574 941407
rect 610642 941351 610698 941407
rect 610766 941351 610822 941407
rect 610890 941351 610946 941407
rect 611014 941351 611070 941407
rect 611138 941351 611194 941407
rect 609278 941227 609334 941283
rect 609402 941227 609458 941283
rect 609526 941227 609582 941283
rect 609650 941227 609706 941283
rect 609774 941227 609830 941283
rect 609898 941227 609954 941283
rect 610022 941227 610078 941283
rect 610146 941227 610202 941283
rect 610270 941227 610326 941283
rect 610394 941227 610450 941283
rect 610518 941227 610574 941283
rect 610642 941227 610698 941283
rect 610766 941227 610822 941283
rect 610890 941227 610946 941283
rect 611014 941227 611070 941283
rect 611138 941227 611194 941283
rect 609278 941103 609334 941159
rect 609402 941103 609458 941159
rect 609526 941103 609582 941159
rect 609650 941103 609706 941159
rect 609774 941103 609830 941159
rect 609898 941103 609954 941159
rect 610022 941103 610078 941159
rect 610146 941103 610202 941159
rect 610270 941103 610326 941159
rect 610394 941103 610450 941159
rect 610518 941103 610574 941159
rect 610642 941103 610698 941159
rect 610766 941103 610822 941159
rect 610890 941103 610946 941159
rect 611014 941103 611070 941159
rect 611138 941103 611194 941159
rect 609278 940979 609334 941035
rect 609402 940979 609458 941035
rect 609526 940979 609582 941035
rect 609650 940979 609706 941035
rect 609774 940979 609830 941035
rect 609898 940979 609954 941035
rect 610022 940979 610078 941035
rect 610146 940979 610202 941035
rect 610270 940979 610326 941035
rect 610394 940979 610450 941035
rect 610518 940979 610574 941035
rect 610642 940979 610698 941035
rect 610766 940979 610822 941035
rect 610890 940979 610946 941035
rect 611014 940979 611070 941035
rect 611138 940979 611194 941035
rect 609278 940855 609334 940911
rect 609402 940855 609458 940911
rect 609526 940855 609582 940911
rect 609650 940855 609706 940911
rect 609774 940855 609830 940911
rect 609898 940855 609954 940911
rect 610022 940855 610078 940911
rect 610146 940855 610202 940911
rect 610270 940855 610326 940911
rect 610394 940855 610450 940911
rect 610518 940855 610574 940911
rect 610642 940855 610698 940911
rect 610766 940855 610822 940911
rect 610890 940855 610946 940911
rect 611014 940855 611070 940911
rect 611138 940855 611194 940911
rect 609278 940731 609334 940787
rect 609402 940731 609458 940787
rect 609526 940731 609582 940787
rect 609650 940731 609706 940787
rect 609774 940731 609830 940787
rect 609898 940731 609954 940787
rect 610022 940731 610078 940787
rect 610146 940731 610202 940787
rect 610270 940731 610326 940787
rect 610394 940731 610450 940787
rect 610518 940731 610574 940787
rect 610642 940731 610698 940787
rect 610766 940731 610822 940787
rect 610890 940731 610946 940787
rect 611014 940731 611070 940787
rect 611138 940731 611194 940787
rect 609278 940607 609334 940663
rect 609402 940607 609458 940663
rect 609526 940607 609582 940663
rect 609650 940607 609706 940663
rect 609774 940607 609830 940663
rect 609898 940607 609954 940663
rect 610022 940607 610078 940663
rect 610146 940607 610202 940663
rect 610270 940607 610326 940663
rect 610394 940607 610450 940663
rect 610518 940607 610574 940663
rect 610642 940607 610698 940663
rect 610766 940607 610822 940663
rect 610890 940607 610946 940663
rect 611014 940607 611070 940663
rect 611138 940607 611194 940663
rect 609278 940483 609334 940539
rect 609402 940483 609458 940539
rect 609526 940483 609582 940539
rect 609650 940483 609706 940539
rect 609774 940483 609830 940539
rect 609898 940483 609954 940539
rect 610022 940483 610078 940539
rect 610146 940483 610202 940539
rect 610270 940483 610326 940539
rect 610394 940483 610450 940539
rect 610518 940483 610574 940539
rect 610642 940483 610698 940539
rect 610766 940483 610822 940539
rect 610890 940483 610946 940539
rect 611014 940483 611070 940539
rect 611138 940483 611194 940539
rect 609278 940359 609334 940415
rect 609402 940359 609458 940415
rect 609526 940359 609582 940415
rect 609650 940359 609706 940415
rect 609774 940359 609830 940415
rect 609898 940359 609954 940415
rect 610022 940359 610078 940415
rect 610146 940359 610202 940415
rect 610270 940359 610326 940415
rect 610394 940359 610450 940415
rect 610518 940359 610574 940415
rect 610642 940359 610698 940415
rect 610766 940359 610822 940415
rect 610890 940359 610946 940415
rect 611014 940359 611070 940415
rect 611138 940359 611194 940415
rect 609278 940235 609334 940291
rect 609402 940235 609458 940291
rect 609526 940235 609582 940291
rect 609650 940235 609706 940291
rect 609774 940235 609830 940291
rect 609898 940235 609954 940291
rect 610022 940235 610078 940291
rect 610146 940235 610202 940291
rect 610270 940235 610326 940291
rect 610394 940235 610450 940291
rect 610518 940235 610574 940291
rect 610642 940235 610698 940291
rect 610766 940235 610822 940291
rect 610890 940235 610946 940291
rect 611014 940235 611070 940291
rect 611138 940235 611194 940291
rect 609278 940111 609334 940167
rect 609402 940111 609458 940167
rect 609526 940111 609582 940167
rect 609650 940111 609706 940167
rect 609774 940111 609830 940167
rect 609898 940111 609954 940167
rect 610022 940111 610078 940167
rect 610146 940111 610202 940167
rect 610270 940111 610326 940167
rect 610394 940111 610450 940167
rect 610518 940111 610574 940167
rect 610642 940111 610698 940167
rect 610766 940111 610822 940167
rect 610890 940111 610946 940167
rect 611014 940111 611070 940167
rect 611138 940111 611194 940167
rect 609278 939987 609334 940043
rect 609402 939987 609458 940043
rect 609526 939987 609582 940043
rect 609650 939987 609706 940043
rect 609774 939987 609830 940043
rect 609898 939987 609954 940043
rect 610022 939987 610078 940043
rect 610146 939987 610202 940043
rect 610270 939987 610326 940043
rect 610394 939987 610450 940043
rect 610518 939987 610574 940043
rect 610642 939987 610698 940043
rect 610766 939987 610822 940043
rect 610890 939987 610946 940043
rect 611014 939987 611070 940043
rect 611138 939987 611194 940043
rect 609278 939863 609334 939919
rect 609402 939863 609458 939919
rect 609526 939863 609582 939919
rect 609650 939863 609706 939919
rect 609774 939863 609830 939919
rect 609898 939863 609954 939919
rect 610022 939863 610078 939919
rect 610146 939863 610202 939919
rect 610270 939863 610326 939919
rect 610394 939863 610450 939919
rect 610518 939863 610574 939919
rect 610642 939863 610698 939919
rect 610766 939863 610822 939919
rect 610890 939863 610946 939919
rect 611014 939863 611070 939919
rect 611138 939863 611194 939919
rect 611882 941599 611938 941655
rect 612006 941599 612062 941655
rect 612130 941599 612186 941655
rect 612254 941599 612310 941655
rect 612378 941599 612434 941655
rect 612502 941599 612558 941655
rect 612626 941599 612682 941655
rect 612750 941599 612806 941655
rect 612874 941599 612930 941655
rect 612998 941599 613054 941655
rect 613122 941599 613178 941655
rect 613246 941599 613302 941655
rect 613370 941599 613426 941655
rect 613494 941599 613550 941655
rect 613618 941599 613674 941655
rect 611882 941475 611938 941531
rect 612006 941475 612062 941531
rect 612130 941475 612186 941531
rect 612254 941475 612310 941531
rect 612378 941475 612434 941531
rect 612502 941475 612558 941531
rect 612626 941475 612682 941531
rect 612750 941475 612806 941531
rect 612874 941475 612930 941531
rect 612998 941475 613054 941531
rect 613122 941475 613178 941531
rect 613246 941475 613302 941531
rect 613370 941475 613426 941531
rect 613494 941475 613550 941531
rect 613618 941475 613674 941531
rect 611882 941351 611938 941407
rect 612006 941351 612062 941407
rect 612130 941351 612186 941407
rect 612254 941351 612310 941407
rect 612378 941351 612434 941407
rect 612502 941351 612558 941407
rect 612626 941351 612682 941407
rect 612750 941351 612806 941407
rect 612874 941351 612930 941407
rect 612998 941351 613054 941407
rect 613122 941351 613178 941407
rect 613246 941351 613302 941407
rect 613370 941351 613426 941407
rect 613494 941351 613550 941407
rect 613618 941351 613674 941407
rect 611882 941227 611938 941283
rect 612006 941227 612062 941283
rect 612130 941227 612186 941283
rect 612254 941227 612310 941283
rect 612378 941227 612434 941283
rect 612502 941227 612558 941283
rect 612626 941227 612682 941283
rect 612750 941227 612806 941283
rect 612874 941227 612930 941283
rect 612998 941227 613054 941283
rect 613122 941227 613178 941283
rect 613246 941227 613302 941283
rect 613370 941227 613426 941283
rect 613494 941227 613550 941283
rect 613618 941227 613674 941283
rect 611882 941103 611938 941159
rect 612006 941103 612062 941159
rect 612130 941103 612186 941159
rect 612254 941103 612310 941159
rect 612378 941103 612434 941159
rect 612502 941103 612558 941159
rect 612626 941103 612682 941159
rect 612750 941103 612806 941159
rect 612874 941103 612930 941159
rect 612998 941103 613054 941159
rect 613122 941103 613178 941159
rect 613246 941103 613302 941159
rect 613370 941103 613426 941159
rect 613494 941103 613550 941159
rect 613618 941103 613674 941159
rect 611882 940979 611938 941035
rect 612006 940979 612062 941035
rect 612130 940979 612186 941035
rect 612254 940979 612310 941035
rect 612378 940979 612434 941035
rect 612502 940979 612558 941035
rect 612626 940979 612682 941035
rect 612750 940979 612806 941035
rect 612874 940979 612930 941035
rect 612998 940979 613054 941035
rect 613122 940979 613178 941035
rect 613246 940979 613302 941035
rect 613370 940979 613426 941035
rect 613494 940979 613550 941035
rect 613618 940979 613674 941035
rect 611882 940855 611938 940911
rect 612006 940855 612062 940911
rect 612130 940855 612186 940911
rect 612254 940855 612310 940911
rect 612378 940855 612434 940911
rect 612502 940855 612558 940911
rect 612626 940855 612682 940911
rect 612750 940855 612806 940911
rect 612874 940855 612930 940911
rect 612998 940855 613054 940911
rect 613122 940855 613178 940911
rect 613246 940855 613302 940911
rect 613370 940855 613426 940911
rect 613494 940855 613550 940911
rect 613618 940855 613674 940911
rect 611882 940731 611938 940787
rect 612006 940731 612062 940787
rect 612130 940731 612186 940787
rect 612254 940731 612310 940787
rect 612378 940731 612434 940787
rect 612502 940731 612558 940787
rect 612626 940731 612682 940787
rect 612750 940731 612806 940787
rect 612874 940731 612930 940787
rect 612998 940731 613054 940787
rect 613122 940731 613178 940787
rect 613246 940731 613302 940787
rect 613370 940731 613426 940787
rect 613494 940731 613550 940787
rect 613618 940731 613674 940787
rect 611882 940607 611938 940663
rect 612006 940607 612062 940663
rect 612130 940607 612186 940663
rect 612254 940607 612310 940663
rect 612378 940607 612434 940663
rect 612502 940607 612558 940663
rect 612626 940607 612682 940663
rect 612750 940607 612806 940663
rect 612874 940607 612930 940663
rect 612998 940607 613054 940663
rect 613122 940607 613178 940663
rect 613246 940607 613302 940663
rect 613370 940607 613426 940663
rect 613494 940607 613550 940663
rect 613618 940607 613674 940663
rect 611882 940483 611938 940539
rect 612006 940483 612062 940539
rect 612130 940483 612186 940539
rect 612254 940483 612310 940539
rect 612378 940483 612434 940539
rect 612502 940483 612558 940539
rect 612626 940483 612682 940539
rect 612750 940483 612806 940539
rect 612874 940483 612930 940539
rect 612998 940483 613054 940539
rect 613122 940483 613178 940539
rect 613246 940483 613302 940539
rect 613370 940483 613426 940539
rect 613494 940483 613550 940539
rect 613618 940483 613674 940539
rect 611882 940359 611938 940415
rect 612006 940359 612062 940415
rect 612130 940359 612186 940415
rect 612254 940359 612310 940415
rect 612378 940359 612434 940415
rect 612502 940359 612558 940415
rect 612626 940359 612682 940415
rect 612750 940359 612806 940415
rect 612874 940359 612930 940415
rect 612998 940359 613054 940415
rect 613122 940359 613178 940415
rect 613246 940359 613302 940415
rect 613370 940359 613426 940415
rect 613494 940359 613550 940415
rect 613618 940359 613674 940415
rect 611882 940235 611938 940291
rect 612006 940235 612062 940291
rect 612130 940235 612186 940291
rect 612254 940235 612310 940291
rect 612378 940235 612434 940291
rect 612502 940235 612558 940291
rect 612626 940235 612682 940291
rect 612750 940235 612806 940291
rect 612874 940235 612930 940291
rect 612998 940235 613054 940291
rect 613122 940235 613178 940291
rect 613246 940235 613302 940291
rect 613370 940235 613426 940291
rect 613494 940235 613550 940291
rect 613618 940235 613674 940291
rect 611882 940111 611938 940167
rect 612006 940111 612062 940167
rect 612130 940111 612186 940167
rect 612254 940111 612310 940167
rect 612378 940111 612434 940167
rect 612502 940111 612558 940167
rect 612626 940111 612682 940167
rect 612750 940111 612806 940167
rect 612874 940111 612930 940167
rect 612998 940111 613054 940167
rect 613122 940111 613178 940167
rect 613246 940111 613302 940167
rect 613370 940111 613426 940167
rect 613494 940111 613550 940167
rect 613618 940111 613674 940167
rect 611882 939987 611938 940043
rect 612006 939987 612062 940043
rect 612130 939987 612186 940043
rect 612254 939987 612310 940043
rect 612378 939987 612434 940043
rect 612502 939987 612558 940043
rect 612626 939987 612682 940043
rect 612750 939987 612806 940043
rect 612874 939987 612930 940043
rect 612998 939987 613054 940043
rect 613122 939987 613178 940043
rect 613246 939987 613302 940043
rect 613370 939987 613426 940043
rect 613494 939987 613550 940043
rect 613618 939987 613674 940043
rect 611882 939863 611938 939919
rect 612006 939863 612062 939919
rect 612130 939863 612186 939919
rect 612254 939863 612310 939919
rect 612378 939863 612434 939919
rect 612502 939863 612558 939919
rect 612626 939863 612682 939919
rect 612750 939863 612806 939919
rect 612874 939863 612930 939919
rect 612998 939863 613054 939919
rect 613122 939863 613178 939919
rect 613246 939863 613302 939919
rect 613370 939863 613426 939919
rect 613494 939863 613550 939919
rect 613618 939863 613674 939919
rect 70047 878605 70103 878661
rect 70171 878605 70227 878661
rect 70295 878605 70351 878661
rect 70419 878605 70475 878661
rect 70047 878481 70103 878537
rect 70171 878481 70227 878537
rect 70295 878481 70351 878537
rect 70419 878481 70475 878537
rect 70047 878357 70103 878413
rect 70171 878357 70227 878413
rect 70295 878357 70351 878413
rect 70419 878357 70475 878413
rect 70047 878233 70103 878289
rect 70171 878233 70227 878289
rect 70295 878233 70351 878289
rect 70419 878233 70475 878289
rect 70047 878109 70103 878165
rect 70171 878109 70227 878165
rect 70295 878109 70351 878165
rect 70419 878109 70475 878165
rect 70047 877985 70103 878041
rect 70171 877985 70227 878041
rect 70295 877985 70351 878041
rect 70419 877985 70475 878041
rect 70047 877861 70103 877917
rect 70171 877861 70227 877917
rect 70295 877861 70351 877917
rect 70419 877861 70475 877917
rect 70047 877737 70103 877793
rect 70171 877737 70227 877793
rect 70295 877737 70351 877793
rect 70419 877737 70475 877793
rect 70047 877613 70103 877669
rect 70171 877613 70227 877669
rect 70295 877613 70351 877669
rect 70419 877613 70475 877669
rect 70047 877489 70103 877545
rect 70171 877489 70227 877545
rect 70295 877489 70351 877545
rect 70419 877489 70475 877545
rect 70047 877365 70103 877421
rect 70171 877365 70227 877421
rect 70295 877365 70351 877421
rect 70419 877365 70475 877421
rect 70047 877241 70103 877297
rect 70171 877241 70227 877297
rect 70295 877241 70351 877297
rect 70419 877241 70475 877297
rect 70047 877117 70103 877173
rect 70171 877117 70227 877173
rect 70295 877117 70351 877173
rect 70419 877117 70475 877173
rect 70047 876993 70103 877049
rect 70171 876993 70227 877049
rect 70295 876993 70351 877049
rect 70419 876993 70475 877049
rect 70047 876869 70103 876925
rect 70171 876869 70227 876925
rect 70295 876869 70351 876925
rect 70419 876869 70475 876925
rect 705525 877631 705581 877687
rect 705649 877631 705705 877687
rect 705773 877631 705829 877687
rect 705897 877631 705953 877687
rect 705525 877507 705581 877563
rect 705649 877507 705705 877563
rect 705773 877507 705829 877563
rect 705897 877507 705953 877563
rect 705525 877383 705581 877439
rect 705649 877383 705705 877439
rect 705773 877383 705829 877439
rect 705897 877383 705953 877439
rect 705525 877259 705581 877315
rect 705649 877259 705705 877315
rect 705773 877259 705829 877315
rect 705897 877259 705953 877315
rect 705525 877135 705581 877191
rect 705649 877135 705705 877191
rect 705773 877135 705829 877191
rect 705897 877135 705953 877191
rect 705525 877011 705581 877067
rect 705649 877011 705705 877067
rect 705773 877011 705829 877067
rect 705897 877011 705953 877067
rect 705525 876887 705581 876943
rect 705649 876887 705705 876943
rect 705773 876887 705829 876943
rect 705897 876887 705953 876943
rect 705525 876763 705581 876819
rect 705649 876763 705705 876819
rect 705773 876763 705829 876819
rect 705897 876763 705953 876819
rect 705525 876639 705581 876695
rect 705649 876639 705705 876695
rect 705773 876639 705829 876695
rect 705897 876639 705953 876695
rect 705525 876515 705581 876571
rect 705649 876515 705705 876571
rect 705773 876515 705829 876571
rect 705897 876515 705953 876571
rect 705525 876391 705581 876447
rect 705649 876391 705705 876447
rect 705773 876391 705829 876447
rect 705897 876391 705953 876447
rect 705525 876267 705581 876323
rect 705649 876267 705705 876323
rect 705773 876267 705829 876323
rect 705897 876267 705953 876323
rect 70047 876125 70103 876181
rect 70171 876125 70227 876181
rect 70295 876125 70351 876181
rect 70419 876125 70475 876181
rect 70047 876001 70103 876057
rect 70171 876001 70227 876057
rect 70295 876001 70351 876057
rect 70419 876001 70475 876057
rect 70047 875877 70103 875933
rect 70171 875877 70227 875933
rect 70295 875877 70351 875933
rect 70419 875877 70475 875933
rect 705525 876143 705581 876199
rect 705649 876143 705705 876199
rect 705773 876143 705829 876199
rect 705897 876143 705953 876199
rect 705525 876019 705581 876075
rect 705649 876019 705705 876075
rect 705773 876019 705829 876075
rect 705897 876019 705953 876075
rect 705525 875895 705581 875951
rect 705649 875895 705705 875951
rect 705773 875895 705829 875951
rect 705897 875895 705953 875951
rect 70047 875753 70103 875809
rect 70171 875753 70227 875809
rect 70295 875753 70351 875809
rect 70419 875753 70475 875809
rect 70047 875629 70103 875685
rect 70171 875629 70227 875685
rect 70295 875629 70351 875685
rect 70419 875629 70475 875685
rect 70047 875505 70103 875561
rect 70171 875505 70227 875561
rect 70295 875505 70351 875561
rect 70419 875505 70475 875561
rect 70047 875381 70103 875437
rect 70171 875381 70227 875437
rect 70295 875381 70351 875437
rect 70419 875381 70475 875437
rect 70047 875257 70103 875313
rect 70171 875257 70227 875313
rect 70295 875257 70351 875313
rect 70419 875257 70475 875313
rect 70047 875133 70103 875189
rect 70171 875133 70227 875189
rect 70295 875133 70351 875189
rect 70419 875133 70475 875189
rect 70047 875009 70103 875065
rect 70171 875009 70227 875065
rect 70295 875009 70351 875065
rect 70419 875009 70475 875065
rect 70047 874885 70103 874941
rect 70171 874885 70227 874941
rect 70295 874885 70351 874941
rect 70419 874885 70475 874941
rect 70047 874761 70103 874817
rect 70171 874761 70227 874817
rect 70295 874761 70351 874817
rect 70419 874761 70475 874817
rect 70047 874637 70103 874693
rect 70171 874637 70227 874693
rect 70295 874637 70351 874693
rect 70419 874637 70475 874693
rect 70047 874513 70103 874569
rect 70171 874513 70227 874569
rect 70295 874513 70351 874569
rect 70419 874513 70475 874569
rect 70047 874389 70103 874445
rect 70171 874389 70227 874445
rect 70295 874389 70351 874445
rect 70419 874389 70475 874445
rect 70047 874265 70103 874321
rect 70171 874265 70227 874321
rect 70295 874265 70351 874321
rect 70419 874265 70475 874321
rect 705525 875125 705581 875181
rect 705649 875125 705705 875181
rect 705773 875125 705829 875181
rect 705897 875125 705953 875181
rect 705525 875001 705581 875057
rect 705649 875001 705705 875057
rect 705773 875001 705829 875057
rect 705897 875001 705953 875057
rect 705525 874877 705581 874933
rect 705649 874877 705705 874933
rect 705773 874877 705829 874933
rect 705897 874877 705953 874933
rect 705525 874753 705581 874809
rect 705649 874753 705705 874809
rect 705773 874753 705829 874809
rect 705897 874753 705953 874809
rect 705525 874629 705581 874685
rect 705649 874629 705705 874685
rect 705773 874629 705829 874685
rect 705897 874629 705953 874685
rect 705525 874505 705581 874561
rect 705649 874505 705705 874561
rect 705773 874505 705829 874561
rect 705897 874505 705953 874561
rect 705525 874381 705581 874437
rect 705649 874381 705705 874437
rect 705773 874381 705829 874437
rect 705897 874381 705953 874437
rect 705525 874257 705581 874313
rect 705649 874257 705705 874313
rect 705773 874257 705829 874313
rect 705897 874257 705953 874313
rect 705525 874133 705581 874189
rect 705649 874133 705705 874189
rect 705773 874133 705829 874189
rect 705897 874133 705953 874189
rect 705525 874009 705581 874065
rect 705649 874009 705705 874065
rect 705773 874009 705829 874065
rect 705897 874009 705953 874065
rect 705525 873885 705581 873941
rect 705649 873885 705705 873941
rect 705773 873885 705829 873941
rect 705897 873885 705953 873941
rect 70047 873755 70103 873811
rect 70171 873755 70227 873811
rect 70295 873755 70351 873811
rect 70419 873755 70475 873811
rect 70047 873631 70103 873687
rect 70171 873631 70227 873687
rect 70295 873631 70351 873687
rect 70419 873631 70475 873687
rect 70047 873507 70103 873563
rect 70171 873507 70227 873563
rect 70295 873507 70351 873563
rect 70419 873507 70475 873563
rect 70047 873383 70103 873439
rect 70171 873383 70227 873439
rect 70295 873383 70351 873439
rect 70419 873383 70475 873439
rect 70047 873259 70103 873315
rect 70171 873259 70227 873315
rect 70295 873259 70351 873315
rect 70419 873259 70475 873315
rect 705525 873761 705581 873817
rect 705649 873761 705705 873817
rect 705773 873761 705829 873817
rect 705897 873761 705953 873817
rect 705525 873637 705581 873693
rect 705649 873637 705705 873693
rect 705773 873637 705829 873693
rect 705897 873637 705953 873693
rect 705525 873513 705581 873569
rect 705649 873513 705705 873569
rect 705773 873513 705829 873569
rect 705897 873513 705953 873569
rect 705525 873389 705581 873445
rect 705649 873389 705705 873445
rect 705773 873389 705829 873445
rect 705897 873389 705953 873445
rect 705525 873265 705581 873321
rect 705649 873265 705705 873321
rect 705773 873265 705829 873321
rect 705897 873265 705953 873321
rect 70047 873135 70103 873191
rect 70171 873135 70227 873191
rect 70295 873135 70351 873191
rect 70419 873135 70475 873191
rect 70047 873011 70103 873067
rect 70171 873011 70227 873067
rect 70295 873011 70351 873067
rect 70419 873011 70475 873067
rect 70047 872887 70103 872943
rect 70171 872887 70227 872943
rect 70295 872887 70351 872943
rect 70419 872887 70475 872943
rect 70047 872763 70103 872819
rect 70171 872763 70227 872819
rect 70295 872763 70351 872819
rect 70419 872763 70475 872819
rect 70047 872639 70103 872695
rect 70171 872639 70227 872695
rect 70295 872639 70351 872695
rect 70419 872639 70475 872695
rect 70047 872515 70103 872571
rect 70171 872515 70227 872571
rect 70295 872515 70351 872571
rect 70419 872515 70475 872571
rect 70047 872391 70103 872447
rect 70171 872391 70227 872447
rect 70295 872391 70351 872447
rect 70419 872391 70475 872447
rect 70047 872267 70103 872323
rect 70171 872267 70227 872323
rect 70295 872267 70351 872323
rect 70419 872267 70475 872323
rect 70047 872143 70103 872199
rect 70171 872143 70227 872199
rect 70295 872143 70351 872199
rect 70419 872143 70475 872199
rect 70047 872019 70103 872075
rect 70171 872019 70227 872075
rect 70295 872019 70351 872075
rect 70419 872019 70475 872075
rect 70047 871895 70103 871951
rect 70171 871895 70227 871951
rect 70295 871895 70351 871951
rect 70419 871895 70475 871951
rect 705525 872755 705581 872811
rect 705649 872755 705705 872811
rect 705773 872755 705829 872811
rect 705897 872755 705953 872811
rect 705525 872631 705581 872687
rect 705649 872631 705705 872687
rect 705773 872631 705829 872687
rect 705897 872631 705953 872687
rect 705525 872507 705581 872563
rect 705649 872507 705705 872563
rect 705773 872507 705829 872563
rect 705897 872507 705953 872563
rect 705525 872383 705581 872439
rect 705649 872383 705705 872439
rect 705773 872383 705829 872439
rect 705897 872383 705953 872439
rect 705525 872259 705581 872315
rect 705649 872259 705705 872315
rect 705773 872259 705829 872315
rect 705897 872259 705953 872315
rect 705525 872135 705581 872191
rect 705649 872135 705705 872191
rect 705773 872135 705829 872191
rect 705897 872135 705953 872191
rect 705525 872011 705581 872067
rect 705649 872011 705705 872067
rect 705773 872011 705829 872067
rect 705897 872011 705953 872067
rect 705525 871887 705581 871943
rect 705649 871887 705705 871943
rect 705773 871887 705829 871943
rect 705897 871887 705953 871943
rect 705525 871763 705581 871819
rect 705649 871763 705705 871819
rect 705773 871763 705829 871819
rect 705897 871763 705953 871819
rect 705525 871639 705581 871695
rect 705649 871639 705705 871695
rect 705773 871639 705829 871695
rect 705897 871639 705953 871695
rect 705525 871515 705581 871571
rect 705649 871515 705705 871571
rect 705773 871515 705829 871571
rect 705897 871515 705953 871571
rect 705525 871391 705581 871447
rect 705649 871391 705705 871447
rect 705773 871391 705829 871447
rect 705897 871391 705953 871447
rect 705525 871267 705581 871323
rect 705649 871267 705705 871323
rect 705773 871267 705829 871323
rect 705897 871267 705953 871323
rect 70047 871049 70103 871105
rect 70171 871049 70227 871105
rect 70295 871049 70351 871105
rect 70419 871049 70475 871105
rect 70047 870925 70103 870981
rect 70171 870925 70227 870981
rect 70295 870925 70351 870981
rect 70419 870925 70475 870981
rect 70047 870801 70103 870857
rect 70171 870801 70227 870857
rect 70295 870801 70351 870857
rect 70419 870801 70475 870857
rect 705525 871143 705581 871199
rect 705649 871143 705705 871199
rect 705773 871143 705829 871199
rect 705897 871143 705953 871199
rect 705525 871019 705581 871075
rect 705649 871019 705705 871075
rect 705773 871019 705829 871075
rect 705897 871019 705953 871075
rect 705525 870895 705581 870951
rect 705649 870895 705705 870951
rect 705773 870895 705829 870951
rect 705897 870895 705953 870951
rect 70047 870677 70103 870733
rect 70171 870677 70227 870733
rect 70295 870677 70351 870733
rect 70419 870677 70475 870733
rect 70047 870553 70103 870609
rect 70171 870553 70227 870609
rect 70295 870553 70351 870609
rect 70419 870553 70475 870609
rect 70047 870429 70103 870485
rect 70171 870429 70227 870485
rect 70295 870429 70351 870485
rect 70419 870429 70475 870485
rect 70047 870305 70103 870361
rect 70171 870305 70227 870361
rect 70295 870305 70351 870361
rect 70419 870305 70475 870361
rect 70047 870181 70103 870237
rect 70171 870181 70227 870237
rect 70295 870181 70351 870237
rect 70419 870181 70475 870237
rect 70047 870057 70103 870113
rect 70171 870057 70227 870113
rect 70295 870057 70351 870113
rect 70419 870057 70475 870113
rect 70047 869933 70103 869989
rect 70171 869933 70227 869989
rect 70295 869933 70351 869989
rect 70419 869933 70475 869989
rect 70047 869809 70103 869865
rect 70171 869809 70227 869865
rect 70295 869809 70351 869865
rect 70419 869809 70475 869865
rect 70047 869685 70103 869741
rect 70171 869685 70227 869741
rect 70295 869685 70351 869741
rect 70419 869685 70475 869741
rect 70047 869561 70103 869617
rect 70171 869561 70227 869617
rect 70295 869561 70351 869617
rect 70419 869561 70475 869617
rect 70047 869437 70103 869493
rect 70171 869437 70227 869493
rect 70295 869437 70351 869493
rect 70419 869437 70475 869493
rect 70047 869313 70103 869369
rect 70171 869313 70227 869369
rect 70295 869313 70351 869369
rect 70419 869313 70475 869369
rect 70047 869189 70103 869245
rect 70171 869189 70227 869245
rect 70295 869189 70351 869245
rect 70419 869189 70475 869245
rect 705525 870049 705581 870105
rect 705649 870049 705705 870105
rect 705773 870049 705829 870105
rect 705897 870049 705953 870105
rect 705525 869925 705581 869981
rect 705649 869925 705705 869981
rect 705773 869925 705829 869981
rect 705897 869925 705953 869981
rect 705525 869801 705581 869857
rect 705649 869801 705705 869857
rect 705773 869801 705829 869857
rect 705897 869801 705953 869857
rect 705525 869677 705581 869733
rect 705649 869677 705705 869733
rect 705773 869677 705829 869733
rect 705897 869677 705953 869733
rect 705525 869553 705581 869609
rect 705649 869553 705705 869609
rect 705773 869553 705829 869609
rect 705897 869553 705953 869609
rect 705525 869429 705581 869485
rect 705649 869429 705705 869485
rect 705773 869429 705829 869485
rect 705897 869429 705953 869485
rect 705525 869305 705581 869361
rect 705649 869305 705705 869361
rect 705773 869305 705829 869361
rect 705897 869305 705953 869361
rect 705525 869181 705581 869237
rect 705649 869181 705705 869237
rect 705773 869181 705829 869237
rect 705897 869181 705953 869237
rect 705525 869057 705581 869113
rect 705649 869057 705705 869113
rect 705773 869057 705829 869113
rect 705897 869057 705953 869113
rect 705525 868933 705581 868989
rect 705649 868933 705705 868989
rect 705773 868933 705829 868989
rect 705897 868933 705953 868989
rect 705525 868809 705581 868865
rect 705649 868809 705705 868865
rect 705773 868809 705829 868865
rect 705897 868809 705953 868865
rect 70047 868679 70103 868735
rect 70171 868679 70227 868735
rect 70295 868679 70351 868735
rect 70419 868679 70475 868735
rect 70047 868555 70103 868611
rect 70171 868555 70227 868611
rect 70295 868555 70351 868611
rect 70419 868555 70475 868611
rect 70047 868431 70103 868487
rect 70171 868431 70227 868487
rect 70295 868431 70351 868487
rect 70419 868431 70475 868487
rect 70047 868307 70103 868363
rect 70171 868307 70227 868363
rect 70295 868307 70351 868363
rect 70419 868307 70475 868363
rect 70047 868183 70103 868239
rect 70171 868183 70227 868239
rect 70295 868183 70351 868239
rect 70419 868183 70475 868239
rect 705525 868685 705581 868741
rect 705649 868685 705705 868741
rect 705773 868685 705829 868741
rect 705897 868685 705953 868741
rect 705525 868561 705581 868617
rect 705649 868561 705705 868617
rect 705773 868561 705829 868617
rect 705897 868561 705953 868617
rect 705525 868437 705581 868493
rect 705649 868437 705705 868493
rect 705773 868437 705829 868493
rect 705897 868437 705953 868493
rect 705525 868313 705581 868369
rect 705649 868313 705705 868369
rect 705773 868313 705829 868369
rect 705897 868313 705953 868369
rect 705525 868189 705581 868245
rect 705649 868189 705705 868245
rect 705773 868189 705829 868245
rect 705897 868189 705953 868245
rect 70047 868059 70103 868115
rect 70171 868059 70227 868115
rect 70295 868059 70351 868115
rect 70419 868059 70475 868115
rect 70047 867935 70103 867991
rect 70171 867935 70227 867991
rect 70295 867935 70351 867991
rect 70419 867935 70475 867991
rect 70047 867811 70103 867867
rect 70171 867811 70227 867867
rect 70295 867811 70351 867867
rect 70419 867811 70475 867867
rect 70047 867687 70103 867743
rect 70171 867687 70227 867743
rect 70295 867687 70351 867743
rect 70419 867687 70475 867743
rect 70047 867563 70103 867619
rect 70171 867563 70227 867619
rect 70295 867563 70351 867619
rect 70419 867563 70475 867619
rect 70047 867439 70103 867495
rect 70171 867439 70227 867495
rect 70295 867439 70351 867495
rect 70419 867439 70475 867495
rect 70047 867315 70103 867371
rect 70171 867315 70227 867371
rect 70295 867315 70351 867371
rect 70419 867315 70475 867371
rect 70047 867191 70103 867247
rect 70171 867191 70227 867247
rect 70295 867191 70351 867247
rect 70419 867191 70475 867247
rect 70047 867067 70103 867123
rect 70171 867067 70227 867123
rect 70295 867067 70351 867123
rect 70419 867067 70475 867123
rect 70047 866943 70103 866999
rect 70171 866943 70227 866999
rect 70295 866943 70351 866999
rect 70419 866943 70475 866999
rect 70047 866819 70103 866875
rect 70171 866819 70227 866875
rect 70295 866819 70351 866875
rect 70419 866819 70475 866875
rect 705525 867679 705581 867735
rect 705649 867679 705705 867735
rect 705773 867679 705829 867735
rect 705897 867679 705953 867735
rect 705525 867555 705581 867611
rect 705649 867555 705705 867611
rect 705773 867555 705829 867611
rect 705897 867555 705953 867611
rect 705525 867431 705581 867487
rect 705649 867431 705705 867487
rect 705773 867431 705829 867487
rect 705897 867431 705953 867487
rect 705525 867307 705581 867363
rect 705649 867307 705705 867363
rect 705773 867307 705829 867363
rect 705897 867307 705953 867363
rect 705525 867183 705581 867239
rect 705649 867183 705705 867239
rect 705773 867183 705829 867239
rect 705897 867183 705953 867239
rect 705525 867059 705581 867115
rect 705649 867059 705705 867115
rect 705773 867059 705829 867115
rect 705897 867059 705953 867115
rect 705525 866935 705581 866991
rect 705649 866935 705705 866991
rect 705773 866935 705829 866991
rect 705897 866935 705953 866991
rect 705525 866811 705581 866867
rect 705649 866811 705705 866867
rect 705773 866811 705829 866867
rect 705897 866811 705953 866867
rect 705525 866687 705581 866743
rect 705649 866687 705705 866743
rect 705773 866687 705829 866743
rect 705897 866687 705953 866743
rect 705525 866563 705581 866619
rect 705649 866563 705705 866619
rect 705773 866563 705829 866619
rect 705897 866563 705953 866619
rect 705525 866439 705581 866495
rect 705649 866439 705705 866495
rect 705773 866439 705829 866495
rect 705897 866439 705953 866495
rect 705525 866315 705581 866371
rect 705649 866315 705705 866371
rect 705773 866315 705829 866371
rect 705897 866315 705953 866371
rect 705525 866191 705581 866247
rect 705649 866191 705705 866247
rect 705773 866191 705829 866247
rect 705897 866191 705953 866247
rect 70047 866049 70103 866105
rect 70171 866049 70227 866105
rect 70295 866049 70351 866105
rect 70419 866049 70475 866105
rect 70047 865925 70103 865981
rect 70171 865925 70227 865981
rect 70295 865925 70351 865981
rect 70419 865925 70475 865981
rect 70047 865801 70103 865857
rect 70171 865801 70227 865857
rect 70295 865801 70351 865857
rect 70419 865801 70475 865857
rect 705525 866067 705581 866123
rect 705649 866067 705705 866123
rect 705773 866067 705829 866123
rect 705897 866067 705953 866123
rect 705525 865943 705581 865999
rect 705649 865943 705705 865999
rect 705773 865943 705829 865999
rect 705897 865943 705953 865999
rect 705525 865819 705581 865875
rect 705649 865819 705705 865875
rect 705773 865819 705829 865875
rect 705897 865819 705953 865875
rect 70047 865677 70103 865733
rect 70171 865677 70227 865733
rect 70295 865677 70351 865733
rect 70419 865677 70475 865733
rect 70047 865553 70103 865609
rect 70171 865553 70227 865609
rect 70295 865553 70351 865609
rect 70419 865553 70475 865609
rect 70047 865429 70103 865485
rect 70171 865429 70227 865485
rect 70295 865429 70351 865485
rect 70419 865429 70475 865485
rect 70047 865305 70103 865361
rect 70171 865305 70227 865361
rect 70295 865305 70351 865361
rect 70419 865305 70475 865361
rect 70047 865181 70103 865237
rect 70171 865181 70227 865237
rect 70295 865181 70351 865237
rect 70419 865181 70475 865237
rect 70047 865057 70103 865113
rect 70171 865057 70227 865113
rect 70295 865057 70351 865113
rect 70419 865057 70475 865113
rect 70047 864933 70103 864989
rect 70171 864933 70227 864989
rect 70295 864933 70351 864989
rect 70419 864933 70475 864989
rect 70047 864809 70103 864865
rect 70171 864809 70227 864865
rect 70295 864809 70351 864865
rect 70419 864809 70475 864865
rect 70047 864685 70103 864741
rect 70171 864685 70227 864741
rect 70295 864685 70351 864741
rect 70419 864685 70475 864741
rect 70047 864561 70103 864617
rect 70171 864561 70227 864617
rect 70295 864561 70351 864617
rect 70419 864561 70475 864617
rect 70047 864437 70103 864493
rect 70171 864437 70227 864493
rect 70295 864437 70351 864493
rect 70419 864437 70475 864493
rect 70047 864313 70103 864369
rect 70171 864313 70227 864369
rect 70295 864313 70351 864369
rect 70419 864313 70475 864369
rect 705525 865075 705581 865131
rect 705649 865075 705705 865131
rect 705773 865075 705829 865131
rect 705897 865075 705953 865131
rect 705525 864951 705581 865007
rect 705649 864951 705705 865007
rect 705773 864951 705829 865007
rect 705897 864951 705953 865007
rect 705525 864827 705581 864883
rect 705649 864827 705705 864883
rect 705773 864827 705829 864883
rect 705897 864827 705953 864883
rect 705525 864703 705581 864759
rect 705649 864703 705705 864759
rect 705773 864703 705829 864759
rect 705897 864703 705953 864759
rect 705525 864579 705581 864635
rect 705649 864579 705705 864635
rect 705773 864579 705829 864635
rect 705897 864579 705953 864635
rect 705525 864455 705581 864511
rect 705649 864455 705705 864511
rect 705773 864455 705829 864511
rect 705897 864455 705953 864511
rect 705525 864331 705581 864387
rect 705649 864331 705705 864387
rect 705773 864331 705829 864387
rect 705897 864331 705953 864387
rect 705525 864207 705581 864263
rect 705649 864207 705705 864263
rect 705773 864207 705829 864263
rect 705897 864207 705953 864263
rect 705525 864083 705581 864139
rect 705649 864083 705705 864139
rect 705773 864083 705829 864139
rect 705897 864083 705953 864139
rect 705525 863959 705581 864015
rect 705649 863959 705705 864015
rect 705773 863959 705829 864015
rect 705897 863959 705953 864015
rect 705525 863835 705581 863891
rect 705649 863835 705705 863891
rect 705773 863835 705829 863891
rect 705897 863835 705953 863891
rect 705525 863711 705581 863767
rect 705649 863711 705705 863767
rect 705773 863711 705829 863767
rect 705897 863711 705953 863767
rect 705525 863587 705581 863643
rect 705649 863587 705705 863643
rect 705773 863587 705829 863643
rect 705897 863587 705953 863643
rect 705525 863463 705581 863519
rect 705649 863463 705705 863519
rect 705773 863463 705829 863519
rect 705897 863463 705953 863519
rect 705525 863339 705581 863395
rect 705649 863339 705705 863395
rect 705773 863339 705829 863395
rect 705897 863339 705953 863395
rect 70047 837605 70103 837661
rect 70171 837605 70227 837661
rect 70295 837605 70351 837661
rect 70419 837605 70475 837661
rect 70047 837481 70103 837537
rect 70171 837481 70227 837537
rect 70295 837481 70351 837537
rect 70419 837481 70475 837537
rect 70047 837357 70103 837413
rect 70171 837357 70227 837413
rect 70295 837357 70351 837413
rect 70419 837357 70475 837413
rect 70047 837233 70103 837289
rect 70171 837233 70227 837289
rect 70295 837233 70351 837289
rect 70419 837233 70475 837289
rect 70047 837109 70103 837165
rect 70171 837109 70227 837165
rect 70295 837109 70351 837165
rect 70419 837109 70475 837165
rect 70047 836985 70103 837041
rect 70171 836985 70227 837041
rect 70295 836985 70351 837041
rect 70419 836985 70475 837041
rect 70047 836861 70103 836917
rect 70171 836861 70227 836917
rect 70295 836861 70351 836917
rect 70419 836861 70475 836917
rect 70047 836737 70103 836793
rect 70171 836737 70227 836793
rect 70295 836737 70351 836793
rect 70419 836737 70475 836793
rect 70047 836613 70103 836669
rect 70171 836613 70227 836669
rect 70295 836613 70351 836669
rect 70419 836613 70475 836669
rect 70047 836489 70103 836545
rect 70171 836489 70227 836545
rect 70295 836489 70351 836545
rect 70419 836489 70475 836545
rect 70047 836365 70103 836421
rect 70171 836365 70227 836421
rect 70295 836365 70351 836421
rect 70419 836365 70475 836421
rect 70047 836241 70103 836297
rect 70171 836241 70227 836297
rect 70295 836241 70351 836297
rect 70419 836241 70475 836297
rect 70047 836117 70103 836173
rect 70171 836117 70227 836173
rect 70295 836117 70351 836173
rect 70419 836117 70475 836173
rect 70047 835993 70103 836049
rect 70171 835993 70227 836049
rect 70295 835993 70351 836049
rect 70419 835993 70475 836049
rect 70047 835869 70103 835925
rect 70171 835869 70227 835925
rect 70295 835869 70351 835925
rect 70419 835869 70475 835925
rect 70047 835125 70103 835181
rect 70171 835125 70227 835181
rect 70295 835125 70351 835181
rect 70419 835125 70475 835181
rect 70047 835001 70103 835057
rect 70171 835001 70227 835057
rect 70295 835001 70351 835057
rect 70419 835001 70475 835057
rect 70047 834877 70103 834933
rect 70171 834877 70227 834933
rect 70295 834877 70351 834933
rect 70419 834877 70475 834933
rect 70047 834753 70103 834809
rect 70171 834753 70227 834809
rect 70295 834753 70351 834809
rect 70419 834753 70475 834809
rect 70047 834629 70103 834685
rect 70171 834629 70227 834685
rect 70295 834629 70351 834685
rect 70419 834629 70475 834685
rect 70047 834505 70103 834561
rect 70171 834505 70227 834561
rect 70295 834505 70351 834561
rect 70419 834505 70475 834561
rect 70047 834381 70103 834437
rect 70171 834381 70227 834437
rect 70295 834381 70351 834437
rect 70419 834381 70475 834437
rect 70047 834257 70103 834313
rect 70171 834257 70227 834313
rect 70295 834257 70351 834313
rect 70419 834257 70475 834313
rect 70047 834133 70103 834189
rect 70171 834133 70227 834189
rect 70295 834133 70351 834189
rect 70419 834133 70475 834189
rect 70047 834009 70103 834065
rect 70171 834009 70227 834065
rect 70295 834009 70351 834065
rect 70419 834009 70475 834065
rect 70047 833885 70103 833941
rect 70171 833885 70227 833941
rect 70295 833885 70351 833941
rect 70419 833885 70475 833941
rect 70047 833761 70103 833817
rect 70171 833761 70227 833817
rect 70295 833761 70351 833817
rect 70419 833761 70475 833817
rect 70047 833637 70103 833693
rect 70171 833637 70227 833693
rect 70295 833637 70351 833693
rect 70419 833637 70475 833693
rect 70047 833513 70103 833569
rect 70171 833513 70227 833569
rect 70295 833513 70351 833569
rect 70419 833513 70475 833569
rect 70047 833389 70103 833445
rect 70171 833389 70227 833445
rect 70295 833389 70351 833445
rect 70419 833389 70475 833445
rect 70047 833265 70103 833321
rect 70171 833265 70227 833321
rect 70295 833265 70351 833321
rect 70419 833265 70475 833321
rect 70047 832755 70103 832811
rect 70171 832755 70227 832811
rect 70295 832755 70351 832811
rect 70419 832755 70475 832811
rect 70047 832631 70103 832687
rect 70171 832631 70227 832687
rect 70295 832631 70351 832687
rect 70419 832631 70475 832687
rect 70047 832507 70103 832563
rect 70171 832507 70227 832563
rect 70295 832507 70351 832563
rect 70419 832507 70475 832563
rect 70047 832383 70103 832439
rect 70171 832383 70227 832439
rect 70295 832383 70351 832439
rect 70419 832383 70475 832439
rect 70047 832259 70103 832315
rect 70171 832259 70227 832315
rect 70295 832259 70351 832315
rect 70419 832259 70475 832315
rect 70047 832135 70103 832191
rect 70171 832135 70227 832191
rect 70295 832135 70351 832191
rect 70419 832135 70475 832191
rect 70047 832011 70103 832067
rect 70171 832011 70227 832067
rect 70295 832011 70351 832067
rect 70419 832011 70475 832067
rect 70047 831887 70103 831943
rect 70171 831887 70227 831943
rect 70295 831887 70351 831943
rect 70419 831887 70475 831943
rect 70047 831763 70103 831819
rect 70171 831763 70227 831819
rect 70295 831763 70351 831819
rect 70419 831763 70475 831819
rect 70047 831639 70103 831695
rect 70171 831639 70227 831695
rect 70295 831639 70351 831695
rect 70419 831639 70475 831695
rect 70047 831515 70103 831571
rect 70171 831515 70227 831571
rect 70295 831515 70351 831571
rect 70419 831515 70475 831571
rect 70047 831391 70103 831447
rect 70171 831391 70227 831447
rect 70295 831391 70351 831447
rect 70419 831391 70475 831447
rect 70047 831267 70103 831323
rect 70171 831267 70227 831323
rect 70295 831267 70351 831323
rect 70419 831267 70475 831323
rect 70047 831143 70103 831199
rect 70171 831143 70227 831199
rect 70295 831143 70351 831199
rect 70419 831143 70475 831199
rect 70047 831019 70103 831075
rect 70171 831019 70227 831075
rect 70295 831019 70351 831075
rect 70419 831019 70475 831075
rect 70047 830895 70103 830951
rect 70171 830895 70227 830951
rect 70295 830895 70351 830951
rect 70419 830895 70475 830951
rect 70047 830049 70103 830105
rect 70171 830049 70227 830105
rect 70295 830049 70351 830105
rect 70419 830049 70475 830105
rect 70047 829925 70103 829981
rect 70171 829925 70227 829981
rect 70295 829925 70351 829981
rect 70419 829925 70475 829981
rect 70047 829801 70103 829857
rect 70171 829801 70227 829857
rect 70295 829801 70351 829857
rect 70419 829801 70475 829857
rect 70047 829677 70103 829733
rect 70171 829677 70227 829733
rect 70295 829677 70351 829733
rect 70419 829677 70475 829733
rect 70047 829553 70103 829609
rect 70171 829553 70227 829609
rect 70295 829553 70351 829609
rect 70419 829553 70475 829609
rect 70047 829429 70103 829485
rect 70171 829429 70227 829485
rect 70295 829429 70351 829485
rect 70419 829429 70475 829485
rect 70047 829305 70103 829361
rect 70171 829305 70227 829361
rect 70295 829305 70351 829361
rect 70419 829305 70475 829361
rect 70047 829181 70103 829237
rect 70171 829181 70227 829237
rect 70295 829181 70351 829237
rect 70419 829181 70475 829237
rect 70047 829057 70103 829113
rect 70171 829057 70227 829113
rect 70295 829057 70351 829113
rect 70419 829057 70475 829113
rect 70047 828933 70103 828989
rect 70171 828933 70227 828989
rect 70295 828933 70351 828989
rect 70419 828933 70475 828989
rect 70047 828809 70103 828865
rect 70171 828809 70227 828865
rect 70295 828809 70351 828865
rect 70419 828809 70475 828865
rect 70047 828685 70103 828741
rect 70171 828685 70227 828741
rect 70295 828685 70351 828741
rect 70419 828685 70475 828741
rect 70047 828561 70103 828617
rect 70171 828561 70227 828617
rect 70295 828561 70351 828617
rect 70419 828561 70475 828617
rect 70047 828437 70103 828493
rect 70171 828437 70227 828493
rect 70295 828437 70351 828493
rect 70419 828437 70475 828493
rect 70047 828313 70103 828369
rect 70171 828313 70227 828369
rect 70295 828313 70351 828369
rect 70419 828313 70475 828369
rect 70047 828189 70103 828245
rect 70171 828189 70227 828245
rect 70295 828189 70351 828245
rect 70419 828189 70475 828245
rect 70047 827679 70103 827735
rect 70171 827679 70227 827735
rect 70295 827679 70351 827735
rect 70419 827679 70475 827735
rect 70047 827555 70103 827611
rect 70171 827555 70227 827611
rect 70295 827555 70351 827611
rect 70419 827555 70475 827611
rect 70047 827431 70103 827487
rect 70171 827431 70227 827487
rect 70295 827431 70351 827487
rect 70419 827431 70475 827487
rect 70047 827307 70103 827363
rect 70171 827307 70227 827363
rect 70295 827307 70351 827363
rect 70419 827307 70475 827363
rect 70047 827183 70103 827239
rect 70171 827183 70227 827239
rect 70295 827183 70351 827239
rect 70419 827183 70475 827239
rect 70047 827059 70103 827115
rect 70171 827059 70227 827115
rect 70295 827059 70351 827115
rect 70419 827059 70475 827115
rect 70047 826935 70103 826991
rect 70171 826935 70227 826991
rect 70295 826935 70351 826991
rect 70419 826935 70475 826991
rect 70047 826811 70103 826867
rect 70171 826811 70227 826867
rect 70295 826811 70351 826867
rect 70419 826811 70475 826867
rect 70047 826687 70103 826743
rect 70171 826687 70227 826743
rect 70295 826687 70351 826743
rect 70419 826687 70475 826743
rect 70047 826563 70103 826619
rect 70171 826563 70227 826619
rect 70295 826563 70351 826619
rect 70419 826563 70475 826619
rect 70047 826439 70103 826495
rect 70171 826439 70227 826495
rect 70295 826439 70351 826495
rect 70419 826439 70475 826495
rect 70047 826315 70103 826371
rect 70171 826315 70227 826371
rect 70295 826315 70351 826371
rect 70419 826315 70475 826371
rect 70047 826191 70103 826247
rect 70171 826191 70227 826247
rect 70295 826191 70351 826247
rect 70419 826191 70475 826247
rect 70047 826067 70103 826123
rect 70171 826067 70227 826123
rect 70295 826067 70351 826123
rect 70419 826067 70475 826123
rect 70047 825943 70103 825999
rect 70171 825943 70227 825999
rect 70295 825943 70351 825999
rect 70419 825943 70475 825999
rect 70047 825819 70103 825875
rect 70171 825819 70227 825875
rect 70295 825819 70351 825875
rect 70419 825819 70475 825875
rect 70047 825049 70103 825105
rect 70171 825049 70227 825105
rect 70295 825049 70351 825105
rect 70419 825049 70475 825105
rect 70047 824925 70103 824981
rect 70171 824925 70227 824981
rect 70295 824925 70351 824981
rect 70419 824925 70475 824981
rect 70047 824801 70103 824857
rect 70171 824801 70227 824857
rect 70295 824801 70351 824857
rect 70419 824801 70475 824857
rect 70047 824677 70103 824733
rect 70171 824677 70227 824733
rect 70295 824677 70351 824733
rect 70419 824677 70475 824733
rect 70047 824553 70103 824609
rect 70171 824553 70227 824609
rect 70295 824553 70351 824609
rect 70419 824553 70475 824609
rect 70047 824429 70103 824485
rect 70171 824429 70227 824485
rect 70295 824429 70351 824485
rect 70419 824429 70475 824485
rect 70047 824305 70103 824361
rect 70171 824305 70227 824361
rect 70295 824305 70351 824361
rect 70419 824305 70475 824361
rect 70047 824181 70103 824237
rect 70171 824181 70227 824237
rect 70295 824181 70351 824237
rect 70419 824181 70475 824237
rect 70047 824057 70103 824113
rect 70171 824057 70227 824113
rect 70295 824057 70351 824113
rect 70419 824057 70475 824113
rect 70047 823933 70103 823989
rect 70171 823933 70227 823989
rect 70295 823933 70351 823989
rect 70419 823933 70475 823989
rect 70047 823809 70103 823865
rect 70171 823809 70227 823865
rect 70295 823809 70351 823865
rect 70419 823809 70475 823865
rect 70047 823685 70103 823741
rect 70171 823685 70227 823741
rect 70295 823685 70351 823741
rect 70419 823685 70475 823741
rect 70047 823561 70103 823617
rect 70171 823561 70227 823617
rect 70295 823561 70351 823617
rect 70419 823561 70475 823617
rect 70047 823437 70103 823493
rect 70171 823437 70227 823493
rect 70295 823437 70351 823493
rect 70419 823437 70475 823493
rect 70047 823313 70103 823369
rect 70171 823313 70227 823369
rect 70295 823313 70351 823369
rect 70419 823313 70475 823369
rect 70047 796605 70103 796661
rect 70171 796605 70227 796661
rect 70295 796605 70351 796661
rect 70419 796605 70475 796661
rect 70047 796481 70103 796537
rect 70171 796481 70227 796537
rect 70295 796481 70351 796537
rect 70419 796481 70475 796537
rect 70047 796357 70103 796413
rect 70171 796357 70227 796413
rect 70295 796357 70351 796413
rect 70419 796357 70475 796413
rect 70047 796233 70103 796289
rect 70171 796233 70227 796289
rect 70295 796233 70351 796289
rect 70419 796233 70475 796289
rect 70047 796109 70103 796165
rect 70171 796109 70227 796165
rect 70295 796109 70351 796165
rect 70419 796109 70475 796165
rect 70047 795985 70103 796041
rect 70171 795985 70227 796041
rect 70295 795985 70351 796041
rect 70419 795985 70475 796041
rect 70047 795861 70103 795917
rect 70171 795861 70227 795917
rect 70295 795861 70351 795917
rect 70419 795861 70475 795917
rect 70047 795737 70103 795793
rect 70171 795737 70227 795793
rect 70295 795737 70351 795793
rect 70419 795737 70475 795793
rect 70047 795613 70103 795669
rect 70171 795613 70227 795669
rect 70295 795613 70351 795669
rect 70419 795613 70475 795669
rect 70047 795489 70103 795545
rect 70171 795489 70227 795545
rect 70295 795489 70351 795545
rect 70419 795489 70475 795545
rect 70047 795365 70103 795421
rect 70171 795365 70227 795421
rect 70295 795365 70351 795421
rect 70419 795365 70475 795421
rect 70047 795241 70103 795297
rect 70171 795241 70227 795297
rect 70295 795241 70351 795297
rect 70419 795241 70475 795297
rect 70047 795117 70103 795173
rect 70171 795117 70227 795173
rect 70295 795117 70351 795173
rect 70419 795117 70475 795173
rect 70047 794993 70103 795049
rect 70171 794993 70227 795049
rect 70295 794993 70351 795049
rect 70419 794993 70475 795049
rect 70047 794869 70103 794925
rect 70171 794869 70227 794925
rect 70295 794869 70351 794925
rect 70419 794869 70475 794925
rect 70047 794125 70103 794181
rect 70171 794125 70227 794181
rect 70295 794125 70351 794181
rect 70419 794125 70475 794181
rect 70047 794001 70103 794057
rect 70171 794001 70227 794057
rect 70295 794001 70351 794057
rect 70419 794001 70475 794057
rect 70047 793877 70103 793933
rect 70171 793877 70227 793933
rect 70295 793877 70351 793933
rect 70419 793877 70475 793933
rect 70047 793753 70103 793809
rect 70171 793753 70227 793809
rect 70295 793753 70351 793809
rect 70419 793753 70475 793809
rect 70047 793629 70103 793685
rect 70171 793629 70227 793685
rect 70295 793629 70351 793685
rect 70419 793629 70475 793685
rect 70047 793505 70103 793561
rect 70171 793505 70227 793561
rect 70295 793505 70351 793561
rect 70419 793505 70475 793561
rect 70047 793381 70103 793437
rect 70171 793381 70227 793437
rect 70295 793381 70351 793437
rect 70419 793381 70475 793437
rect 70047 793257 70103 793313
rect 70171 793257 70227 793313
rect 70295 793257 70351 793313
rect 70419 793257 70475 793313
rect 70047 793133 70103 793189
rect 70171 793133 70227 793189
rect 70295 793133 70351 793189
rect 70419 793133 70475 793189
rect 70047 793009 70103 793065
rect 70171 793009 70227 793065
rect 70295 793009 70351 793065
rect 70419 793009 70475 793065
rect 70047 792885 70103 792941
rect 70171 792885 70227 792941
rect 70295 792885 70351 792941
rect 70419 792885 70475 792941
rect 70047 792761 70103 792817
rect 70171 792761 70227 792817
rect 70295 792761 70351 792817
rect 70419 792761 70475 792817
rect 70047 792637 70103 792693
rect 70171 792637 70227 792693
rect 70295 792637 70351 792693
rect 70419 792637 70475 792693
rect 70047 792513 70103 792569
rect 70171 792513 70227 792569
rect 70295 792513 70351 792569
rect 70419 792513 70475 792569
rect 70047 792389 70103 792445
rect 70171 792389 70227 792445
rect 70295 792389 70351 792445
rect 70419 792389 70475 792445
rect 70047 792265 70103 792321
rect 70171 792265 70227 792321
rect 70295 792265 70351 792321
rect 70419 792265 70475 792321
rect 70047 791755 70103 791811
rect 70171 791755 70227 791811
rect 70295 791755 70351 791811
rect 70419 791755 70475 791811
rect 70047 791631 70103 791687
rect 70171 791631 70227 791687
rect 70295 791631 70351 791687
rect 70419 791631 70475 791687
rect 70047 791507 70103 791563
rect 70171 791507 70227 791563
rect 70295 791507 70351 791563
rect 70419 791507 70475 791563
rect 70047 791383 70103 791439
rect 70171 791383 70227 791439
rect 70295 791383 70351 791439
rect 70419 791383 70475 791439
rect 70047 791259 70103 791315
rect 70171 791259 70227 791315
rect 70295 791259 70351 791315
rect 70419 791259 70475 791315
rect 70047 791135 70103 791191
rect 70171 791135 70227 791191
rect 70295 791135 70351 791191
rect 70419 791135 70475 791191
rect 70047 791011 70103 791067
rect 70171 791011 70227 791067
rect 70295 791011 70351 791067
rect 70419 791011 70475 791067
rect 70047 790887 70103 790943
rect 70171 790887 70227 790943
rect 70295 790887 70351 790943
rect 70419 790887 70475 790943
rect 70047 790763 70103 790819
rect 70171 790763 70227 790819
rect 70295 790763 70351 790819
rect 70419 790763 70475 790819
rect 70047 790639 70103 790695
rect 70171 790639 70227 790695
rect 70295 790639 70351 790695
rect 70419 790639 70475 790695
rect 70047 790515 70103 790571
rect 70171 790515 70227 790571
rect 70295 790515 70351 790571
rect 70419 790515 70475 790571
rect 70047 790391 70103 790447
rect 70171 790391 70227 790447
rect 70295 790391 70351 790447
rect 70419 790391 70475 790447
rect 70047 790267 70103 790323
rect 70171 790267 70227 790323
rect 70295 790267 70351 790323
rect 70419 790267 70475 790323
rect 70047 790143 70103 790199
rect 70171 790143 70227 790199
rect 70295 790143 70351 790199
rect 70419 790143 70475 790199
rect 70047 790019 70103 790075
rect 70171 790019 70227 790075
rect 70295 790019 70351 790075
rect 70419 790019 70475 790075
rect 70047 789895 70103 789951
rect 70171 789895 70227 789951
rect 70295 789895 70351 789951
rect 70419 789895 70475 789951
rect 705525 791631 705581 791687
rect 705649 791631 705705 791687
rect 705773 791631 705829 791687
rect 705897 791631 705953 791687
rect 705525 791507 705581 791563
rect 705649 791507 705705 791563
rect 705773 791507 705829 791563
rect 705897 791507 705953 791563
rect 705525 791383 705581 791439
rect 705649 791383 705705 791439
rect 705773 791383 705829 791439
rect 705897 791383 705953 791439
rect 705525 791259 705581 791315
rect 705649 791259 705705 791315
rect 705773 791259 705829 791315
rect 705897 791259 705953 791315
rect 705525 791135 705581 791191
rect 705649 791135 705705 791191
rect 705773 791135 705829 791191
rect 705897 791135 705953 791191
rect 705525 791011 705581 791067
rect 705649 791011 705705 791067
rect 705773 791011 705829 791067
rect 705897 791011 705953 791067
rect 705525 790887 705581 790943
rect 705649 790887 705705 790943
rect 705773 790887 705829 790943
rect 705897 790887 705953 790943
rect 705525 790763 705581 790819
rect 705649 790763 705705 790819
rect 705773 790763 705829 790819
rect 705897 790763 705953 790819
rect 705525 790639 705581 790695
rect 705649 790639 705705 790695
rect 705773 790639 705829 790695
rect 705897 790639 705953 790695
rect 705525 790515 705581 790571
rect 705649 790515 705705 790571
rect 705773 790515 705829 790571
rect 705897 790515 705953 790571
rect 705525 790391 705581 790447
rect 705649 790391 705705 790447
rect 705773 790391 705829 790447
rect 705897 790391 705953 790447
rect 705525 790267 705581 790323
rect 705649 790267 705705 790323
rect 705773 790267 705829 790323
rect 705897 790267 705953 790323
rect 705525 790143 705581 790199
rect 705649 790143 705705 790199
rect 705773 790143 705829 790199
rect 705897 790143 705953 790199
rect 705525 790019 705581 790075
rect 705649 790019 705705 790075
rect 705773 790019 705829 790075
rect 705897 790019 705953 790075
rect 705525 789895 705581 789951
rect 705649 789895 705705 789951
rect 705773 789895 705829 789951
rect 705897 789895 705953 789951
rect 70047 789049 70103 789105
rect 70171 789049 70227 789105
rect 70295 789049 70351 789105
rect 70419 789049 70475 789105
rect 70047 788925 70103 788981
rect 70171 788925 70227 788981
rect 70295 788925 70351 788981
rect 70419 788925 70475 788981
rect 70047 788801 70103 788857
rect 70171 788801 70227 788857
rect 70295 788801 70351 788857
rect 70419 788801 70475 788857
rect 70047 788677 70103 788733
rect 70171 788677 70227 788733
rect 70295 788677 70351 788733
rect 70419 788677 70475 788733
rect 70047 788553 70103 788609
rect 70171 788553 70227 788609
rect 70295 788553 70351 788609
rect 70419 788553 70475 788609
rect 70047 788429 70103 788485
rect 70171 788429 70227 788485
rect 70295 788429 70351 788485
rect 70419 788429 70475 788485
rect 70047 788305 70103 788361
rect 70171 788305 70227 788361
rect 70295 788305 70351 788361
rect 70419 788305 70475 788361
rect 70047 788181 70103 788237
rect 70171 788181 70227 788237
rect 70295 788181 70351 788237
rect 70419 788181 70475 788237
rect 70047 788057 70103 788113
rect 70171 788057 70227 788113
rect 70295 788057 70351 788113
rect 70419 788057 70475 788113
rect 70047 787933 70103 787989
rect 70171 787933 70227 787989
rect 70295 787933 70351 787989
rect 70419 787933 70475 787989
rect 70047 787809 70103 787865
rect 70171 787809 70227 787865
rect 70295 787809 70351 787865
rect 70419 787809 70475 787865
rect 70047 787685 70103 787741
rect 70171 787685 70227 787741
rect 70295 787685 70351 787741
rect 70419 787685 70475 787741
rect 70047 787561 70103 787617
rect 70171 787561 70227 787617
rect 70295 787561 70351 787617
rect 70419 787561 70475 787617
rect 70047 787437 70103 787493
rect 70171 787437 70227 787493
rect 70295 787437 70351 787493
rect 70419 787437 70475 787493
rect 70047 787313 70103 787369
rect 70171 787313 70227 787369
rect 70295 787313 70351 787369
rect 70419 787313 70475 787369
rect 70047 787189 70103 787245
rect 70171 787189 70227 787245
rect 70295 787189 70351 787245
rect 70419 787189 70475 787245
rect 705525 789125 705581 789181
rect 705649 789125 705705 789181
rect 705773 789125 705829 789181
rect 705897 789125 705953 789181
rect 705525 789001 705581 789057
rect 705649 789001 705705 789057
rect 705773 789001 705829 789057
rect 705897 789001 705953 789057
rect 705525 788877 705581 788933
rect 705649 788877 705705 788933
rect 705773 788877 705829 788933
rect 705897 788877 705953 788933
rect 705525 788753 705581 788809
rect 705649 788753 705705 788809
rect 705773 788753 705829 788809
rect 705897 788753 705953 788809
rect 705525 788629 705581 788685
rect 705649 788629 705705 788685
rect 705773 788629 705829 788685
rect 705897 788629 705953 788685
rect 705525 788505 705581 788561
rect 705649 788505 705705 788561
rect 705773 788505 705829 788561
rect 705897 788505 705953 788561
rect 705525 788381 705581 788437
rect 705649 788381 705705 788437
rect 705773 788381 705829 788437
rect 705897 788381 705953 788437
rect 705525 788257 705581 788313
rect 705649 788257 705705 788313
rect 705773 788257 705829 788313
rect 705897 788257 705953 788313
rect 705525 788133 705581 788189
rect 705649 788133 705705 788189
rect 705773 788133 705829 788189
rect 705897 788133 705953 788189
rect 705525 788009 705581 788065
rect 705649 788009 705705 788065
rect 705773 788009 705829 788065
rect 705897 788009 705953 788065
rect 705525 787885 705581 787941
rect 705649 787885 705705 787941
rect 705773 787885 705829 787941
rect 705897 787885 705953 787941
rect 705525 787761 705581 787817
rect 705649 787761 705705 787817
rect 705773 787761 705829 787817
rect 705897 787761 705953 787817
rect 705525 787637 705581 787693
rect 705649 787637 705705 787693
rect 705773 787637 705829 787693
rect 705897 787637 705953 787693
rect 705525 787513 705581 787569
rect 705649 787513 705705 787569
rect 705773 787513 705829 787569
rect 705897 787513 705953 787569
rect 705525 787389 705581 787445
rect 705649 787389 705705 787445
rect 705773 787389 705829 787445
rect 705897 787389 705953 787445
rect 705525 787265 705581 787321
rect 705649 787265 705705 787321
rect 705773 787265 705829 787321
rect 705897 787265 705953 787321
rect 70047 786679 70103 786735
rect 70171 786679 70227 786735
rect 70295 786679 70351 786735
rect 70419 786679 70475 786735
rect 70047 786555 70103 786611
rect 70171 786555 70227 786611
rect 70295 786555 70351 786611
rect 70419 786555 70475 786611
rect 70047 786431 70103 786487
rect 70171 786431 70227 786487
rect 70295 786431 70351 786487
rect 70419 786431 70475 786487
rect 70047 786307 70103 786363
rect 70171 786307 70227 786363
rect 70295 786307 70351 786363
rect 70419 786307 70475 786363
rect 70047 786183 70103 786239
rect 70171 786183 70227 786239
rect 70295 786183 70351 786239
rect 70419 786183 70475 786239
rect 70047 786059 70103 786115
rect 70171 786059 70227 786115
rect 70295 786059 70351 786115
rect 70419 786059 70475 786115
rect 70047 785935 70103 785991
rect 70171 785935 70227 785991
rect 70295 785935 70351 785991
rect 70419 785935 70475 785991
rect 70047 785811 70103 785867
rect 70171 785811 70227 785867
rect 70295 785811 70351 785867
rect 70419 785811 70475 785867
rect 70047 785687 70103 785743
rect 70171 785687 70227 785743
rect 70295 785687 70351 785743
rect 70419 785687 70475 785743
rect 70047 785563 70103 785619
rect 70171 785563 70227 785619
rect 70295 785563 70351 785619
rect 70419 785563 70475 785619
rect 70047 785439 70103 785495
rect 70171 785439 70227 785495
rect 70295 785439 70351 785495
rect 70419 785439 70475 785495
rect 70047 785315 70103 785371
rect 70171 785315 70227 785371
rect 70295 785315 70351 785371
rect 70419 785315 70475 785371
rect 70047 785191 70103 785247
rect 70171 785191 70227 785247
rect 70295 785191 70351 785247
rect 70419 785191 70475 785247
rect 70047 785067 70103 785123
rect 70171 785067 70227 785123
rect 70295 785067 70351 785123
rect 70419 785067 70475 785123
rect 70047 784943 70103 784999
rect 70171 784943 70227 784999
rect 70295 784943 70351 784999
rect 70419 784943 70475 784999
rect 70047 784819 70103 784875
rect 70171 784819 70227 784875
rect 70295 784819 70351 784875
rect 70419 784819 70475 784875
rect 705525 786755 705581 786811
rect 705649 786755 705705 786811
rect 705773 786755 705829 786811
rect 705897 786755 705953 786811
rect 705525 786631 705581 786687
rect 705649 786631 705705 786687
rect 705773 786631 705829 786687
rect 705897 786631 705953 786687
rect 705525 786507 705581 786563
rect 705649 786507 705705 786563
rect 705773 786507 705829 786563
rect 705897 786507 705953 786563
rect 705525 786383 705581 786439
rect 705649 786383 705705 786439
rect 705773 786383 705829 786439
rect 705897 786383 705953 786439
rect 705525 786259 705581 786315
rect 705649 786259 705705 786315
rect 705773 786259 705829 786315
rect 705897 786259 705953 786315
rect 705525 786135 705581 786191
rect 705649 786135 705705 786191
rect 705773 786135 705829 786191
rect 705897 786135 705953 786191
rect 705525 786011 705581 786067
rect 705649 786011 705705 786067
rect 705773 786011 705829 786067
rect 705897 786011 705953 786067
rect 705525 785887 705581 785943
rect 705649 785887 705705 785943
rect 705773 785887 705829 785943
rect 705897 785887 705953 785943
rect 705525 785763 705581 785819
rect 705649 785763 705705 785819
rect 705773 785763 705829 785819
rect 705897 785763 705953 785819
rect 705525 785639 705581 785695
rect 705649 785639 705705 785695
rect 705773 785639 705829 785695
rect 705897 785639 705953 785695
rect 705525 785515 705581 785571
rect 705649 785515 705705 785571
rect 705773 785515 705829 785571
rect 705897 785515 705953 785571
rect 705525 785391 705581 785447
rect 705649 785391 705705 785447
rect 705773 785391 705829 785447
rect 705897 785391 705953 785447
rect 705525 785267 705581 785323
rect 705649 785267 705705 785323
rect 705773 785267 705829 785323
rect 705897 785267 705953 785323
rect 705525 785143 705581 785199
rect 705649 785143 705705 785199
rect 705773 785143 705829 785199
rect 705897 785143 705953 785199
rect 705525 785019 705581 785075
rect 705649 785019 705705 785075
rect 705773 785019 705829 785075
rect 705897 785019 705953 785075
rect 705525 784895 705581 784951
rect 705649 784895 705705 784951
rect 705773 784895 705829 784951
rect 705897 784895 705953 784951
rect 70047 784049 70103 784105
rect 70171 784049 70227 784105
rect 70295 784049 70351 784105
rect 70419 784049 70475 784105
rect 70047 783925 70103 783981
rect 70171 783925 70227 783981
rect 70295 783925 70351 783981
rect 70419 783925 70475 783981
rect 70047 783801 70103 783857
rect 70171 783801 70227 783857
rect 70295 783801 70351 783857
rect 70419 783801 70475 783857
rect 70047 783677 70103 783733
rect 70171 783677 70227 783733
rect 70295 783677 70351 783733
rect 70419 783677 70475 783733
rect 70047 783553 70103 783609
rect 70171 783553 70227 783609
rect 70295 783553 70351 783609
rect 70419 783553 70475 783609
rect 70047 783429 70103 783485
rect 70171 783429 70227 783485
rect 70295 783429 70351 783485
rect 70419 783429 70475 783485
rect 70047 783305 70103 783361
rect 70171 783305 70227 783361
rect 70295 783305 70351 783361
rect 70419 783305 70475 783361
rect 70047 783181 70103 783237
rect 70171 783181 70227 783237
rect 70295 783181 70351 783237
rect 70419 783181 70475 783237
rect 70047 783057 70103 783113
rect 70171 783057 70227 783113
rect 70295 783057 70351 783113
rect 70419 783057 70475 783113
rect 70047 782933 70103 782989
rect 70171 782933 70227 782989
rect 70295 782933 70351 782989
rect 70419 782933 70475 782989
rect 70047 782809 70103 782865
rect 70171 782809 70227 782865
rect 70295 782809 70351 782865
rect 70419 782809 70475 782865
rect 70047 782685 70103 782741
rect 70171 782685 70227 782741
rect 70295 782685 70351 782741
rect 70419 782685 70475 782741
rect 70047 782561 70103 782617
rect 70171 782561 70227 782617
rect 70295 782561 70351 782617
rect 70419 782561 70475 782617
rect 70047 782437 70103 782493
rect 70171 782437 70227 782493
rect 70295 782437 70351 782493
rect 70419 782437 70475 782493
rect 70047 782313 70103 782369
rect 70171 782313 70227 782369
rect 70295 782313 70351 782369
rect 70419 782313 70475 782369
rect 705525 784049 705581 784105
rect 705649 784049 705705 784105
rect 705773 784049 705829 784105
rect 705897 784049 705953 784105
rect 705525 783925 705581 783981
rect 705649 783925 705705 783981
rect 705773 783925 705829 783981
rect 705897 783925 705953 783981
rect 705525 783801 705581 783857
rect 705649 783801 705705 783857
rect 705773 783801 705829 783857
rect 705897 783801 705953 783857
rect 705525 783677 705581 783733
rect 705649 783677 705705 783733
rect 705773 783677 705829 783733
rect 705897 783677 705953 783733
rect 705525 783553 705581 783609
rect 705649 783553 705705 783609
rect 705773 783553 705829 783609
rect 705897 783553 705953 783609
rect 705525 783429 705581 783485
rect 705649 783429 705705 783485
rect 705773 783429 705829 783485
rect 705897 783429 705953 783485
rect 705525 783305 705581 783361
rect 705649 783305 705705 783361
rect 705773 783305 705829 783361
rect 705897 783305 705953 783361
rect 705525 783181 705581 783237
rect 705649 783181 705705 783237
rect 705773 783181 705829 783237
rect 705897 783181 705953 783237
rect 705525 783057 705581 783113
rect 705649 783057 705705 783113
rect 705773 783057 705829 783113
rect 705897 783057 705953 783113
rect 705525 782933 705581 782989
rect 705649 782933 705705 782989
rect 705773 782933 705829 782989
rect 705897 782933 705953 782989
rect 705525 782809 705581 782865
rect 705649 782809 705705 782865
rect 705773 782809 705829 782865
rect 705897 782809 705953 782865
rect 705525 782685 705581 782741
rect 705649 782685 705705 782741
rect 705773 782685 705829 782741
rect 705897 782685 705953 782741
rect 705525 782561 705581 782617
rect 705649 782561 705705 782617
rect 705773 782561 705829 782617
rect 705897 782561 705953 782617
rect 705525 782437 705581 782493
rect 705649 782437 705705 782493
rect 705773 782437 705829 782493
rect 705897 782437 705953 782493
rect 705525 782313 705581 782369
rect 705649 782313 705705 782369
rect 705773 782313 705829 782369
rect 705897 782313 705953 782369
rect 705525 782189 705581 782245
rect 705649 782189 705705 782245
rect 705773 782189 705829 782245
rect 705897 782189 705953 782245
rect 705525 781679 705581 781735
rect 705649 781679 705705 781735
rect 705773 781679 705829 781735
rect 705897 781679 705953 781735
rect 705525 781555 705581 781611
rect 705649 781555 705705 781611
rect 705773 781555 705829 781611
rect 705897 781555 705953 781611
rect 705525 781431 705581 781487
rect 705649 781431 705705 781487
rect 705773 781431 705829 781487
rect 705897 781431 705953 781487
rect 705525 781307 705581 781363
rect 705649 781307 705705 781363
rect 705773 781307 705829 781363
rect 705897 781307 705953 781363
rect 705525 781183 705581 781239
rect 705649 781183 705705 781239
rect 705773 781183 705829 781239
rect 705897 781183 705953 781239
rect 705525 781059 705581 781115
rect 705649 781059 705705 781115
rect 705773 781059 705829 781115
rect 705897 781059 705953 781115
rect 705525 780935 705581 780991
rect 705649 780935 705705 780991
rect 705773 780935 705829 780991
rect 705897 780935 705953 780991
rect 705525 780811 705581 780867
rect 705649 780811 705705 780867
rect 705773 780811 705829 780867
rect 705897 780811 705953 780867
rect 705525 780687 705581 780743
rect 705649 780687 705705 780743
rect 705773 780687 705829 780743
rect 705897 780687 705953 780743
rect 705525 780563 705581 780619
rect 705649 780563 705705 780619
rect 705773 780563 705829 780619
rect 705897 780563 705953 780619
rect 705525 780439 705581 780495
rect 705649 780439 705705 780495
rect 705773 780439 705829 780495
rect 705897 780439 705953 780495
rect 705525 780315 705581 780371
rect 705649 780315 705705 780371
rect 705773 780315 705829 780371
rect 705897 780315 705953 780371
rect 705525 780191 705581 780247
rect 705649 780191 705705 780247
rect 705773 780191 705829 780247
rect 705897 780191 705953 780247
rect 705525 780067 705581 780123
rect 705649 780067 705705 780123
rect 705773 780067 705829 780123
rect 705897 780067 705953 780123
rect 705525 779943 705581 779999
rect 705649 779943 705705 779999
rect 705773 779943 705829 779999
rect 705897 779943 705953 779999
rect 705525 779819 705581 779875
rect 705649 779819 705705 779875
rect 705773 779819 705829 779875
rect 705897 779819 705953 779875
rect 705525 779075 705581 779131
rect 705649 779075 705705 779131
rect 705773 779075 705829 779131
rect 705897 779075 705953 779131
rect 705525 778951 705581 779007
rect 705649 778951 705705 779007
rect 705773 778951 705829 779007
rect 705897 778951 705953 779007
rect 705525 778827 705581 778883
rect 705649 778827 705705 778883
rect 705773 778827 705829 778883
rect 705897 778827 705953 778883
rect 705525 778703 705581 778759
rect 705649 778703 705705 778759
rect 705773 778703 705829 778759
rect 705897 778703 705953 778759
rect 705525 778579 705581 778635
rect 705649 778579 705705 778635
rect 705773 778579 705829 778635
rect 705897 778579 705953 778635
rect 705525 778455 705581 778511
rect 705649 778455 705705 778511
rect 705773 778455 705829 778511
rect 705897 778455 705953 778511
rect 705525 778331 705581 778387
rect 705649 778331 705705 778387
rect 705773 778331 705829 778387
rect 705897 778331 705953 778387
rect 705525 778207 705581 778263
rect 705649 778207 705705 778263
rect 705773 778207 705829 778263
rect 705897 778207 705953 778263
rect 705525 778083 705581 778139
rect 705649 778083 705705 778139
rect 705773 778083 705829 778139
rect 705897 778083 705953 778139
rect 705525 777959 705581 778015
rect 705649 777959 705705 778015
rect 705773 777959 705829 778015
rect 705897 777959 705953 778015
rect 705525 777835 705581 777891
rect 705649 777835 705705 777891
rect 705773 777835 705829 777891
rect 705897 777835 705953 777891
rect 705525 777711 705581 777767
rect 705649 777711 705705 777767
rect 705773 777711 705829 777767
rect 705897 777711 705953 777767
rect 705525 777587 705581 777643
rect 705649 777587 705705 777643
rect 705773 777587 705829 777643
rect 705897 777587 705953 777643
rect 705525 777463 705581 777519
rect 705649 777463 705705 777519
rect 705773 777463 705829 777519
rect 705897 777463 705953 777519
rect 705525 777339 705581 777395
rect 705649 777339 705705 777395
rect 705773 777339 705829 777395
rect 705897 777339 705953 777395
rect 705525 490631 705581 490687
rect 705649 490631 705705 490687
rect 705773 490631 705829 490687
rect 705897 490631 705953 490687
rect 705525 490507 705581 490563
rect 705649 490507 705705 490563
rect 705773 490507 705829 490563
rect 705897 490507 705953 490563
rect 705525 490383 705581 490439
rect 705649 490383 705705 490439
rect 705773 490383 705829 490439
rect 705897 490383 705953 490439
rect 705525 490259 705581 490315
rect 705649 490259 705705 490315
rect 705773 490259 705829 490315
rect 705897 490259 705953 490315
rect 705525 490135 705581 490191
rect 705649 490135 705705 490191
rect 705773 490135 705829 490191
rect 705897 490135 705953 490191
rect 705525 490011 705581 490067
rect 705649 490011 705705 490067
rect 705773 490011 705829 490067
rect 705897 490011 705953 490067
rect 705525 489887 705581 489943
rect 705649 489887 705705 489943
rect 705773 489887 705829 489943
rect 705897 489887 705953 489943
rect 705525 489763 705581 489819
rect 705649 489763 705705 489819
rect 705773 489763 705829 489819
rect 705897 489763 705953 489819
rect 705525 489639 705581 489695
rect 705649 489639 705705 489695
rect 705773 489639 705829 489695
rect 705897 489639 705953 489695
rect 705525 489515 705581 489571
rect 705649 489515 705705 489571
rect 705773 489515 705829 489571
rect 705897 489515 705953 489571
rect 705525 489391 705581 489447
rect 705649 489391 705705 489447
rect 705773 489391 705829 489447
rect 705897 489391 705953 489447
rect 705525 489267 705581 489323
rect 705649 489267 705705 489323
rect 705773 489267 705829 489323
rect 705897 489267 705953 489323
rect 705525 489143 705581 489199
rect 705649 489143 705705 489199
rect 705773 489143 705829 489199
rect 705897 489143 705953 489199
rect 705525 489019 705581 489075
rect 705649 489019 705705 489075
rect 705773 489019 705829 489075
rect 705897 489019 705953 489075
rect 705525 488895 705581 488951
rect 705649 488895 705705 488951
rect 705773 488895 705829 488951
rect 705897 488895 705953 488951
rect 705525 488125 705581 488181
rect 705649 488125 705705 488181
rect 705773 488125 705829 488181
rect 705897 488125 705953 488181
rect 705525 488001 705581 488057
rect 705649 488001 705705 488057
rect 705773 488001 705829 488057
rect 705897 488001 705953 488057
rect 705525 487877 705581 487933
rect 705649 487877 705705 487933
rect 705773 487877 705829 487933
rect 705897 487877 705953 487933
rect 705525 487753 705581 487809
rect 705649 487753 705705 487809
rect 705773 487753 705829 487809
rect 705897 487753 705953 487809
rect 705525 487629 705581 487685
rect 705649 487629 705705 487685
rect 705773 487629 705829 487685
rect 705897 487629 705953 487685
rect 705525 487505 705581 487561
rect 705649 487505 705705 487561
rect 705773 487505 705829 487561
rect 705897 487505 705953 487561
rect 705525 487381 705581 487437
rect 705649 487381 705705 487437
rect 705773 487381 705829 487437
rect 705897 487381 705953 487437
rect 705525 487257 705581 487313
rect 705649 487257 705705 487313
rect 705773 487257 705829 487313
rect 705897 487257 705953 487313
rect 705525 487133 705581 487189
rect 705649 487133 705705 487189
rect 705773 487133 705829 487189
rect 705897 487133 705953 487189
rect 705525 487009 705581 487065
rect 705649 487009 705705 487065
rect 705773 487009 705829 487065
rect 705897 487009 705953 487065
rect 705525 486885 705581 486941
rect 705649 486885 705705 486941
rect 705773 486885 705829 486941
rect 705897 486885 705953 486941
rect 705525 486761 705581 486817
rect 705649 486761 705705 486817
rect 705773 486761 705829 486817
rect 705897 486761 705953 486817
rect 705525 486637 705581 486693
rect 705649 486637 705705 486693
rect 705773 486637 705829 486693
rect 705897 486637 705953 486693
rect 705525 486513 705581 486569
rect 705649 486513 705705 486569
rect 705773 486513 705829 486569
rect 705897 486513 705953 486569
rect 705525 486389 705581 486445
rect 705649 486389 705705 486445
rect 705773 486389 705829 486445
rect 705897 486389 705953 486445
rect 705525 486265 705581 486321
rect 705649 486265 705705 486321
rect 705773 486265 705829 486321
rect 705897 486265 705953 486321
rect 705525 485755 705581 485811
rect 705649 485755 705705 485811
rect 705773 485755 705829 485811
rect 705897 485755 705953 485811
rect 705525 485631 705581 485687
rect 705649 485631 705705 485687
rect 705773 485631 705829 485687
rect 705897 485631 705953 485687
rect 705525 485507 705581 485563
rect 705649 485507 705705 485563
rect 705773 485507 705829 485563
rect 705897 485507 705953 485563
rect 705525 485383 705581 485439
rect 705649 485383 705705 485439
rect 705773 485383 705829 485439
rect 705897 485383 705953 485439
rect 705525 485259 705581 485315
rect 705649 485259 705705 485315
rect 705773 485259 705829 485315
rect 705897 485259 705953 485315
rect 705525 485135 705581 485191
rect 705649 485135 705705 485191
rect 705773 485135 705829 485191
rect 705897 485135 705953 485191
rect 705525 485011 705581 485067
rect 705649 485011 705705 485067
rect 705773 485011 705829 485067
rect 705897 485011 705953 485067
rect 705525 484887 705581 484943
rect 705649 484887 705705 484943
rect 705773 484887 705829 484943
rect 705897 484887 705953 484943
rect 705525 484763 705581 484819
rect 705649 484763 705705 484819
rect 705773 484763 705829 484819
rect 705897 484763 705953 484819
rect 705525 484639 705581 484695
rect 705649 484639 705705 484695
rect 705773 484639 705829 484695
rect 705897 484639 705953 484695
rect 705525 484515 705581 484571
rect 705649 484515 705705 484571
rect 705773 484515 705829 484571
rect 705897 484515 705953 484571
rect 705525 484391 705581 484447
rect 705649 484391 705705 484447
rect 705773 484391 705829 484447
rect 705897 484391 705953 484447
rect 705525 484267 705581 484323
rect 705649 484267 705705 484323
rect 705773 484267 705829 484323
rect 705897 484267 705953 484323
rect 705525 484143 705581 484199
rect 705649 484143 705705 484199
rect 705773 484143 705829 484199
rect 705897 484143 705953 484199
rect 705525 484019 705581 484075
rect 705649 484019 705705 484075
rect 705773 484019 705829 484075
rect 705897 484019 705953 484075
rect 705525 483895 705581 483951
rect 705649 483895 705705 483951
rect 705773 483895 705829 483951
rect 705897 483895 705953 483951
rect 705525 483049 705581 483105
rect 705649 483049 705705 483105
rect 705773 483049 705829 483105
rect 705897 483049 705953 483105
rect 705525 482925 705581 482981
rect 705649 482925 705705 482981
rect 705773 482925 705829 482981
rect 705897 482925 705953 482981
rect 705525 482801 705581 482857
rect 705649 482801 705705 482857
rect 705773 482801 705829 482857
rect 705897 482801 705953 482857
rect 705525 482677 705581 482733
rect 705649 482677 705705 482733
rect 705773 482677 705829 482733
rect 705897 482677 705953 482733
rect 705525 482553 705581 482609
rect 705649 482553 705705 482609
rect 705773 482553 705829 482609
rect 705897 482553 705953 482609
rect 705525 482429 705581 482485
rect 705649 482429 705705 482485
rect 705773 482429 705829 482485
rect 705897 482429 705953 482485
rect 705525 482305 705581 482361
rect 705649 482305 705705 482361
rect 705773 482305 705829 482361
rect 705897 482305 705953 482361
rect 705525 482181 705581 482237
rect 705649 482181 705705 482237
rect 705773 482181 705829 482237
rect 705897 482181 705953 482237
rect 705525 482057 705581 482113
rect 705649 482057 705705 482113
rect 705773 482057 705829 482113
rect 705897 482057 705953 482113
rect 705525 481933 705581 481989
rect 705649 481933 705705 481989
rect 705773 481933 705829 481989
rect 705897 481933 705953 481989
rect 705525 481809 705581 481865
rect 705649 481809 705705 481865
rect 705773 481809 705829 481865
rect 705897 481809 705953 481865
rect 705525 481685 705581 481741
rect 705649 481685 705705 481741
rect 705773 481685 705829 481741
rect 705897 481685 705953 481741
rect 705525 481561 705581 481617
rect 705649 481561 705705 481617
rect 705773 481561 705829 481617
rect 705897 481561 705953 481617
rect 705525 481437 705581 481493
rect 705649 481437 705705 481493
rect 705773 481437 705829 481493
rect 705897 481437 705953 481493
rect 705525 481313 705581 481369
rect 705649 481313 705705 481369
rect 705773 481313 705829 481369
rect 705897 481313 705953 481369
rect 705525 481189 705581 481245
rect 705649 481189 705705 481245
rect 705773 481189 705829 481245
rect 705897 481189 705953 481245
rect 705525 480679 705581 480735
rect 705649 480679 705705 480735
rect 705773 480679 705829 480735
rect 705897 480679 705953 480735
rect 705525 480555 705581 480611
rect 705649 480555 705705 480611
rect 705773 480555 705829 480611
rect 705897 480555 705953 480611
rect 705525 480431 705581 480487
rect 705649 480431 705705 480487
rect 705773 480431 705829 480487
rect 705897 480431 705953 480487
rect 705525 480307 705581 480363
rect 705649 480307 705705 480363
rect 705773 480307 705829 480363
rect 705897 480307 705953 480363
rect 705525 480183 705581 480239
rect 705649 480183 705705 480239
rect 705773 480183 705829 480239
rect 705897 480183 705953 480239
rect 705525 480059 705581 480115
rect 705649 480059 705705 480115
rect 705773 480059 705829 480115
rect 705897 480059 705953 480115
rect 705525 479935 705581 479991
rect 705649 479935 705705 479991
rect 705773 479935 705829 479991
rect 705897 479935 705953 479991
rect 705525 479811 705581 479867
rect 705649 479811 705705 479867
rect 705773 479811 705829 479867
rect 705897 479811 705953 479867
rect 705525 479687 705581 479743
rect 705649 479687 705705 479743
rect 705773 479687 705829 479743
rect 705897 479687 705953 479743
rect 705525 479563 705581 479619
rect 705649 479563 705705 479619
rect 705773 479563 705829 479619
rect 705897 479563 705953 479619
rect 705525 479439 705581 479495
rect 705649 479439 705705 479495
rect 705773 479439 705829 479495
rect 705897 479439 705953 479495
rect 705525 479315 705581 479371
rect 705649 479315 705705 479371
rect 705773 479315 705829 479371
rect 705897 479315 705953 479371
rect 705525 479191 705581 479247
rect 705649 479191 705705 479247
rect 705773 479191 705829 479247
rect 705897 479191 705953 479247
rect 705525 479067 705581 479123
rect 705649 479067 705705 479123
rect 705773 479067 705829 479123
rect 705897 479067 705953 479123
rect 705525 478943 705581 478999
rect 705649 478943 705705 478999
rect 705773 478943 705829 478999
rect 705897 478943 705953 478999
rect 705525 478819 705581 478875
rect 705649 478819 705705 478875
rect 705773 478819 705829 478875
rect 705897 478819 705953 478875
rect 705525 478075 705581 478131
rect 705649 478075 705705 478131
rect 705773 478075 705829 478131
rect 705897 478075 705953 478131
rect 705525 477951 705581 478007
rect 705649 477951 705705 478007
rect 705773 477951 705829 478007
rect 705897 477951 705953 478007
rect 705525 477827 705581 477883
rect 705649 477827 705705 477883
rect 705773 477827 705829 477883
rect 705897 477827 705953 477883
rect 705525 477703 705581 477759
rect 705649 477703 705705 477759
rect 705773 477703 705829 477759
rect 705897 477703 705953 477759
rect 705525 477579 705581 477635
rect 705649 477579 705705 477635
rect 705773 477579 705829 477635
rect 705897 477579 705953 477635
rect 705525 477455 705581 477511
rect 705649 477455 705705 477511
rect 705773 477455 705829 477511
rect 705897 477455 705953 477511
rect 705525 477331 705581 477387
rect 705649 477331 705705 477387
rect 705773 477331 705829 477387
rect 705897 477331 705953 477387
rect 705525 477207 705581 477263
rect 705649 477207 705705 477263
rect 705773 477207 705829 477263
rect 705897 477207 705953 477263
rect 705525 477083 705581 477139
rect 705649 477083 705705 477139
rect 705773 477083 705829 477139
rect 705897 477083 705953 477139
rect 705525 476959 705581 477015
rect 705649 476959 705705 477015
rect 705773 476959 705829 477015
rect 705897 476959 705953 477015
rect 705525 476835 705581 476891
rect 705649 476835 705705 476891
rect 705773 476835 705829 476891
rect 705897 476835 705953 476891
rect 705525 476711 705581 476767
rect 705649 476711 705705 476767
rect 705773 476711 705829 476767
rect 705897 476711 705953 476767
rect 705525 476587 705581 476643
rect 705649 476587 705705 476643
rect 705773 476587 705829 476643
rect 705897 476587 705953 476643
rect 705525 476463 705581 476519
rect 705649 476463 705705 476519
rect 705773 476463 705829 476519
rect 705897 476463 705953 476519
rect 705525 476339 705581 476395
rect 705649 476339 705705 476395
rect 705773 476339 705829 476395
rect 705897 476339 705953 476395
rect 70047 468605 70103 468661
rect 70171 468605 70227 468661
rect 70295 468605 70351 468661
rect 70419 468605 70475 468661
rect 70047 468481 70103 468537
rect 70171 468481 70227 468537
rect 70295 468481 70351 468537
rect 70419 468481 70475 468537
rect 70047 468357 70103 468413
rect 70171 468357 70227 468413
rect 70295 468357 70351 468413
rect 70419 468357 70475 468413
rect 70047 468233 70103 468289
rect 70171 468233 70227 468289
rect 70295 468233 70351 468289
rect 70419 468233 70475 468289
rect 70047 468109 70103 468165
rect 70171 468109 70227 468165
rect 70295 468109 70351 468165
rect 70419 468109 70475 468165
rect 70047 467985 70103 468041
rect 70171 467985 70227 468041
rect 70295 467985 70351 468041
rect 70419 467985 70475 468041
rect 70047 467861 70103 467917
rect 70171 467861 70227 467917
rect 70295 467861 70351 467917
rect 70419 467861 70475 467917
rect 70047 467737 70103 467793
rect 70171 467737 70227 467793
rect 70295 467737 70351 467793
rect 70419 467737 70475 467793
rect 70047 467613 70103 467669
rect 70171 467613 70227 467669
rect 70295 467613 70351 467669
rect 70419 467613 70475 467669
rect 70047 467489 70103 467545
rect 70171 467489 70227 467545
rect 70295 467489 70351 467545
rect 70419 467489 70475 467545
rect 70047 467365 70103 467421
rect 70171 467365 70227 467421
rect 70295 467365 70351 467421
rect 70419 467365 70475 467421
rect 70047 467241 70103 467297
rect 70171 467241 70227 467297
rect 70295 467241 70351 467297
rect 70419 467241 70475 467297
rect 70047 467117 70103 467173
rect 70171 467117 70227 467173
rect 70295 467117 70351 467173
rect 70419 467117 70475 467173
rect 70047 466993 70103 467049
rect 70171 466993 70227 467049
rect 70295 466993 70351 467049
rect 70419 466993 70475 467049
rect 70047 466869 70103 466925
rect 70171 466869 70227 466925
rect 70295 466869 70351 466925
rect 70419 466869 70475 466925
rect 70047 466125 70103 466181
rect 70171 466125 70227 466181
rect 70295 466125 70351 466181
rect 70419 466125 70475 466181
rect 70047 466001 70103 466057
rect 70171 466001 70227 466057
rect 70295 466001 70351 466057
rect 70419 466001 70475 466057
rect 70047 465877 70103 465933
rect 70171 465877 70227 465933
rect 70295 465877 70351 465933
rect 70419 465877 70475 465933
rect 70047 465753 70103 465809
rect 70171 465753 70227 465809
rect 70295 465753 70351 465809
rect 70419 465753 70475 465809
rect 70047 465629 70103 465685
rect 70171 465629 70227 465685
rect 70295 465629 70351 465685
rect 70419 465629 70475 465685
rect 70047 465505 70103 465561
rect 70171 465505 70227 465561
rect 70295 465505 70351 465561
rect 70419 465505 70475 465561
rect 70047 465381 70103 465437
rect 70171 465381 70227 465437
rect 70295 465381 70351 465437
rect 70419 465381 70475 465437
rect 70047 465257 70103 465313
rect 70171 465257 70227 465313
rect 70295 465257 70351 465313
rect 70419 465257 70475 465313
rect 70047 465133 70103 465189
rect 70171 465133 70227 465189
rect 70295 465133 70351 465189
rect 70419 465133 70475 465189
rect 70047 465009 70103 465065
rect 70171 465009 70227 465065
rect 70295 465009 70351 465065
rect 70419 465009 70475 465065
rect 70047 464885 70103 464941
rect 70171 464885 70227 464941
rect 70295 464885 70351 464941
rect 70419 464885 70475 464941
rect 70047 464761 70103 464817
rect 70171 464761 70227 464817
rect 70295 464761 70351 464817
rect 70419 464761 70475 464817
rect 70047 464637 70103 464693
rect 70171 464637 70227 464693
rect 70295 464637 70351 464693
rect 70419 464637 70475 464693
rect 70047 464513 70103 464569
rect 70171 464513 70227 464569
rect 70295 464513 70351 464569
rect 70419 464513 70475 464569
rect 70047 464389 70103 464445
rect 70171 464389 70227 464445
rect 70295 464389 70351 464445
rect 70419 464389 70475 464445
rect 70047 464265 70103 464321
rect 70171 464265 70227 464321
rect 70295 464265 70351 464321
rect 70419 464265 70475 464321
rect 70047 463755 70103 463811
rect 70171 463755 70227 463811
rect 70295 463755 70351 463811
rect 70419 463755 70475 463811
rect 70047 463631 70103 463687
rect 70171 463631 70227 463687
rect 70295 463631 70351 463687
rect 70419 463631 70475 463687
rect 70047 463507 70103 463563
rect 70171 463507 70227 463563
rect 70295 463507 70351 463563
rect 70419 463507 70475 463563
rect 70047 463383 70103 463439
rect 70171 463383 70227 463439
rect 70295 463383 70351 463439
rect 70419 463383 70475 463439
rect 70047 463259 70103 463315
rect 70171 463259 70227 463315
rect 70295 463259 70351 463315
rect 70419 463259 70475 463315
rect 70047 463135 70103 463191
rect 70171 463135 70227 463191
rect 70295 463135 70351 463191
rect 70419 463135 70475 463191
rect 70047 463011 70103 463067
rect 70171 463011 70227 463067
rect 70295 463011 70351 463067
rect 70419 463011 70475 463067
rect 70047 462887 70103 462943
rect 70171 462887 70227 462943
rect 70295 462887 70351 462943
rect 70419 462887 70475 462943
rect 70047 462763 70103 462819
rect 70171 462763 70227 462819
rect 70295 462763 70351 462819
rect 70419 462763 70475 462819
rect 70047 462639 70103 462695
rect 70171 462639 70227 462695
rect 70295 462639 70351 462695
rect 70419 462639 70475 462695
rect 70047 462515 70103 462571
rect 70171 462515 70227 462571
rect 70295 462515 70351 462571
rect 70419 462515 70475 462571
rect 70047 462391 70103 462447
rect 70171 462391 70227 462447
rect 70295 462391 70351 462447
rect 70419 462391 70475 462447
rect 70047 462267 70103 462323
rect 70171 462267 70227 462323
rect 70295 462267 70351 462323
rect 70419 462267 70475 462323
rect 70047 462143 70103 462199
rect 70171 462143 70227 462199
rect 70295 462143 70351 462199
rect 70419 462143 70475 462199
rect 70047 462019 70103 462075
rect 70171 462019 70227 462075
rect 70295 462019 70351 462075
rect 70419 462019 70475 462075
rect 70047 461895 70103 461951
rect 70171 461895 70227 461951
rect 70295 461895 70351 461951
rect 70419 461895 70475 461951
rect 70047 461049 70103 461105
rect 70171 461049 70227 461105
rect 70295 461049 70351 461105
rect 70419 461049 70475 461105
rect 70047 460925 70103 460981
rect 70171 460925 70227 460981
rect 70295 460925 70351 460981
rect 70419 460925 70475 460981
rect 70047 460801 70103 460857
rect 70171 460801 70227 460857
rect 70295 460801 70351 460857
rect 70419 460801 70475 460857
rect 70047 460677 70103 460733
rect 70171 460677 70227 460733
rect 70295 460677 70351 460733
rect 70419 460677 70475 460733
rect 70047 460553 70103 460609
rect 70171 460553 70227 460609
rect 70295 460553 70351 460609
rect 70419 460553 70475 460609
rect 70047 460429 70103 460485
rect 70171 460429 70227 460485
rect 70295 460429 70351 460485
rect 70419 460429 70475 460485
rect 70047 460305 70103 460361
rect 70171 460305 70227 460361
rect 70295 460305 70351 460361
rect 70419 460305 70475 460361
rect 70047 460181 70103 460237
rect 70171 460181 70227 460237
rect 70295 460181 70351 460237
rect 70419 460181 70475 460237
rect 70047 460057 70103 460113
rect 70171 460057 70227 460113
rect 70295 460057 70351 460113
rect 70419 460057 70475 460113
rect 70047 459933 70103 459989
rect 70171 459933 70227 459989
rect 70295 459933 70351 459989
rect 70419 459933 70475 459989
rect 70047 459809 70103 459865
rect 70171 459809 70227 459865
rect 70295 459809 70351 459865
rect 70419 459809 70475 459865
rect 70047 459685 70103 459741
rect 70171 459685 70227 459741
rect 70295 459685 70351 459741
rect 70419 459685 70475 459741
rect 70047 459561 70103 459617
rect 70171 459561 70227 459617
rect 70295 459561 70351 459617
rect 70419 459561 70475 459617
rect 70047 459437 70103 459493
rect 70171 459437 70227 459493
rect 70295 459437 70351 459493
rect 70419 459437 70475 459493
rect 70047 459313 70103 459369
rect 70171 459313 70227 459369
rect 70295 459313 70351 459369
rect 70419 459313 70475 459369
rect 70047 459189 70103 459245
rect 70171 459189 70227 459245
rect 70295 459189 70351 459245
rect 70419 459189 70475 459245
rect 70047 458679 70103 458735
rect 70171 458679 70227 458735
rect 70295 458679 70351 458735
rect 70419 458679 70475 458735
rect 70047 458555 70103 458611
rect 70171 458555 70227 458611
rect 70295 458555 70351 458611
rect 70419 458555 70475 458611
rect 70047 458431 70103 458487
rect 70171 458431 70227 458487
rect 70295 458431 70351 458487
rect 70419 458431 70475 458487
rect 70047 458307 70103 458363
rect 70171 458307 70227 458363
rect 70295 458307 70351 458363
rect 70419 458307 70475 458363
rect 70047 458183 70103 458239
rect 70171 458183 70227 458239
rect 70295 458183 70351 458239
rect 70419 458183 70475 458239
rect 70047 458059 70103 458115
rect 70171 458059 70227 458115
rect 70295 458059 70351 458115
rect 70419 458059 70475 458115
rect 70047 457935 70103 457991
rect 70171 457935 70227 457991
rect 70295 457935 70351 457991
rect 70419 457935 70475 457991
rect 70047 457811 70103 457867
rect 70171 457811 70227 457867
rect 70295 457811 70351 457867
rect 70419 457811 70475 457867
rect 70047 457687 70103 457743
rect 70171 457687 70227 457743
rect 70295 457687 70351 457743
rect 70419 457687 70475 457743
rect 70047 457563 70103 457619
rect 70171 457563 70227 457619
rect 70295 457563 70351 457619
rect 70419 457563 70475 457619
rect 70047 457439 70103 457495
rect 70171 457439 70227 457495
rect 70295 457439 70351 457495
rect 70419 457439 70475 457495
rect 70047 457315 70103 457371
rect 70171 457315 70227 457371
rect 70295 457315 70351 457371
rect 70419 457315 70475 457371
rect 70047 457191 70103 457247
rect 70171 457191 70227 457247
rect 70295 457191 70351 457247
rect 70419 457191 70475 457247
rect 70047 457067 70103 457123
rect 70171 457067 70227 457123
rect 70295 457067 70351 457123
rect 70419 457067 70475 457123
rect 70047 456943 70103 456999
rect 70171 456943 70227 456999
rect 70295 456943 70351 456999
rect 70419 456943 70475 456999
rect 70047 456819 70103 456875
rect 70171 456819 70227 456875
rect 70295 456819 70351 456875
rect 70419 456819 70475 456875
rect 70047 456049 70103 456105
rect 70171 456049 70227 456105
rect 70295 456049 70351 456105
rect 70419 456049 70475 456105
rect 70047 455925 70103 455981
rect 70171 455925 70227 455981
rect 70295 455925 70351 455981
rect 70419 455925 70475 455981
rect 70047 455801 70103 455857
rect 70171 455801 70227 455857
rect 70295 455801 70351 455857
rect 70419 455801 70475 455857
rect 70047 455677 70103 455733
rect 70171 455677 70227 455733
rect 70295 455677 70351 455733
rect 70419 455677 70475 455733
rect 70047 455553 70103 455609
rect 70171 455553 70227 455609
rect 70295 455553 70351 455609
rect 70419 455553 70475 455609
rect 70047 455429 70103 455485
rect 70171 455429 70227 455485
rect 70295 455429 70351 455485
rect 70419 455429 70475 455485
rect 70047 455305 70103 455361
rect 70171 455305 70227 455361
rect 70295 455305 70351 455361
rect 70419 455305 70475 455361
rect 70047 455181 70103 455237
rect 70171 455181 70227 455237
rect 70295 455181 70351 455237
rect 70419 455181 70475 455237
rect 70047 455057 70103 455113
rect 70171 455057 70227 455113
rect 70295 455057 70351 455113
rect 70419 455057 70475 455113
rect 70047 454933 70103 454989
rect 70171 454933 70227 454989
rect 70295 454933 70351 454989
rect 70419 454933 70475 454989
rect 70047 454809 70103 454865
rect 70171 454809 70227 454865
rect 70295 454809 70351 454865
rect 70419 454809 70475 454865
rect 70047 454685 70103 454741
rect 70171 454685 70227 454741
rect 70295 454685 70351 454741
rect 70419 454685 70475 454741
rect 70047 454561 70103 454617
rect 70171 454561 70227 454617
rect 70295 454561 70351 454617
rect 70419 454561 70475 454617
rect 70047 454437 70103 454493
rect 70171 454437 70227 454493
rect 70295 454437 70351 454493
rect 70419 454437 70475 454493
rect 70047 454313 70103 454369
rect 70171 454313 70227 454369
rect 70295 454313 70351 454369
rect 70419 454313 70475 454369
rect 705525 447631 705581 447687
rect 705649 447631 705705 447687
rect 705773 447631 705829 447687
rect 705897 447631 705953 447687
rect 705525 447507 705581 447563
rect 705649 447507 705705 447563
rect 705773 447507 705829 447563
rect 705897 447507 705953 447563
rect 705525 447383 705581 447439
rect 705649 447383 705705 447439
rect 705773 447383 705829 447439
rect 705897 447383 705953 447439
rect 705525 447259 705581 447315
rect 705649 447259 705705 447315
rect 705773 447259 705829 447315
rect 705897 447259 705953 447315
rect 705525 447135 705581 447191
rect 705649 447135 705705 447191
rect 705773 447135 705829 447191
rect 705897 447135 705953 447191
rect 705525 447011 705581 447067
rect 705649 447011 705705 447067
rect 705773 447011 705829 447067
rect 705897 447011 705953 447067
rect 705525 446887 705581 446943
rect 705649 446887 705705 446943
rect 705773 446887 705829 446943
rect 705897 446887 705953 446943
rect 705525 446763 705581 446819
rect 705649 446763 705705 446819
rect 705773 446763 705829 446819
rect 705897 446763 705953 446819
rect 705525 446639 705581 446695
rect 705649 446639 705705 446695
rect 705773 446639 705829 446695
rect 705897 446639 705953 446695
rect 705525 446515 705581 446571
rect 705649 446515 705705 446571
rect 705773 446515 705829 446571
rect 705897 446515 705953 446571
rect 705525 446391 705581 446447
rect 705649 446391 705705 446447
rect 705773 446391 705829 446447
rect 705897 446391 705953 446447
rect 705525 446267 705581 446323
rect 705649 446267 705705 446323
rect 705773 446267 705829 446323
rect 705897 446267 705953 446323
rect 705525 446143 705581 446199
rect 705649 446143 705705 446199
rect 705773 446143 705829 446199
rect 705897 446143 705953 446199
rect 705525 446019 705581 446075
rect 705649 446019 705705 446075
rect 705773 446019 705829 446075
rect 705897 446019 705953 446075
rect 705525 445895 705581 445951
rect 705649 445895 705705 445951
rect 705773 445895 705829 445951
rect 705897 445895 705953 445951
rect 705525 445125 705581 445181
rect 705649 445125 705705 445181
rect 705773 445125 705829 445181
rect 705897 445125 705953 445181
rect 705525 445001 705581 445057
rect 705649 445001 705705 445057
rect 705773 445001 705829 445057
rect 705897 445001 705953 445057
rect 705525 444877 705581 444933
rect 705649 444877 705705 444933
rect 705773 444877 705829 444933
rect 705897 444877 705953 444933
rect 705525 444753 705581 444809
rect 705649 444753 705705 444809
rect 705773 444753 705829 444809
rect 705897 444753 705953 444809
rect 705525 444629 705581 444685
rect 705649 444629 705705 444685
rect 705773 444629 705829 444685
rect 705897 444629 705953 444685
rect 705525 444505 705581 444561
rect 705649 444505 705705 444561
rect 705773 444505 705829 444561
rect 705897 444505 705953 444561
rect 705525 444381 705581 444437
rect 705649 444381 705705 444437
rect 705773 444381 705829 444437
rect 705897 444381 705953 444437
rect 705525 444257 705581 444313
rect 705649 444257 705705 444313
rect 705773 444257 705829 444313
rect 705897 444257 705953 444313
rect 705525 444133 705581 444189
rect 705649 444133 705705 444189
rect 705773 444133 705829 444189
rect 705897 444133 705953 444189
rect 705525 444009 705581 444065
rect 705649 444009 705705 444065
rect 705773 444009 705829 444065
rect 705897 444009 705953 444065
rect 705525 443885 705581 443941
rect 705649 443885 705705 443941
rect 705773 443885 705829 443941
rect 705897 443885 705953 443941
rect 705525 443761 705581 443817
rect 705649 443761 705705 443817
rect 705773 443761 705829 443817
rect 705897 443761 705953 443817
rect 705525 443637 705581 443693
rect 705649 443637 705705 443693
rect 705773 443637 705829 443693
rect 705897 443637 705953 443693
rect 705525 443513 705581 443569
rect 705649 443513 705705 443569
rect 705773 443513 705829 443569
rect 705897 443513 705953 443569
rect 705525 443389 705581 443445
rect 705649 443389 705705 443445
rect 705773 443389 705829 443445
rect 705897 443389 705953 443445
rect 705525 443265 705581 443321
rect 705649 443265 705705 443321
rect 705773 443265 705829 443321
rect 705897 443265 705953 443321
rect 705525 442755 705581 442811
rect 705649 442755 705705 442811
rect 705773 442755 705829 442811
rect 705897 442755 705953 442811
rect 705525 442631 705581 442687
rect 705649 442631 705705 442687
rect 705773 442631 705829 442687
rect 705897 442631 705953 442687
rect 705525 442507 705581 442563
rect 705649 442507 705705 442563
rect 705773 442507 705829 442563
rect 705897 442507 705953 442563
rect 705525 442383 705581 442439
rect 705649 442383 705705 442439
rect 705773 442383 705829 442439
rect 705897 442383 705953 442439
rect 705525 442259 705581 442315
rect 705649 442259 705705 442315
rect 705773 442259 705829 442315
rect 705897 442259 705953 442315
rect 705525 442135 705581 442191
rect 705649 442135 705705 442191
rect 705773 442135 705829 442191
rect 705897 442135 705953 442191
rect 705525 442011 705581 442067
rect 705649 442011 705705 442067
rect 705773 442011 705829 442067
rect 705897 442011 705953 442067
rect 705525 441887 705581 441943
rect 705649 441887 705705 441943
rect 705773 441887 705829 441943
rect 705897 441887 705953 441943
rect 705525 441763 705581 441819
rect 705649 441763 705705 441819
rect 705773 441763 705829 441819
rect 705897 441763 705953 441819
rect 705525 441639 705581 441695
rect 705649 441639 705705 441695
rect 705773 441639 705829 441695
rect 705897 441639 705953 441695
rect 705525 441515 705581 441571
rect 705649 441515 705705 441571
rect 705773 441515 705829 441571
rect 705897 441515 705953 441571
rect 705525 441391 705581 441447
rect 705649 441391 705705 441447
rect 705773 441391 705829 441447
rect 705897 441391 705953 441447
rect 705525 441267 705581 441323
rect 705649 441267 705705 441323
rect 705773 441267 705829 441323
rect 705897 441267 705953 441323
rect 705525 441143 705581 441199
rect 705649 441143 705705 441199
rect 705773 441143 705829 441199
rect 705897 441143 705953 441199
rect 705525 441019 705581 441075
rect 705649 441019 705705 441075
rect 705773 441019 705829 441075
rect 705897 441019 705953 441075
rect 705525 440895 705581 440951
rect 705649 440895 705705 440951
rect 705773 440895 705829 440951
rect 705897 440895 705953 440951
rect 705525 440049 705581 440105
rect 705649 440049 705705 440105
rect 705773 440049 705829 440105
rect 705897 440049 705953 440105
rect 705525 439925 705581 439981
rect 705649 439925 705705 439981
rect 705773 439925 705829 439981
rect 705897 439925 705953 439981
rect 705525 439801 705581 439857
rect 705649 439801 705705 439857
rect 705773 439801 705829 439857
rect 705897 439801 705953 439857
rect 705525 439677 705581 439733
rect 705649 439677 705705 439733
rect 705773 439677 705829 439733
rect 705897 439677 705953 439733
rect 705525 439553 705581 439609
rect 705649 439553 705705 439609
rect 705773 439553 705829 439609
rect 705897 439553 705953 439609
rect 705525 439429 705581 439485
rect 705649 439429 705705 439485
rect 705773 439429 705829 439485
rect 705897 439429 705953 439485
rect 705525 439305 705581 439361
rect 705649 439305 705705 439361
rect 705773 439305 705829 439361
rect 705897 439305 705953 439361
rect 705525 439181 705581 439237
rect 705649 439181 705705 439237
rect 705773 439181 705829 439237
rect 705897 439181 705953 439237
rect 705525 439057 705581 439113
rect 705649 439057 705705 439113
rect 705773 439057 705829 439113
rect 705897 439057 705953 439113
rect 705525 438933 705581 438989
rect 705649 438933 705705 438989
rect 705773 438933 705829 438989
rect 705897 438933 705953 438989
rect 705525 438809 705581 438865
rect 705649 438809 705705 438865
rect 705773 438809 705829 438865
rect 705897 438809 705953 438865
rect 705525 438685 705581 438741
rect 705649 438685 705705 438741
rect 705773 438685 705829 438741
rect 705897 438685 705953 438741
rect 705525 438561 705581 438617
rect 705649 438561 705705 438617
rect 705773 438561 705829 438617
rect 705897 438561 705953 438617
rect 705525 438437 705581 438493
rect 705649 438437 705705 438493
rect 705773 438437 705829 438493
rect 705897 438437 705953 438493
rect 705525 438313 705581 438369
rect 705649 438313 705705 438369
rect 705773 438313 705829 438369
rect 705897 438313 705953 438369
rect 705525 438189 705581 438245
rect 705649 438189 705705 438245
rect 705773 438189 705829 438245
rect 705897 438189 705953 438245
rect 705525 437679 705581 437735
rect 705649 437679 705705 437735
rect 705773 437679 705829 437735
rect 705897 437679 705953 437735
rect 705525 437555 705581 437611
rect 705649 437555 705705 437611
rect 705773 437555 705829 437611
rect 705897 437555 705953 437611
rect 705525 437431 705581 437487
rect 705649 437431 705705 437487
rect 705773 437431 705829 437487
rect 705897 437431 705953 437487
rect 705525 437307 705581 437363
rect 705649 437307 705705 437363
rect 705773 437307 705829 437363
rect 705897 437307 705953 437363
rect 705525 437183 705581 437239
rect 705649 437183 705705 437239
rect 705773 437183 705829 437239
rect 705897 437183 705953 437239
rect 705525 437059 705581 437115
rect 705649 437059 705705 437115
rect 705773 437059 705829 437115
rect 705897 437059 705953 437115
rect 705525 436935 705581 436991
rect 705649 436935 705705 436991
rect 705773 436935 705829 436991
rect 705897 436935 705953 436991
rect 705525 436811 705581 436867
rect 705649 436811 705705 436867
rect 705773 436811 705829 436867
rect 705897 436811 705953 436867
rect 705525 436687 705581 436743
rect 705649 436687 705705 436743
rect 705773 436687 705829 436743
rect 705897 436687 705953 436743
rect 705525 436563 705581 436619
rect 705649 436563 705705 436619
rect 705773 436563 705829 436619
rect 705897 436563 705953 436619
rect 705525 436439 705581 436495
rect 705649 436439 705705 436495
rect 705773 436439 705829 436495
rect 705897 436439 705953 436495
rect 705525 436315 705581 436371
rect 705649 436315 705705 436371
rect 705773 436315 705829 436371
rect 705897 436315 705953 436371
rect 705525 436191 705581 436247
rect 705649 436191 705705 436247
rect 705773 436191 705829 436247
rect 705897 436191 705953 436247
rect 705525 435075 705581 435131
rect 705649 435075 705705 435131
rect 705773 435075 705829 435131
rect 705897 435075 705953 435131
rect 705525 434951 705581 435007
rect 705649 434951 705705 435007
rect 705773 434951 705829 435007
rect 705897 434951 705953 435007
rect 705525 434827 705581 434883
rect 705649 434827 705705 434883
rect 705773 434827 705829 434883
rect 705897 434827 705953 434883
rect 705525 434703 705581 434759
rect 705649 434703 705705 434759
rect 705773 434703 705829 434759
rect 705897 434703 705953 434759
rect 705525 434579 705581 434635
rect 705649 434579 705705 434635
rect 705773 434579 705829 434635
rect 705897 434579 705953 434635
rect 705525 434455 705581 434511
rect 705649 434455 705705 434511
rect 705773 434455 705829 434511
rect 705897 434455 705953 434511
rect 705525 434331 705581 434387
rect 705649 434331 705705 434387
rect 705773 434331 705829 434387
rect 705897 434331 705953 434387
rect 705525 434207 705581 434263
rect 705649 434207 705705 434263
rect 705773 434207 705829 434263
rect 705897 434207 705953 434263
rect 705525 434083 705581 434139
rect 705649 434083 705705 434139
rect 705773 434083 705829 434139
rect 705897 434083 705953 434139
rect 705525 433959 705581 434015
rect 705649 433959 705705 434015
rect 705773 433959 705829 434015
rect 705897 433959 705953 434015
rect 705525 433835 705581 433891
rect 705649 433835 705705 433891
rect 705773 433835 705829 433891
rect 705897 433835 705953 433891
rect 705525 433711 705581 433767
rect 705649 433711 705705 433767
rect 705773 433711 705829 433767
rect 705897 433711 705953 433767
rect 705525 433587 705581 433643
rect 705649 433587 705705 433643
rect 705773 433587 705829 433643
rect 705897 433587 705953 433643
rect 705525 433463 705581 433519
rect 705649 433463 705705 433519
rect 705773 433463 705829 433519
rect 705897 433463 705953 433519
rect 705525 433339 705581 433395
rect 705649 433339 705705 433395
rect 705773 433339 705829 433395
rect 705897 433339 705953 433395
rect 70047 427605 70103 427661
rect 70171 427605 70227 427661
rect 70295 427605 70351 427661
rect 70419 427605 70475 427661
rect 70047 427481 70103 427537
rect 70171 427481 70227 427537
rect 70295 427481 70351 427537
rect 70419 427481 70475 427537
rect 70047 427357 70103 427413
rect 70171 427357 70227 427413
rect 70295 427357 70351 427413
rect 70419 427357 70475 427413
rect 70047 427233 70103 427289
rect 70171 427233 70227 427289
rect 70295 427233 70351 427289
rect 70419 427233 70475 427289
rect 70047 427109 70103 427165
rect 70171 427109 70227 427165
rect 70295 427109 70351 427165
rect 70419 427109 70475 427165
rect 70047 426985 70103 427041
rect 70171 426985 70227 427041
rect 70295 426985 70351 427041
rect 70419 426985 70475 427041
rect 70047 426861 70103 426917
rect 70171 426861 70227 426917
rect 70295 426861 70351 426917
rect 70419 426861 70475 426917
rect 70047 426737 70103 426793
rect 70171 426737 70227 426793
rect 70295 426737 70351 426793
rect 70419 426737 70475 426793
rect 70047 426613 70103 426669
rect 70171 426613 70227 426669
rect 70295 426613 70351 426669
rect 70419 426613 70475 426669
rect 70047 426489 70103 426545
rect 70171 426489 70227 426545
rect 70295 426489 70351 426545
rect 70419 426489 70475 426545
rect 70047 426365 70103 426421
rect 70171 426365 70227 426421
rect 70295 426365 70351 426421
rect 70419 426365 70475 426421
rect 70047 426241 70103 426297
rect 70171 426241 70227 426297
rect 70295 426241 70351 426297
rect 70419 426241 70475 426297
rect 70047 426117 70103 426173
rect 70171 426117 70227 426173
rect 70295 426117 70351 426173
rect 70419 426117 70475 426173
rect 70047 425993 70103 426049
rect 70171 425993 70227 426049
rect 70295 425993 70351 426049
rect 70419 425993 70475 426049
rect 70047 425869 70103 425925
rect 70171 425869 70227 425925
rect 70295 425869 70351 425925
rect 70419 425869 70475 425925
rect 70047 425125 70103 425181
rect 70171 425125 70227 425181
rect 70295 425125 70351 425181
rect 70419 425125 70475 425181
rect 70047 425001 70103 425057
rect 70171 425001 70227 425057
rect 70295 425001 70351 425057
rect 70419 425001 70475 425057
rect 70047 424877 70103 424933
rect 70171 424877 70227 424933
rect 70295 424877 70351 424933
rect 70419 424877 70475 424933
rect 70047 424753 70103 424809
rect 70171 424753 70227 424809
rect 70295 424753 70351 424809
rect 70419 424753 70475 424809
rect 70047 424629 70103 424685
rect 70171 424629 70227 424685
rect 70295 424629 70351 424685
rect 70419 424629 70475 424685
rect 70047 424505 70103 424561
rect 70171 424505 70227 424561
rect 70295 424505 70351 424561
rect 70419 424505 70475 424561
rect 70047 424381 70103 424437
rect 70171 424381 70227 424437
rect 70295 424381 70351 424437
rect 70419 424381 70475 424437
rect 70047 424257 70103 424313
rect 70171 424257 70227 424313
rect 70295 424257 70351 424313
rect 70419 424257 70475 424313
rect 70047 424133 70103 424189
rect 70171 424133 70227 424189
rect 70295 424133 70351 424189
rect 70419 424133 70475 424189
rect 70047 424009 70103 424065
rect 70171 424009 70227 424065
rect 70295 424009 70351 424065
rect 70419 424009 70475 424065
rect 70047 423885 70103 423941
rect 70171 423885 70227 423941
rect 70295 423885 70351 423941
rect 70419 423885 70475 423941
rect 70047 423761 70103 423817
rect 70171 423761 70227 423817
rect 70295 423761 70351 423817
rect 70419 423761 70475 423817
rect 70047 423637 70103 423693
rect 70171 423637 70227 423693
rect 70295 423637 70351 423693
rect 70419 423637 70475 423693
rect 70047 423513 70103 423569
rect 70171 423513 70227 423569
rect 70295 423513 70351 423569
rect 70419 423513 70475 423569
rect 70047 423389 70103 423445
rect 70171 423389 70227 423445
rect 70295 423389 70351 423445
rect 70419 423389 70475 423445
rect 70047 423265 70103 423321
rect 70171 423265 70227 423321
rect 70295 423265 70351 423321
rect 70419 423265 70475 423321
rect 70047 422755 70103 422811
rect 70171 422755 70227 422811
rect 70295 422755 70351 422811
rect 70419 422755 70475 422811
rect 70047 422631 70103 422687
rect 70171 422631 70227 422687
rect 70295 422631 70351 422687
rect 70419 422631 70475 422687
rect 70047 422507 70103 422563
rect 70171 422507 70227 422563
rect 70295 422507 70351 422563
rect 70419 422507 70475 422563
rect 70047 422383 70103 422439
rect 70171 422383 70227 422439
rect 70295 422383 70351 422439
rect 70419 422383 70475 422439
rect 70047 422259 70103 422315
rect 70171 422259 70227 422315
rect 70295 422259 70351 422315
rect 70419 422259 70475 422315
rect 70047 422135 70103 422191
rect 70171 422135 70227 422191
rect 70295 422135 70351 422191
rect 70419 422135 70475 422191
rect 70047 422011 70103 422067
rect 70171 422011 70227 422067
rect 70295 422011 70351 422067
rect 70419 422011 70475 422067
rect 70047 421887 70103 421943
rect 70171 421887 70227 421943
rect 70295 421887 70351 421943
rect 70419 421887 70475 421943
rect 70047 421763 70103 421819
rect 70171 421763 70227 421819
rect 70295 421763 70351 421819
rect 70419 421763 70475 421819
rect 70047 421639 70103 421695
rect 70171 421639 70227 421695
rect 70295 421639 70351 421695
rect 70419 421639 70475 421695
rect 70047 421515 70103 421571
rect 70171 421515 70227 421571
rect 70295 421515 70351 421571
rect 70419 421515 70475 421571
rect 70047 421391 70103 421447
rect 70171 421391 70227 421447
rect 70295 421391 70351 421447
rect 70419 421391 70475 421447
rect 70047 421267 70103 421323
rect 70171 421267 70227 421323
rect 70295 421267 70351 421323
rect 70419 421267 70475 421323
rect 70047 421143 70103 421199
rect 70171 421143 70227 421199
rect 70295 421143 70351 421199
rect 70419 421143 70475 421199
rect 70047 421019 70103 421075
rect 70171 421019 70227 421075
rect 70295 421019 70351 421075
rect 70419 421019 70475 421075
rect 70047 420895 70103 420951
rect 70171 420895 70227 420951
rect 70295 420895 70351 420951
rect 70419 420895 70475 420951
rect 70047 420049 70103 420105
rect 70171 420049 70227 420105
rect 70295 420049 70351 420105
rect 70419 420049 70475 420105
rect 70047 419925 70103 419981
rect 70171 419925 70227 419981
rect 70295 419925 70351 419981
rect 70419 419925 70475 419981
rect 70047 419801 70103 419857
rect 70171 419801 70227 419857
rect 70295 419801 70351 419857
rect 70419 419801 70475 419857
rect 70047 419677 70103 419733
rect 70171 419677 70227 419733
rect 70295 419677 70351 419733
rect 70419 419677 70475 419733
rect 70047 419553 70103 419609
rect 70171 419553 70227 419609
rect 70295 419553 70351 419609
rect 70419 419553 70475 419609
rect 70047 419429 70103 419485
rect 70171 419429 70227 419485
rect 70295 419429 70351 419485
rect 70419 419429 70475 419485
rect 70047 419305 70103 419361
rect 70171 419305 70227 419361
rect 70295 419305 70351 419361
rect 70419 419305 70475 419361
rect 70047 419181 70103 419237
rect 70171 419181 70227 419237
rect 70295 419181 70351 419237
rect 70419 419181 70475 419237
rect 70047 419057 70103 419113
rect 70171 419057 70227 419113
rect 70295 419057 70351 419113
rect 70419 419057 70475 419113
rect 70047 418933 70103 418989
rect 70171 418933 70227 418989
rect 70295 418933 70351 418989
rect 70419 418933 70475 418989
rect 70047 418809 70103 418865
rect 70171 418809 70227 418865
rect 70295 418809 70351 418865
rect 70419 418809 70475 418865
rect 70047 418685 70103 418741
rect 70171 418685 70227 418741
rect 70295 418685 70351 418741
rect 70419 418685 70475 418741
rect 70047 418561 70103 418617
rect 70171 418561 70227 418617
rect 70295 418561 70351 418617
rect 70419 418561 70475 418617
rect 70047 418437 70103 418493
rect 70171 418437 70227 418493
rect 70295 418437 70351 418493
rect 70419 418437 70475 418493
rect 70047 418313 70103 418369
rect 70171 418313 70227 418369
rect 70295 418313 70351 418369
rect 70419 418313 70475 418369
rect 70047 418189 70103 418245
rect 70171 418189 70227 418245
rect 70295 418189 70351 418245
rect 70419 418189 70475 418245
rect 70047 417679 70103 417735
rect 70171 417679 70227 417735
rect 70295 417679 70351 417735
rect 70419 417679 70475 417735
rect 70047 417555 70103 417611
rect 70171 417555 70227 417611
rect 70295 417555 70351 417611
rect 70419 417555 70475 417611
rect 70047 417431 70103 417487
rect 70171 417431 70227 417487
rect 70295 417431 70351 417487
rect 70419 417431 70475 417487
rect 70047 417307 70103 417363
rect 70171 417307 70227 417363
rect 70295 417307 70351 417363
rect 70419 417307 70475 417363
rect 70047 417183 70103 417239
rect 70171 417183 70227 417239
rect 70295 417183 70351 417239
rect 70419 417183 70475 417239
rect 70047 417059 70103 417115
rect 70171 417059 70227 417115
rect 70295 417059 70351 417115
rect 70419 417059 70475 417115
rect 70047 416935 70103 416991
rect 70171 416935 70227 416991
rect 70295 416935 70351 416991
rect 70419 416935 70475 416991
rect 70047 416811 70103 416867
rect 70171 416811 70227 416867
rect 70295 416811 70351 416867
rect 70419 416811 70475 416867
rect 70047 416687 70103 416743
rect 70171 416687 70227 416743
rect 70295 416687 70351 416743
rect 70419 416687 70475 416743
rect 70047 416563 70103 416619
rect 70171 416563 70227 416619
rect 70295 416563 70351 416619
rect 70419 416563 70475 416619
rect 70047 416439 70103 416495
rect 70171 416439 70227 416495
rect 70295 416439 70351 416495
rect 70419 416439 70475 416495
rect 70047 416315 70103 416371
rect 70171 416315 70227 416371
rect 70295 416315 70351 416371
rect 70419 416315 70475 416371
rect 70047 416191 70103 416247
rect 70171 416191 70227 416247
rect 70295 416191 70351 416247
rect 70419 416191 70475 416247
rect 70047 416067 70103 416123
rect 70171 416067 70227 416123
rect 70295 416067 70351 416123
rect 70419 416067 70475 416123
rect 70047 415943 70103 415999
rect 70171 415943 70227 415999
rect 70295 415943 70351 415999
rect 70419 415943 70475 415999
rect 70047 415819 70103 415875
rect 70171 415819 70227 415875
rect 70295 415819 70351 415875
rect 70419 415819 70475 415875
rect 70047 415049 70103 415105
rect 70171 415049 70227 415105
rect 70295 415049 70351 415105
rect 70419 415049 70475 415105
rect 70047 414925 70103 414981
rect 70171 414925 70227 414981
rect 70295 414925 70351 414981
rect 70419 414925 70475 414981
rect 70047 414801 70103 414857
rect 70171 414801 70227 414857
rect 70295 414801 70351 414857
rect 70419 414801 70475 414857
rect 70047 414677 70103 414733
rect 70171 414677 70227 414733
rect 70295 414677 70351 414733
rect 70419 414677 70475 414733
rect 70047 414553 70103 414609
rect 70171 414553 70227 414609
rect 70295 414553 70351 414609
rect 70419 414553 70475 414609
rect 70047 414429 70103 414485
rect 70171 414429 70227 414485
rect 70295 414429 70351 414485
rect 70419 414429 70475 414485
rect 70047 414305 70103 414361
rect 70171 414305 70227 414361
rect 70295 414305 70351 414361
rect 70419 414305 70475 414361
rect 70047 414181 70103 414237
rect 70171 414181 70227 414237
rect 70295 414181 70351 414237
rect 70419 414181 70475 414237
rect 70047 414057 70103 414113
rect 70171 414057 70227 414113
rect 70295 414057 70351 414113
rect 70419 414057 70475 414113
rect 70047 413933 70103 413989
rect 70171 413933 70227 413989
rect 70295 413933 70351 413989
rect 70419 413933 70475 413989
rect 70047 413809 70103 413865
rect 70171 413809 70227 413865
rect 70295 413809 70351 413865
rect 70419 413809 70475 413865
rect 70047 413685 70103 413741
rect 70171 413685 70227 413741
rect 70295 413685 70351 413741
rect 70419 413685 70475 413741
rect 70047 413561 70103 413617
rect 70171 413561 70227 413617
rect 70295 413561 70351 413617
rect 70419 413561 70475 413617
rect 70047 413437 70103 413493
rect 70171 413437 70227 413493
rect 70295 413437 70351 413493
rect 70419 413437 70475 413493
rect 70047 413313 70103 413369
rect 70171 413313 70227 413369
rect 70295 413313 70351 413369
rect 70419 413313 70475 413369
rect 705525 404631 705581 404687
rect 705649 404631 705705 404687
rect 705773 404631 705829 404687
rect 705897 404631 705953 404687
rect 705525 404507 705581 404563
rect 705649 404507 705705 404563
rect 705773 404507 705829 404563
rect 705897 404507 705953 404563
rect 705525 404383 705581 404439
rect 705649 404383 705705 404439
rect 705773 404383 705829 404439
rect 705897 404383 705953 404439
rect 705525 404259 705581 404315
rect 705649 404259 705705 404315
rect 705773 404259 705829 404315
rect 705897 404259 705953 404315
rect 705525 404135 705581 404191
rect 705649 404135 705705 404191
rect 705773 404135 705829 404191
rect 705897 404135 705953 404191
rect 705525 404011 705581 404067
rect 705649 404011 705705 404067
rect 705773 404011 705829 404067
rect 705897 404011 705953 404067
rect 705525 403887 705581 403943
rect 705649 403887 705705 403943
rect 705773 403887 705829 403943
rect 705897 403887 705953 403943
rect 705525 403763 705581 403819
rect 705649 403763 705705 403819
rect 705773 403763 705829 403819
rect 705897 403763 705953 403819
rect 705525 403639 705581 403695
rect 705649 403639 705705 403695
rect 705773 403639 705829 403695
rect 705897 403639 705953 403695
rect 705525 403515 705581 403571
rect 705649 403515 705705 403571
rect 705773 403515 705829 403571
rect 705897 403515 705953 403571
rect 705525 403391 705581 403447
rect 705649 403391 705705 403447
rect 705773 403391 705829 403447
rect 705897 403391 705953 403447
rect 705525 403267 705581 403323
rect 705649 403267 705705 403323
rect 705773 403267 705829 403323
rect 705897 403267 705953 403323
rect 705525 403143 705581 403199
rect 705649 403143 705705 403199
rect 705773 403143 705829 403199
rect 705897 403143 705953 403199
rect 705525 403019 705581 403075
rect 705649 403019 705705 403075
rect 705773 403019 705829 403075
rect 705897 403019 705953 403075
rect 705525 402895 705581 402951
rect 705649 402895 705705 402951
rect 705773 402895 705829 402951
rect 705897 402895 705953 402951
rect 705525 402125 705581 402181
rect 705649 402125 705705 402181
rect 705773 402125 705829 402181
rect 705897 402125 705953 402181
rect 705525 402001 705581 402057
rect 705649 402001 705705 402057
rect 705773 402001 705829 402057
rect 705897 402001 705953 402057
rect 705525 401877 705581 401933
rect 705649 401877 705705 401933
rect 705773 401877 705829 401933
rect 705897 401877 705953 401933
rect 705525 401753 705581 401809
rect 705649 401753 705705 401809
rect 705773 401753 705829 401809
rect 705897 401753 705953 401809
rect 705525 401629 705581 401685
rect 705649 401629 705705 401685
rect 705773 401629 705829 401685
rect 705897 401629 705953 401685
rect 705525 401505 705581 401561
rect 705649 401505 705705 401561
rect 705773 401505 705829 401561
rect 705897 401505 705953 401561
rect 705525 401381 705581 401437
rect 705649 401381 705705 401437
rect 705773 401381 705829 401437
rect 705897 401381 705953 401437
rect 705525 401257 705581 401313
rect 705649 401257 705705 401313
rect 705773 401257 705829 401313
rect 705897 401257 705953 401313
rect 705525 401133 705581 401189
rect 705649 401133 705705 401189
rect 705773 401133 705829 401189
rect 705897 401133 705953 401189
rect 705525 401009 705581 401065
rect 705649 401009 705705 401065
rect 705773 401009 705829 401065
rect 705897 401009 705953 401065
rect 705525 400885 705581 400941
rect 705649 400885 705705 400941
rect 705773 400885 705829 400941
rect 705897 400885 705953 400941
rect 705525 400761 705581 400817
rect 705649 400761 705705 400817
rect 705773 400761 705829 400817
rect 705897 400761 705953 400817
rect 705525 400637 705581 400693
rect 705649 400637 705705 400693
rect 705773 400637 705829 400693
rect 705897 400637 705953 400693
rect 705525 400513 705581 400569
rect 705649 400513 705705 400569
rect 705773 400513 705829 400569
rect 705897 400513 705953 400569
rect 705525 400389 705581 400445
rect 705649 400389 705705 400445
rect 705773 400389 705829 400445
rect 705897 400389 705953 400445
rect 705525 400265 705581 400321
rect 705649 400265 705705 400321
rect 705773 400265 705829 400321
rect 705897 400265 705953 400321
rect 705525 399755 705581 399811
rect 705649 399755 705705 399811
rect 705773 399755 705829 399811
rect 705897 399755 705953 399811
rect 705525 399631 705581 399687
rect 705649 399631 705705 399687
rect 705773 399631 705829 399687
rect 705897 399631 705953 399687
rect 705525 399507 705581 399563
rect 705649 399507 705705 399563
rect 705773 399507 705829 399563
rect 705897 399507 705953 399563
rect 705525 399383 705581 399439
rect 705649 399383 705705 399439
rect 705773 399383 705829 399439
rect 705897 399383 705953 399439
rect 705525 399259 705581 399315
rect 705649 399259 705705 399315
rect 705773 399259 705829 399315
rect 705897 399259 705953 399315
rect 705525 399135 705581 399191
rect 705649 399135 705705 399191
rect 705773 399135 705829 399191
rect 705897 399135 705953 399191
rect 705525 399011 705581 399067
rect 705649 399011 705705 399067
rect 705773 399011 705829 399067
rect 705897 399011 705953 399067
rect 705525 398887 705581 398943
rect 705649 398887 705705 398943
rect 705773 398887 705829 398943
rect 705897 398887 705953 398943
rect 705525 398763 705581 398819
rect 705649 398763 705705 398819
rect 705773 398763 705829 398819
rect 705897 398763 705953 398819
rect 705525 398639 705581 398695
rect 705649 398639 705705 398695
rect 705773 398639 705829 398695
rect 705897 398639 705953 398695
rect 705525 398515 705581 398571
rect 705649 398515 705705 398571
rect 705773 398515 705829 398571
rect 705897 398515 705953 398571
rect 705525 398391 705581 398447
rect 705649 398391 705705 398447
rect 705773 398391 705829 398447
rect 705897 398391 705953 398447
rect 705525 398267 705581 398323
rect 705649 398267 705705 398323
rect 705773 398267 705829 398323
rect 705897 398267 705953 398323
rect 705525 398143 705581 398199
rect 705649 398143 705705 398199
rect 705773 398143 705829 398199
rect 705897 398143 705953 398199
rect 705525 398019 705581 398075
rect 705649 398019 705705 398075
rect 705773 398019 705829 398075
rect 705897 398019 705953 398075
rect 705525 397895 705581 397951
rect 705649 397895 705705 397951
rect 705773 397895 705829 397951
rect 705897 397895 705953 397951
rect 705525 397049 705581 397105
rect 705649 397049 705705 397105
rect 705773 397049 705829 397105
rect 705897 397049 705953 397105
rect 705525 396925 705581 396981
rect 705649 396925 705705 396981
rect 705773 396925 705829 396981
rect 705897 396925 705953 396981
rect 705525 396801 705581 396857
rect 705649 396801 705705 396857
rect 705773 396801 705829 396857
rect 705897 396801 705953 396857
rect 705525 396677 705581 396733
rect 705649 396677 705705 396733
rect 705773 396677 705829 396733
rect 705897 396677 705953 396733
rect 705525 396553 705581 396609
rect 705649 396553 705705 396609
rect 705773 396553 705829 396609
rect 705897 396553 705953 396609
rect 705525 396429 705581 396485
rect 705649 396429 705705 396485
rect 705773 396429 705829 396485
rect 705897 396429 705953 396485
rect 705525 396305 705581 396361
rect 705649 396305 705705 396361
rect 705773 396305 705829 396361
rect 705897 396305 705953 396361
rect 705525 396181 705581 396237
rect 705649 396181 705705 396237
rect 705773 396181 705829 396237
rect 705897 396181 705953 396237
rect 705525 396057 705581 396113
rect 705649 396057 705705 396113
rect 705773 396057 705829 396113
rect 705897 396057 705953 396113
rect 705525 395933 705581 395989
rect 705649 395933 705705 395989
rect 705773 395933 705829 395989
rect 705897 395933 705953 395989
rect 705525 395809 705581 395865
rect 705649 395809 705705 395865
rect 705773 395809 705829 395865
rect 705897 395809 705953 395865
rect 705525 395685 705581 395741
rect 705649 395685 705705 395741
rect 705773 395685 705829 395741
rect 705897 395685 705953 395741
rect 705525 395561 705581 395617
rect 705649 395561 705705 395617
rect 705773 395561 705829 395617
rect 705897 395561 705953 395617
rect 705525 395437 705581 395493
rect 705649 395437 705705 395493
rect 705773 395437 705829 395493
rect 705897 395437 705953 395493
rect 705525 395313 705581 395369
rect 705649 395313 705705 395369
rect 705773 395313 705829 395369
rect 705897 395313 705953 395369
rect 705525 395189 705581 395245
rect 705649 395189 705705 395245
rect 705773 395189 705829 395245
rect 705897 395189 705953 395245
rect 705525 394679 705581 394735
rect 705649 394679 705705 394735
rect 705773 394679 705829 394735
rect 705897 394679 705953 394735
rect 705525 394555 705581 394611
rect 705649 394555 705705 394611
rect 705773 394555 705829 394611
rect 705897 394555 705953 394611
rect 705525 394431 705581 394487
rect 705649 394431 705705 394487
rect 705773 394431 705829 394487
rect 705897 394431 705953 394487
rect 705525 394307 705581 394363
rect 705649 394307 705705 394363
rect 705773 394307 705829 394363
rect 705897 394307 705953 394363
rect 705525 394183 705581 394239
rect 705649 394183 705705 394239
rect 705773 394183 705829 394239
rect 705897 394183 705953 394239
rect 705525 394059 705581 394115
rect 705649 394059 705705 394115
rect 705773 394059 705829 394115
rect 705897 394059 705953 394115
rect 705525 393935 705581 393991
rect 705649 393935 705705 393991
rect 705773 393935 705829 393991
rect 705897 393935 705953 393991
rect 705525 393811 705581 393867
rect 705649 393811 705705 393867
rect 705773 393811 705829 393867
rect 705897 393811 705953 393867
rect 705525 393687 705581 393743
rect 705649 393687 705705 393743
rect 705773 393687 705829 393743
rect 705897 393687 705953 393743
rect 705525 393563 705581 393619
rect 705649 393563 705705 393619
rect 705773 393563 705829 393619
rect 705897 393563 705953 393619
rect 705525 393439 705581 393495
rect 705649 393439 705705 393495
rect 705773 393439 705829 393495
rect 705897 393439 705953 393495
rect 705525 393315 705581 393371
rect 705649 393315 705705 393371
rect 705773 393315 705829 393371
rect 705897 393315 705953 393371
rect 705525 393191 705581 393247
rect 705649 393191 705705 393247
rect 705773 393191 705829 393247
rect 705897 393191 705953 393247
rect 705525 393067 705581 393123
rect 705649 393067 705705 393123
rect 705773 393067 705829 393123
rect 705897 393067 705953 393123
rect 705525 392943 705581 392999
rect 705649 392943 705705 392999
rect 705773 392943 705829 392999
rect 705897 392943 705953 392999
rect 705525 392819 705581 392875
rect 705649 392819 705705 392875
rect 705773 392819 705829 392875
rect 705897 392819 705953 392875
rect 705525 392075 705581 392131
rect 705649 392075 705705 392131
rect 705773 392075 705829 392131
rect 705897 392075 705953 392131
rect 705525 391951 705581 392007
rect 705649 391951 705705 392007
rect 705773 391951 705829 392007
rect 705897 391951 705953 392007
rect 705525 391827 705581 391883
rect 705649 391827 705705 391883
rect 705773 391827 705829 391883
rect 705897 391827 705953 391883
rect 705525 391703 705581 391759
rect 705649 391703 705705 391759
rect 705773 391703 705829 391759
rect 705897 391703 705953 391759
rect 705525 391579 705581 391635
rect 705649 391579 705705 391635
rect 705773 391579 705829 391635
rect 705897 391579 705953 391635
rect 705525 391455 705581 391511
rect 705649 391455 705705 391511
rect 705773 391455 705829 391511
rect 705897 391455 705953 391511
rect 705525 391331 705581 391387
rect 705649 391331 705705 391387
rect 705773 391331 705829 391387
rect 705897 391331 705953 391387
rect 705525 391207 705581 391263
rect 705649 391207 705705 391263
rect 705773 391207 705829 391263
rect 705897 391207 705953 391263
rect 705525 391083 705581 391139
rect 705649 391083 705705 391139
rect 705773 391083 705829 391139
rect 705897 391083 705953 391139
rect 705525 390959 705581 391015
rect 705649 390959 705705 391015
rect 705773 390959 705829 391015
rect 705897 390959 705953 391015
rect 705525 390835 705581 390891
rect 705649 390835 705705 390891
rect 705773 390835 705829 390891
rect 705897 390835 705953 390891
rect 705525 390711 705581 390767
rect 705649 390711 705705 390767
rect 705773 390711 705829 390767
rect 705897 390711 705953 390767
rect 705525 390587 705581 390643
rect 705649 390587 705705 390643
rect 705773 390587 705829 390643
rect 705897 390587 705953 390643
rect 705525 390463 705581 390519
rect 705649 390463 705705 390519
rect 705773 390463 705829 390519
rect 705897 390463 705953 390519
rect 705525 390339 705581 390395
rect 705649 390339 705705 390395
rect 705773 390339 705829 390395
rect 705897 390339 705953 390395
rect 70047 140605 70103 140661
rect 70171 140605 70227 140661
rect 70295 140605 70351 140661
rect 70419 140605 70475 140661
rect 70047 140481 70103 140537
rect 70171 140481 70227 140537
rect 70295 140481 70351 140537
rect 70419 140481 70475 140537
rect 70047 140357 70103 140413
rect 70171 140357 70227 140413
rect 70295 140357 70351 140413
rect 70419 140357 70475 140413
rect 70047 140233 70103 140289
rect 70171 140233 70227 140289
rect 70295 140233 70351 140289
rect 70419 140233 70475 140289
rect 70047 140109 70103 140165
rect 70171 140109 70227 140165
rect 70295 140109 70351 140165
rect 70419 140109 70475 140165
rect 70047 139985 70103 140041
rect 70171 139985 70227 140041
rect 70295 139985 70351 140041
rect 70419 139985 70475 140041
rect 70047 139861 70103 139917
rect 70171 139861 70227 139917
rect 70295 139861 70351 139917
rect 70419 139861 70475 139917
rect 70047 139737 70103 139793
rect 70171 139737 70227 139793
rect 70295 139737 70351 139793
rect 70419 139737 70475 139793
rect 70047 139613 70103 139669
rect 70171 139613 70227 139669
rect 70295 139613 70351 139669
rect 70419 139613 70475 139669
rect 70047 139489 70103 139545
rect 70171 139489 70227 139545
rect 70295 139489 70351 139545
rect 70419 139489 70475 139545
rect 70047 139365 70103 139421
rect 70171 139365 70227 139421
rect 70295 139365 70351 139421
rect 70419 139365 70475 139421
rect 70047 139241 70103 139297
rect 70171 139241 70227 139297
rect 70295 139241 70351 139297
rect 70419 139241 70475 139297
rect 70047 139117 70103 139173
rect 70171 139117 70227 139173
rect 70295 139117 70351 139173
rect 70419 139117 70475 139173
rect 70047 138993 70103 139049
rect 70171 138993 70227 139049
rect 70295 138993 70351 139049
rect 70419 138993 70475 139049
rect 70047 138869 70103 138925
rect 70171 138869 70227 138925
rect 70295 138869 70351 138925
rect 70419 138869 70475 138925
rect 70047 138125 70103 138181
rect 70171 138125 70227 138181
rect 70295 138125 70351 138181
rect 70419 138125 70475 138181
rect 70047 138001 70103 138057
rect 70171 138001 70227 138057
rect 70295 138001 70351 138057
rect 70419 138001 70475 138057
rect 70047 137877 70103 137933
rect 70171 137877 70227 137933
rect 70295 137877 70351 137933
rect 70419 137877 70475 137933
rect 70047 137753 70103 137809
rect 70171 137753 70227 137809
rect 70295 137753 70351 137809
rect 70419 137753 70475 137809
rect 70047 137629 70103 137685
rect 70171 137629 70227 137685
rect 70295 137629 70351 137685
rect 70419 137629 70475 137685
rect 70047 137505 70103 137561
rect 70171 137505 70227 137561
rect 70295 137505 70351 137561
rect 70419 137505 70475 137561
rect 70047 137381 70103 137437
rect 70171 137381 70227 137437
rect 70295 137381 70351 137437
rect 70419 137381 70475 137437
rect 70047 137257 70103 137313
rect 70171 137257 70227 137313
rect 70295 137257 70351 137313
rect 70419 137257 70475 137313
rect 70047 137133 70103 137189
rect 70171 137133 70227 137189
rect 70295 137133 70351 137189
rect 70419 137133 70475 137189
rect 70047 137009 70103 137065
rect 70171 137009 70227 137065
rect 70295 137009 70351 137065
rect 70419 137009 70475 137065
rect 70047 136885 70103 136941
rect 70171 136885 70227 136941
rect 70295 136885 70351 136941
rect 70419 136885 70475 136941
rect 70047 136761 70103 136817
rect 70171 136761 70227 136817
rect 70295 136761 70351 136817
rect 70419 136761 70475 136817
rect 70047 136637 70103 136693
rect 70171 136637 70227 136693
rect 70295 136637 70351 136693
rect 70419 136637 70475 136693
rect 70047 136513 70103 136569
rect 70171 136513 70227 136569
rect 70295 136513 70351 136569
rect 70419 136513 70475 136569
rect 70047 136389 70103 136445
rect 70171 136389 70227 136445
rect 70295 136389 70351 136445
rect 70419 136389 70475 136445
rect 70047 136265 70103 136321
rect 70171 136265 70227 136321
rect 70295 136265 70351 136321
rect 70419 136265 70475 136321
rect 70047 135755 70103 135811
rect 70171 135755 70227 135811
rect 70295 135755 70351 135811
rect 70419 135755 70475 135811
rect 70047 135631 70103 135687
rect 70171 135631 70227 135687
rect 70295 135631 70351 135687
rect 70419 135631 70475 135687
rect 70047 135507 70103 135563
rect 70171 135507 70227 135563
rect 70295 135507 70351 135563
rect 70419 135507 70475 135563
rect 70047 135383 70103 135439
rect 70171 135383 70227 135439
rect 70295 135383 70351 135439
rect 70419 135383 70475 135439
rect 70047 135259 70103 135315
rect 70171 135259 70227 135315
rect 70295 135259 70351 135315
rect 70419 135259 70475 135315
rect 70047 135135 70103 135191
rect 70171 135135 70227 135191
rect 70295 135135 70351 135191
rect 70419 135135 70475 135191
rect 70047 135011 70103 135067
rect 70171 135011 70227 135067
rect 70295 135011 70351 135067
rect 70419 135011 70475 135067
rect 70047 134887 70103 134943
rect 70171 134887 70227 134943
rect 70295 134887 70351 134943
rect 70419 134887 70475 134943
rect 70047 134763 70103 134819
rect 70171 134763 70227 134819
rect 70295 134763 70351 134819
rect 70419 134763 70475 134819
rect 70047 134639 70103 134695
rect 70171 134639 70227 134695
rect 70295 134639 70351 134695
rect 70419 134639 70475 134695
rect 70047 134515 70103 134571
rect 70171 134515 70227 134571
rect 70295 134515 70351 134571
rect 70419 134515 70475 134571
rect 70047 134391 70103 134447
rect 70171 134391 70227 134447
rect 70295 134391 70351 134447
rect 70419 134391 70475 134447
rect 70047 134267 70103 134323
rect 70171 134267 70227 134323
rect 70295 134267 70351 134323
rect 70419 134267 70475 134323
rect 70047 134143 70103 134199
rect 70171 134143 70227 134199
rect 70295 134143 70351 134199
rect 70419 134143 70475 134199
rect 70047 134019 70103 134075
rect 70171 134019 70227 134075
rect 70295 134019 70351 134075
rect 70419 134019 70475 134075
rect 70047 133895 70103 133951
rect 70171 133895 70227 133951
rect 70295 133895 70351 133951
rect 70419 133895 70475 133951
rect 70047 133049 70103 133105
rect 70171 133049 70227 133105
rect 70295 133049 70351 133105
rect 70419 133049 70475 133105
rect 70047 132925 70103 132981
rect 70171 132925 70227 132981
rect 70295 132925 70351 132981
rect 70419 132925 70475 132981
rect 70047 132801 70103 132857
rect 70171 132801 70227 132857
rect 70295 132801 70351 132857
rect 70419 132801 70475 132857
rect 70047 132677 70103 132733
rect 70171 132677 70227 132733
rect 70295 132677 70351 132733
rect 70419 132677 70475 132733
rect 70047 132553 70103 132609
rect 70171 132553 70227 132609
rect 70295 132553 70351 132609
rect 70419 132553 70475 132609
rect 70047 132429 70103 132485
rect 70171 132429 70227 132485
rect 70295 132429 70351 132485
rect 70419 132429 70475 132485
rect 70047 132305 70103 132361
rect 70171 132305 70227 132361
rect 70295 132305 70351 132361
rect 70419 132305 70475 132361
rect 70047 132181 70103 132237
rect 70171 132181 70227 132237
rect 70295 132181 70351 132237
rect 70419 132181 70475 132237
rect 70047 132057 70103 132113
rect 70171 132057 70227 132113
rect 70295 132057 70351 132113
rect 70419 132057 70475 132113
rect 70047 131933 70103 131989
rect 70171 131933 70227 131989
rect 70295 131933 70351 131989
rect 70419 131933 70475 131989
rect 70047 131809 70103 131865
rect 70171 131809 70227 131865
rect 70295 131809 70351 131865
rect 70419 131809 70475 131865
rect 70047 131685 70103 131741
rect 70171 131685 70227 131741
rect 70295 131685 70351 131741
rect 70419 131685 70475 131741
rect 70047 131561 70103 131617
rect 70171 131561 70227 131617
rect 70295 131561 70351 131617
rect 70419 131561 70475 131617
rect 70047 131437 70103 131493
rect 70171 131437 70227 131493
rect 70295 131437 70351 131493
rect 70419 131437 70475 131493
rect 70047 131313 70103 131369
rect 70171 131313 70227 131369
rect 70295 131313 70351 131369
rect 70419 131313 70475 131369
rect 70047 131189 70103 131245
rect 70171 131189 70227 131245
rect 70295 131189 70351 131245
rect 70419 131189 70475 131245
rect 70047 130679 70103 130735
rect 70171 130679 70227 130735
rect 70295 130679 70351 130735
rect 70419 130679 70475 130735
rect 70047 130555 70103 130611
rect 70171 130555 70227 130611
rect 70295 130555 70351 130611
rect 70419 130555 70475 130611
rect 70047 130431 70103 130487
rect 70171 130431 70227 130487
rect 70295 130431 70351 130487
rect 70419 130431 70475 130487
rect 70047 130307 70103 130363
rect 70171 130307 70227 130363
rect 70295 130307 70351 130363
rect 70419 130307 70475 130363
rect 70047 130183 70103 130239
rect 70171 130183 70227 130239
rect 70295 130183 70351 130239
rect 70419 130183 70475 130239
rect 70047 130059 70103 130115
rect 70171 130059 70227 130115
rect 70295 130059 70351 130115
rect 70419 130059 70475 130115
rect 70047 129935 70103 129991
rect 70171 129935 70227 129991
rect 70295 129935 70351 129991
rect 70419 129935 70475 129991
rect 70047 129811 70103 129867
rect 70171 129811 70227 129867
rect 70295 129811 70351 129867
rect 70419 129811 70475 129867
rect 70047 129687 70103 129743
rect 70171 129687 70227 129743
rect 70295 129687 70351 129743
rect 70419 129687 70475 129743
rect 70047 129563 70103 129619
rect 70171 129563 70227 129619
rect 70295 129563 70351 129619
rect 70419 129563 70475 129619
rect 70047 129439 70103 129495
rect 70171 129439 70227 129495
rect 70295 129439 70351 129495
rect 70419 129439 70475 129495
rect 70047 129315 70103 129371
rect 70171 129315 70227 129371
rect 70295 129315 70351 129371
rect 70419 129315 70475 129371
rect 70047 129191 70103 129247
rect 70171 129191 70227 129247
rect 70295 129191 70351 129247
rect 70419 129191 70475 129247
rect 70047 129067 70103 129123
rect 70171 129067 70227 129123
rect 70295 129067 70351 129123
rect 70419 129067 70475 129123
rect 70047 128943 70103 128999
rect 70171 128943 70227 128999
rect 70295 128943 70351 128999
rect 70419 128943 70475 128999
rect 70047 128819 70103 128875
rect 70171 128819 70227 128875
rect 70295 128819 70351 128875
rect 70419 128819 70475 128875
rect 70047 128049 70103 128105
rect 70171 128049 70227 128105
rect 70295 128049 70351 128105
rect 70419 128049 70475 128105
rect 70047 127925 70103 127981
rect 70171 127925 70227 127981
rect 70295 127925 70351 127981
rect 70419 127925 70475 127981
rect 70047 127801 70103 127857
rect 70171 127801 70227 127857
rect 70295 127801 70351 127857
rect 70419 127801 70475 127857
rect 70047 127677 70103 127733
rect 70171 127677 70227 127733
rect 70295 127677 70351 127733
rect 70419 127677 70475 127733
rect 70047 127553 70103 127609
rect 70171 127553 70227 127609
rect 70295 127553 70351 127609
rect 70419 127553 70475 127609
rect 70047 127429 70103 127485
rect 70171 127429 70227 127485
rect 70295 127429 70351 127485
rect 70419 127429 70475 127485
rect 70047 127305 70103 127361
rect 70171 127305 70227 127361
rect 70295 127305 70351 127361
rect 70419 127305 70475 127361
rect 70047 127181 70103 127237
rect 70171 127181 70227 127237
rect 70295 127181 70351 127237
rect 70419 127181 70475 127237
rect 70047 127057 70103 127113
rect 70171 127057 70227 127113
rect 70295 127057 70351 127113
rect 70419 127057 70475 127113
rect 70047 126933 70103 126989
rect 70171 126933 70227 126989
rect 70295 126933 70351 126989
rect 70419 126933 70475 126989
rect 70047 126809 70103 126865
rect 70171 126809 70227 126865
rect 70295 126809 70351 126865
rect 70419 126809 70475 126865
rect 70047 126685 70103 126741
rect 70171 126685 70227 126741
rect 70295 126685 70351 126741
rect 70419 126685 70475 126741
rect 70047 126561 70103 126617
rect 70171 126561 70227 126617
rect 70295 126561 70351 126617
rect 70419 126561 70475 126617
rect 70047 126437 70103 126493
rect 70171 126437 70227 126493
rect 70295 126437 70351 126493
rect 70419 126437 70475 126493
rect 70047 126313 70103 126369
rect 70171 126313 70227 126369
rect 70295 126313 70351 126369
rect 70419 126313 70475 126369
rect 70047 99605 70103 99661
rect 70171 99605 70227 99661
rect 70295 99605 70351 99661
rect 70419 99605 70475 99661
rect 70047 99481 70103 99537
rect 70171 99481 70227 99537
rect 70295 99481 70351 99537
rect 70419 99481 70475 99537
rect 70047 99357 70103 99413
rect 70171 99357 70227 99413
rect 70295 99357 70351 99413
rect 70419 99357 70475 99413
rect 70047 99233 70103 99289
rect 70171 99233 70227 99289
rect 70295 99233 70351 99289
rect 70419 99233 70475 99289
rect 70047 99109 70103 99165
rect 70171 99109 70227 99165
rect 70295 99109 70351 99165
rect 70419 99109 70475 99165
rect 70047 98985 70103 99041
rect 70171 98985 70227 99041
rect 70295 98985 70351 99041
rect 70419 98985 70475 99041
rect 70047 98861 70103 98917
rect 70171 98861 70227 98917
rect 70295 98861 70351 98917
rect 70419 98861 70475 98917
rect 70047 98737 70103 98793
rect 70171 98737 70227 98793
rect 70295 98737 70351 98793
rect 70419 98737 70475 98793
rect 70047 98613 70103 98669
rect 70171 98613 70227 98669
rect 70295 98613 70351 98669
rect 70419 98613 70475 98669
rect 70047 98489 70103 98545
rect 70171 98489 70227 98545
rect 70295 98489 70351 98545
rect 70419 98489 70475 98545
rect 70047 98365 70103 98421
rect 70171 98365 70227 98421
rect 70295 98365 70351 98421
rect 70419 98365 70475 98421
rect 70047 98241 70103 98297
rect 70171 98241 70227 98297
rect 70295 98241 70351 98297
rect 70419 98241 70475 98297
rect 70047 98117 70103 98173
rect 70171 98117 70227 98173
rect 70295 98117 70351 98173
rect 70419 98117 70475 98173
rect 70047 97993 70103 98049
rect 70171 97993 70227 98049
rect 70295 97993 70351 98049
rect 70419 97993 70475 98049
rect 70047 97869 70103 97925
rect 70171 97869 70227 97925
rect 70295 97869 70351 97925
rect 70419 97869 70475 97925
rect 70047 97125 70103 97181
rect 70171 97125 70227 97181
rect 70295 97125 70351 97181
rect 70419 97125 70475 97181
rect 70047 97001 70103 97057
rect 70171 97001 70227 97057
rect 70295 97001 70351 97057
rect 70419 97001 70475 97057
rect 70047 96877 70103 96933
rect 70171 96877 70227 96933
rect 70295 96877 70351 96933
rect 70419 96877 70475 96933
rect 70047 96753 70103 96809
rect 70171 96753 70227 96809
rect 70295 96753 70351 96809
rect 70419 96753 70475 96809
rect 70047 96629 70103 96685
rect 70171 96629 70227 96685
rect 70295 96629 70351 96685
rect 70419 96629 70475 96685
rect 70047 96505 70103 96561
rect 70171 96505 70227 96561
rect 70295 96505 70351 96561
rect 70419 96505 70475 96561
rect 70047 96381 70103 96437
rect 70171 96381 70227 96437
rect 70295 96381 70351 96437
rect 70419 96381 70475 96437
rect 70047 96257 70103 96313
rect 70171 96257 70227 96313
rect 70295 96257 70351 96313
rect 70419 96257 70475 96313
rect 70047 96133 70103 96189
rect 70171 96133 70227 96189
rect 70295 96133 70351 96189
rect 70419 96133 70475 96189
rect 70047 96009 70103 96065
rect 70171 96009 70227 96065
rect 70295 96009 70351 96065
rect 70419 96009 70475 96065
rect 70047 95885 70103 95941
rect 70171 95885 70227 95941
rect 70295 95885 70351 95941
rect 70419 95885 70475 95941
rect 70047 95761 70103 95817
rect 70171 95761 70227 95817
rect 70295 95761 70351 95817
rect 70419 95761 70475 95817
rect 70047 95637 70103 95693
rect 70171 95637 70227 95693
rect 70295 95637 70351 95693
rect 70419 95637 70475 95693
rect 70047 95513 70103 95569
rect 70171 95513 70227 95569
rect 70295 95513 70351 95569
rect 70419 95513 70475 95569
rect 70047 95389 70103 95445
rect 70171 95389 70227 95445
rect 70295 95389 70351 95445
rect 70419 95389 70475 95445
rect 70047 95265 70103 95321
rect 70171 95265 70227 95321
rect 70295 95265 70351 95321
rect 70419 95265 70475 95321
rect 70047 94755 70103 94811
rect 70171 94755 70227 94811
rect 70295 94755 70351 94811
rect 70419 94755 70475 94811
rect 70047 94631 70103 94687
rect 70171 94631 70227 94687
rect 70295 94631 70351 94687
rect 70419 94631 70475 94687
rect 70047 94507 70103 94563
rect 70171 94507 70227 94563
rect 70295 94507 70351 94563
rect 70419 94507 70475 94563
rect 70047 94383 70103 94439
rect 70171 94383 70227 94439
rect 70295 94383 70351 94439
rect 70419 94383 70475 94439
rect 70047 94259 70103 94315
rect 70171 94259 70227 94315
rect 70295 94259 70351 94315
rect 70419 94259 70475 94315
rect 70047 94135 70103 94191
rect 70171 94135 70227 94191
rect 70295 94135 70351 94191
rect 70419 94135 70475 94191
rect 70047 94011 70103 94067
rect 70171 94011 70227 94067
rect 70295 94011 70351 94067
rect 70419 94011 70475 94067
rect 70047 93887 70103 93943
rect 70171 93887 70227 93943
rect 70295 93887 70351 93943
rect 70419 93887 70475 93943
rect 70047 93763 70103 93819
rect 70171 93763 70227 93819
rect 70295 93763 70351 93819
rect 70419 93763 70475 93819
rect 70047 93639 70103 93695
rect 70171 93639 70227 93695
rect 70295 93639 70351 93695
rect 70419 93639 70475 93695
rect 70047 93515 70103 93571
rect 70171 93515 70227 93571
rect 70295 93515 70351 93571
rect 70419 93515 70475 93571
rect 70047 93391 70103 93447
rect 70171 93391 70227 93447
rect 70295 93391 70351 93447
rect 70419 93391 70475 93447
rect 70047 93267 70103 93323
rect 70171 93267 70227 93323
rect 70295 93267 70351 93323
rect 70419 93267 70475 93323
rect 70047 93143 70103 93199
rect 70171 93143 70227 93199
rect 70295 93143 70351 93199
rect 70419 93143 70475 93199
rect 70047 93019 70103 93075
rect 70171 93019 70227 93075
rect 70295 93019 70351 93075
rect 70419 93019 70475 93075
rect 70047 92895 70103 92951
rect 70171 92895 70227 92951
rect 70295 92895 70351 92951
rect 70419 92895 70475 92951
rect 70047 92049 70103 92105
rect 70171 92049 70227 92105
rect 70295 92049 70351 92105
rect 70419 92049 70475 92105
rect 70047 91925 70103 91981
rect 70171 91925 70227 91981
rect 70295 91925 70351 91981
rect 70419 91925 70475 91981
rect 70047 91801 70103 91857
rect 70171 91801 70227 91857
rect 70295 91801 70351 91857
rect 70419 91801 70475 91857
rect 70047 91677 70103 91733
rect 70171 91677 70227 91733
rect 70295 91677 70351 91733
rect 70419 91677 70475 91733
rect 70047 91553 70103 91609
rect 70171 91553 70227 91609
rect 70295 91553 70351 91609
rect 70419 91553 70475 91609
rect 70047 91429 70103 91485
rect 70171 91429 70227 91485
rect 70295 91429 70351 91485
rect 70419 91429 70475 91485
rect 70047 91305 70103 91361
rect 70171 91305 70227 91361
rect 70295 91305 70351 91361
rect 70419 91305 70475 91361
rect 70047 91181 70103 91237
rect 70171 91181 70227 91237
rect 70295 91181 70351 91237
rect 70419 91181 70475 91237
rect 70047 91057 70103 91113
rect 70171 91057 70227 91113
rect 70295 91057 70351 91113
rect 70419 91057 70475 91113
rect 70047 90933 70103 90989
rect 70171 90933 70227 90989
rect 70295 90933 70351 90989
rect 70419 90933 70475 90989
rect 70047 90809 70103 90865
rect 70171 90809 70227 90865
rect 70295 90809 70351 90865
rect 70419 90809 70475 90865
rect 70047 90685 70103 90741
rect 70171 90685 70227 90741
rect 70295 90685 70351 90741
rect 70419 90685 70475 90741
rect 70047 90561 70103 90617
rect 70171 90561 70227 90617
rect 70295 90561 70351 90617
rect 70419 90561 70475 90617
rect 70047 90437 70103 90493
rect 70171 90437 70227 90493
rect 70295 90437 70351 90493
rect 70419 90437 70475 90493
rect 70047 90313 70103 90369
rect 70171 90313 70227 90369
rect 70295 90313 70351 90369
rect 70419 90313 70475 90369
rect 70047 90189 70103 90245
rect 70171 90189 70227 90245
rect 70295 90189 70351 90245
rect 70419 90189 70475 90245
rect 70047 89679 70103 89735
rect 70171 89679 70227 89735
rect 70295 89679 70351 89735
rect 70419 89679 70475 89735
rect 70047 89555 70103 89611
rect 70171 89555 70227 89611
rect 70295 89555 70351 89611
rect 70419 89555 70475 89611
rect 70047 89431 70103 89487
rect 70171 89431 70227 89487
rect 70295 89431 70351 89487
rect 70419 89431 70475 89487
rect 70047 89307 70103 89363
rect 70171 89307 70227 89363
rect 70295 89307 70351 89363
rect 70419 89307 70475 89363
rect 70047 89183 70103 89239
rect 70171 89183 70227 89239
rect 70295 89183 70351 89239
rect 70419 89183 70475 89239
rect 70047 89059 70103 89115
rect 70171 89059 70227 89115
rect 70295 89059 70351 89115
rect 70419 89059 70475 89115
rect 70047 88935 70103 88991
rect 70171 88935 70227 88991
rect 70295 88935 70351 88991
rect 70419 88935 70475 88991
rect 70047 88811 70103 88867
rect 70171 88811 70227 88867
rect 70295 88811 70351 88867
rect 70419 88811 70475 88867
rect 70047 88687 70103 88743
rect 70171 88687 70227 88743
rect 70295 88687 70351 88743
rect 70419 88687 70475 88743
rect 70047 88563 70103 88619
rect 70171 88563 70227 88619
rect 70295 88563 70351 88619
rect 70419 88563 70475 88619
rect 70047 88439 70103 88495
rect 70171 88439 70227 88495
rect 70295 88439 70351 88495
rect 70419 88439 70475 88495
rect 70047 88315 70103 88371
rect 70171 88315 70227 88371
rect 70295 88315 70351 88371
rect 70419 88315 70475 88371
rect 70047 88191 70103 88247
rect 70171 88191 70227 88247
rect 70295 88191 70351 88247
rect 70419 88191 70475 88247
rect 70047 88067 70103 88123
rect 70171 88067 70227 88123
rect 70295 88067 70351 88123
rect 70419 88067 70475 88123
rect 70047 87943 70103 87999
rect 70171 87943 70227 87999
rect 70295 87943 70351 87999
rect 70419 87943 70475 87999
rect 70047 87819 70103 87875
rect 70171 87819 70227 87875
rect 70295 87819 70351 87875
rect 70419 87819 70475 87875
rect 70047 87049 70103 87105
rect 70171 87049 70227 87105
rect 70295 87049 70351 87105
rect 70419 87049 70475 87105
rect 70047 86925 70103 86981
rect 70171 86925 70227 86981
rect 70295 86925 70351 86981
rect 70419 86925 70475 86981
rect 70047 86801 70103 86857
rect 70171 86801 70227 86857
rect 70295 86801 70351 86857
rect 70419 86801 70475 86857
rect 70047 86677 70103 86733
rect 70171 86677 70227 86733
rect 70295 86677 70351 86733
rect 70419 86677 70475 86733
rect 70047 86553 70103 86609
rect 70171 86553 70227 86609
rect 70295 86553 70351 86609
rect 70419 86553 70475 86609
rect 70047 86429 70103 86485
rect 70171 86429 70227 86485
rect 70295 86429 70351 86485
rect 70419 86429 70475 86485
rect 70047 86305 70103 86361
rect 70171 86305 70227 86361
rect 70295 86305 70351 86361
rect 70419 86305 70475 86361
rect 70047 86181 70103 86237
rect 70171 86181 70227 86237
rect 70295 86181 70351 86237
rect 70419 86181 70475 86237
rect 70047 86057 70103 86113
rect 70171 86057 70227 86113
rect 70295 86057 70351 86113
rect 70419 86057 70475 86113
rect 70047 85933 70103 85989
rect 70171 85933 70227 85989
rect 70295 85933 70351 85989
rect 70419 85933 70475 85989
rect 70047 85809 70103 85865
rect 70171 85809 70227 85865
rect 70295 85809 70351 85865
rect 70419 85809 70475 85865
rect 70047 85685 70103 85741
rect 70171 85685 70227 85741
rect 70295 85685 70351 85741
rect 70419 85685 70475 85741
rect 70047 85561 70103 85617
rect 70171 85561 70227 85617
rect 70295 85561 70351 85617
rect 70419 85561 70475 85617
rect 70047 85437 70103 85493
rect 70171 85437 70227 85493
rect 70295 85437 70351 85493
rect 70419 85437 70475 85493
rect 70047 85313 70103 85369
rect 70171 85313 70227 85369
rect 70295 85313 70351 85369
rect 70419 85313 70475 85369
rect 655326 75889 655382 75945
rect 655450 75889 655506 75945
rect 655574 75889 655630 75945
rect 655698 75889 655754 75945
rect 655822 75889 655878 75945
rect 655946 75889 656002 75945
rect 656070 75889 656126 75945
rect 656194 75889 656250 75945
rect 656318 75889 656374 75945
rect 655326 75765 655382 75821
rect 655450 75765 655506 75821
rect 655574 75765 655630 75821
rect 655698 75765 655754 75821
rect 655822 75765 655878 75821
rect 655946 75765 656002 75821
rect 656070 75765 656126 75821
rect 656194 75765 656250 75821
rect 656318 75765 656374 75821
rect 655326 75641 655382 75697
rect 655450 75641 655506 75697
rect 655574 75641 655630 75697
rect 655698 75641 655754 75697
rect 655822 75641 655878 75697
rect 655946 75641 656002 75697
rect 656070 75641 656126 75697
rect 656194 75641 656250 75697
rect 656318 75641 656374 75697
rect 655326 75517 655382 75573
rect 655450 75517 655506 75573
rect 655574 75517 655630 75573
rect 655698 75517 655754 75573
rect 655822 75517 655878 75573
rect 655946 75517 656002 75573
rect 656070 75517 656126 75573
rect 656194 75517 656250 75573
rect 656318 75517 656374 75573
rect 655326 75393 655382 75449
rect 655450 75393 655506 75449
rect 655574 75393 655630 75449
rect 655698 75393 655754 75449
rect 655822 75393 655878 75449
rect 655946 75393 656002 75449
rect 656070 75393 656126 75449
rect 656194 75393 656250 75449
rect 656318 75393 656374 75449
rect 655326 75269 655382 75325
rect 655450 75269 655506 75325
rect 655574 75269 655630 75325
rect 655698 75269 655754 75325
rect 655822 75269 655878 75325
rect 655946 75269 656002 75325
rect 656070 75269 656126 75325
rect 656194 75269 656250 75325
rect 656318 75269 656374 75325
rect 655326 75145 655382 75201
rect 655450 75145 655506 75201
rect 655574 75145 655630 75201
rect 655698 75145 655754 75201
rect 655822 75145 655878 75201
rect 655946 75145 656002 75201
rect 656070 75145 656126 75201
rect 656194 75145 656250 75201
rect 656318 75145 656374 75201
rect 655326 75021 655382 75077
rect 655450 75021 655506 75077
rect 655574 75021 655630 75077
rect 655698 75021 655754 75077
rect 655822 75021 655878 75077
rect 655946 75021 656002 75077
rect 656070 75021 656126 75077
rect 656194 75021 656250 75077
rect 656318 75021 656374 75077
rect 655326 74897 655382 74953
rect 655450 74897 655506 74953
rect 655574 74897 655630 74953
rect 655698 74897 655754 74953
rect 655822 74897 655878 74953
rect 655946 74897 656002 74953
rect 656070 74897 656126 74953
rect 656194 74897 656250 74953
rect 656318 74897 656374 74953
rect 655326 74773 655382 74829
rect 655450 74773 655506 74829
rect 655574 74773 655630 74829
rect 655698 74773 655754 74829
rect 655822 74773 655878 74829
rect 655946 74773 656002 74829
rect 656070 74773 656126 74829
rect 656194 74773 656250 74829
rect 656318 74773 656374 74829
rect 655326 74649 655382 74705
rect 655450 74649 655506 74705
rect 655574 74649 655630 74705
rect 655698 74649 655754 74705
rect 655822 74649 655878 74705
rect 655946 74649 656002 74705
rect 656070 74649 656126 74705
rect 656194 74649 656250 74705
rect 656318 74649 656374 74705
rect 655326 74525 655382 74581
rect 655450 74525 655506 74581
rect 655574 74525 655630 74581
rect 655698 74525 655754 74581
rect 655822 74525 655878 74581
rect 655946 74525 656002 74581
rect 656070 74525 656126 74581
rect 656194 74525 656250 74581
rect 656318 74525 656374 74581
rect 105326 73889 105382 73945
rect 105450 73889 105506 73945
rect 105574 73889 105630 73945
rect 105698 73889 105754 73945
rect 105822 73889 105878 73945
rect 105946 73889 106002 73945
rect 106070 73889 106126 73945
rect 106194 73889 106250 73945
rect 106318 73889 106374 73945
rect 106442 73889 106498 73945
rect 106566 73889 106622 73945
rect 106690 73889 106746 73945
rect 106814 73889 106870 73945
rect 106938 73889 106994 73945
rect 107062 73889 107118 73945
rect 105326 73765 105382 73821
rect 105450 73765 105506 73821
rect 105574 73765 105630 73821
rect 105698 73765 105754 73821
rect 105822 73765 105878 73821
rect 105946 73765 106002 73821
rect 106070 73765 106126 73821
rect 106194 73765 106250 73821
rect 106318 73765 106374 73821
rect 106442 73765 106498 73821
rect 106566 73765 106622 73821
rect 106690 73765 106746 73821
rect 106814 73765 106870 73821
rect 106938 73765 106994 73821
rect 107062 73765 107118 73821
rect 105326 73641 105382 73697
rect 105450 73641 105506 73697
rect 105574 73641 105630 73697
rect 105698 73641 105754 73697
rect 105822 73641 105878 73697
rect 105946 73641 106002 73697
rect 106070 73641 106126 73697
rect 106194 73641 106250 73697
rect 106318 73641 106374 73697
rect 106442 73641 106498 73697
rect 106566 73641 106622 73697
rect 106690 73641 106746 73697
rect 106814 73641 106870 73697
rect 106938 73641 106994 73697
rect 107062 73641 107118 73697
rect 105326 73517 105382 73573
rect 105450 73517 105506 73573
rect 105574 73517 105630 73573
rect 105698 73517 105754 73573
rect 105822 73517 105878 73573
rect 105946 73517 106002 73573
rect 106070 73517 106126 73573
rect 106194 73517 106250 73573
rect 106318 73517 106374 73573
rect 106442 73517 106498 73573
rect 106566 73517 106622 73573
rect 106690 73517 106746 73573
rect 106814 73517 106870 73573
rect 106938 73517 106994 73573
rect 107062 73517 107118 73573
rect 105326 73393 105382 73449
rect 105450 73393 105506 73449
rect 105574 73393 105630 73449
rect 105698 73393 105754 73449
rect 105822 73393 105878 73449
rect 105946 73393 106002 73449
rect 106070 73393 106126 73449
rect 106194 73393 106250 73449
rect 106318 73393 106374 73449
rect 106442 73393 106498 73449
rect 106566 73393 106622 73449
rect 106690 73393 106746 73449
rect 106814 73393 106870 73449
rect 106938 73393 106994 73449
rect 107062 73393 107118 73449
rect 105326 73269 105382 73325
rect 105450 73269 105506 73325
rect 105574 73269 105630 73325
rect 105698 73269 105754 73325
rect 105822 73269 105878 73325
rect 105946 73269 106002 73325
rect 106070 73269 106126 73325
rect 106194 73269 106250 73325
rect 106318 73269 106374 73325
rect 106442 73269 106498 73325
rect 106566 73269 106622 73325
rect 106690 73269 106746 73325
rect 106814 73269 106870 73325
rect 106938 73269 106994 73325
rect 107062 73269 107118 73325
rect 105326 73145 105382 73201
rect 105450 73145 105506 73201
rect 105574 73145 105630 73201
rect 105698 73145 105754 73201
rect 105822 73145 105878 73201
rect 105946 73145 106002 73201
rect 106070 73145 106126 73201
rect 106194 73145 106250 73201
rect 106318 73145 106374 73201
rect 106442 73145 106498 73201
rect 106566 73145 106622 73201
rect 106690 73145 106746 73201
rect 106814 73145 106870 73201
rect 106938 73145 106994 73201
rect 107062 73145 107118 73201
rect 105326 73021 105382 73077
rect 105450 73021 105506 73077
rect 105574 73021 105630 73077
rect 105698 73021 105754 73077
rect 105822 73021 105878 73077
rect 105946 73021 106002 73077
rect 106070 73021 106126 73077
rect 106194 73021 106250 73077
rect 106318 73021 106374 73077
rect 106442 73021 106498 73077
rect 106566 73021 106622 73077
rect 106690 73021 106746 73077
rect 106814 73021 106870 73077
rect 106938 73021 106994 73077
rect 107062 73021 107118 73077
rect 105326 72897 105382 72953
rect 105450 72897 105506 72953
rect 105574 72897 105630 72953
rect 105698 72897 105754 72953
rect 105822 72897 105878 72953
rect 105946 72897 106002 72953
rect 106070 72897 106126 72953
rect 106194 72897 106250 72953
rect 106318 72897 106374 72953
rect 106442 72897 106498 72953
rect 106566 72897 106622 72953
rect 106690 72897 106746 72953
rect 106814 72897 106870 72953
rect 106938 72897 106994 72953
rect 107062 72897 107118 72953
rect 105326 72773 105382 72829
rect 105450 72773 105506 72829
rect 105574 72773 105630 72829
rect 105698 72773 105754 72829
rect 105822 72773 105878 72829
rect 105946 72773 106002 72829
rect 106070 72773 106126 72829
rect 106194 72773 106250 72829
rect 106318 72773 106374 72829
rect 106442 72773 106498 72829
rect 106566 72773 106622 72829
rect 106690 72773 106746 72829
rect 106814 72773 106870 72829
rect 106938 72773 106994 72829
rect 107062 72773 107118 72829
rect 105326 72649 105382 72705
rect 105450 72649 105506 72705
rect 105574 72649 105630 72705
rect 105698 72649 105754 72705
rect 105822 72649 105878 72705
rect 105946 72649 106002 72705
rect 106070 72649 106126 72705
rect 106194 72649 106250 72705
rect 106318 72649 106374 72705
rect 106442 72649 106498 72705
rect 106566 72649 106622 72705
rect 106690 72649 106746 72705
rect 106814 72649 106870 72705
rect 106938 72649 106994 72705
rect 107062 72649 107118 72705
rect 105326 72525 105382 72581
rect 105450 72525 105506 72581
rect 105574 72525 105630 72581
rect 105698 72525 105754 72581
rect 105822 72525 105878 72581
rect 105946 72525 106002 72581
rect 106070 72525 106126 72581
rect 106194 72525 106250 72581
rect 106318 72525 106374 72581
rect 106442 72525 106498 72581
rect 106566 72525 106622 72581
rect 106690 72525 106746 72581
rect 106814 72525 106870 72581
rect 106938 72525 106994 72581
rect 107062 72525 107118 72581
rect 105326 72401 105382 72457
rect 105450 72401 105506 72457
rect 105574 72401 105630 72457
rect 105698 72401 105754 72457
rect 105822 72401 105878 72457
rect 105946 72401 106002 72457
rect 106070 72401 106126 72457
rect 106194 72401 106250 72457
rect 106318 72401 106374 72457
rect 106442 72401 106498 72457
rect 106566 72401 106622 72457
rect 106690 72401 106746 72457
rect 106814 72401 106870 72457
rect 106938 72401 106994 72457
rect 107062 72401 107118 72457
rect 105326 72277 105382 72333
rect 105450 72277 105506 72333
rect 105574 72277 105630 72333
rect 105698 72277 105754 72333
rect 105822 72277 105878 72333
rect 105946 72277 106002 72333
rect 106070 72277 106126 72333
rect 106194 72277 106250 72333
rect 106318 72277 106374 72333
rect 106442 72277 106498 72333
rect 106566 72277 106622 72333
rect 106690 72277 106746 72333
rect 106814 72277 106870 72333
rect 106938 72277 106994 72333
rect 107062 72277 107118 72333
rect 105326 72153 105382 72209
rect 105450 72153 105506 72209
rect 105574 72153 105630 72209
rect 105698 72153 105754 72209
rect 105822 72153 105878 72209
rect 105946 72153 106002 72209
rect 106070 72153 106126 72209
rect 106194 72153 106250 72209
rect 106318 72153 106374 72209
rect 106442 72153 106498 72209
rect 106566 72153 106622 72209
rect 106690 72153 106746 72209
rect 106814 72153 106870 72209
rect 106938 72153 106994 72209
rect 107062 72153 107118 72209
rect 109046 73889 109102 73945
rect 109170 73889 109226 73945
rect 109294 73889 109350 73945
rect 109418 73889 109474 73945
rect 109542 73889 109598 73945
rect 109666 73889 109722 73945
rect 109046 73765 109102 73821
rect 109170 73765 109226 73821
rect 109294 73765 109350 73821
rect 109418 73765 109474 73821
rect 109542 73765 109598 73821
rect 109666 73765 109722 73821
rect 109046 73641 109102 73697
rect 109170 73641 109226 73697
rect 109294 73641 109350 73697
rect 109418 73641 109474 73697
rect 109542 73641 109598 73697
rect 109666 73641 109722 73697
rect 109046 73517 109102 73573
rect 109170 73517 109226 73573
rect 109294 73517 109350 73573
rect 109418 73517 109474 73573
rect 109542 73517 109598 73573
rect 109666 73517 109722 73573
rect 109046 73393 109102 73449
rect 109170 73393 109226 73449
rect 109294 73393 109350 73449
rect 109418 73393 109474 73449
rect 109542 73393 109598 73449
rect 109666 73393 109722 73449
rect 109046 73269 109102 73325
rect 109170 73269 109226 73325
rect 109294 73269 109350 73325
rect 109418 73269 109474 73325
rect 109542 73269 109598 73325
rect 109666 73269 109722 73325
rect 109046 73145 109102 73201
rect 109170 73145 109226 73201
rect 109294 73145 109350 73201
rect 109418 73145 109474 73201
rect 109542 73145 109598 73201
rect 109666 73145 109722 73201
rect 109046 73021 109102 73077
rect 109170 73021 109226 73077
rect 109294 73021 109350 73077
rect 109418 73021 109474 73077
rect 109542 73021 109598 73077
rect 109666 73021 109722 73077
rect 109046 72897 109102 72953
rect 109170 72897 109226 72953
rect 109294 72897 109350 72953
rect 109418 72897 109474 72953
rect 109542 72897 109598 72953
rect 109666 72897 109722 72953
rect 109046 72773 109102 72829
rect 109170 72773 109226 72829
rect 109294 72773 109350 72829
rect 109418 72773 109474 72829
rect 109542 72773 109598 72829
rect 109666 72773 109722 72829
rect 109046 72649 109102 72705
rect 109170 72649 109226 72705
rect 109294 72649 109350 72705
rect 109418 72649 109474 72705
rect 109542 72649 109598 72705
rect 109666 72649 109722 72705
rect 109046 72525 109102 72581
rect 109170 72525 109226 72581
rect 109294 72525 109350 72581
rect 109418 72525 109474 72581
rect 109542 72525 109598 72581
rect 109666 72525 109722 72581
rect 109046 72401 109102 72457
rect 109170 72401 109226 72457
rect 109294 72401 109350 72457
rect 109418 72401 109474 72457
rect 109542 72401 109598 72457
rect 109666 72401 109722 72457
rect 109046 72277 109102 72333
rect 109170 72277 109226 72333
rect 109294 72277 109350 72333
rect 109418 72277 109474 72333
rect 109542 72277 109598 72333
rect 109666 72277 109722 72333
rect 109046 72153 109102 72209
rect 109170 72153 109226 72209
rect 109294 72153 109350 72209
rect 109418 72153 109474 72209
rect 109542 72153 109598 72209
rect 109666 72153 109722 72209
rect 110176 73889 110232 73945
rect 110300 73889 110356 73945
rect 110424 73889 110480 73945
rect 110548 73889 110604 73945
rect 110672 73889 110728 73945
rect 110796 73889 110852 73945
rect 110920 73889 110976 73945
rect 111044 73889 111100 73945
rect 111168 73889 111224 73945
rect 111292 73889 111348 73945
rect 111416 73889 111472 73945
rect 111540 73889 111596 73945
rect 111664 73889 111720 73945
rect 111788 73889 111844 73945
rect 111912 73889 111968 73945
rect 112036 73889 112092 73945
rect 110176 73765 110232 73821
rect 110300 73765 110356 73821
rect 110424 73765 110480 73821
rect 110548 73765 110604 73821
rect 110672 73765 110728 73821
rect 110796 73765 110852 73821
rect 110920 73765 110976 73821
rect 111044 73765 111100 73821
rect 111168 73765 111224 73821
rect 111292 73765 111348 73821
rect 111416 73765 111472 73821
rect 111540 73765 111596 73821
rect 111664 73765 111720 73821
rect 111788 73765 111844 73821
rect 111912 73765 111968 73821
rect 112036 73765 112092 73821
rect 110176 73641 110232 73697
rect 110300 73641 110356 73697
rect 110424 73641 110480 73697
rect 110548 73641 110604 73697
rect 110672 73641 110728 73697
rect 110796 73641 110852 73697
rect 110920 73641 110976 73697
rect 111044 73641 111100 73697
rect 111168 73641 111224 73697
rect 111292 73641 111348 73697
rect 111416 73641 111472 73697
rect 111540 73641 111596 73697
rect 111664 73641 111720 73697
rect 111788 73641 111844 73697
rect 111912 73641 111968 73697
rect 112036 73641 112092 73697
rect 110176 73517 110232 73573
rect 110300 73517 110356 73573
rect 110424 73517 110480 73573
rect 110548 73517 110604 73573
rect 110672 73517 110728 73573
rect 110796 73517 110852 73573
rect 110920 73517 110976 73573
rect 111044 73517 111100 73573
rect 111168 73517 111224 73573
rect 111292 73517 111348 73573
rect 111416 73517 111472 73573
rect 111540 73517 111596 73573
rect 111664 73517 111720 73573
rect 111788 73517 111844 73573
rect 111912 73517 111968 73573
rect 112036 73517 112092 73573
rect 110176 73393 110232 73449
rect 110300 73393 110356 73449
rect 110424 73393 110480 73449
rect 110548 73393 110604 73449
rect 110672 73393 110728 73449
rect 110796 73393 110852 73449
rect 110920 73393 110976 73449
rect 111044 73393 111100 73449
rect 111168 73393 111224 73449
rect 111292 73393 111348 73449
rect 111416 73393 111472 73449
rect 111540 73393 111596 73449
rect 111664 73393 111720 73449
rect 111788 73393 111844 73449
rect 111912 73393 111968 73449
rect 112036 73393 112092 73449
rect 110176 73269 110232 73325
rect 110300 73269 110356 73325
rect 110424 73269 110480 73325
rect 110548 73269 110604 73325
rect 110672 73269 110728 73325
rect 110796 73269 110852 73325
rect 110920 73269 110976 73325
rect 111044 73269 111100 73325
rect 111168 73269 111224 73325
rect 111292 73269 111348 73325
rect 111416 73269 111472 73325
rect 111540 73269 111596 73325
rect 111664 73269 111720 73325
rect 111788 73269 111844 73325
rect 111912 73269 111968 73325
rect 112036 73269 112092 73325
rect 110176 73145 110232 73201
rect 110300 73145 110356 73201
rect 110424 73145 110480 73201
rect 110548 73145 110604 73201
rect 110672 73145 110728 73201
rect 110796 73145 110852 73201
rect 110920 73145 110976 73201
rect 111044 73145 111100 73201
rect 111168 73145 111224 73201
rect 111292 73145 111348 73201
rect 111416 73145 111472 73201
rect 111540 73145 111596 73201
rect 111664 73145 111720 73201
rect 111788 73145 111844 73201
rect 111912 73145 111968 73201
rect 112036 73145 112092 73201
rect 110176 73021 110232 73077
rect 110300 73021 110356 73077
rect 110424 73021 110480 73077
rect 110548 73021 110604 73077
rect 110672 73021 110728 73077
rect 110796 73021 110852 73077
rect 110920 73021 110976 73077
rect 111044 73021 111100 73077
rect 111168 73021 111224 73077
rect 111292 73021 111348 73077
rect 111416 73021 111472 73077
rect 111540 73021 111596 73077
rect 111664 73021 111720 73077
rect 111788 73021 111844 73077
rect 111912 73021 111968 73077
rect 112036 73021 112092 73077
rect 110176 72897 110232 72953
rect 110300 72897 110356 72953
rect 110424 72897 110480 72953
rect 110548 72897 110604 72953
rect 110672 72897 110728 72953
rect 110796 72897 110852 72953
rect 110920 72897 110976 72953
rect 111044 72897 111100 72953
rect 111168 72897 111224 72953
rect 111292 72897 111348 72953
rect 111416 72897 111472 72953
rect 111540 72897 111596 72953
rect 111664 72897 111720 72953
rect 111788 72897 111844 72953
rect 111912 72897 111968 72953
rect 112036 72897 112092 72953
rect 110176 72773 110232 72829
rect 110300 72773 110356 72829
rect 110424 72773 110480 72829
rect 110548 72773 110604 72829
rect 110672 72773 110728 72829
rect 110796 72773 110852 72829
rect 110920 72773 110976 72829
rect 111044 72773 111100 72829
rect 111168 72773 111224 72829
rect 111292 72773 111348 72829
rect 111416 72773 111472 72829
rect 111540 72773 111596 72829
rect 111664 72773 111720 72829
rect 111788 72773 111844 72829
rect 111912 72773 111968 72829
rect 112036 72773 112092 72829
rect 110176 72649 110232 72705
rect 110300 72649 110356 72705
rect 110424 72649 110480 72705
rect 110548 72649 110604 72705
rect 110672 72649 110728 72705
rect 110796 72649 110852 72705
rect 110920 72649 110976 72705
rect 111044 72649 111100 72705
rect 111168 72649 111224 72705
rect 111292 72649 111348 72705
rect 111416 72649 111472 72705
rect 111540 72649 111596 72705
rect 111664 72649 111720 72705
rect 111788 72649 111844 72705
rect 111912 72649 111968 72705
rect 112036 72649 112092 72705
rect 110176 72525 110232 72581
rect 110300 72525 110356 72581
rect 110424 72525 110480 72581
rect 110548 72525 110604 72581
rect 110672 72525 110728 72581
rect 110796 72525 110852 72581
rect 110920 72525 110976 72581
rect 111044 72525 111100 72581
rect 111168 72525 111224 72581
rect 111292 72525 111348 72581
rect 111416 72525 111472 72581
rect 111540 72525 111596 72581
rect 111664 72525 111720 72581
rect 111788 72525 111844 72581
rect 111912 72525 111968 72581
rect 112036 72525 112092 72581
rect 110176 72401 110232 72457
rect 110300 72401 110356 72457
rect 110424 72401 110480 72457
rect 110548 72401 110604 72457
rect 110672 72401 110728 72457
rect 110796 72401 110852 72457
rect 110920 72401 110976 72457
rect 111044 72401 111100 72457
rect 111168 72401 111224 72457
rect 111292 72401 111348 72457
rect 111416 72401 111472 72457
rect 111540 72401 111596 72457
rect 111664 72401 111720 72457
rect 111788 72401 111844 72457
rect 111912 72401 111968 72457
rect 112036 72401 112092 72457
rect 110176 72277 110232 72333
rect 110300 72277 110356 72333
rect 110424 72277 110480 72333
rect 110548 72277 110604 72333
rect 110672 72277 110728 72333
rect 110796 72277 110852 72333
rect 110920 72277 110976 72333
rect 111044 72277 111100 72333
rect 111168 72277 111224 72333
rect 111292 72277 111348 72333
rect 111416 72277 111472 72333
rect 111540 72277 111596 72333
rect 111664 72277 111720 72333
rect 111788 72277 111844 72333
rect 111912 72277 111968 72333
rect 112036 72277 112092 72333
rect 110176 72153 110232 72209
rect 110300 72153 110356 72209
rect 110424 72153 110480 72209
rect 110548 72153 110604 72209
rect 110672 72153 110728 72209
rect 110796 72153 110852 72209
rect 110920 72153 110976 72209
rect 111044 72153 111100 72209
rect 111168 72153 111224 72209
rect 111292 72153 111348 72209
rect 111416 72153 111472 72209
rect 111540 72153 111596 72209
rect 111664 72153 111720 72209
rect 111788 72153 111844 72209
rect 111912 72153 111968 72209
rect 112036 72153 112092 72209
rect 112882 73889 112938 73945
rect 113006 73889 113062 73945
rect 113130 73889 113186 73945
rect 113254 73889 113310 73945
rect 113378 73889 113434 73945
rect 113502 73889 113558 73945
rect 113626 73889 113682 73945
rect 113750 73889 113806 73945
rect 113874 73889 113930 73945
rect 113998 73889 114054 73945
rect 114122 73889 114178 73945
rect 114246 73889 114302 73945
rect 114370 73889 114426 73945
rect 114494 73889 114550 73945
rect 114618 73889 114674 73945
rect 114742 73889 114798 73945
rect 112882 73765 112938 73821
rect 113006 73765 113062 73821
rect 113130 73765 113186 73821
rect 113254 73765 113310 73821
rect 113378 73765 113434 73821
rect 113502 73765 113558 73821
rect 113626 73765 113682 73821
rect 113750 73765 113806 73821
rect 113874 73765 113930 73821
rect 113998 73765 114054 73821
rect 114122 73765 114178 73821
rect 114246 73765 114302 73821
rect 114370 73765 114426 73821
rect 114494 73765 114550 73821
rect 114618 73765 114674 73821
rect 114742 73765 114798 73821
rect 112882 73641 112938 73697
rect 113006 73641 113062 73697
rect 113130 73641 113186 73697
rect 113254 73641 113310 73697
rect 113378 73641 113434 73697
rect 113502 73641 113558 73697
rect 113626 73641 113682 73697
rect 113750 73641 113806 73697
rect 113874 73641 113930 73697
rect 113998 73641 114054 73697
rect 114122 73641 114178 73697
rect 114246 73641 114302 73697
rect 114370 73641 114426 73697
rect 114494 73641 114550 73697
rect 114618 73641 114674 73697
rect 114742 73641 114798 73697
rect 112882 73517 112938 73573
rect 113006 73517 113062 73573
rect 113130 73517 113186 73573
rect 113254 73517 113310 73573
rect 113378 73517 113434 73573
rect 113502 73517 113558 73573
rect 113626 73517 113682 73573
rect 113750 73517 113806 73573
rect 113874 73517 113930 73573
rect 113998 73517 114054 73573
rect 114122 73517 114178 73573
rect 114246 73517 114302 73573
rect 114370 73517 114426 73573
rect 114494 73517 114550 73573
rect 114618 73517 114674 73573
rect 114742 73517 114798 73573
rect 112882 73393 112938 73449
rect 113006 73393 113062 73449
rect 113130 73393 113186 73449
rect 113254 73393 113310 73449
rect 113378 73393 113434 73449
rect 113502 73393 113558 73449
rect 113626 73393 113682 73449
rect 113750 73393 113806 73449
rect 113874 73393 113930 73449
rect 113998 73393 114054 73449
rect 114122 73393 114178 73449
rect 114246 73393 114302 73449
rect 114370 73393 114426 73449
rect 114494 73393 114550 73449
rect 114618 73393 114674 73449
rect 114742 73393 114798 73449
rect 112882 73269 112938 73325
rect 113006 73269 113062 73325
rect 113130 73269 113186 73325
rect 113254 73269 113310 73325
rect 113378 73269 113434 73325
rect 113502 73269 113558 73325
rect 113626 73269 113682 73325
rect 113750 73269 113806 73325
rect 113874 73269 113930 73325
rect 113998 73269 114054 73325
rect 114122 73269 114178 73325
rect 114246 73269 114302 73325
rect 114370 73269 114426 73325
rect 114494 73269 114550 73325
rect 114618 73269 114674 73325
rect 114742 73269 114798 73325
rect 112882 73145 112938 73201
rect 113006 73145 113062 73201
rect 113130 73145 113186 73201
rect 113254 73145 113310 73201
rect 113378 73145 113434 73201
rect 113502 73145 113558 73201
rect 113626 73145 113682 73201
rect 113750 73145 113806 73201
rect 113874 73145 113930 73201
rect 113998 73145 114054 73201
rect 114122 73145 114178 73201
rect 114246 73145 114302 73201
rect 114370 73145 114426 73201
rect 114494 73145 114550 73201
rect 114618 73145 114674 73201
rect 114742 73145 114798 73201
rect 112882 73021 112938 73077
rect 113006 73021 113062 73077
rect 113130 73021 113186 73077
rect 113254 73021 113310 73077
rect 113378 73021 113434 73077
rect 113502 73021 113558 73077
rect 113626 73021 113682 73077
rect 113750 73021 113806 73077
rect 113874 73021 113930 73077
rect 113998 73021 114054 73077
rect 114122 73021 114178 73077
rect 114246 73021 114302 73077
rect 114370 73021 114426 73077
rect 114494 73021 114550 73077
rect 114618 73021 114674 73077
rect 114742 73021 114798 73077
rect 112882 72897 112938 72953
rect 113006 72897 113062 72953
rect 113130 72897 113186 72953
rect 113254 72897 113310 72953
rect 113378 72897 113434 72953
rect 113502 72897 113558 72953
rect 113626 72897 113682 72953
rect 113750 72897 113806 72953
rect 113874 72897 113930 72953
rect 113998 72897 114054 72953
rect 114122 72897 114178 72953
rect 114246 72897 114302 72953
rect 114370 72897 114426 72953
rect 114494 72897 114550 72953
rect 114618 72897 114674 72953
rect 114742 72897 114798 72953
rect 112882 72773 112938 72829
rect 113006 72773 113062 72829
rect 113130 72773 113186 72829
rect 113254 72773 113310 72829
rect 113378 72773 113434 72829
rect 113502 72773 113558 72829
rect 113626 72773 113682 72829
rect 113750 72773 113806 72829
rect 113874 72773 113930 72829
rect 113998 72773 114054 72829
rect 114122 72773 114178 72829
rect 114246 72773 114302 72829
rect 114370 72773 114426 72829
rect 114494 72773 114550 72829
rect 114618 72773 114674 72829
rect 114742 72773 114798 72829
rect 112882 72649 112938 72705
rect 113006 72649 113062 72705
rect 113130 72649 113186 72705
rect 113254 72649 113310 72705
rect 113378 72649 113434 72705
rect 113502 72649 113558 72705
rect 113626 72649 113682 72705
rect 113750 72649 113806 72705
rect 113874 72649 113930 72705
rect 113998 72649 114054 72705
rect 114122 72649 114178 72705
rect 114246 72649 114302 72705
rect 114370 72649 114426 72705
rect 114494 72649 114550 72705
rect 114618 72649 114674 72705
rect 114742 72649 114798 72705
rect 112882 72525 112938 72581
rect 113006 72525 113062 72581
rect 113130 72525 113186 72581
rect 113254 72525 113310 72581
rect 113378 72525 113434 72581
rect 113502 72525 113558 72581
rect 113626 72525 113682 72581
rect 113750 72525 113806 72581
rect 113874 72525 113930 72581
rect 113998 72525 114054 72581
rect 114122 72525 114178 72581
rect 114246 72525 114302 72581
rect 114370 72525 114426 72581
rect 114494 72525 114550 72581
rect 114618 72525 114674 72581
rect 114742 72525 114798 72581
rect 112882 72401 112938 72457
rect 113006 72401 113062 72457
rect 113130 72401 113186 72457
rect 113254 72401 113310 72457
rect 113378 72401 113434 72457
rect 113502 72401 113558 72457
rect 113626 72401 113682 72457
rect 113750 72401 113806 72457
rect 113874 72401 113930 72457
rect 113998 72401 114054 72457
rect 114122 72401 114178 72457
rect 114246 72401 114302 72457
rect 114370 72401 114426 72457
rect 114494 72401 114550 72457
rect 114618 72401 114674 72457
rect 114742 72401 114798 72457
rect 112882 72277 112938 72333
rect 113006 72277 113062 72333
rect 113130 72277 113186 72333
rect 113254 72277 113310 72333
rect 113378 72277 113434 72333
rect 113502 72277 113558 72333
rect 113626 72277 113682 72333
rect 113750 72277 113806 72333
rect 113874 72277 113930 72333
rect 113998 72277 114054 72333
rect 114122 72277 114178 72333
rect 114246 72277 114302 72333
rect 114370 72277 114426 72333
rect 114494 72277 114550 72333
rect 114618 72277 114674 72333
rect 114742 72277 114798 72333
rect 112882 72153 112938 72209
rect 113006 72153 113062 72209
rect 113130 72153 113186 72209
rect 113254 72153 113310 72209
rect 113378 72153 113434 72209
rect 113502 72153 113558 72209
rect 113626 72153 113682 72209
rect 113750 72153 113806 72209
rect 113874 72153 113930 72209
rect 113998 72153 114054 72209
rect 114122 72153 114178 72209
rect 114246 72153 114302 72209
rect 114370 72153 114426 72209
rect 114494 72153 114550 72209
rect 114618 72153 114674 72209
rect 114742 72153 114798 72209
rect 115252 73889 115308 73945
rect 115376 73889 115432 73945
rect 115500 73889 115556 73945
rect 115624 73889 115680 73945
rect 115748 73889 115804 73945
rect 115872 73889 115928 73945
rect 115996 73889 116052 73945
rect 116120 73889 116176 73945
rect 116244 73889 116300 73945
rect 116368 73889 116424 73945
rect 116492 73889 116548 73945
rect 116616 73889 116672 73945
rect 116740 73889 116796 73945
rect 116864 73889 116920 73945
rect 116988 73889 117044 73945
rect 117112 73889 117168 73945
rect 115252 73765 115308 73821
rect 115376 73765 115432 73821
rect 115500 73765 115556 73821
rect 115624 73765 115680 73821
rect 115748 73765 115804 73821
rect 115872 73765 115928 73821
rect 115996 73765 116052 73821
rect 116120 73765 116176 73821
rect 116244 73765 116300 73821
rect 116368 73765 116424 73821
rect 116492 73765 116548 73821
rect 116616 73765 116672 73821
rect 116740 73765 116796 73821
rect 116864 73765 116920 73821
rect 116988 73765 117044 73821
rect 117112 73765 117168 73821
rect 115252 73641 115308 73697
rect 115376 73641 115432 73697
rect 115500 73641 115556 73697
rect 115624 73641 115680 73697
rect 115748 73641 115804 73697
rect 115872 73641 115928 73697
rect 115996 73641 116052 73697
rect 116120 73641 116176 73697
rect 116244 73641 116300 73697
rect 116368 73641 116424 73697
rect 116492 73641 116548 73697
rect 116616 73641 116672 73697
rect 116740 73641 116796 73697
rect 116864 73641 116920 73697
rect 116988 73641 117044 73697
rect 117112 73641 117168 73697
rect 115252 73517 115308 73573
rect 115376 73517 115432 73573
rect 115500 73517 115556 73573
rect 115624 73517 115680 73573
rect 115748 73517 115804 73573
rect 115872 73517 115928 73573
rect 115996 73517 116052 73573
rect 116120 73517 116176 73573
rect 116244 73517 116300 73573
rect 116368 73517 116424 73573
rect 116492 73517 116548 73573
rect 116616 73517 116672 73573
rect 116740 73517 116796 73573
rect 116864 73517 116920 73573
rect 116988 73517 117044 73573
rect 117112 73517 117168 73573
rect 115252 73393 115308 73449
rect 115376 73393 115432 73449
rect 115500 73393 115556 73449
rect 115624 73393 115680 73449
rect 115748 73393 115804 73449
rect 115872 73393 115928 73449
rect 115996 73393 116052 73449
rect 116120 73393 116176 73449
rect 116244 73393 116300 73449
rect 116368 73393 116424 73449
rect 116492 73393 116548 73449
rect 116616 73393 116672 73449
rect 116740 73393 116796 73449
rect 116864 73393 116920 73449
rect 116988 73393 117044 73449
rect 117112 73393 117168 73449
rect 115252 73269 115308 73325
rect 115376 73269 115432 73325
rect 115500 73269 115556 73325
rect 115624 73269 115680 73325
rect 115748 73269 115804 73325
rect 115872 73269 115928 73325
rect 115996 73269 116052 73325
rect 116120 73269 116176 73325
rect 116244 73269 116300 73325
rect 116368 73269 116424 73325
rect 116492 73269 116548 73325
rect 116616 73269 116672 73325
rect 116740 73269 116796 73325
rect 116864 73269 116920 73325
rect 116988 73269 117044 73325
rect 117112 73269 117168 73325
rect 115252 73145 115308 73201
rect 115376 73145 115432 73201
rect 115500 73145 115556 73201
rect 115624 73145 115680 73201
rect 115748 73145 115804 73201
rect 115872 73145 115928 73201
rect 115996 73145 116052 73201
rect 116120 73145 116176 73201
rect 116244 73145 116300 73201
rect 116368 73145 116424 73201
rect 116492 73145 116548 73201
rect 116616 73145 116672 73201
rect 116740 73145 116796 73201
rect 116864 73145 116920 73201
rect 116988 73145 117044 73201
rect 117112 73145 117168 73201
rect 115252 73021 115308 73077
rect 115376 73021 115432 73077
rect 115500 73021 115556 73077
rect 115624 73021 115680 73077
rect 115748 73021 115804 73077
rect 115872 73021 115928 73077
rect 115996 73021 116052 73077
rect 116120 73021 116176 73077
rect 116244 73021 116300 73077
rect 116368 73021 116424 73077
rect 116492 73021 116548 73077
rect 116616 73021 116672 73077
rect 116740 73021 116796 73077
rect 116864 73021 116920 73077
rect 116988 73021 117044 73077
rect 117112 73021 117168 73077
rect 115252 72897 115308 72953
rect 115376 72897 115432 72953
rect 115500 72897 115556 72953
rect 115624 72897 115680 72953
rect 115748 72897 115804 72953
rect 115872 72897 115928 72953
rect 115996 72897 116052 72953
rect 116120 72897 116176 72953
rect 116244 72897 116300 72953
rect 116368 72897 116424 72953
rect 116492 72897 116548 72953
rect 116616 72897 116672 72953
rect 116740 72897 116796 72953
rect 116864 72897 116920 72953
rect 116988 72897 117044 72953
rect 117112 72897 117168 72953
rect 115252 72773 115308 72829
rect 115376 72773 115432 72829
rect 115500 72773 115556 72829
rect 115624 72773 115680 72829
rect 115748 72773 115804 72829
rect 115872 72773 115928 72829
rect 115996 72773 116052 72829
rect 116120 72773 116176 72829
rect 116244 72773 116300 72829
rect 116368 72773 116424 72829
rect 116492 72773 116548 72829
rect 116616 72773 116672 72829
rect 116740 72773 116796 72829
rect 116864 72773 116920 72829
rect 116988 72773 117044 72829
rect 117112 72773 117168 72829
rect 115252 72649 115308 72705
rect 115376 72649 115432 72705
rect 115500 72649 115556 72705
rect 115624 72649 115680 72705
rect 115748 72649 115804 72705
rect 115872 72649 115928 72705
rect 115996 72649 116052 72705
rect 116120 72649 116176 72705
rect 116244 72649 116300 72705
rect 116368 72649 116424 72705
rect 116492 72649 116548 72705
rect 116616 72649 116672 72705
rect 116740 72649 116796 72705
rect 116864 72649 116920 72705
rect 116988 72649 117044 72705
rect 117112 72649 117168 72705
rect 115252 72525 115308 72581
rect 115376 72525 115432 72581
rect 115500 72525 115556 72581
rect 115624 72525 115680 72581
rect 115748 72525 115804 72581
rect 115872 72525 115928 72581
rect 115996 72525 116052 72581
rect 116120 72525 116176 72581
rect 116244 72525 116300 72581
rect 116368 72525 116424 72581
rect 116492 72525 116548 72581
rect 116616 72525 116672 72581
rect 116740 72525 116796 72581
rect 116864 72525 116920 72581
rect 116988 72525 117044 72581
rect 117112 72525 117168 72581
rect 115252 72401 115308 72457
rect 115376 72401 115432 72457
rect 115500 72401 115556 72457
rect 115624 72401 115680 72457
rect 115748 72401 115804 72457
rect 115872 72401 115928 72457
rect 115996 72401 116052 72457
rect 116120 72401 116176 72457
rect 116244 72401 116300 72457
rect 116368 72401 116424 72457
rect 116492 72401 116548 72457
rect 116616 72401 116672 72457
rect 116740 72401 116796 72457
rect 116864 72401 116920 72457
rect 116988 72401 117044 72457
rect 117112 72401 117168 72457
rect 115252 72277 115308 72333
rect 115376 72277 115432 72333
rect 115500 72277 115556 72333
rect 115624 72277 115680 72333
rect 115748 72277 115804 72333
rect 115872 72277 115928 72333
rect 115996 72277 116052 72333
rect 116120 72277 116176 72333
rect 116244 72277 116300 72333
rect 116368 72277 116424 72333
rect 116492 72277 116548 72333
rect 116616 72277 116672 72333
rect 116740 72277 116796 72333
rect 116864 72277 116920 72333
rect 116988 72277 117044 72333
rect 117112 72277 117168 72333
rect 115252 72153 115308 72209
rect 115376 72153 115432 72209
rect 115500 72153 115556 72209
rect 115624 72153 115680 72209
rect 115748 72153 115804 72209
rect 115872 72153 115928 72209
rect 115996 72153 116052 72209
rect 116120 72153 116176 72209
rect 116244 72153 116300 72209
rect 116368 72153 116424 72209
rect 116492 72153 116548 72209
rect 116616 72153 116672 72209
rect 116740 72153 116796 72209
rect 116864 72153 116920 72209
rect 116988 72153 117044 72209
rect 117112 72153 117168 72209
rect 117882 73889 117938 73945
rect 118006 73889 118062 73945
rect 118130 73889 118186 73945
rect 118254 73889 118310 73945
rect 118378 73889 118434 73945
rect 118502 73889 118558 73945
rect 118626 73889 118682 73945
rect 118750 73889 118806 73945
rect 118874 73889 118930 73945
rect 118998 73889 119054 73945
rect 119122 73889 119178 73945
rect 119246 73889 119302 73945
rect 119370 73889 119426 73945
rect 119494 73889 119550 73945
rect 119618 73889 119674 73945
rect 117882 73765 117938 73821
rect 118006 73765 118062 73821
rect 118130 73765 118186 73821
rect 118254 73765 118310 73821
rect 118378 73765 118434 73821
rect 118502 73765 118558 73821
rect 118626 73765 118682 73821
rect 118750 73765 118806 73821
rect 118874 73765 118930 73821
rect 118998 73765 119054 73821
rect 119122 73765 119178 73821
rect 119246 73765 119302 73821
rect 119370 73765 119426 73821
rect 119494 73765 119550 73821
rect 119618 73765 119674 73821
rect 117882 73641 117938 73697
rect 118006 73641 118062 73697
rect 118130 73641 118186 73697
rect 118254 73641 118310 73697
rect 118378 73641 118434 73697
rect 118502 73641 118558 73697
rect 118626 73641 118682 73697
rect 118750 73641 118806 73697
rect 118874 73641 118930 73697
rect 118998 73641 119054 73697
rect 119122 73641 119178 73697
rect 119246 73641 119302 73697
rect 119370 73641 119426 73697
rect 119494 73641 119550 73697
rect 119618 73641 119674 73697
rect 117882 73517 117938 73573
rect 118006 73517 118062 73573
rect 118130 73517 118186 73573
rect 118254 73517 118310 73573
rect 118378 73517 118434 73573
rect 118502 73517 118558 73573
rect 118626 73517 118682 73573
rect 118750 73517 118806 73573
rect 118874 73517 118930 73573
rect 118998 73517 119054 73573
rect 119122 73517 119178 73573
rect 119246 73517 119302 73573
rect 119370 73517 119426 73573
rect 119494 73517 119550 73573
rect 119618 73517 119674 73573
rect 117882 73393 117938 73449
rect 118006 73393 118062 73449
rect 118130 73393 118186 73449
rect 118254 73393 118310 73449
rect 118378 73393 118434 73449
rect 118502 73393 118558 73449
rect 118626 73393 118682 73449
rect 118750 73393 118806 73449
rect 118874 73393 118930 73449
rect 118998 73393 119054 73449
rect 119122 73393 119178 73449
rect 119246 73393 119302 73449
rect 119370 73393 119426 73449
rect 119494 73393 119550 73449
rect 119618 73393 119674 73449
rect 117882 73269 117938 73325
rect 118006 73269 118062 73325
rect 118130 73269 118186 73325
rect 118254 73269 118310 73325
rect 118378 73269 118434 73325
rect 118502 73269 118558 73325
rect 118626 73269 118682 73325
rect 118750 73269 118806 73325
rect 118874 73269 118930 73325
rect 118998 73269 119054 73325
rect 119122 73269 119178 73325
rect 119246 73269 119302 73325
rect 119370 73269 119426 73325
rect 119494 73269 119550 73325
rect 119618 73269 119674 73325
rect 117882 73145 117938 73201
rect 118006 73145 118062 73201
rect 118130 73145 118186 73201
rect 118254 73145 118310 73201
rect 118378 73145 118434 73201
rect 118502 73145 118558 73201
rect 118626 73145 118682 73201
rect 118750 73145 118806 73201
rect 118874 73145 118930 73201
rect 118998 73145 119054 73201
rect 119122 73145 119178 73201
rect 119246 73145 119302 73201
rect 119370 73145 119426 73201
rect 119494 73145 119550 73201
rect 119618 73145 119674 73201
rect 117882 73021 117938 73077
rect 118006 73021 118062 73077
rect 118130 73021 118186 73077
rect 118254 73021 118310 73077
rect 118378 73021 118434 73077
rect 118502 73021 118558 73077
rect 118626 73021 118682 73077
rect 118750 73021 118806 73077
rect 118874 73021 118930 73077
rect 118998 73021 119054 73077
rect 119122 73021 119178 73077
rect 119246 73021 119302 73077
rect 119370 73021 119426 73077
rect 119494 73021 119550 73077
rect 119618 73021 119674 73077
rect 117882 72897 117938 72953
rect 118006 72897 118062 72953
rect 118130 72897 118186 72953
rect 118254 72897 118310 72953
rect 118378 72897 118434 72953
rect 118502 72897 118558 72953
rect 118626 72897 118682 72953
rect 118750 72897 118806 72953
rect 118874 72897 118930 72953
rect 118998 72897 119054 72953
rect 119122 72897 119178 72953
rect 119246 72897 119302 72953
rect 119370 72897 119426 72953
rect 119494 72897 119550 72953
rect 119618 72897 119674 72953
rect 117882 72773 117938 72829
rect 118006 72773 118062 72829
rect 118130 72773 118186 72829
rect 118254 72773 118310 72829
rect 118378 72773 118434 72829
rect 118502 72773 118558 72829
rect 118626 72773 118682 72829
rect 118750 72773 118806 72829
rect 118874 72773 118930 72829
rect 118998 72773 119054 72829
rect 119122 72773 119178 72829
rect 119246 72773 119302 72829
rect 119370 72773 119426 72829
rect 119494 72773 119550 72829
rect 119618 72773 119674 72829
rect 117882 72649 117938 72705
rect 118006 72649 118062 72705
rect 118130 72649 118186 72705
rect 118254 72649 118310 72705
rect 118378 72649 118434 72705
rect 118502 72649 118558 72705
rect 118626 72649 118682 72705
rect 118750 72649 118806 72705
rect 118874 72649 118930 72705
rect 118998 72649 119054 72705
rect 119122 72649 119178 72705
rect 119246 72649 119302 72705
rect 119370 72649 119426 72705
rect 119494 72649 119550 72705
rect 119618 72649 119674 72705
rect 117882 72525 117938 72581
rect 118006 72525 118062 72581
rect 118130 72525 118186 72581
rect 118254 72525 118310 72581
rect 118378 72525 118434 72581
rect 118502 72525 118558 72581
rect 118626 72525 118682 72581
rect 118750 72525 118806 72581
rect 118874 72525 118930 72581
rect 118998 72525 119054 72581
rect 119122 72525 119178 72581
rect 119246 72525 119302 72581
rect 119370 72525 119426 72581
rect 119494 72525 119550 72581
rect 119618 72525 119674 72581
rect 117882 72401 117938 72457
rect 118006 72401 118062 72457
rect 118130 72401 118186 72457
rect 118254 72401 118310 72457
rect 118378 72401 118434 72457
rect 118502 72401 118558 72457
rect 118626 72401 118682 72457
rect 118750 72401 118806 72457
rect 118874 72401 118930 72457
rect 118998 72401 119054 72457
rect 119122 72401 119178 72457
rect 119246 72401 119302 72457
rect 119370 72401 119426 72457
rect 119494 72401 119550 72457
rect 119618 72401 119674 72457
rect 117882 72277 117938 72333
rect 118006 72277 118062 72333
rect 118130 72277 118186 72333
rect 118254 72277 118310 72333
rect 118378 72277 118434 72333
rect 118502 72277 118558 72333
rect 118626 72277 118682 72333
rect 118750 72277 118806 72333
rect 118874 72277 118930 72333
rect 118998 72277 119054 72333
rect 119122 72277 119178 72333
rect 119246 72277 119302 72333
rect 119370 72277 119426 72333
rect 119494 72277 119550 72333
rect 119618 72277 119674 72333
rect 117882 72153 117938 72209
rect 118006 72153 118062 72209
rect 118130 72153 118186 72209
rect 118254 72153 118310 72209
rect 118378 72153 118434 72209
rect 118502 72153 118558 72209
rect 118626 72153 118682 72209
rect 118750 72153 118806 72209
rect 118874 72153 118930 72209
rect 118998 72153 119054 72209
rect 119122 72153 119178 72209
rect 119246 72153 119302 72209
rect 119370 72153 119426 72209
rect 119494 72153 119550 72209
rect 119618 72153 119674 72209
rect 270326 73889 270382 73945
rect 270450 73889 270506 73945
rect 270574 73889 270630 73945
rect 270698 73889 270754 73945
rect 270822 73889 270878 73945
rect 270946 73889 271002 73945
rect 271070 73889 271126 73945
rect 271194 73889 271250 73945
rect 271318 73889 271374 73945
rect 271442 73889 271498 73945
rect 271566 73889 271622 73945
rect 271690 73889 271746 73945
rect 271814 73889 271870 73945
rect 271938 73889 271994 73945
rect 272062 73889 272118 73945
rect 270326 73765 270382 73821
rect 270450 73765 270506 73821
rect 270574 73765 270630 73821
rect 270698 73765 270754 73821
rect 270822 73765 270878 73821
rect 270946 73765 271002 73821
rect 271070 73765 271126 73821
rect 271194 73765 271250 73821
rect 271318 73765 271374 73821
rect 271442 73765 271498 73821
rect 271566 73765 271622 73821
rect 271690 73765 271746 73821
rect 271814 73765 271870 73821
rect 271938 73765 271994 73821
rect 272062 73765 272118 73821
rect 270326 73641 270382 73697
rect 270450 73641 270506 73697
rect 270574 73641 270630 73697
rect 270698 73641 270754 73697
rect 270822 73641 270878 73697
rect 270946 73641 271002 73697
rect 271070 73641 271126 73697
rect 271194 73641 271250 73697
rect 271318 73641 271374 73697
rect 271442 73641 271498 73697
rect 271566 73641 271622 73697
rect 271690 73641 271746 73697
rect 271814 73641 271870 73697
rect 271938 73641 271994 73697
rect 272062 73641 272118 73697
rect 270326 73517 270382 73573
rect 270450 73517 270506 73573
rect 270574 73517 270630 73573
rect 270698 73517 270754 73573
rect 270822 73517 270878 73573
rect 270946 73517 271002 73573
rect 271070 73517 271126 73573
rect 271194 73517 271250 73573
rect 271318 73517 271374 73573
rect 271442 73517 271498 73573
rect 271566 73517 271622 73573
rect 271690 73517 271746 73573
rect 271814 73517 271870 73573
rect 271938 73517 271994 73573
rect 272062 73517 272118 73573
rect 270326 73393 270382 73449
rect 270450 73393 270506 73449
rect 270574 73393 270630 73449
rect 270698 73393 270754 73449
rect 270822 73393 270878 73449
rect 270946 73393 271002 73449
rect 271070 73393 271126 73449
rect 271194 73393 271250 73449
rect 271318 73393 271374 73449
rect 271442 73393 271498 73449
rect 271566 73393 271622 73449
rect 271690 73393 271746 73449
rect 271814 73393 271870 73449
rect 271938 73393 271994 73449
rect 272062 73393 272118 73449
rect 270326 73269 270382 73325
rect 270450 73269 270506 73325
rect 270574 73269 270630 73325
rect 270698 73269 270754 73325
rect 270822 73269 270878 73325
rect 270946 73269 271002 73325
rect 271070 73269 271126 73325
rect 271194 73269 271250 73325
rect 271318 73269 271374 73325
rect 271442 73269 271498 73325
rect 271566 73269 271622 73325
rect 271690 73269 271746 73325
rect 271814 73269 271870 73325
rect 271938 73269 271994 73325
rect 272062 73269 272118 73325
rect 270326 73145 270382 73201
rect 270450 73145 270506 73201
rect 270574 73145 270630 73201
rect 270698 73145 270754 73201
rect 270822 73145 270878 73201
rect 270946 73145 271002 73201
rect 271070 73145 271126 73201
rect 271194 73145 271250 73201
rect 271318 73145 271374 73201
rect 271442 73145 271498 73201
rect 271566 73145 271622 73201
rect 271690 73145 271746 73201
rect 271814 73145 271870 73201
rect 271938 73145 271994 73201
rect 272062 73145 272118 73201
rect 270326 73021 270382 73077
rect 270450 73021 270506 73077
rect 270574 73021 270630 73077
rect 270698 73021 270754 73077
rect 270822 73021 270878 73077
rect 270946 73021 271002 73077
rect 271070 73021 271126 73077
rect 271194 73021 271250 73077
rect 271318 73021 271374 73077
rect 271442 73021 271498 73077
rect 271566 73021 271622 73077
rect 271690 73021 271746 73077
rect 271814 73021 271870 73077
rect 271938 73021 271994 73077
rect 272062 73021 272118 73077
rect 270326 72897 270382 72953
rect 270450 72897 270506 72953
rect 270574 72897 270630 72953
rect 270698 72897 270754 72953
rect 270822 72897 270878 72953
rect 270946 72897 271002 72953
rect 271070 72897 271126 72953
rect 271194 72897 271250 72953
rect 271318 72897 271374 72953
rect 271442 72897 271498 72953
rect 271566 72897 271622 72953
rect 271690 72897 271746 72953
rect 271814 72897 271870 72953
rect 271938 72897 271994 72953
rect 272062 72897 272118 72953
rect 270326 72773 270382 72829
rect 270450 72773 270506 72829
rect 270574 72773 270630 72829
rect 270698 72773 270754 72829
rect 270822 72773 270878 72829
rect 270946 72773 271002 72829
rect 271070 72773 271126 72829
rect 271194 72773 271250 72829
rect 271318 72773 271374 72829
rect 271442 72773 271498 72829
rect 271566 72773 271622 72829
rect 271690 72773 271746 72829
rect 271814 72773 271870 72829
rect 271938 72773 271994 72829
rect 272062 72773 272118 72829
rect 270326 72649 270382 72705
rect 270450 72649 270506 72705
rect 270574 72649 270630 72705
rect 270698 72649 270754 72705
rect 270822 72649 270878 72705
rect 270946 72649 271002 72705
rect 271070 72649 271126 72705
rect 271194 72649 271250 72705
rect 271318 72649 271374 72705
rect 271442 72649 271498 72705
rect 271566 72649 271622 72705
rect 271690 72649 271746 72705
rect 271814 72649 271870 72705
rect 271938 72649 271994 72705
rect 272062 72649 272118 72705
rect 270326 72525 270382 72581
rect 270450 72525 270506 72581
rect 270574 72525 270630 72581
rect 270698 72525 270754 72581
rect 270822 72525 270878 72581
rect 270946 72525 271002 72581
rect 271070 72525 271126 72581
rect 271194 72525 271250 72581
rect 271318 72525 271374 72581
rect 271442 72525 271498 72581
rect 271566 72525 271622 72581
rect 271690 72525 271746 72581
rect 271814 72525 271870 72581
rect 271938 72525 271994 72581
rect 272062 72525 272118 72581
rect 270326 72401 270382 72457
rect 270450 72401 270506 72457
rect 270574 72401 270630 72457
rect 270698 72401 270754 72457
rect 270822 72401 270878 72457
rect 270946 72401 271002 72457
rect 271070 72401 271126 72457
rect 271194 72401 271250 72457
rect 271318 72401 271374 72457
rect 271442 72401 271498 72457
rect 271566 72401 271622 72457
rect 271690 72401 271746 72457
rect 271814 72401 271870 72457
rect 271938 72401 271994 72457
rect 272062 72401 272118 72457
rect 270326 72277 270382 72333
rect 270450 72277 270506 72333
rect 270574 72277 270630 72333
rect 270698 72277 270754 72333
rect 270822 72277 270878 72333
rect 270946 72277 271002 72333
rect 271070 72277 271126 72333
rect 271194 72277 271250 72333
rect 271318 72277 271374 72333
rect 271442 72277 271498 72333
rect 271566 72277 271622 72333
rect 271690 72277 271746 72333
rect 271814 72277 271870 72333
rect 271938 72277 271994 72333
rect 272062 72277 272118 72333
rect 270326 72153 270382 72209
rect 270450 72153 270506 72209
rect 270574 72153 270630 72209
rect 270698 72153 270754 72209
rect 270822 72153 270878 72209
rect 270946 72153 271002 72209
rect 271070 72153 271126 72209
rect 271194 72153 271250 72209
rect 271318 72153 271374 72209
rect 271442 72153 271498 72209
rect 271566 72153 271622 72209
rect 271690 72153 271746 72209
rect 271814 72153 271870 72209
rect 271938 72153 271994 72209
rect 272062 72153 272118 72209
rect 272806 73889 272862 73945
rect 272930 73889 272986 73945
rect 273054 73889 273110 73945
rect 273178 73889 273234 73945
rect 273302 73889 273358 73945
rect 273426 73889 273482 73945
rect 273550 73889 273606 73945
rect 273674 73889 273730 73945
rect 273798 73889 273854 73945
rect 273922 73889 273978 73945
rect 274046 73889 274102 73945
rect 274170 73889 274226 73945
rect 274294 73889 274350 73945
rect 274418 73889 274474 73945
rect 274542 73889 274598 73945
rect 274666 73889 274722 73945
rect 272806 73765 272862 73821
rect 272930 73765 272986 73821
rect 273054 73765 273110 73821
rect 273178 73765 273234 73821
rect 273302 73765 273358 73821
rect 273426 73765 273482 73821
rect 273550 73765 273606 73821
rect 273674 73765 273730 73821
rect 273798 73765 273854 73821
rect 273922 73765 273978 73821
rect 274046 73765 274102 73821
rect 274170 73765 274226 73821
rect 274294 73765 274350 73821
rect 274418 73765 274474 73821
rect 274542 73765 274598 73821
rect 274666 73765 274722 73821
rect 272806 73641 272862 73697
rect 272930 73641 272986 73697
rect 273054 73641 273110 73697
rect 273178 73641 273234 73697
rect 273302 73641 273358 73697
rect 273426 73641 273482 73697
rect 273550 73641 273606 73697
rect 273674 73641 273730 73697
rect 273798 73641 273854 73697
rect 273922 73641 273978 73697
rect 274046 73641 274102 73697
rect 274170 73641 274226 73697
rect 274294 73641 274350 73697
rect 274418 73641 274474 73697
rect 274542 73641 274598 73697
rect 274666 73641 274722 73697
rect 272806 73517 272862 73573
rect 272930 73517 272986 73573
rect 273054 73517 273110 73573
rect 273178 73517 273234 73573
rect 273302 73517 273358 73573
rect 273426 73517 273482 73573
rect 273550 73517 273606 73573
rect 273674 73517 273730 73573
rect 273798 73517 273854 73573
rect 273922 73517 273978 73573
rect 274046 73517 274102 73573
rect 274170 73517 274226 73573
rect 274294 73517 274350 73573
rect 274418 73517 274474 73573
rect 274542 73517 274598 73573
rect 274666 73517 274722 73573
rect 272806 73393 272862 73449
rect 272930 73393 272986 73449
rect 273054 73393 273110 73449
rect 273178 73393 273234 73449
rect 273302 73393 273358 73449
rect 273426 73393 273482 73449
rect 273550 73393 273606 73449
rect 273674 73393 273730 73449
rect 273798 73393 273854 73449
rect 273922 73393 273978 73449
rect 274046 73393 274102 73449
rect 274170 73393 274226 73449
rect 274294 73393 274350 73449
rect 274418 73393 274474 73449
rect 274542 73393 274598 73449
rect 274666 73393 274722 73449
rect 272806 73269 272862 73325
rect 272930 73269 272986 73325
rect 273054 73269 273110 73325
rect 273178 73269 273234 73325
rect 273302 73269 273358 73325
rect 273426 73269 273482 73325
rect 273550 73269 273606 73325
rect 273674 73269 273730 73325
rect 273798 73269 273854 73325
rect 273922 73269 273978 73325
rect 274046 73269 274102 73325
rect 274170 73269 274226 73325
rect 274294 73269 274350 73325
rect 274418 73269 274474 73325
rect 274542 73269 274598 73325
rect 274666 73269 274722 73325
rect 272806 73145 272862 73201
rect 272930 73145 272986 73201
rect 273054 73145 273110 73201
rect 273178 73145 273234 73201
rect 273302 73145 273358 73201
rect 273426 73145 273482 73201
rect 273550 73145 273606 73201
rect 273674 73145 273730 73201
rect 273798 73145 273854 73201
rect 273922 73145 273978 73201
rect 274046 73145 274102 73201
rect 274170 73145 274226 73201
rect 274294 73145 274350 73201
rect 274418 73145 274474 73201
rect 274542 73145 274598 73201
rect 274666 73145 274722 73201
rect 272806 73021 272862 73077
rect 272930 73021 272986 73077
rect 273054 73021 273110 73077
rect 273178 73021 273234 73077
rect 273302 73021 273358 73077
rect 273426 73021 273482 73077
rect 273550 73021 273606 73077
rect 273674 73021 273730 73077
rect 273798 73021 273854 73077
rect 273922 73021 273978 73077
rect 274046 73021 274102 73077
rect 274170 73021 274226 73077
rect 274294 73021 274350 73077
rect 274418 73021 274474 73077
rect 274542 73021 274598 73077
rect 274666 73021 274722 73077
rect 272806 72897 272862 72953
rect 272930 72897 272986 72953
rect 273054 72897 273110 72953
rect 273178 72897 273234 72953
rect 273302 72897 273358 72953
rect 273426 72897 273482 72953
rect 273550 72897 273606 72953
rect 273674 72897 273730 72953
rect 273798 72897 273854 72953
rect 273922 72897 273978 72953
rect 274046 72897 274102 72953
rect 274170 72897 274226 72953
rect 274294 72897 274350 72953
rect 274418 72897 274474 72953
rect 274542 72897 274598 72953
rect 274666 72897 274722 72953
rect 272806 72773 272862 72829
rect 272930 72773 272986 72829
rect 273054 72773 273110 72829
rect 273178 72773 273234 72829
rect 273302 72773 273358 72829
rect 273426 72773 273482 72829
rect 273550 72773 273606 72829
rect 273674 72773 273730 72829
rect 273798 72773 273854 72829
rect 273922 72773 273978 72829
rect 274046 72773 274102 72829
rect 274170 72773 274226 72829
rect 274294 72773 274350 72829
rect 274418 72773 274474 72829
rect 274542 72773 274598 72829
rect 274666 72773 274722 72829
rect 272806 72649 272862 72705
rect 272930 72649 272986 72705
rect 273054 72649 273110 72705
rect 273178 72649 273234 72705
rect 273302 72649 273358 72705
rect 273426 72649 273482 72705
rect 273550 72649 273606 72705
rect 273674 72649 273730 72705
rect 273798 72649 273854 72705
rect 273922 72649 273978 72705
rect 274046 72649 274102 72705
rect 274170 72649 274226 72705
rect 274294 72649 274350 72705
rect 274418 72649 274474 72705
rect 274542 72649 274598 72705
rect 274666 72649 274722 72705
rect 272806 72525 272862 72581
rect 272930 72525 272986 72581
rect 273054 72525 273110 72581
rect 273178 72525 273234 72581
rect 273302 72525 273358 72581
rect 273426 72525 273482 72581
rect 273550 72525 273606 72581
rect 273674 72525 273730 72581
rect 273798 72525 273854 72581
rect 273922 72525 273978 72581
rect 274046 72525 274102 72581
rect 274170 72525 274226 72581
rect 274294 72525 274350 72581
rect 274418 72525 274474 72581
rect 274542 72525 274598 72581
rect 274666 72525 274722 72581
rect 272806 72401 272862 72457
rect 272930 72401 272986 72457
rect 273054 72401 273110 72457
rect 273178 72401 273234 72457
rect 273302 72401 273358 72457
rect 273426 72401 273482 72457
rect 273550 72401 273606 72457
rect 273674 72401 273730 72457
rect 273798 72401 273854 72457
rect 273922 72401 273978 72457
rect 274046 72401 274102 72457
rect 274170 72401 274226 72457
rect 274294 72401 274350 72457
rect 274418 72401 274474 72457
rect 274542 72401 274598 72457
rect 274666 72401 274722 72457
rect 272806 72277 272862 72333
rect 272930 72277 272986 72333
rect 273054 72277 273110 72333
rect 273178 72277 273234 72333
rect 273302 72277 273358 72333
rect 273426 72277 273482 72333
rect 273550 72277 273606 72333
rect 273674 72277 273730 72333
rect 273798 72277 273854 72333
rect 273922 72277 273978 72333
rect 274046 72277 274102 72333
rect 274170 72277 274226 72333
rect 274294 72277 274350 72333
rect 274418 72277 274474 72333
rect 274542 72277 274598 72333
rect 274666 72277 274722 72333
rect 272806 72153 272862 72209
rect 272930 72153 272986 72209
rect 273054 72153 273110 72209
rect 273178 72153 273234 72209
rect 273302 72153 273358 72209
rect 273426 72153 273482 72209
rect 273550 72153 273606 72209
rect 273674 72153 273730 72209
rect 273798 72153 273854 72209
rect 273922 72153 273978 72209
rect 274046 72153 274102 72209
rect 274170 72153 274226 72209
rect 274294 72153 274350 72209
rect 274418 72153 274474 72209
rect 274542 72153 274598 72209
rect 274666 72153 274722 72209
rect 275176 73889 275232 73945
rect 275300 73889 275356 73945
rect 275424 73889 275480 73945
rect 275548 73889 275604 73945
rect 275672 73889 275728 73945
rect 275796 73889 275852 73945
rect 275920 73889 275976 73945
rect 276044 73889 276100 73945
rect 276168 73889 276224 73945
rect 276292 73889 276348 73945
rect 276416 73889 276472 73945
rect 276540 73889 276596 73945
rect 276664 73889 276720 73945
rect 276788 73889 276844 73945
rect 276912 73889 276968 73945
rect 277036 73889 277092 73945
rect 275176 73765 275232 73821
rect 275300 73765 275356 73821
rect 275424 73765 275480 73821
rect 275548 73765 275604 73821
rect 275672 73765 275728 73821
rect 275796 73765 275852 73821
rect 275920 73765 275976 73821
rect 276044 73765 276100 73821
rect 276168 73765 276224 73821
rect 276292 73765 276348 73821
rect 276416 73765 276472 73821
rect 276540 73765 276596 73821
rect 276664 73765 276720 73821
rect 276788 73765 276844 73821
rect 276912 73765 276968 73821
rect 277036 73765 277092 73821
rect 275176 73641 275232 73697
rect 275300 73641 275356 73697
rect 275424 73641 275480 73697
rect 275548 73641 275604 73697
rect 275672 73641 275728 73697
rect 275796 73641 275852 73697
rect 275920 73641 275976 73697
rect 276044 73641 276100 73697
rect 276168 73641 276224 73697
rect 276292 73641 276348 73697
rect 276416 73641 276472 73697
rect 276540 73641 276596 73697
rect 276664 73641 276720 73697
rect 276788 73641 276844 73697
rect 276912 73641 276968 73697
rect 277036 73641 277092 73697
rect 275176 73517 275232 73573
rect 275300 73517 275356 73573
rect 275424 73517 275480 73573
rect 275548 73517 275604 73573
rect 275672 73517 275728 73573
rect 275796 73517 275852 73573
rect 275920 73517 275976 73573
rect 276044 73517 276100 73573
rect 276168 73517 276224 73573
rect 276292 73517 276348 73573
rect 276416 73517 276472 73573
rect 276540 73517 276596 73573
rect 276664 73517 276720 73573
rect 276788 73517 276844 73573
rect 276912 73517 276968 73573
rect 277036 73517 277092 73573
rect 275176 73393 275232 73449
rect 275300 73393 275356 73449
rect 275424 73393 275480 73449
rect 275548 73393 275604 73449
rect 275672 73393 275728 73449
rect 275796 73393 275852 73449
rect 275920 73393 275976 73449
rect 276044 73393 276100 73449
rect 276168 73393 276224 73449
rect 276292 73393 276348 73449
rect 276416 73393 276472 73449
rect 276540 73393 276596 73449
rect 276664 73393 276720 73449
rect 276788 73393 276844 73449
rect 276912 73393 276968 73449
rect 277036 73393 277092 73449
rect 275176 73269 275232 73325
rect 275300 73269 275356 73325
rect 275424 73269 275480 73325
rect 275548 73269 275604 73325
rect 275672 73269 275728 73325
rect 275796 73269 275852 73325
rect 275920 73269 275976 73325
rect 276044 73269 276100 73325
rect 276168 73269 276224 73325
rect 276292 73269 276348 73325
rect 276416 73269 276472 73325
rect 276540 73269 276596 73325
rect 276664 73269 276720 73325
rect 276788 73269 276844 73325
rect 276912 73269 276968 73325
rect 277036 73269 277092 73325
rect 275176 73145 275232 73201
rect 275300 73145 275356 73201
rect 275424 73145 275480 73201
rect 275548 73145 275604 73201
rect 275672 73145 275728 73201
rect 275796 73145 275852 73201
rect 275920 73145 275976 73201
rect 276044 73145 276100 73201
rect 276168 73145 276224 73201
rect 276292 73145 276348 73201
rect 276416 73145 276472 73201
rect 276540 73145 276596 73201
rect 276664 73145 276720 73201
rect 276788 73145 276844 73201
rect 276912 73145 276968 73201
rect 277036 73145 277092 73201
rect 275176 73021 275232 73077
rect 275300 73021 275356 73077
rect 275424 73021 275480 73077
rect 275548 73021 275604 73077
rect 275672 73021 275728 73077
rect 275796 73021 275852 73077
rect 275920 73021 275976 73077
rect 276044 73021 276100 73077
rect 276168 73021 276224 73077
rect 276292 73021 276348 73077
rect 276416 73021 276472 73077
rect 276540 73021 276596 73077
rect 276664 73021 276720 73077
rect 276788 73021 276844 73077
rect 276912 73021 276968 73077
rect 277036 73021 277092 73077
rect 275176 72897 275232 72953
rect 275300 72897 275356 72953
rect 275424 72897 275480 72953
rect 275548 72897 275604 72953
rect 275672 72897 275728 72953
rect 275796 72897 275852 72953
rect 275920 72897 275976 72953
rect 276044 72897 276100 72953
rect 276168 72897 276224 72953
rect 276292 72897 276348 72953
rect 276416 72897 276472 72953
rect 276540 72897 276596 72953
rect 276664 72897 276720 72953
rect 276788 72897 276844 72953
rect 276912 72897 276968 72953
rect 277036 72897 277092 72953
rect 275176 72773 275232 72829
rect 275300 72773 275356 72829
rect 275424 72773 275480 72829
rect 275548 72773 275604 72829
rect 275672 72773 275728 72829
rect 275796 72773 275852 72829
rect 275920 72773 275976 72829
rect 276044 72773 276100 72829
rect 276168 72773 276224 72829
rect 276292 72773 276348 72829
rect 276416 72773 276472 72829
rect 276540 72773 276596 72829
rect 276664 72773 276720 72829
rect 276788 72773 276844 72829
rect 276912 72773 276968 72829
rect 277036 72773 277092 72829
rect 275176 72649 275232 72705
rect 275300 72649 275356 72705
rect 275424 72649 275480 72705
rect 275548 72649 275604 72705
rect 275672 72649 275728 72705
rect 275796 72649 275852 72705
rect 275920 72649 275976 72705
rect 276044 72649 276100 72705
rect 276168 72649 276224 72705
rect 276292 72649 276348 72705
rect 276416 72649 276472 72705
rect 276540 72649 276596 72705
rect 276664 72649 276720 72705
rect 276788 72649 276844 72705
rect 276912 72649 276968 72705
rect 277036 72649 277092 72705
rect 275176 72525 275232 72581
rect 275300 72525 275356 72581
rect 275424 72525 275480 72581
rect 275548 72525 275604 72581
rect 275672 72525 275728 72581
rect 275796 72525 275852 72581
rect 275920 72525 275976 72581
rect 276044 72525 276100 72581
rect 276168 72525 276224 72581
rect 276292 72525 276348 72581
rect 276416 72525 276472 72581
rect 276540 72525 276596 72581
rect 276664 72525 276720 72581
rect 276788 72525 276844 72581
rect 276912 72525 276968 72581
rect 277036 72525 277092 72581
rect 275176 72401 275232 72457
rect 275300 72401 275356 72457
rect 275424 72401 275480 72457
rect 275548 72401 275604 72457
rect 275672 72401 275728 72457
rect 275796 72401 275852 72457
rect 275920 72401 275976 72457
rect 276044 72401 276100 72457
rect 276168 72401 276224 72457
rect 276292 72401 276348 72457
rect 276416 72401 276472 72457
rect 276540 72401 276596 72457
rect 276664 72401 276720 72457
rect 276788 72401 276844 72457
rect 276912 72401 276968 72457
rect 277036 72401 277092 72457
rect 275176 72277 275232 72333
rect 275300 72277 275356 72333
rect 275424 72277 275480 72333
rect 275548 72277 275604 72333
rect 275672 72277 275728 72333
rect 275796 72277 275852 72333
rect 275920 72277 275976 72333
rect 276044 72277 276100 72333
rect 276168 72277 276224 72333
rect 276292 72277 276348 72333
rect 276416 72277 276472 72333
rect 276540 72277 276596 72333
rect 276664 72277 276720 72333
rect 276788 72277 276844 72333
rect 276912 72277 276968 72333
rect 277036 72277 277092 72333
rect 275176 72153 275232 72209
rect 275300 72153 275356 72209
rect 275424 72153 275480 72209
rect 275548 72153 275604 72209
rect 275672 72153 275728 72209
rect 275796 72153 275852 72209
rect 275920 72153 275976 72209
rect 276044 72153 276100 72209
rect 276168 72153 276224 72209
rect 276292 72153 276348 72209
rect 276416 72153 276472 72209
rect 276540 72153 276596 72209
rect 276664 72153 276720 72209
rect 276788 72153 276844 72209
rect 276912 72153 276968 72209
rect 277036 72153 277092 72209
rect 277882 73889 277938 73945
rect 278006 73889 278062 73945
rect 278130 73889 278186 73945
rect 278254 73889 278310 73945
rect 278378 73889 278434 73945
rect 278502 73889 278558 73945
rect 278626 73889 278682 73945
rect 278750 73889 278806 73945
rect 278874 73889 278930 73945
rect 278998 73889 279054 73945
rect 279122 73889 279178 73945
rect 279246 73889 279302 73945
rect 279370 73889 279426 73945
rect 279494 73889 279550 73945
rect 279618 73889 279674 73945
rect 279742 73889 279798 73945
rect 277882 73765 277938 73821
rect 278006 73765 278062 73821
rect 278130 73765 278186 73821
rect 278254 73765 278310 73821
rect 278378 73765 278434 73821
rect 278502 73765 278558 73821
rect 278626 73765 278682 73821
rect 278750 73765 278806 73821
rect 278874 73765 278930 73821
rect 278998 73765 279054 73821
rect 279122 73765 279178 73821
rect 279246 73765 279302 73821
rect 279370 73765 279426 73821
rect 279494 73765 279550 73821
rect 279618 73765 279674 73821
rect 279742 73765 279798 73821
rect 277882 73641 277938 73697
rect 278006 73641 278062 73697
rect 278130 73641 278186 73697
rect 278254 73641 278310 73697
rect 278378 73641 278434 73697
rect 278502 73641 278558 73697
rect 278626 73641 278682 73697
rect 278750 73641 278806 73697
rect 278874 73641 278930 73697
rect 278998 73641 279054 73697
rect 279122 73641 279178 73697
rect 279246 73641 279302 73697
rect 279370 73641 279426 73697
rect 279494 73641 279550 73697
rect 279618 73641 279674 73697
rect 279742 73641 279798 73697
rect 277882 73517 277938 73573
rect 278006 73517 278062 73573
rect 278130 73517 278186 73573
rect 278254 73517 278310 73573
rect 278378 73517 278434 73573
rect 278502 73517 278558 73573
rect 278626 73517 278682 73573
rect 278750 73517 278806 73573
rect 278874 73517 278930 73573
rect 278998 73517 279054 73573
rect 279122 73517 279178 73573
rect 279246 73517 279302 73573
rect 279370 73517 279426 73573
rect 279494 73517 279550 73573
rect 279618 73517 279674 73573
rect 279742 73517 279798 73573
rect 277882 73393 277938 73449
rect 278006 73393 278062 73449
rect 278130 73393 278186 73449
rect 278254 73393 278310 73449
rect 278378 73393 278434 73449
rect 278502 73393 278558 73449
rect 278626 73393 278682 73449
rect 278750 73393 278806 73449
rect 278874 73393 278930 73449
rect 278998 73393 279054 73449
rect 279122 73393 279178 73449
rect 279246 73393 279302 73449
rect 279370 73393 279426 73449
rect 279494 73393 279550 73449
rect 279618 73393 279674 73449
rect 279742 73393 279798 73449
rect 277882 73269 277938 73325
rect 278006 73269 278062 73325
rect 278130 73269 278186 73325
rect 278254 73269 278310 73325
rect 278378 73269 278434 73325
rect 278502 73269 278558 73325
rect 278626 73269 278682 73325
rect 278750 73269 278806 73325
rect 278874 73269 278930 73325
rect 278998 73269 279054 73325
rect 279122 73269 279178 73325
rect 279246 73269 279302 73325
rect 279370 73269 279426 73325
rect 279494 73269 279550 73325
rect 279618 73269 279674 73325
rect 279742 73269 279798 73325
rect 277882 73145 277938 73201
rect 278006 73145 278062 73201
rect 278130 73145 278186 73201
rect 278254 73145 278310 73201
rect 278378 73145 278434 73201
rect 278502 73145 278558 73201
rect 278626 73145 278682 73201
rect 278750 73145 278806 73201
rect 278874 73145 278930 73201
rect 278998 73145 279054 73201
rect 279122 73145 279178 73201
rect 279246 73145 279302 73201
rect 279370 73145 279426 73201
rect 279494 73145 279550 73201
rect 279618 73145 279674 73201
rect 279742 73145 279798 73201
rect 277882 73021 277938 73077
rect 278006 73021 278062 73077
rect 278130 73021 278186 73077
rect 278254 73021 278310 73077
rect 278378 73021 278434 73077
rect 278502 73021 278558 73077
rect 278626 73021 278682 73077
rect 278750 73021 278806 73077
rect 278874 73021 278930 73077
rect 278998 73021 279054 73077
rect 279122 73021 279178 73077
rect 279246 73021 279302 73077
rect 279370 73021 279426 73077
rect 279494 73021 279550 73077
rect 279618 73021 279674 73077
rect 279742 73021 279798 73077
rect 277882 72897 277938 72953
rect 278006 72897 278062 72953
rect 278130 72897 278186 72953
rect 278254 72897 278310 72953
rect 278378 72897 278434 72953
rect 278502 72897 278558 72953
rect 278626 72897 278682 72953
rect 278750 72897 278806 72953
rect 278874 72897 278930 72953
rect 278998 72897 279054 72953
rect 279122 72897 279178 72953
rect 279246 72897 279302 72953
rect 279370 72897 279426 72953
rect 279494 72897 279550 72953
rect 279618 72897 279674 72953
rect 279742 72897 279798 72953
rect 277882 72773 277938 72829
rect 278006 72773 278062 72829
rect 278130 72773 278186 72829
rect 278254 72773 278310 72829
rect 278378 72773 278434 72829
rect 278502 72773 278558 72829
rect 278626 72773 278682 72829
rect 278750 72773 278806 72829
rect 278874 72773 278930 72829
rect 278998 72773 279054 72829
rect 279122 72773 279178 72829
rect 279246 72773 279302 72829
rect 279370 72773 279426 72829
rect 279494 72773 279550 72829
rect 279618 72773 279674 72829
rect 279742 72773 279798 72829
rect 277882 72649 277938 72705
rect 278006 72649 278062 72705
rect 278130 72649 278186 72705
rect 278254 72649 278310 72705
rect 278378 72649 278434 72705
rect 278502 72649 278558 72705
rect 278626 72649 278682 72705
rect 278750 72649 278806 72705
rect 278874 72649 278930 72705
rect 278998 72649 279054 72705
rect 279122 72649 279178 72705
rect 279246 72649 279302 72705
rect 279370 72649 279426 72705
rect 279494 72649 279550 72705
rect 279618 72649 279674 72705
rect 279742 72649 279798 72705
rect 277882 72525 277938 72581
rect 278006 72525 278062 72581
rect 278130 72525 278186 72581
rect 278254 72525 278310 72581
rect 278378 72525 278434 72581
rect 278502 72525 278558 72581
rect 278626 72525 278682 72581
rect 278750 72525 278806 72581
rect 278874 72525 278930 72581
rect 278998 72525 279054 72581
rect 279122 72525 279178 72581
rect 279246 72525 279302 72581
rect 279370 72525 279426 72581
rect 279494 72525 279550 72581
rect 279618 72525 279674 72581
rect 279742 72525 279798 72581
rect 277882 72401 277938 72457
rect 278006 72401 278062 72457
rect 278130 72401 278186 72457
rect 278254 72401 278310 72457
rect 278378 72401 278434 72457
rect 278502 72401 278558 72457
rect 278626 72401 278682 72457
rect 278750 72401 278806 72457
rect 278874 72401 278930 72457
rect 278998 72401 279054 72457
rect 279122 72401 279178 72457
rect 279246 72401 279302 72457
rect 279370 72401 279426 72457
rect 279494 72401 279550 72457
rect 279618 72401 279674 72457
rect 279742 72401 279798 72457
rect 277882 72277 277938 72333
rect 278006 72277 278062 72333
rect 278130 72277 278186 72333
rect 278254 72277 278310 72333
rect 278378 72277 278434 72333
rect 278502 72277 278558 72333
rect 278626 72277 278682 72333
rect 278750 72277 278806 72333
rect 278874 72277 278930 72333
rect 278998 72277 279054 72333
rect 279122 72277 279178 72333
rect 279246 72277 279302 72333
rect 279370 72277 279426 72333
rect 279494 72277 279550 72333
rect 279618 72277 279674 72333
rect 279742 72277 279798 72333
rect 277882 72153 277938 72209
rect 278006 72153 278062 72209
rect 278130 72153 278186 72209
rect 278254 72153 278310 72209
rect 278378 72153 278434 72209
rect 278502 72153 278558 72209
rect 278626 72153 278682 72209
rect 278750 72153 278806 72209
rect 278874 72153 278930 72209
rect 278998 72153 279054 72209
rect 279122 72153 279178 72209
rect 279246 72153 279302 72209
rect 279370 72153 279426 72209
rect 279494 72153 279550 72209
rect 279618 72153 279674 72209
rect 279742 72153 279798 72209
rect 280252 73889 280308 73945
rect 280376 73889 280432 73945
rect 280500 73889 280556 73945
rect 280624 73889 280680 73945
rect 280748 73889 280804 73945
rect 280872 73889 280928 73945
rect 280996 73889 281052 73945
rect 281120 73889 281176 73945
rect 281244 73889 281300 73945
rect 281368 73889 281424 73945
rect 281492 73889 281548 73945
rect 281616 73889 281672 73945
rect 281740 73889 281796 73945
rect 281864 73889 281920 73945
rect 281988 73889 282044 73945
rect 282112 73889 282168 73945
rect 280252 73765 280308 73821
rect 280376 73765 280432 73821
rect 280500 73765 280556 73821
rect 280624 73765 280680 73821
rect 280748 73765 280804 73821
rect 280872 73765 280928 73821
rect 280996 73765 281052 73821
rect 281120 73765 281176 73821
rect 281244 73765 281300 73821
rect 281368 73765 281424 73821
rect 281492 73765 281548 73821
rect 281616 73765 281672 73821
rect 281740 73765 281796 73821
rect 281864 73765 281920 73821
rect 281988 73765 282044 73821
rect 282112 73765 282168 73821
rect 280252 73641 280308 73697
rect 280376 73641 280432 73697
rect 280500 73641 280556 73697
rect 280624 73641 280680 73697
rect 280748 73641 280804 73697
rect 280872 73641 280928 73697
rect 280996 73641 281052 73697
rect 281120 73641 281176 73697
rect 281244 73641 281300 73697
rect 281368 73641 281424 73697
rect 281492 73641 281548 73697
rect 281616 73641 281672 73697
rect 281740 73641 281796 73697
rect 281864 73641 281920 73697
rect 281988 73641 282044 73697
rect 282112 73641 282168 73697
rect 280252 73517 280308 73573
rect 280376 73517 280432 73573
rect 280500 73517 280556 73573
rect 280624 73517 280680 73573
rect 280748 73517 280804 73573
rect 280872 73517 280928 73573
rect 280996 73517 281052 73573
rect 281120 73517 281176 73573
rect 281244 73517 281300 73573
rect 281368 73517 281424 73573
rect 281492 73517 281548 73573
rect 281616 73517 281672 73573
rect 281740 73517 281796 73573
rect 281864 73517 281920 73573
rect 281988 73517 282044 73573
rect 282112 73517 282168 73573
rect 280252 73393 280308 73449
rect 280376 73393 280432 73449
rect 280500 73393 280556 73449
rect 280624 73393 280680 73449
rect 280748 73393 280804 73449
rect 280872 73393 280928 73449
rect 280996 73393 281052 73449
rect 281120 73393 281176 73449
rect 281244 73393 281300 73449
rect 281368 73393 281424 73449
rect 281492 73393 281548 73449
rect 281616 73393 281672 73449
rect 281740 73393 281796 73449
rect 281864 73393 281920 73449
rect 281988 73393 282044 73449
rect 282112 73393 282168 73449
rect 280252 73269 280308 73325
rect 280376 73269 280432 73325
rect 280500 73269 280556 73325
rect 280624 73269 280680 73325
rect 280748 73269 280804 73325
rect 280872 73269 280928 73325
rect 280996 73269 281052 73325
rect 281120 73269 281176 73325
rect 281244 73269 281300 73325
rect 281368 73269 281424 73325
rect 281492 73269 281548 73325
rect 281616 73269 281672 73325
rect 281740 73269 281796 73325
rect 281864 73269 281920 73325
rect 281988 73269 282044 73325
rect 282112 73269 282168 73325
rect 280252 73145 280308 73201
rect 280376 73145 280432 73201
rect 280500 73145 280556 73201
rect 280624 73145 280680 73201
rect 280748 73145 280804 73201
rect 280872 73145 280928 73201
rect 280996 73145 281052 73201
rect 281120 73145 281176 73201
rect 281244 73145 281300 73201
rect 281368 73145 281424 73201
rect 281492 73145 281548 73201
rect 281616 73145 281672 73201
rect 281740 73145 281796 73201
rect 281864 73145 281920 73201
rect 281988 73145 282044 73201
rect 282112 73145 282168 73201
rect 280252 73021 280308 73077
rect 280376 73021 280432 73077
rect 280500 73021 280556 73077
rect 280624 73021 280680 73077
rect 280748 73021 280804 73077
rect 280872 73021 280928 73077
rect 280996 73021 281052 73077
rect 281120 73021 281176 73077
rect 281244 73021 281300 73077
rect 281368 73021 281424 73077
rect 281492 73021 281548 73077
rect 281616 73021 281672 73077
rect 281740 73021 281796 73077
rect 281864 73021 281920 73077
rect 281988 73021 282044 73077
rect 282112 73021 282168 73077
rect 280252 72897 280308 72953
rect 280376 72897 280432 72953
rect 280500 72897 280556 72953
rect 280624 72897 280680 72953
rect 280748 72897 280804 72953
rect 280872 72897 280928 72953
rect 280996 72897 281052 72953
rect 281120 72897 281176 72953
rect 281244 72897 281300 72953
rect 281368 72897 281424 72953
rect 281492 72897 281548 72953
rect 281616 72897 281672 72953
rect 281740 72897 281796 72953
rect 281864 72897 281920 72953
rect 281988 72897 282044 72953
rect 282112 72897 282168 72953
rect 280252 72773 280308 72829
rect 280376 72773 280432 72829
rect 280500 72773 280556 72829
rect 280624 72773 280680 72829
rect 280748 72773 280804 72829
rect 280872 72773 280928 72829
rect 280996 72773 281052 72829
rect 281120 72773 281176 72829
rect 281244 72773 281300 72829
rect 281368 72773 281424 72829
rect 281492 72773 281548 72829
rect 281616 72773 281672 72829
rect 281740 72773 281796 72829
rect 281864 72773 281920 72829
rect 281988 72773 282044 72829
rect 282112 72773 282168 72829
rect 280252 72649 280308 72705
rect 280376 72649 280432 72705
rect 280500 72649 280556 72705
rect 280624 72649 280680 72705
rect 280748 72649 280804 72705
rect 280872 72649 280928 72705
rect 280996 72649 281052 72705
rect 281120 72649 281176 72705
rect 281244 72649 281300 72705
rect 281368 72649 281424 72705
rect 281492 72649 281548 72705
rect 281616 72649 281672 72705
rect 281740 72649 281796 72705
rect 281864 72649 281920 72705
rect 281988 72649 282044 72705
rect 282112 72649 282168 72705
rect 280252 72525 280308 72581
rect 280376 72525 280432 72581
rect 280500 72525 280556 72581
rect 280624 72525 280680 72581
rect 280748 72525 280804 72581
rect 280872 72525 280928 72581
rect 280996 72525 281052 72581
rect 281120 72525 281176 72581
rect 281244 72525 281300 72581
rect 281368 72525 281424 72581
rect 281492 72525 281548 72581
rect 281616 72525 281672 72581
rect 281740 72525 281796 72581
rect 281864 72525 281920 72581
rect 281988 72525 282044 72581
rect 282112 72525 282168 72581
rect 280252 72401 280308 72457
rect 280376 72401 280432 72457
rect 280500 72401 280556 72457
rect 280624 72401 280680 72457
rect 280748 72401 280804 72457
rect 280872 72401 280928 72457
rect 280996 72401 281052 72457
rect 281120 72401 281176 72457
rect 281244 72401 281300 72457
rect 281368 72401 281424 72457
rect 281492 72401 281548 72457
rect 281616 72401 281672 72457
rect 281740 72401 281796 72457
rect 281864 72401 281920 72457
rect 281988 72401 282044 72457
rect 282112 72401 282168 72457
rect 280252 72277 280308 72333
rect 280376 72277 280432 72333
rect 280500 72277 280556 72333
rect 280624 72277 280680 72333
rect 280748 72277 280804 72333
rect 280872 72277 280928 72333
rect 280996 72277 281052 72333
rect 281120 72277 281176 72333
rect 281244 72277 281300 72333
rect 281368 72277 281424 72333
rect 281492 72277 281548 72333
rect 281616 72277 281672 72333
rect 281740 72277 281796 72333
rect 281864 72277 281920 72333
rect 281988 72277 282044 72333
rect 282112 72277 282168 72333
rect 280252 72153 280308 72209
rect 280376 72153 280432 72209
rect 280500 72153 280556 72209
rect 280624 72153 280680 72209
rect 280748 72153 280804 72209
rect 280872 72153 280928 72209
rect 280996 72153 281052 72209
rect 281120 72153 281176 72209
rect 281244 72153 281300 72209
rect 281368 72153 281424 72209
rect 281492 72153 281548 72209
rect 281616 72153 281672 72209
rect 281740 72153 281796 72209
rect 281864 72153 281920 72209
rect 281988 72153 282044 72209
rect 282112 72153 282168 72209
rect 282882 73889 282938 73945
rect 283006 73889 283062 73945
rect 283130 73889 283186 73945
rect 283254 73889 283310 73945
rect 283378 73889 283434 73945
rect 283502 73889 283558 73945
rect 283626 73889 283682 73945
rect 283750 73889 283806 73945
rect 283874 73889 283930 73945
rect 282882 73765 282938 73821
rect 283006 73765 283062 73821
rect 283130 73765 283186 73821
rect 283254 73765 283310 73821
rect 283378 73765 283434 73821
rect 283502 73765 283558 73821
rect 283626 73765 283682 73821
rect 283750 73765 283806 73821
rect 283874 73765 283930 73821
rect 282882 73641 282938 73697
rect 283006 73641 283062 73697
rect 283130 73641 283186 73697
rect 283254 73641 283310 73697
rect 283378 73641 283434 73697
rect 283502 73641 283558 73697
rect 283626 73641 283682 73697
rect 283750 73641 283806 73697
rect 283874 73641 283930 73697
rect 282882 73517 282938 73573
rect 283006 73517 283062 73573
rect 283130 73517 283186 73573
rect 283254 73517 283310 73573
rect 283378 73517 283434 73573
rect 283502 73517 283558 73573
rect 283626 73517 283682 73573
rect 283750 73517 283806 73573
rect 283874 73517 283930 73573
rect 282882 73393 282938 73449
rect 283006 73393 283062 73449
rect 283130 73393 283186 73449
rect 283254 73393 283310 73449
rect 283378 73393 283434 73449
rect 283502 73393 283558 73449
rect 283626 73393 283682 73449
rect 283750 73393 283806 73449
rect 283874 73393 283930 73449
rect 282882 73269 282938 73325
rect 283006 73269 283062 73325
rect 283130 73269 283186 73325
rect 283254 73269 283310 73325
rect 283378 73269 283434 73325
rect 283502 73269 283558 73325
rect 283626 73269 283682 73325
rect 283750 73269 283806 73325
rect 283874 73269 283930 73325
rect 282882 73145 282938 73201
rect 283006 73145 283062 73201
rect 283130 73145 283186 73201
rect 283254 73145 283310 73201
rect 283378 73145 283434 73201
rect 283502 73145 283558 73201
rect 283626 73145 283682 73201
rect 283750 73145 283806 73201
rect 283874 73145 283930 73201
rect 282882 73021 282938 73077
rect 283006 73021 283062 73077
rect 283130 73021 283186 73077
rect 283254 73021 283310 73077
rect 283378 73021 283434 73077
rect 283502 73021 283558 73077
rect 283626 73021 283682 73077
rect 283750 73021 283806 73077
rect 283874 73021 283930 73077
rect 282882 72897 282938 72953
rect 283006 72897 283062 72953
rect 283130 72897 283186 72953
rect 283254 72897 283310 72953
rect 283378 72897 283434 72953
rect 283502 72897 283558 72953
rect 283626 72897 283682 72953
rect 283750 72897 283806 72953
rect 283874 72897 283930 72953
rect 282882 72773 282938 72829
rect 283006 72773 283062 72829
rect 283130 72773 283186 72829
rect 283254 72773 283310 72829
rect 283378 72773 283434 72829
rect 283502 72773 283558 72829
rect 283626 72773 283682 72829
rect 283750 72773 283806 72829
rect 283874 72773 283930 72829
rect 282882 72649 282938 72705
rect 283006 72649 283062 72705
rect 283130 72649 283186 72705
rect 283254 72649 283310 72705
rect 283378 72649 283434 72705
rect 283502 72649 283558 72705
rect 283626 72649 283682 72705
rect 283750 72649 283806 72705
rect 283874 72649 283930 72705
rect 282882 72525 282938 72581
rect 283006 72525 283062 72581
rect 283130 72525 283186 72581
rect 283254 72525 283310 72581
rect 283378 72525 283434 72581
rect 283502 72525 283558 72581
rect 283626 72525 283682 72581
rect 283750 72525 283806 72581
rect 283874 72525 283930 72581
rect 282882 72401 282938 72457
rect 283006 72401 283062 72457
rect 283130 72401 283186 72457
rect 283254 72401 283310 72457
rect 283378 72401 283434 72457
rect 283502 72401 283558 72457
rect 283626 72401 283682 72457
rect 283750 72401 283806 72457
rect 283874 72401 283930 72457
rect 282882 72277 282938 72333
rect 283006 72277 283062 72333
rect 283130 72277 283186 72333
rect 283254 72277 283310 72333
rect 283378 72277 283434 72333
rect 283502 72277 283558 72333
rect 283626 72277 283682 72333
rect 283750 72277 283806 72333
rect 283874 72277 283930 72333
rect 282882 72153 282938 72209
rect 283006 72153 283062 72209
rect 283130 72153 283186 72209
rect 283254 72153 283310 72209
rect 283378 72153 283434 72209
rect 283502 72153 283558 72209
rect 283626 72153 283682 72209
rect 283750 72153 283806 72209
rect 283874 72153 283930 72209
rect 600326 73889 600382 73945
rect 600450 73889 600506 73945
rect 600574 73889 600630 73945
rect 600698 73889 600754 73945
rect 600822 73889 600878 73945
rect 600946 73889 601002 73945
rect 601070 73889 601126 73945
rect 601194 73889 601250 73945
rect 601318 73889 601374 73945
rect 601442 73889 601498 73945
rect 601566 73889 601622 73945
rect 601690 73889 601746 73945
rect 601814 73889 601870 73945
rect 601938 73889 601994 73945
rect 602062 73889 602118 73945
rect 600326 73765 600382 73821
rect 600450 73765 600506 73821
rect 600574 73765 600630 73821
rect 600698 73765 600754 73821
rect 600822 73765 600878 73821
rect 600946 73765 601002 73821
rect 601070 73765 601126 73821
rect 601194 73765 601250 73821
rect 601318 73765 601374 73821
rect 601442 73765 601498 73821
rect 601566 73765 601622 73821
rect 601690 73765 601746 73821
rect 601814 73765 601870 73821
rect 601938 73765 601994 73821
rect 602062 73765 602118 73821
rect 600326 73641 600382 73697
rect 600450 73641 600506 73697
rect 600574 73641 600630 73697
rect 600698 73641 600754 73697
rect 600822 73641 600878 73697
rect 600946 73641 601002 73697
rect 601070 73641 601126 73697
rect 601194 73641 601250 73697
rect 601318 73641 601374 73697
rect 601442 73641 601498 73697
rect 601566 73641 601622 73697
rect 601690 73641 601746 73697
rect 601814 73641 601870 73697
rect 601938 73641 601994 73697
rect 602062 73641 602118 73697
rect 600326 73517 600382 73573
rect 600450 73517 600506 73573
rect 600574 73517 600630 73573
rect 600698 73517 600754 73573
rect 600822 73517 600878 73573
rect 600946 73517 601002 73573
rect 601070 73517 601126 73573
rect 601194 73517 601250 73573
rect 601318 73517 601374 73573
rect 601442 73517 601498 73573
rect 601566 73517 601622 73573
rect 601690 73517 601746 73573
rect 601814 73517 601870 73573
rect 601938 73517 601994 73573
rect 602062 73517 602118 73573
rect 600326 73393 600382 73449
rect 600450 73393 600506 73449
rect 600574 73393 600630 73449
rect 600698 73393 600754 73449
rect 600822 73393 600878 73449
rect 600946 73393 601002 73449
rect 601070 73393 601126 73449
rect 601194 73393 601250 73449
rect 601318 73393 601374 73449
rect 601442 73393 601498 73449
rect 601566 73393 601622 73449
rect 601690 73393 601746 73449
rect 601814 73393 601870 73449
rect 601938 73393 601994 73449
rect 602062 73393 602118 73449
rect 600326 73269 600382 73325
rect 600450 73269 600506 73325
rect 600574 73269 600630 73325
rect 600698 73269 600754 73325
rect 600822 73269 600878 73325
rect 600946 73269 601002 73325
rect 601070 73269 601126 73325
rect 601194 73269 601250 73325
rect 601318 73269 601374 73325
rect 601442 73269 601498 73325
rect 601566 73269 601622 73325
rect 601690 73269 601746 73325
rect 601814 73269 601870 73325
rect 601938 73269 601994 73325
rect 602062 73269 602118 73325
rect 600326 73145 600382 73201
rect 600450 73145 600506 73201
rect 600574 73145 600630 73201
rect 600698 73145 600754 73201
rect 600822 73145 600878 73201
rect 600946 73145 601002 73201
rect 601070 73145 601126 73201
rect 601194 73145 601250 73201
rect 601318 73145 601374 73201
rect 601442 73145 601498 73201
rect 601566 73145 601622 73201
rect 601690 73145 601746 73201
rect 601814 73145 601870 73201
rect 601938 73145 601994 73201
rect 602062 73145 602118 73201
rect 600326 73021 600382 73077
rect 600450 73021 600506 73077
rect 600574 73021 600630 73077
rect 600698 73021 600754 73077
rect 600822 73021 600878 73077
rect 600946 73021 601002 73077
rect 601070 73021 601126 73077
rect 601194 73021 601250 73077
rect 601318 73021 601374 73077
rect 601442 73021 601498 73077
rect 601566 73021 601622 73077
rect 601690 73021 601746 73077
rect 601814 73021 601870 73077
rect 601938 73021 601994 73077
rect 602062 73021 602118 73077
rect 600326 72897 600382 72953
rect 600450 72897 600506 72953
rect 600574 72897 600630 72953
rect 600698 72897 600754 72953
rect 600822 72897 600878 72953
rect 600946 72897 601002 72953
rect 601070 72897 601126 72953
rect 601194 72897 601250 72953
rect 601318 72897 601374 72953
rect 601442 72897 601498 72953
rect 601566 72897 601622 72953
rect 601690 72897 601746 72953
rect 601814 72897 601870 72953
rect 601938 72897 601994 72953
rect 602062 72897 602118 72953
rect 600326 72773 600382 72829
rect 600450 72773 600506 72829
rect 600574 72773 600630 72829
rect 600698 72773 600754 72829
rect 600822 72773 600878 72829
rect 600946 72773 601002 72829
rect 601070 72773 601126 72829
rect 601194 72773 601250 72829
rect 601318 72773 601374 72829
rect 601442 72773 601498 72829
rect 601566 72773 601622 72829
rect 601690 72773 601746 72829
rect 601814 72773 601870 72829
rect 601938 72773 601994 72829
rect 602062 72773 602118 72829
rect 600326 72649 600382 72705
rect 600450 72649 600506 72705
rect 600574 72649 600630 72705
rect 600698 72649 600754 72705
rect 600822 72649 600878 72705
rect 600946 72649 601002 72705
rect 601070 72649 601126 72705
rect 601194 72649 601250 72705
rect 601318 72649 601374 72705
rect 601442 72649 601498 72705
rect 601566 72649 601622 72705
rect 601690 72649 601746 72705
rect 601814 72649 601870 72705
rect 601938 72649 601994 72705
rect 602062 72649 602118 72705
rect 600326 72525 600382 72581
rect 600450 72525 600506 72581
rect 600574 72525 600630 72581
rect 600698 72525 600754 72581
rect 600822 72525 600878 72581
rect 600946 72525 601002 72581
rect 601070 72525 601126 72581
rect 601194 72525 601250 72581
rect 601318 72525 601374 72581
rect 601442 72525 601498 72581
rect 601566 72525 601622 72581
rect 601690 72525 601746 72581
rect 601814 72525 601870 72581
rect 601938 72525 601994 72581
rect 602062 72525 602118 72581
rect 600326 72401 600382 72457
rect 600450 72401 600506 72457
rect 600574 72401 600630 72457
rect 600698 72401 600754 72457
rect 600822 72401 600878 72457
rect 600946 72401 601002 72457
rect 601070 72401 601126 72457
rect 601194 72401 601250 72457
rect 601318 72401 601374 72457
rect 601442 72401 601498 72457
rect 601566 72401 601622 72457
rect 601690 72401 601746 72457
rect 601814 72401 601870 72457
rect 601938 72401 601994 72457
rect 602062 72401 602118 72457
rect 600326 72277 600382 72333
rect 600450 72277 600506 72333
rect 600574 72277 600630 72333
rect 600698 72277 600754 72333
rect 600822 72277 600878 72333
rect 600946 72277 601002 72333
rect 601070 72277 601126 72333
rect 601194 72277 601250 72333
rect 601318 72277 601374 72333
rect 601442 72277 601498 72333
rect 601566 72277 601622 72333
rect 601690 72277 601746 72333
rect 601814 72277 601870 72333
rect 601938 72277 601994 72333
rect 602062 72277 602118 72333
rect 600326 72153 600382 72209
rect 600450 72153 600506 72209
rect 600574 72153 600630 72209
rect 600698 72153 600754 72209
rect 600822 72153 600878 72209
rect 600946 72153 601002 72209
rect 601070 72153 601126 72209
rect 601194 72153 601250 72209
rect 601318 72153 601374 72209
rect 601442 72153 601498 72209
rect 601566 72153 601622 72209
rect 601690 72153 601746 72209
rect 601814 72153 601870 72209
rect 601938 72153 601994 72209
rect 602062 72153 602118 72209
rect 602806 73889 602862 73945
rect 602930 73889 602986 73945
rect 603054 73889 603110 73945
rect 603178 73889 603234 73945
rect 603302 73889 603358 73945
rect 603426 73889 603482 73945
rect 603550 73889 603606 73945
rect 603674 73889 603730 73945
rect 603798 73889 603854 73945
rect 603922 73889 603978 73945
rect 602806 73765 602862 73821
rect 602930 73765 602986 73821
rect 603054 73765 603110 73821
rect 603178 73765 603234 73821
rect 603302 73765 603358 73821
rect 603426 73765 603482 73821
rect 603550 73765 603606 73821
rect 603674 73765 603730 73821
rect 603798 73765 603854 73821
rect 603922 73765 603978 73821
rect 602806 73641 602862 73697
rect 602930 73641 602986 73697
rect 603054 73641 603110 73697
rect 603178 73641 603234 73697
rect 603302 73641 603358 73697
rect 603426 73641 603482 73697
rect 603550 73641 603606 73697
rect 603674 73641 603730 73697
rect 603798 73641 603854 73697
rect 603922 73641 603978 73697
rect 602806 73517 602862 73573
rect 602930 73517 602986 73573
rect 603054 73517 603110 73573
rect 603178 73517 603234 73573
rect 603302 73517 603358 73573
rect 603426 73517 603482 73573
rect 603550 73517 603606 73573
rect 603674 73517 603730 73573
rect 603798 73517 603854 73573
rect 603922 73517 603978 73573
rect 602806 73393 602862 73449
rect 602930 73393 602986 73449
rect 603054 73393 603110 73449
rect 603178 73393 603234 73449
rect 603302 73393 603358 73449
rect 603426 73393 603482 73449
rect 603550 73393 603606 73449
rect 603674 73393 603730 73449
rect 603798 73393 603854 73449
rect 603922 73393 603978 73449
rect 602806 73269 602862 73325
rect 602930 73269 602986 73325
rect 603054 73269 603110 73325
rect 603178 73269 603234 73325
rect 603302 73269 603358 73325
rect 603426 73269 603482 73325
rect 603550 73269 603606 73325
rect 603674 73269 603730 73325
rect 603798 73269 603854 73325
rect 603922 73269 603978 73325
rect 602806 73145 602862 73201
rect 602930 73145 602986 73201
rect 603054 73145 603110 73201
rect 603178 73145 603234 73201
rect 603302 73145 603358 73201
rect 603426 73145 603482 73201
rect 603550 73145 603606 73201
rect 603674 73145 603730 73201
rect 603798 73145 603854 73201
rect 603922 73145 603978 73201
rect 602806 73021 602862 73077
rect 602930 73021 602986 73077
rect 603054 73021 603110 73077
rect 603178 73021 603234 73077
rect 603302 73021 603358 73077
rect 603426 73021 603482 73077
rect 603550 73021 603606 73077
rect 603674 73021 603730 73077
rect 603798 73021 603854 73077
rect 603922 73021 603978 73077
rect 602806 72897 602862 72953
rect 602930 72897 602986 72953
rect 603054 72897 603110 72953
rect 603178 72897 603234 72953
rect 603302 72897 603358 72953
rect 603426 72897 603482 72953
rect 603550 72897 603606 72953
rect 603674 72897 603730 72953
rect 603798 72897 603854 72953
rect 603922 72897 603978 72953
rect 602806 72773 602862 72829
rect 602930 72773 602986 72829
rect 603054 72773 603110 72829
rect 603178 72773 603234 72829
rect 603302 72773 603358 72829
rect 603426 72773 603482 72829
rect 603550 72773 603606 72829
rect 603674 72773 603730 72829
rect 603798 72773 603854 72829
rect 603922 72773 603978 72829
rect 602806 72649 602862 72705
rect 602930 72649 602986 72705
rect 603054 72649 603110 72705
rect 603178 72649 603234 72705
rect 603302 72649 603358 72705
rect 603426 72649 603482 72705
rect 603550 72649 603606 72705
rect 603674 72649 603730 72705
rect 603798 72649 603854 72705
rect 603922 72649 603978 72705
rect 602806 72525 602862 72581
rect 602930 72525 602986 72581
rect 603054 72525 603110 72581
rect 603178 72525 603234 72581
rect 603302 72525 603358 72581
rect 603426 72525 603482 72581
rect 603550 72525 603606 72581
rect 603674 72525 603730 72581
rect 603798 72525 603854 72581
rect 603922 72525 603978 72581
rect 602806 72401 602862 72457
rect 602930 72401 602986 72457
rect 603054 72401 603110 72457
rect 603178 72401 603234 72457
rect 603302 72401 603358 72457
rect 603426 72401 603482 72457
rect 603550 72401 603606 72457
rect 603674 72401 603730 72457
rect 603798 72401 603854 72457
rect 603922 72401 603978 72457
rect 602806 72277 602862 72333
rect 602930 72277 602986 72333
rect 603054 72277 603110 72333
rect 603178 72277 603234 72333
rect 603302 72277 603358 72333
rect 603426 72277 603482 72333
rect 603550 72277 603606 72333
rect 603674 72277 603730 72333
rect 603798 72277 603854 72333
rect 603922 72277 603978 72333
rect 602806 72153 602862 72209
rect 602930 72153 602986 72209
rect 603054 72153 603110 72209
rect 603178 72153 603234 72209
rect 603302 72153 603358 72209
rect 603426 72153 603482 72209
rect 603550 72153 603606 72209
rect 603674 72153 603730 72209
rect 603798 72153 603854 72209
rect 603922 72153 603978 72209
rect 605176 73889 605232 73945
rect 605300 73889 605356 73945
rect 605424 73889 605480 73945
rect 605548 73889 605604 73945
rect 605672 73889 605728 73945
rect 605796 73889 605852 73945
rect 605920 73889 605976 73945
rect 606044 73889 606100 73945
rect 606168 73889 606224 73945
rect 606292 73889 606348 73945
rect 606416 73889 606472 73945
rect 606540 73889 606596 73945
rect 606664 73889 606720 73945
rect 606788 73889 606844 73945
rect 606912 73889 606968 73945
rect 607036 73889 607092 73945
rect 605176 73765 605232 73821
rect 605300 73765 605356 73821
rect 605424 73765 605480 73821
rect 605548 73765 605604 73821
rect 605672 73765 605728 73821
rect 605796 73765 605852 73821
rect 605920 73765 605976 73821
rect 606044 73765 606100 73821
rect 606168 73765 606224 73821
rect 606292 73765 606348 73821
rect 606416 73765 606472 73821
rect 606540 73765 606596 73821
rect 606664 73765 606720 73821
rect 606788 73765 606844 73821
rect 606912 73765 606968 73821
rect 607036 73765 607092 73821
rect 605176 73641 605232 73697
rect 605300 73641 605356 73697
rect 605424 73641 605480 73697
rect 605548 73641 605604 73697
rect 605672 73641 605728 73697
rect 605796 73641 605852 73697
rect 605920 73641 605976 73697
rect 606044 73641 606100 73697
rect 606168 73641 606224 73697
rect 606292 73641 606348 73697
rect 606416 73641 606472 73697
rect 606540 73641 606596 73697
rect 606664 73641 606720 73697
rect 606788 73641 606844 73697
rect 606912 73641 606968 73697
rect 607036 73641 607092 73697
rect 605176 73517 605232 73573
rect 605300 73517 605356 73573
rect 605424 73517 605480 73573
rect 605548 73517 605604 73573
rect 605672 73517 605728 73573
rect 605796 73517 605852 73573
rect 605920 73517 605976 73573
rect 606044 73517 606100 73573
rect 606168 73517 606224 73573
rect 606292 73517 606348 73573
rect 606416 73517 606472 73573
rect 606540 73517 606596 73573
rect 606664 73517 606720 73573
rect 606788 73517 606844 73573
rect 606912 73517 606968 73573
rect 607036 73517 607092 73573
rect 605176 73393 605232 73449
rect 605300 73393 605356 73449
rect 605424 73393 605480 73449
rect 605548 73393 605604 73449
rect 605672 73393 605728 73449
rect 605796 73393 605852 73449
rect 605920 73393 605976 73449
rect 606044 73393 606100 73449
rect 606168 73393 606224 73449
rect 606292 73393 606348 73449
rect 606416 73393 606472 73449
rect 606540 73393 606596 73449
rect 606664 73393 606720 73449
rect 606788 73393 606844 73449
rect 606912 73393 606968 73449
rect 607036 73393 607092 73449
rect 605176 73269 605232 73325
rect 605300 73269 605356 73325
rect 605424 73269 605480 73325
rect 605548 73269 605604 73325
rect 605672 73269 605728 73325
rect 605796 73269 605852 73325
rect 605920 73269 605976 73325
rect 606044 73269 606100 73325
rect 606168 73269 606224 73325
rect 606292 73269 606348 73325
rect 606416 73269 606472 73325
rect 606540 73269 606596 73325
rect 606664 73269 606720 73325
rect 606788 73269 606844 73325
rect 606912 73269 606968 73325
rect 607036 73269 607092 73325
rect 605176 73145 605232 73201
rect 605300 73145 605356 73201
rect 605424 73145 605480 73201
rect 605548 73145 605604 73201
rect 605672 73145 605728 73201
rect 605796 73145 605852 73201
rect 605920 73145 605976 73201
rect 606044 73145 606100 73201
rect 606168 73145 606224 73201
rect 606292 73145 606348 73201
rect 606416 73145 606472 73201
rect 606540 73145 606596 73201
rect 606664 73145 606720 73201
rect 606788 73145 606844 73201
rect 606912 73145 606968 73201
rect 607036 73145 607092 73201
rect 605176 73021 605232 73077
rect 605300 73021 605356 73077
rect 605424 73021 605480 73077
rect 605548 73021 605604 73077
rect 605672 73021 605728 73077
rect 605796 73021 605852 73077
rect 605920 73021 605976 73077
rect 606044 73021 606100 73077
rect 606168 73021 606224 73077
rect 606292 73021 606348 73077
rect 606416 73021 606472 73077
rect 606540 73021 606596 73077
rect 606664 73021 606720 73077
rect 606788 73021 606844 73077
rect 606912 73021 606968 73077
rect 607036 73021 607092 73077
rect 605176 72897 605232 72953
rect 605300 72897 605356 72953
rect 605424 72897 605480 72953
rect 605548 72897 605604 72953
rect 605672 72897 605728 72953
rect 605796 72897 605852 72953
rect 605920 72897 605976 72953
rect 606044 72897 606100 72953
rect 606168 72897 606224 72953
rect 606292 72897 606348 72953
rect 606416 72897 606472 72953
rect 606540 72897 606596 72953
rect 606664 72897 606720 72953
rect 606788 72897 606844 72953
rect 606912 72897 606968 72953
rect 607036 72897 607092 72953
rect 605176 72773 605232 72829
rect 605300 72773 605356 72829
rect 605424 72773 605480 72829
rect 605548 72773 605604 72829
rect 605672 72773 605728 72829
rect 605796 72773 605852 72829
rect 605920 72773 605976 72829
rect 606044 72773 606100 72829
rect 606168 72773 606224 72829
rect 606292 72773 606348 72829
rect 606416 72773 606472 72829
rect 606540 72773 606596 72829
rect 606664 72773 606720 72829
rect 606788 72773 606844 72829
rect 606912 72773 606968 72829
rect 607036 72773 607092 72829
rect 605176 72649 605232 72705
rect 605300 72649 605356 72705
rect 605424 72649 605480 72705
rect 605548 72649 605604 72705
rect 605672 72649 605728 72705
rect 605796 72649 605852 72705
rect 605920 72649 605976 72705
rect 606044 72649 606100 72705
rect 606168 72649 606224 72705
rect 606292 72649 606348 72705
rect 606416 72649 606472 72705
rect 606540 72649 606596 72705
rect 606664 72649 606720 72705
rect 606788 72649 606844 72705
rect 606912 72649 606968 72705
rect 607036 72649 607092 72705
rect 605176 72525 605232 72581
rect 605300 72525 605356 72581
rect 605424 72525 605480 72581
rect 605548 72525 605604 72581
rect 605672 72525 605728 72581
rect 605796 72525 605852 72581
rect 605920 72525 605976 72581
rect 606044 72525 606100 72581
rect 606168 72525 606224 72581
rect 606292 72525 606348 72581
rect 606416 72525 606472 72581
rect 606540 72525 606596 72581
rect 606664 72525 606720 72581
rect 606788 72525 606844 72581
rect 606912 72525 606968 72581
rect 607036 72525 607092 72581
rect 605176 72401 605232 72457
rect 605300 72401 605356 72457
rect 605424 72401 605480 72457
rect 605548 72401 605604 72457
rect 605672 72401 605728 72457
rect 605796 72401 605852 72457
rect 605920 72401 605976 72457
rect 606044 72401 606100 72457
rect 606168 72401 606224 72457
rect 606292 72401 606348 72457
rect 606416 72401 606472 72457
rect 606540 72401 606596 72457
rect 606664 72401 606720 72457
rect 606788 72401 606844 72457
rect 606912 72401 606968 72457
rect 607036 72401 607092 72457
rect 605176 72277 605232 72333
rect 605300 72277 605356 72333
rect 605424 72277 605480 72333
rect 605548 72277 605604 72333
rect 605672 72277 605728 72333
rect 605796 72277 605852 72333
rect 605920 72277 605976 72333
rect 606044 72277 606100 72333
rect 606168 72277 606224 72333
rect 606292 72277 606348 72333
rect 606416 72277 606472 72333
rect 606540 72277 606596 72333
rect 606664 72277 606720 72333
rect 606788 72277 606844 72333
rect 606912 72277 606968 72333
rect 607036 72277 607092 72333
rect 605176 72153 605232 72209
rect 605300 72153 605356 72209
rect 605424 72153 605480 72209
rect 605548 72153 605604 72209
rect 605672 72153 605728 72209
rect 605796 72153 605852 72209
rect 605920 72153 605976 72209
rect 606044 72153 606100 72209
rect 606168 72153 606224 72209
rect 606292 72153 606348 72209
rect 606416 72153 606472 72209
rect 606540 72153 606596 72209
rect 606664 72153 606720 72209
rect 606788 72153 606844 72209
rect 606912 72153 606968 72209
rect 607036 72153 607092 72209
rect 607882 73889 607938 73945
rect 608006 73889 608062 73945
rect 608130 73889 608186 73945
rect 608254 73889 608310 73945
rect 608378 73889 608434 73945
rect 608502 73889 608558 73945
rect 608626 73889 608682 73945
rect 608750 73889 608806 73945
rect 608874 73889 608930 73945
rect 608998 73889 609054 73945
rect 609122 73889 609178 73945
rect 609246 73889 609302 73945
rect 609370 73889 609426 73945
rect 609494 73889 609550 73945
rect 609618 73889 609674 73945
rect 609742 73889 609798 73945
rect 607882 73765 607938 73821
rect 608006 73765 608062 73821
rect 608130 73765 608186 73821
rect 608254 73765 608310 73821
rect 608378 73765 608434 73821
rect 608502 73765 608558 73821
rect 608626 73765 608682 73821
rect 608750 73765 608806 73821
rect 608874 73765 608930 73821
rect 608998 73765 609054 73821
rect 609122 73765 609178 73821
rect 609246 73765 609302 73821
rect 609370 73765 609426 73821
rect 609494 73765 609550 73821
rect 609618 73765 609674 73821
rect 609742 73765 609798 73821
rect 607882 73641 607938 73697
rect 608006 73641 608062 73697
rect 608130 73641 608186 73697
rect 608254 73641 608310 73697
rect 608378 73641 608434 73697
rect 608502 73641 608558 73697
rect 608626 73641 608682 73697
rect 608750 73641 608806 73697
rect 608874 73641 608930 73697
rect 608998 73641 609054 73697
rect 609122 73641 609178 73697
rect 609246 73641 609302 73697
rect 609370 73641 609426 73697
rect 609494 73641 609550 73697
rect 609618 73641 609674 73697
rect 609742 73641 609798 73697
rect 607882 73517 607938 73573
rect 608006 73517 608062 73573
rect 608130 73517 608186 73573
rect 608254 73517 608310 73573
rect 608378 73517 608434 73573
rect 608502 73517 608558 73573
rect 608626 73517 608682 73573
rect 608750 73517 608806 73573
rect 608874 73517 608930 73573
rect 608998 73517 609054 73573
rect 609122 73517 609178 73573
rect 609246 73517 609302 73573
rect 609370 73517 609426 73573
rect 609494 73517 609550 73573
rect 609618 73517 609674 73573
rect 609742 73517 609798 73573
rect 607882 73393 607938 73449
rect 608006 73393 608062 73449
rect 608130 73393 608186 73449
rect 608254 73393 608310 73449
rect 608378 73393 608434 73449
rect 608502 73393 608558 73449
rect 608626 73393 608682 73449
rect 608750 73393 608806 73449
rect 608874 73393 608930 73449
rect 608998 73393 609054 73449
rect 609122 73393 609178 73449
rect 609246 73393 609302 73449
rect 609370 73393 609426 73449
rect 609494 73393 609550 73449
rect 609618 73393 609674 73449
rect 609742 73393 609798 73449
rect 607882 73269 607938 73325
rect 608006 73269 608062 73325
rect 608130 73269 608186 73325
rect 608254 73269 608310 73325
rect 608378 73269 608434 73325
rect 608502 73269 608558 73325
rect 608626 73269 608682 73325
rect 608750 73269 608806 73325
rect 608874 73269 608930 73325
rect 608998 73269 609054 73325
rect 609122 73269 609178 73325
rect 609246 73269 609302 73325
rect 609370 73269 609426 73325
rect 609494 73269 609550 73325
rect 609618 73269 609674 73325
rect 609742 73269 609798 73325
rect 607882 73145 607938 73201
rect 608006 73145 608062 73201
rect 608130 73145 608186 73201
rect 608254 73145 608310 73201
rect 608378 73145 608434 73201
rect 608502 73145 608558 73201
rect 608626 73145 608682 73201
rect 608750 73145 608806 73201
rect 608874 73145 608930 73201
rect 608998 73145 609054 73201
rect 609122 73145 609178 73201
rect 609246 73145 609302 73201
rect 609370 73145 609426 73201
rect 609494 73145 609550 73201
rect 609618 73145 609674 73201
rect 609742 73145 609798 73201
rect 607882 73021 607938 73077
rect 608006 73021 608062 73077
rect 608130 73021 608186 73077
rect 608254 73021 608310 73077
rect 608378 73021 608434 73077
rect 608502 73021 608558 73077
rect 608626 73021 608682 73077
rect 608750 73021 608806 73077
rect 608874 73021 608930 73077
rect 608998 73021 609054 73077
rect 609122 73021 609178 73077
rect 609246 73021 609302 73077
rect 609370 73021 609426 73077
rect 609494 73021 609550 73077
rect 609618 73021 609674 73077
rect 609742 73021 609798 73077
rect 607882 72897 607938 72953
rect 608006 72897 608062 72953
rect 608130 72897 608186 72953
rect 608254 72897 608310 72953
rect 608378 72897 608434 72953
rect 608502 72897 608558 72953
rect 608626 72897 608682 72953
rect 608750 72897 608806 72953
rect 608874 72897 608930 72953
rect 608998 72897 609054 72953
rect 609122 72897 609178 72953
rect 609246 72897 609302 72953
rect 609370 72897 609426 72953
rect 609494 72897 609550 72953
rect 609618 72897 609674 72953
rect 609742 72897 609798 72953
rect 607882 72773 607938 72829
rect 608006 72773 608062 72829
rect 608130 72773 608186 72829
rect 608254 72773 608310 72829
rect 608378 72773 608434 72829
rect 608502 72773 608558 72829
rect 608626 72773 608682 72829
rect 608750 72773 608806 72829
rect 608874 72773 608930 72829
rect 608998 72773 609054 72829
rect 609122 72773 609178 72829
rect 609246 72773 609302 72829
rect 609370 72773 609426 72829
rect 609494 72773 609550 72829
rect 609618 72773 609674 72829
rect 609742 72773 609798 72829
rect 607882 72649 607938 72705
rect 608006 72649 608062 72705
rect 608130 72649 608186 72705
rect 608254 72649 608310 72705
rect 608378 72649 608434 72705
rect 608502 72649 608558 72705
rect 608626 72649 608682 72705
rect 608750 72649 608806 72705
rect 608874 72649 608930 72705
rect 608998 72649 609054 72705
rect 609122 72649 609178 72705
rect 609246 72649 609302 72705
rect 609370 72649 609426 72705
rect 609494 72649 609550 72705
rect 609618 72649 609674 72705
rect 609742 72649 609798 72705
rect 607882 72525 607938 72581
rect 608006 72525 608062 72581
rect 608130 72525 608186 72581
rect 608254 72525 608310 72581
rect 608378 72525 608434 72581
rect 608502 72525 608558 72581
rect 608626 72525 608682 72581
rect 608750 72525 608806 72581
rect 608874 72525 608930 72581
rect 608998 72525 609054 72581
rect 609122 72525 609178 72581
rect 609246 72525 609302 72581
rect 609370 72525 609426 72581
rect 609494 72525 609550 72581
rect 609618 72525 609674 72581
rect 609742 72525 609798 72581
rect 607882 72401 607938 72457
rect 608006 72401 608062 72457
rect 608130 72401 608186 72457
rect 608254 72401 608310 72457
rect 608378 72401 608434 72457
rect 608502 72401 608558 72457
rect 608626 72401 608682 72457
rect 608750 72401 608806 72457
rect 608874 72401 608930 72457
rect 608998 72401 609054 72457
rect 609122 72401 609178 72457
rect 609246 72401 609302 72457
rect 609370 72401 609426 72457
rect 609494 72401 609550 72457
rect 609618 72401 609674 72457
rect 609742 72401 609798 72457
rect 607882 72277 607938 72333
rect 608006 72277 608062 72333
rect 608130 72277 608186 72333
rect 608254 72277 608310 72333
rect 608378 72277 608434 72333
rect 608502 72277 608558 72333
rect 608626 72277 608682 72333
rect 608750 72277 608806 72333
rect 608874 72277 608930 72333
rect 608998 72277 609054 72333
rect 609122 72277 609178 72333
rect 609246 72277 609302 72333
rect 609370 72277 609426 72333
rect 609494 72277 609550 72333
rect 609618 72277 609674 72333
rect 609742 72277 609798 72333
rect 607882 72153 607938 72209
rect 608006 72153 608062 72209
rect 608130 72153 608186 72209
rect 608254 72153 608310 72209
rect 608378 72153 608434 72209
rect 608502 72153 608558 72209
rect 608626 72153 608682 72209
rect 608750 72153 608806 72209
rect 608874 72153 608930 72209
rect 608998 72153 609054 72209
rect 609122 72153 609178 72209
rect 609246 72153 609302 72209
rect 609370 72153 609426 72209
rect 609494 72153 609550 72209
rect 609618 72153 609674 72209
rect 609742 72153 609798 72209
rect 610252 73889 610308 73945
rect 610376 73889 610432 73945
rect 610500 73889 610556 73945
rect 610624 73889 610680 73945
rect 610748 73889 610804 73945
rect 610872 73889 610928 73945
rect 610996 73889 611052 73945
rect 611120 73889 611176 73945
rect 611244 73889 611300 73945
rect 611368 73889 611424 73945
rect 611492 73889 611548 73945
rect 611616 73889 611672 73945
rect 611740 73889 611796 73945
rect 611864 73889 611920 73945
rect 611988 73889 612044 73945
rect 612112 73889 612168 73945
rect 610252 73765 610308 73821
rect 610376 73765 610432 73821
rect 610500 73765 610556 73821
rect 610624 73765 610680 73821
rect 610748 73765 610804 73821
rect 610872 73765 610928 73821
rect 610996 73765 611052 73821
rect 611120 73765 611176 73821
rect 611244 73765 611300 73821
rect 611368 73765 611424 73821
rect 611492 73765 611548 73821
rect 611616 73765 611672 73821
rect 611740 73765 611796 73821
rect 611864 73765 611920 73821
rect 611988 73765 612044 73821
rect 612112 73765 612168 73821
rect 610252 73641 610308 73697
rect 610376 73641 610432 73697
rect 610500 73641 610556 73697
rect 610624 73641 610680 73697
rect 610748 73641 610804 73697
rect 610872 73641 610928 73697
rect 610996 73641 611052 73697
rect 611120 73641 611176 73697
rect 611244 73641 611300 73697
rect 611368 73641 611424 73697
rect 611492 73641 611548 73697
rect 611616 73641 611672 73697
rect 611740 73641 611796 73697
rect 611864 73641 611920 73697
rect 611988 73641 612044 73697
rect 612112 73641 612168 73697
rect 610252 73517 610308 73573
rect 610376 73517 610432 73573
rect 610500 73517 610556 73573
rect 610624 73517 610680 73573
rect 610748 73517 610804 73573
rect 610872 73517 610928 73573
rect 610996 73517 611052 73573
rect 611120 73517 611176 73573
rect 611244 73517 611300 73573
rect 611368 73517 611424 73573
rect 611492 73517 611548 73573
rect 611616 73517 611672 73573
rect 611740 73517 611796 73573
rect 611864 73517 611920 73573
rect 611988 73517 612044 73573
rect 612112 73517 612168 73573
rect 610252 73393 610308 73449
rect 610376 73393 610432 73449
rect 610500 73393 610556 73449
rect 610624 73393 610680 73449
rect 610748 73393 610804 73449
rect 610872 73393 610928 73449
rect 610996 73393 611052 73449
rect 611120 73393 611176 73449
rect 611244 73393 611300 73449
rect 611368 73393 611424 73449
rect 611492 73393 611548 73449
rect 611616 73393 611672 73449
rect 611740 73393 611796 73449
rect 611864 73393 611920 73449
rect 611988 73393 612044 73449
rect 612112 73393 612168 73449
rect 610252 73269 610308 73325
rect 610376 73269 610432 73325
rect 610500 73269 610556 73325
rect 610624 73269 610680 73325
rect 610748 73269 610804 73325
rect 610872 73269 610928 73325
rect 610996 73269 611052 73325
rect 611120 73269 611176 73325
rect 611244 73269 611300 73325
rect 611368 73269 611424 73325
rect 611492 73269 611548 73325
rect 611616 73269 611672 73325
rect 611740 73269 611796 73325
rect 611864 73269 611920 73325
rect 611988 73269 612044 73325
rect 612112 73269 612168 73325
rect 610252 73145 610308 73201
rect 610376 73145 610432 73201
rect 610500 73145 610556 73201
rect 610624 73145 610680 73201
rect 610748 73145 610804 73201
rect 610872 73145 610928 73201
rect 610996 73145 611052 73201
rect 611120 73145 611176 73201
rect 611244 73145 611300 73201
rect 611368 73145 611424 73201
rect 611492 73145 611548 73201
rect 611616 73145 611672 73201
rect 611740 73145 611796 73201
rect 611864 73145 611920 73201
rect 611988 73145 612044 73201
rect 612112 73145 612168 73201
rect 610252 73021 610308 73077
rect 610376 73021 610432 73077
rect 610500 73021 610556 73077
rect 610624 73021 610680 73077
rect 610748 73021 610804 73077
rect 610872 73021 610928 73077
rect 610996 73021 611052 73077
rect 611120 73021 611176 73077
rect 611244 73021 611300 73077
rect 611368 73021 611424 73077
rect 611492 73021 611548 73077
rect 611616 73021 611672 73077
rect 611740 73021 611796 73077
rect 611864 73021 611920 73077
rect 611988 73021 612044 73077
rect 612112 73021 612168 73077
rect 610252 72897 610308 72953
rect 610376 72897 610432 72953
rect 610500 72897 610556 72953
rect 610624 72897 610680 72953
rect 610748 72897 610804 72953
rect 610872 72897 610928 72953
rect 610996 72897 611052 72953
rect 611120 72897 611176 72953
rect 611244 72897 611300 72953
rect 611368 72897 611424 72953
rect 611492 72897 611548 72953
rect 611616 72897 611672 72953
rect 611740 72897 611796 72953
rect 611864 72897 611920 72953
rect 611988 72897 612044 72953
rect 612112 72897 612168 72953
rect 610252 72773 610308 72829
rect 610376 72773 610432 72829
rect 610500 72773 610556 72829
rect 610624 72773 610680 72829
rect 610748 72773 610804 72829
rect 610872 72773 610928 72829
rect 610996 72773 611052 72829
rect 611120 72773 611176 72829
rect 611244 72773 611300 72829
rect 611368 72773 611424 72829
rect 611492 72773 611548 72829
rect 611616 72773 611672 72829
rect 611740 72773 611796 72829
rect 611864 72773 611920 72829
rect 611988 72773 612044 72829
rect 612112 72773 612168 72829
rect 610252 72649 610308 72705
rect 610376 72649 610432 72705
rect 610500 72649 610556 72705
rect 610624 72649 610680 72705
rect 610748 72649 610804 72705
rect 610872 72649 610928 72705
rect 610996 72649 611052 72705
rect 611120 72649 611176 72705
rect 611244 72649 611300 72705
rect 611368 72649 611424 72705
rect 611492 72649 611548 72705
rect 611616 72649 611672 72705
rect 611740 72649 611796 72705
rect 611864 72649 611920 72705
rect 611988 72649 612044 72705
rect 612112 72649 612168 72705
rect 610252 72525 610308 72581
rect 610376 72525 610432 72581
rect 610500 72525 610556 72581
rect 610624 72525 610680 72581
rect 610748 72525 610804 72581
rect 610872 72525 610928 72581
rect 610996 72525 611052 72581
rect 611120 72525 611176 72581
rect 611244 72525 611300 72581
rect 611368 72525 611424 72581
rect 611492 72525 611548 72581
rect 611616 72525 611672 72581
rect 611740 72525 611796 72581
rect 611864 72525 611920 72581
rect 611988 72525 612044 72581
rect 612112 72525 612168 72581
rect 610252 72401 610308 72457
rect 610376 72401 610432 72457
rect 610500 72401 610556 72457
rect 610624 72401 610680 72457
rect 610748 72401 610804 72457
rect 610872 72401 610928 72457
rect 610996 72401 611052 72457
rect 611120 72401 611176 72457
rect 611244 72401 611300 72457
rect 611368 72401 611424 72457
rect 611492 72401 611548 72457
rect 611616 72401 611672 72457
rect 611740 72401 611796 72457
rect 611864 72401 611920 72457
rect 611988 72401 612044 72457
rect 612112 72401 612168 72457
rect 610252 72277 610308 72333
rect 610376 72277 610432 72333
rect 610500 72277 610556 72333
rect 610624 72277 610680 72333
rect 610748 72277 610804 72333
rect 610872 72277 610928 72333
rect 610996 72277 611052 72333
rect 611120 72277 611176 72333
rect 611244 72277 611300 72333
rect 611368 72277 611424 72333
rect 611492 72277 611548 72333
rect 611616 72277 611672 72333
rect 611740 72277 611796 72333
rect 611864 72277 611920 72333
rect 611988 72277 612044 72333
rect 612112 72277 612168 72333
rect 610252 72153 610308 72209
rect 610376 72153 610432 72209
rect 610500 72153 610556 72209
rect 610624 72153 610680 72209
rect 610748 72153 610804 72209
rect 610872 72153 610928 72209
rect 610996 72153 611052 72209
rect 611120 72153 611176 72209
rect 611244 72153 611300 72209
rect 611368 72153 611424 72209
rect 611492 72153 611548 72209
rect 611616 72153 611672 72209
rect 611740 72153 611796 72209
rect 611864 72153 611920 72209
rect 611988 72153 612044 72209
rect 612112 72153 612168 72209
rect 612882 73889 612938 73945
rect 613006 73889 613062 73945
rect 613130 73889 613186 73945
rect 613254 73889 613310 73945
rect 613378 73889 613434 73945
rect 613502 73889 613558 73945
rect 613626 73889 613682 73945
rect 613750 73889 613806 73945
rect 613874 73889 613930 73945
rect 613998 73889 614054 73945
rect 614122 73889 614178 73945
rect 614246 73889 614302 73945
rect 614370 73889 614426 73945
rect 614494 73889 614550 73945
rect 614618 73889 614674 73945
rect 612882 73765 612938 73821
rect 613006 73765 613062 73821
rect 613130 73765 613186 73821
rect 613254 73765 613310 73821
rect 613378 73765 613434 73821
rect 613502 73765 613558 73821
rect 613626 73765 613682 73821
rect 613750 73765 613806 73821
rect 613874 73765 613930 73821
rect 613998 73765 614054 73821
rect 614122 73765 614178 73821
rect 614246 73765 614302 73821
rect 614370 73765 614426 73821
rect 614494 73765 614550 73821
rect 614618 73765 614674 73821
rect 612882 73641 612938 73697
rect 613006 73641 613062 73697
rect 613130 73641 613186 73697
rect 613254 73641 613310 73697
rect 613378 73641 613434 73697
rect 613502 73641 613558 73697
rect 613626 73641 613682 73697
rect 613750 73641 613806 73697
rect 613874 73641 613930 73697
rect 613998 73641 614054 73697
rect 614122 73641 614178 73697
rect 614246 73641 614302 73697
rect 614370 73641 614426 73697
rect 614494 73641 614550 73697
rect 614618 73641 614674 73697
rect 612882 73517 612938 73573
rect 613006 73517 613062 73573
rect 613130 73517 613186 73573
rect 613254 73517 613310 73573
rect 613378 73517 613434 73573
rect 613502 73517 613558 73573
rect 613626 73517 613682 73573
rect 613750 73517 613806 73573
rect 613874 73517 613930 73573
rect 613998 73517 614054 73573
rect 614122 73517 614178 73573
rect 614246 73517 614302 73573
rect 614370 73517 614426 73573
rect 614494 73517 614550 73573
rect 614618 73517 614674 73573
rect 612882 73393 612938 73449
rect 613006 73393 613062 73449
rect 613130 73393 613186 73449
rect 613254 73393 613310 73449
rect 613378 73393 613434 73449
rect 613502 73393 613558 73449
rect 613626 73393 613682 73449
rect 613750 73393 613806 73449
rect 613874 73393 613930 73449
rect 613998 73393 614054 73449
rect 614122 73393 614178 73449
rect 614246 73393 614302 73449
rect 614370 73393 614426 73449
rect 614494 73393 614550 73449
rect 614618 73393 614674 73449
rect 612882 73269 612938 73325
rect 613006 73269 613062 73325
rect 613130 73269 613186 73325
rect 613254 73269 613310 73325
rect 613378 73269 613434 73325
rect 613502 73269 613558 73325
rect 613626 73269 613682 73325
rect 613750 73269 613806 73325
rect 613874 73269 613930 73325
rect 613998 73269 614054 73325
rect 614122 73269 614178 73325
rect 614246 73269 614302 73325
rect 614370 73269 614426 73325
rect 614494 73269 614550 73325
rect 614618 73269 614674 73325
rect 612882 73145 612938 73201
rect 613006 73145 613062 73201
rect 613130 73145 613186 73201
rect 613254 73145 613310 73201
rect 613378 73145 613434 73201
rect 613502 73145 613558 73201
rect 613626 73145 613682 73201
rect 613750 73145 613806 73201
rect 613874 73145 613930 73201
rect 613998 73145 614054 73201
rect 614122 73145 614178 73201
rect 614246 73145 614302 73201
rect 614370 73145 614426 73201
rect 614494 73145 614550 73201
rect 614618 73145 614674 73201
rect 612882 73021 612938 73077
rect 613006 73021 613062 73077
rect 613130 73021 613186 73077
rect 613254 73021 613310 73077
rect 613378 73021 613434 73077
rect 613502 73021 613558 73077
rect 613626 73021 613682 73077
rect 613750 73021 613806 73077
rect 613874 73021 613930 73077
rect 613998 73021 614054 73077
rect 614122 73021 614178 73077
rect 614246 73021 614302 73077
rect 614370 73021 614426 73077
rect 614494 73021 614550 73077
rect 614618 73021 614674 73077
rect 612882 72897 612938 72953
rect 613006 72897 613062 72953
rect 613130 72897 613186 72953
rect 613254 72897 613310 72953
rect 613378 72897 613434 72953
rect 613502 72897 613558 72953
rect 613626 72897 613682 72953
rect 613750 72897 613806 72953
rect 613874 72897 613930 72953
rect 613998 72897 614054 72953
rect 614122 72897 614178 72953
rect 614246 72897 614302 72953
rect 614370 72897 614426 72953
rect 614494 72897 614550 72953
rect 614618 72897 614674 72953
rect 612882 72773 612938 72829
rect 613006 72773 613062 72829
rect 613130 72773 613186 72829
rect 613254 72773 613310 72829
rect 613378 72773 613434 72829
rect 613502 72773 613558 72829
rect 613626 72773 613682 72829
rect 613750 72773 613806 72829
rect 613874 72773 613930 72829
rect 613998 72773 614054 72829
rect 614122 72773 614178 72829
rect 614246 72773 614302 72829
rect 614370 72773 614426 72829
rect 614494 72773 614550 72829
rect 614618 72773 614674 72829
rect 612882 72649 612938 72705
rect 613006 72649 613062 72705
rect 613130 72649 613186 72705
rect 613254 72649 613310 72705
rect 613378 72649 613434 72705
rect 613502 72649 613558 72705
rect 613626 72649 613682 72705
rect 613750 72649 613806 72705
rect 613874 72649 613930 72705
rect 613998 72649 614054 72705
rect 614122 72649 614178 72705
rect 614246 72649 614302 72705
rect 614370 72649 614426 72705
rect 614494 72649 614550 72705
rect 614618 72649 614674 72705
rect 612882 72525 612938 72581
rect 613006 72525 613062 72581
rect 613130 72525 613186 72581
rect 613254 72525 613310 72581
rect 613378 72525 613434 72581
rect 613502 72525 613558 72581
rect 613626 72525 613682 72581
rect 613750 72525 613806 72581
rect 613874 72525 613930 72581
rect 613998 72525 614054 72581
rect 614122 72525 614178 72581
rect 614246 72525 614302 72581
rect 614370 72525 614426 72581
rect 614494 72525 614550 72581
rect 614618 72525 614674 72581
rect 612882 72401 612938 72457
rect 613006 72401 613062 72457
rect 613130 72401 613186 72457
rect 613254 72401 613310 72457
rect 613378 72401 613434 72457
rect 613502 72401 613558 72457
rect 613626 72401 613682 72457
rect 613750 72401 613806 72457
rect 613874 72401 613930 72457
rect 613998 72401 614054 72457
rect 614122 72401 614178 72457
rect 614246 72401 614302 72457
rect 614370 72401 614426 72457
rect 614494 72401 614550 72457
rect 614618 72401 614674 72457
rect 612882 72277 612938 72333
rect 613006 72277 613062 72333
rect 613130 72277 613186 72333
rect 613254 72277 613310 72333
rect 613378 72277 613434 72333
rect 613502 72277 613558 72333
rect 613626 72277 613682 72333
rect 613750 72277 613806 72333
rect 613874 72277 613930 72333
rect 613998 72277 614054 72333
rect 614122 72277 614178 72333
rect 614246 72277 614302 72333
rect 614370 72277 614426 72333
rect 614494 72277 614550 72333
rect 614618 72277 614674 72333
rect 612882 72153 612938 72209
rect 613006 72153 613062 72209
rect 613130 72153 613186 72209
rect 613254 72153 613310 72209
rect 613378 72153 613434 72209
rect 613502 72153 613558 72209
rect 613626 72153 613682 72209
rect 613750 72153 613806 72209
rect 613874 72153 613930 72209
rect 613998 72153 614054 72209
rect 614122 72153 614178 72209
rect 614246 72153 614302 72209
rect 614370 72153 614426 72209
rect 614494 72153 614550 72209
rect 614618 72153 614674 72209
rect 657806 75889 657862 75945
rect 657930 75889 657986 75945
rect 658054 75889 658110 75945
rect 658178 75889 658234 75945
rect 658302 75889 658358 75945
rect 658426 75889 658482 75945
rect 658550 75889 658606 75945
rect 658674 75889 658730 75945
rect 658798 75889 658854 75945
rect 658922 75889 658978 75945
rect 659046 75889 659102 75945
rect 659170 75889 659226 75945
rect 659294 75889 659350 75945
rect 659418 75889 659474 75945
rect 659542 75889 659598 75945
rect 659666 75889 659722 75945
rect 657806 75765 657862 75821
rect 657930 75765 657986 75821
rect 658054 75765 658110 75821
rect 658178 75765 658234 75821
rect 658302 75765 658358 75821
rect 658426 75765 658482 75821
rect 658550 75765 658606 75821
rect 658674 75765 658730 75821
rect 658798 75765 658854 75821
rect 658922 75765 658978 75821
rect 659046 75765 659102 75821
rect 659170 75765 659226 75821
rect 659294 75765 659350 75821
rect 659418 75765 659474 75821
rect 659542 75765 659598 75821
rect 659666 75765 659722 75821
rect 657806 75641 657862 75697
rect 657930 75641 657986 75697
rect 658054 75641 658110 75697
rect 658178 75641 658234 75697
rect 658302 75641 658358 75697
rect 658426 75641 658482 75697
rect 658550 75641 658606 75697
rect 658674 75641 658730 75697
rect 658798 75641 658854 75697
rect 658922 75641 658978 75697
rect 659046 75641 659102 75697
rect 659170 75641 659226 75697
rect 659294 75641 659350 75697
rect 659418 75641 659474 75697
rect 659542 75641 659598 75697
rect 659666 75641 659722 75697
rect 657806 75517 657862 75573
rect 657930 75517 657986 75573
rect 658054 75517 658110 75573
rect 658178 75517 658234 75573
rect 658302 75517 658358 75573
rect 658426 75517 658482 75573
rect 658550 75517 658606 75573
rect 658674 75517 658730 75573
rect 658798 75517 658854 75573
rect 658922 75517 658978 75573
rect 659046 75517 659102 75573
rect 659170 75517 659226 75573
rect 659294 75517 659350 75573
rect 659418 75517 659474 75573
rect 659542 75517 659598 75573
rect 659666 75517 659722 75573
rect 657806 75393 657862 75449
rect 657930 75393 657986 75449
rect 658054 75393 658110 75449
rect 658178 75393 658234 75449
rect 658302 75393 658358 75449
rect 658426 75393 658482 75449
rect 658550 75393 658606 75449
rect 658674 75393 658730 75449
rect 658798 75393 658854 75449
rect 658922 75393 658978 75449
rect 659046 75393 659102 75449
rect 659170 75393 659226 75449
rect 659294 75393 659350 75449
rect 659418 75393 659474 75449
rect 659542 75393 659598 75449
rect 659666 75393 659722 75449
rect 657806 75269 657862 75325
rect 657930 75269 657986 75325
rect 658054 75269 658110 75325
rect 658178 75269 658234 75325
rect 658302 75269 658358 75325
rect 658426 75269 658482 75325
rect 658550 75269 658606 75325
rect 658674 75269 658730 75325
rect 658798 75269 658854 75325
rect 658922 75269 658978 75325
rect 659046 75269 659102 75325
rect 659170 75269 659226 75325
rect 659294 75269 659350 75325
rect 659418 75269 659474 75325
rect 659542 75269 659598 75325
rect 659666 75269 659722 75325
rect 657806 75145 657862 75201
rect 657930 75145 657986 75201
rect 658054 75145 658110 75201
rect 658178 75145 658234 75201
rect 658302 75145 658358 75201
rect 658426 75145 658482 75201
rect 658550 75145 658606 75201
rect 658674 75145 658730 75201
rect 658798 75145 658854 75201
rect 658922 75145 658978 75201
rect 659046 75145 659102 75201
rect 659170 75145 659226 75201
rect 659294 75145 659350 75201
rect 659418 75145 659474 75201
rect 659542 75145 659598 75201
rect 659666 75145 659722 75201
rect 657806 75021 657862 75077
rect 657930 75021 657986 75077
rect 658054 75021 658110 75077
rect 658178 75021 658234 75077
rect 658302 75021 658358 75077
rect 658426 75021 658482 75077
rect 658550 75021 658606 75077
rect 658674 75021 658730 75077
rect 658798 75021 658854 75077
rect 658922 75021 658978 75077
rect 659046 75021 659102 75077
rect 659170 75021 659226 75077
rect 659294 75021 659350 75077
rect 659418 75021 659474 75077
rect 659542 75021 659598 75077
rect 659666 75021 659722 75077
rect 657806 74897 657862 74953
rect 657930 74897 657986 74953
rect 658054 74897 658110 74953
rect 658178 74897 658234 74953
rect 658302 74897 658358 74953
rect 658426 74897 658482 74953
rect 658550 74897 658606 74953
rect 658674 74897 658730 74953
rect 658798 74897 658854 74953
rect 658922 74897 658978 74953
rect 659046 74897 659102 74953
rect 659170 74897 659226 74953
rect 659294 74897 659350 74953
rect 659418 74897 659474 74953
rect 659542 74897 659598 74953
rect 659666 74897 659722 74953
rect 657806 74773 657862 74829
rect 657930 74773 657986 74829
rect 658054 74773 658110 74829
rect 658178 74773 658234 74829
rect 658302 74773 658358 74829
rect 658426 74773 658482 74829
rect 658550 74773 658606 74829
rect 658674 74773 658730 74829
rect 658798 74773 658854 74829
rect 658922 74773 658978 74829
rect 659046 74773 659102 74829
rect 659170 74773 659226 74829
rect 659294 74773 659350 74829
rect 659418 74773 659474 74829
rect 659542 74773 659598 74829
rect 659666 74773 659722 74829
rect 657806 74649 657862 74705
rect 657930 74649 657986 74705
rect 658054 74649 658110 74705
rect 658178 74649 658234 74705
rect 658302 74649 658358 74705
rect 658426 74649 658482 74705
rect 658550 74649 658606 74705
rect 658674 74649 658730 74705
rect 658798 74649 658854 74705
rect 658922 74649 658978 74705
rect 659046 74649 659102 74705
rect 659170 74649 659226 74705
rect 659294 74649 659350 74705
rect 659418 74649 659474 74705
rect 659542 74649 659598 74705
rect 659666 74649 659722 74705
rect 657806 74525 657862 74581
rect 657930 74525 657986 74581
rect 658054 74525 658110 74581
rect 658178 74525 658234 74581
rect 658302 74525 658358 74581
rect 658426 74525 658482 74581
rect 658550 74525 658606 74581
rect 658674 74525 658730 74581
rect 658798 74525 658854 74581
rect 658922 74525 658978 74581
rect 659046 74525 659102 74581
rect 659170 74525 659226 74581
rect 659294 74525 659350 74581
rect 659418 74525 659474 74581
rect 659542 74525 659598 74581
rect 659666 74525 659722 74581
rect 660176 75889 660232 75945
rect 660300 75889 660356 75945
rect 660424 75889 660480 75945
rect 660548 75889 660604 75945
rect 660672 75889 660728 75945
rect 660796 75889 660852 75945
rect 660920 75889 660976 75945
rect 661044 75889 661100 75945
rect 661168 75889 661224 75945
rect 661292 75889 661348 75945
rect 661416 75889 661472 75945
rect 661540 75889 661596 75945
rect 661664 75889 661720 75945
rect 661788 75889 661844 75945
rect 661912 75889 661968 75945
rect 662036 75889 662092 75945
rect 660176 75765 660232 75821
rect 660300 75765 660356 75821
rect 660424 75765 660480 75821
rect 660548 75765 660604 75821
rect 660672 75765 660728 75821
rect 660796 75765 660852 75821
rect 660920 75765 660976 75821
rect 661044 75765 661100 75821
rect 661168 75765 661224 75821
rect 661292 75765 661348 75821
rect 661416 75765 661472 75821
rect 661540 75765 661596 75821
rect 661664 75765 661720 75821
rect 661788 75765 661844 75821
rect 661912 75765 661968 75821
rect 662036 75765 662092 75821
rect 660176 75641 660232 75697
rect 660300 75641 660356 75697
rect 660424 75641 660480 75697
rect 660548 75641 660604 75697
rect 660672 75641 660728 75697
rect 660796 75641 660852 75697
rect 660920 75641 660976 75697
rect 661044 75641 661100 75697
rect 661168 75641 661224 75697
rect 661292 75641 661348 75697
rect 661416 75641 661472 75697
rect 661540 75641 661596 75697
rect 661664 75641 661720 75697
rect 661788 75641 661844 75697
rect 661912 75641 661968 75697
rect 662036 75641 662092 75697
rect 660176 75517 660232 75573
rect 660300 75517 660356 75573
rect 660424 75517 660480 75573
rect 660548 75517 660604 75573
rect 660672 75517 660728 75573
rect 660796 75517 660852 75573
rect 660920 75517 660976 75573
rect 661044 75517 661100 75573
rect 661168 75517 661224 75573
rect 661292 75517 661348 75573
rect 661416 75517 661472 75573
rect 661540 75517 661596 75573
rect 661664 75517 661720 75573
rect 661788 75517 661844 75573
rect 661912 75517 661968 75573
rect 662036 75517 662092 75573
rect 660176 75393 660232 75449
rect 660300 75393 660356 75449
rect 660424 75393 660480 75449
rect 660548 75393 660604 75449
rect 660672 75393 660728 75449
rect 660796 75393 660852 75449
rect 660920 75393 660976 75449
rect 661044 75393 661100 75449
rect 661168 75393 661224 75449
rect 661292 75393 661348 75449
rect 661416 75393 661472 75449
rect 661540 75393 661596 75449
rect 661664 75393 661720 75449
rect 661788 75393 661844 75449
rect 661912 75393 661968 75449
rect 662036 75393 662092 75449
rect 660176 75269 660232 75325
rect 660300 75269 660356 75325
rect 660424 75269 660480 75325
rect 660548 75269 660604 75325
rect 660672 75269 660728 75325
rect 660796 75269 660852 75325
rect 660920 75269 660976 75325
rect 661044 75269 661100 75325
rect 661168 75269 661224 75325
rect 661292 75269 661348 75325
rect 661416 75269 661472 75325
rect 661540 75269 661596 75325
rect 661664 75269 661720 75325
rect 661788 75269 661844 75325
rect 661912 75269 661968 75325
rect 662036 75269 662092 75325
rect 660176 75145 660232 75201
rect 660300 75145 660356 75201
rect 660424 75145 660480 75201
rect 660548 75145 660604 75201
rect 660672 75145 660728 75201
rect 660796 75145 660852 75201
rect 660920 75145 660976 75201
rect 661044 75145 661100 75201
rect 661168 75145 661224 75201
rect 661292 75145 661348 75201
rect 661416 75145 661472 75201
rect 661540 75145 661596 75201
rect 661664 75145 661720 75201
rect 661788 75145 661844 75201
rect 661912 75145 661968 75201
rect 662036 75145 662092 75201
rect 660176 75021 660232 75077
rect 660300 75021 660356 75077
rect 660424 75021 660480 75077
rect 660548 75021 660604 75077
rect 660672 75021 660728 75077
rect 660796 75021 660852 75077
rect 660920 75021 660976 75077
rect 661044 75021 661100 75077
rect 661168 75021 661224 75077
rect 661292 75021 661348 75077
rect 661416 75021 661472 75077
rect 661540 75021 661596 75077
rect 661664 75021 661720 75077
rect 661788 75021 661844 75077
rect 661912 75021 661968 75077
rect 662036 75021 662092 75077
rect 660176 74897 660232 74953
rect 660300 74897 660356 74953
rect 660424 74897 660480 74953
rect 660548 74897 660604 74953
rect 660672 74897 660728 74953
rect 660796 74897 660852 74953
rect 660920 74897 660976 74953
rect 661044 74897 661100 74953
rect 661168 74897 661224 74953
rect 661292 74897 661348 74953
rect 661416 74897 661472 74953
rect 661540 74897 661596 74953
rect 661664 74897 661720 74953
rect 661788 74897 661844 74953
rect 661912 74897 661968 74953
rect 662036 74897 662092 74953
rect 660176 74773 660232 74829
rect 660300 74773 660356 74829
rect 660424 74773 660480 74829
rect 660548 74773 660604 74829
rect 660672 74773 660728 74829
rect 660796 74773 660852 74829
rect 660920 74773 660976 74829
rect 661044 74773 661100 74829
rect 661168 74773 661224 74829
rect 661292 74773 661348 74829
rect 661416 74773 661472 74829
rect 661540 74773 661596 74829
rect 661664 74773 661720 74829
rect 661788 74773 661844 74829
rect 661912 74773 661968 74829
rect 662036 74773 662092 74829
rect 660176 74649 660232 74705
rect 660300 74649 660356 74705
rect 660424 74649 660480 74705
rect 660548 74649 660604 74705
rect 660672 74649 660728 74705
rect 660796 74649 660852 74705
rect 660920 74649 660976 74705
rect 661044 74649 661100 74705
rect 661168 74649 661224 74705
rect 661292 74649 661348 74705
rect 661416 74649 661472 74705
rect 661540 74649 661596 74705
rect 661664 74649 661720 74705
rect 661788 74649 661844 74705
rect 661912 74649 661968 74705
rect 662036 74649 662092 74705
rect 660176 74525 660232 74581
rect 660300 74525 660356 74581
rect 660424 74525 660480 74581
rect 660548 74525 660604 74581
rect 660672 74525 660728 74581
rect 660796 74525 660852 74581
rect 660920 74525 660976 74581
rect 661044 74525 661100 74581
rect 661168 74525 661224 74581
rect 661292 74525 661348 74581
rect 661416 74525 661472 74581
rect 661540 74525 661596 74581
rect 661664 74525 661720 74581
rect 661788 74525 661844 74581
rect 661912 74525 661968 74581
rect 662036 74525 662092 74581
rect 662882 75889 662938 75945
rect 663006 75889 663062 75945
rect 663130 75889 663186 75945
rect 663254 75889 663310 75945
rect 663378 75889 663434 75945
rect 663502 75889 663558 75945
rect 663626 75889 663682 75945
rect 663750 75889 663806 75945
rect 663874 75889 663930 75945
rect 663998 75889 664054 75945
rect 664122 75889 664178 75945
rect 664246 75889 664302 75945
rect 664370 75889 664426 75945
rect 664494 75889 664550 75945
rect 664618 75889 664674 75945
rect 664742 75889 664798 75945
rect 662882 75765 662938 75821
rect 663006 75765 663062 75821
rect 663130 75765 663186 75821
rect 663254 75765 663310 75821
rect 663378 75765 663434 75821
rect 663502 75765 663558 75821
rect 663626 75765 663682 75821
rect 663750 75765 663806 75821
rect 663874 75765 663930 75821
rect 663998 75765 664054 75821
rect 664122 75765 664178 75821
rect 664246 75765 664302 75821
rect 664370 75765 664426 75821
rect 664494 75765 664550 75821
rect 664618 75765 664674 75821
rect 664742 75765 664798 75821
rect 662882 75641 662938 75697
rect 663006 75641 663062 75697
rect 663130 75641 663186 75697
rect 663254 75641 663310 75697
rect 663378 75641 663434 75697
rect 663502 75641 663558 75697
rect 663626 75641 663682 75697
rect 663750 75641 663806 75697
rect 663874 75641 663930 75697
rect 663998 75641 664054 75697
rect 664122 75641 664178 75697
rect 664246 75641 664302 75697
rect 664370 75641 664426 75697
rect 664494 75641 664550 75697
rect 664618 75641 664674 75697
rect 664742 75641 664798 75697
rect 662882 75517 662938 75573
rect 663006 75517 663062 75573
rect 663130 75517 663186 75573
rect 663254 75517 663310 75573
rect 663378 75517 663434 75573
rect 663502 75517 663558 75573
rect 663626 75517 663682 75573
rect 663750 75517 663806 75573
rect 663874 75517 663930 75573
rect 663998 75517 664054 75573
rect 664122 75517 664178 75573
rect 664246 75517 664302 75573
rect 664370 75517 664426 75573
rect 664494 75517 664550 75573
rect 664618 75517 664674 75573
rect 664742 75517 664798 75573
rect 662882 75393 662938 75449
rect 663006 75393 663062 75449
rect 663130 75393 663186 75449
rect 663254 75393 663310 75449
rect 663378 75393 663434 75449
rect 663502 75393 663558 75449
rect 663626 75393 663682 75449
rect 663750 75393 663806 75449
rect 663874 75393 663930 75449
rect 663998 75393 664054 75449
rect 664122 75393 664178 75449
rect 664246 75393 664302 75449
rect 664370 75393 664426 75449
rect 664494 75393 664550 75449
rect 664618 75393 664674 75449
rect 664742 75393 664798 75449
rect 662882 75269 662938 75325
rect 663006 75269 663062 75325
rect 663130 75269 663186 75325
rect 663254 75269 663310 75325
rect 663378 75269 663434 75325
rect 663502 75269 663558 75325
rect 663626 75269 663682 75325
rect 663750 75269 663806 75325
rect 663874 75269 663930 75325
rect 663998 75269 664054 75325
rect 664122 75269 664178 75325
rect 664246 75269 664302 75325
rect 664370 75269 664426 75325
rect 664494 75269 664550 75325
rect 664618 75269 664674 75325
rect 664742 75269 664798 75325
rect 662882 75145 662938 75201
rect 663006 75145 663062 75201
rect 663130 75145 663186 75201
rect 663254 75145 663310 75201
rect 663378 75145 663434 75201
rect 663502 75145 663558 75201
rect 663626 75145 663682 75201
rect 663750 75145 663806 75201
rect 663874 75145 663930 75201
rect 663998 75145 664054 75201
rect 664122 75145 664178 75201
rect 664246 75145 664302 75201
rect 664370 75145 664426 75201
rect 664494 75145 664550 75201
rect 664618 75145 664674 75201
rect 664742 75145 664798 75201
rect 662882 75021 662938 75077
rect 663006 75021 663062 75077
rect 663130 75021 663186 75077
rect 663254 75021 663310 75077
rect 663378 75021 663434 75077
rect 663502 75021 663558 75077
rect 663626 75021 663682 75077
rect 663750 75021 663806 75077
rect 663874 75021 663930 75077
rect 663998 75021 664054 75077
rect 664122 75021 664178 75077
rect 664246 75021 664302 75077
rect 664370 75021 664426 75077
rect 664494 75021 664550 75077
rect 664618 75021 664674 75077
rect 664742 75021 664798 75077
rect 662882 74897 662938 74953
rect 663006 74897 663062 74953
rect 663130 74897 663186 74953
rect 663254 74897 663310 74953
rect 663378 74897 663434 74953
rect 663502 74897 663558 74953
rect 663626 74897 663682 74953
rect 663750 74897 663806 74953
rect 663874 74897 663930 74953
rect 663998 74897 664054 74953
rect 664122 74897 664178 74953
rect 664246 74897 664302 74953
rect 664370 74897 664426 74953
rect 664494 74897 664550 74953
rect 664618 74897 664674 74953
rect 664742 74897 664798 74953
rect 662882 74773 662938 74829
rect 663006 74773 663062 74829
rect 663130 74773 663186 74829
rect 663254 74773 663310 74829
rect 663378 74773 663434 74829
rect 663502 74773 663558 74829
rect 663626 74773 663682 74829
rect 663750 74773 663806 74829
rect 663874 74773 663930 74829
rect 663998 74773 664054 74829
rect 664122 74773 664178 74829
rect 664246 74773 664302 74829
rect 664370 74773 664426 74829
rect 664494 74773 664550 74829
rect 664618 74773 664674 74829
rect 664742 74773 664798 74829
rect 662882 74649 662938 74705
rect 663006 74649 663062 74705
rect 663130 74649 663186 74705
rect 663254 74649 663310 74705
rect 663378 74649 663434 74705
rect 663502 74649 663558 74705
rect 663626 74649 663682 74705
rect 663750 74649 663806 74705
rect 663874 74649 663930 74705
rect 663998 74649 664054 74705
rect 664122 74649 664178 74705
rect 664246 74649 664302 74705
rect 664370 74649 664426 74705
rect 664494 74649 664550 74705
rect 664618 74649 664674 74705
rect 664742 74649 664798 74705
rect 662882 74525 662938 74581
rect 663006 74525 663062 74581
rect 663130 74525 663186 74581
rect 663254 74525 663310 74581
rect 663378 74525 663434 74581
rect 663502 74525 663558 74581
rect 663626 74525 663682 74581
rect 663750 74525 663806 74581
rect 663874 74525 663930 74581
rect 663998 74525 664054 74581
rect 664122 74525 664178 74581
rect 664246 74525 664302 74581
rect 664370 74525 664426 74581
rect 664494 74525 664550 74581
rect 664618 74525 664674 74581
rect 664742 74525 664798 74581
rect 665252 75889 665308 75945
rect 665376 75889 665432 75945
rect 665500 75889 665556 75945
rect 665624 75889 665680 75945
rect 665748 75889 665804 75945
rect 665872 75889 665928 75945
rect 665996 75889 666052 75945
rect 666120 75889 666176 75945
rect 666244 75889 666300 75945
rect 666368 75889 666424 75945
rect 666492 75889 666548 75945
rect 666616 75889 666672 75945
rect 666740 75889 666796 75945
rect 666864 75889 666920 75945
rect 666988 75889 667044 75945
rect 667112 75889 667168 75945
rect 665252 75765 665308 75821
rect 665376 75765 665432 75821
rect 665500 75765 665556 75821
rect 665624 75765 665680 75821
rect 665748 75765 665804 75821
rect 665872 75765 665928 75821
rect 665996 75765 666052 75821
rect 666120 75765 666176 75821
rect 666244 75765 666300 75821
rect 666368 75765 666424 75821
rect 666492 75765 666548 75821
rect 666616 75765 666672 75821
rect 666740 75765 666796 75821
rect 666864 75765 666920 75821
rect 666988 75765 667044 75821
rect 667112 75765 667168 75821
rect 665252 75641 665308 75697
rect 665376 75641 665432 75697
rect 665500 75641 665556 75697
rect 665624 75641 665680 75697
rect 665748 75641 665804 75697
rect 665872 75641 665928 75697
rect 665996 75641 666052 75697
rect 666120 75641 666176 75697
rect 666244 75641 666300 75697
rect 666368 75641 666424 75697
rect 666492 75641 666548 75697
rect 666616 75641 666672 75697
rect 666740 75641 666796 75697
rect 666864 75641 666920 75697
rect 666988 75641 667044 75697
rect 667112 75641 667168 75697
rect 665252 75517 665308 75573
rect 665376 75517 665432 75573
rect 665500 75517 665556 75573
rect 665624 75517 665680 75573
rect 665748 75517 665804 75573
rect 665872 75517 665928 75573
rect 665996 75517 666052 75573
rect 666120 75517 666176 75573
rect 666244 75517 666300 75573
rect 666368 75517 666424 75573
rect 666492 75517 666548 75573
rect 666616 75517 666672 75573
rect 666740 75517 666796 75573
rect 666864 75517 666920 75573
rect 666988 75517 667044 75573
rect 667112 75517 667168 75573
rect 665252 75393 665308 75449
rect 665376 75393 665432 75449
rect 665500 75393 665556 75449
rect 665624 75393 665680 75449
rect 665748 75393 665804 75449
rect 665872 75393 665928 75449
rect 665996 75393 666052 75449
rect 666120 75393 666176 75449
rect 666244 75393 666300 75449
rect 666368 75393 666424 75449
rect 666492 75393 666548 75449
rect 666616 75393 666672 75449
rect 666740 75393 666796 75449
rect 666864 75393 666920 75449
rect 666988 75393 667044 75449
rect 667112 75393 667168 75449
rect 665252 75269 665308 75325
rect 665376 75269 665432 75325
rect 665500 75269 665556 75325
rect 665624 75269 665680 75325
rect 665748 75269 665804 75325
rect 665872 75269 665928 75325
rect 665996 75269 666052 75325
rect 666120 75269 666176 75325
rect 666244 75269 666300 75325
rect 666368 75269 666424 75325
rect 666492 75269 666548 75325
rect 666616 75269 666672 75325
rect 666740 75269 666796 75325
rect 666864 75269 666920 75325
rect 666988 75269 667044 75325
rect 667112 75269 667168 75325
rect 665252 75145 665308 75201
rect 665376 75145 665432 75201
rect 665500 75145 665556 75201
rect 665624 75145 665680 75201
rect 665748 75145 665804 75201
rect 665872 75145 665928 75201
rect 665996 75145 666052 75201
rect 666120 75145 666176 75201
rect 666244 75145 666300 75201
rect 666368 75145 666424 75201
rect 666492 75145 666548 75201
rect 666616 75145 666672 75201
rect 666740 75145 666796 75201
rect 666864 75145 666920 75201
rect 666988 75145 667044 75201
rect 667112 75145 667168 75201
rect 665252 75021 665308 75077
rect 665376 75021 665432 75077
rect 665500 75021 665556 75077
rect 665624 75021 665680 75077
rect 665748 75021 665804 75077
rect 665872 75021 665928 75077
rect 665996 75021 666052 75077
rect 666120 75021 666176 75077
rect 666244 75021 666300 75077
rect 666368 75021 666424 75077
rect 666492 75021 666548 75077
rect 666616 75021 666672 75077
rect 666740 75021 666796 75077
rect 666864 75021 666920 75077
rect 666988 75021 667044 75077
rect 667112 75021 667168 75077
rect 665252 74897 665308 74953
rect 665376 74897 665432 74953
rect 665500 74897 665556 74953
rect 665624 74897 665680 74953
rect 665748 74897 665804 74953
rect 665872 74897 665928 74953
rect 665996 74897 666052 74953
rect 666120 74897 666176 74953
rect 666244 74897 666300 74953
rect 666368 74897 666424 74953
rect 666492 74897 666548 74953
rect 666616 74897 666672 74953
rect 666740 74897 666796 74953
rect 666864 74897 666920 74953
rect 666988 74897 667044 74953
rect 667112 74897 667168 74953
rect 665252 74773 665308 74829
rect 665376 74773 665432 74829
rect 665500 74773 665556 74829
rect 665624 74773 665680 74829
rect 665748 74773 665804 74829
rect 665872 74773 665928 74829
rect 665996 74773 666052 74829
rect 666120 74773 666176 74829
rect 666244 74773 666300 74829
rect 666368 74773 666424 74829
rect 666492 74773 666548 74829
rect 666616 74773 666672 74829
rect 666740 74773 666796 74829
rect 666864 74773 666920 74829
rect 666988 74773 667044 74829
rect 667112 74773 667168 74829
rect 665252 74649 665308 74705
rect 665376 74649 665432 74705
rect 665500 74649 665556 74705
rect 665624 74649 665680 74705
rect 665748 74649 665804 74705
rect 665872 74649 665928 74705
rect 665996 74649 666052 74705
rect 666120 74649 666176 74705
rect 666244 74649 666300 74705
rect 666368 74649 666424 74705
rect 666492 74649 666548 74705
rect 666616 74649 666672 74705
rect 666740 74649 666796 74705
rect 666864 74649 666920 74705
rect 666988 74649 667044 74705
rect 667112 74649 667168 74705
rect 665252 74525 665308 74581
rect 665376 74525 665432 74581
rect 665500 74525 665556 74581
rect 665624 74525 665680 74581
rect 665748 74525 665804 74581
rect 665872 74525 665928 74581
rect 665996 74525 666052 74581
rect 666120 74525 666176 74581
rect 666244 74525 666300 74581
rect 666368 74525 666424 74581
rect 666492 74525 666548 74581
rect 666616 74525 666672 74581
rect 666740 74525 666796 74581
rect 666864 74525 666920 74581
rect 666988 74525 667044 74581
rect 667112 74525 667168 74581
rect 667882 75889 667938 75945
rect 668006 75889 668062 75945
rect 668130 75889 668186 75945
rect 668254 75889 668310 75945
rect 668378 75889 668434 75945
rect 668502 75889 668558 75945
rect 668626 75889 668682 75945
rect 668750 75889 668806 75945
rect 668874 75889 668930 75945
rect 668998 75889 669054 75945
rect 669122 75889 669178 75945
rect 669246 75889 669302 75945
rect 669370 75889 669426 75945
rect 669494 75889 669550 75945
rect 669618 75889 669674 75945
rect 667882 75765 667938 75821
rect 668006 75765 668062 75821
rect 668130 75765 668186 75821
rect 668254 75765 668310 75821
rect 668378 75765 668434 75821
rect 668502 75765 668558 75821
rect 668626 75765 668682 75821
rect 668750 75765 668806 75821
rect 668874 75765 668930 75821
rect 668998 75765 669054 75821
rect 669122 75765 669178 75821
rect 669246 75765 669302 75821
rect 669370 75765 669426 75821
rect 669494 75765 669550 75821
rect 669618 75765 669674 75821
rect 667882 75641 667938 75697
rect 668006 75641 668062 75697
rect 668130 75641 668186 75697
rect 668254 75641 668310 75697
rect 668378 75641 668434 75697
rect 668502 75641 668558 75697
rect 668626 75641 668682 75697
rect 668750 75641 668806 75697
rect 668874 75641 668930 75697
rect 668998 75641 669054 75697
rect 669122 75641 669178 75697
rect 669246 75641 669302 75697
rect 669370 75641 669426 75697
rect 669494 75641 669550 75697
rect 669618 75641 669674 75697
rect 667882 75517 667938 75573
rect 668006 75517 668062 75573
rect 668130 75517 668186 75573
rect 668254 75517 668310 75573
rect 668378 75517 668434 75573
rect 668502 75517 668558 75573
rect 668626 75517 668682 75573
rect 668750 75517 668806 75573
rect 668874 75517 668930 75573
rect 668998 75517 669054 75573
rect 669122 75517 669178 75573
rect 669246 75517 669302 75573
rect 669370 75517 669426 75573
rect 669494 75517 669550 75573
rect 669618 75517 669674 75573
rect 667882 75393 667938 75449
rect 668006 75393 668062 75449
rect 668130 75393 668186 75449
rect 668254 75393 668310 75449
rect 668378 75393 668434 75449
rect 668502 75393 668558 75449
rect 668626 75393 668682 75449
rect 668750 75393 668806 75449
rect 668874 75393 668930 75449
rect 668998 75393 669054 75449
rect 669122 75393 669178 75449
rect 669246 75393 669302 75449
rect 669370 75393 669426 75449
rect 669494 75393 669550 75449
rect 669618 75393 669674 75449
rect 667882 75269 667938 75325
rect 668006 75269 668062 75325
rect 668130 75269 668186 75325
rect 668254 75269 668310 75325
rect 668378 75269 668434 75325
rect 668502 75269 668558 75325
rect 668626 75269 668682 75325
rect 668750 75269 668806 75325
rect 668874 75269 668930 75325
rect 668998 75269 669054 75325
rect 669122 75269 669178 75325
rect 669246 75269 669302 75325
rect 669370 75269 669426 75325
rect 669494 75269 669550 75325
rect 669618 75269 669674 75325
rect 667882 75145 667938 75201
rect 668006 75145 668062 75201
rect 668130 75145 668186 75201
rect 668254 75145 668310 75201
rect 668378 75145 668434 75201
rect 668502 75145 668558 75201
rect 668626 75145 668682 75201
rect 668750 75145 668806 75201
rect 668874 75145 668930 75201
rect 668998 75145 669054 75201
rect 669122 75145 669178 75201
rect 669246 75145 669302 75201
rect 669370 75145 669426 75201
rect 669494 75145 669550 75201
rect 669618 75145 669674 75201
rect 667882 75021 667938 75077
rect 668006 75021 668062 75077
rect 668130 75021 668186 75077
rect 668254 75021 668310 75077
rect 668378 75021 668434 75077
rect 668502 75021 668558 75077
rect 668626 75021 668682 75077
rect 668750 75021 668806 75077
rect 668874 75021 668930 75077
rect 668998 75021 669054 75077
rect 669122 75021 669178 75077
rect 669246 75021 669302 75077
rect 669370 75021 669426 75077
rect 669494 75021 669550 75077
rect 669618 75021 669674 75077
rect 667882 74897 667938 74953
rect 668006 74897 668062 74953
rect 668130 74897 668186 74953
rect 668254 74897 668310 74953
rect 668378 74897 668434 74953
rect 668502 74897 668558 74953
rect 668626 74897 668682 74953
rect 668750 74897 668806 74953
rect 668874 74897 668930 74953
rect 668998 74897 669054 74953
rect 669122 74897 669178 74953
rect 669246 74897 669302 74953
rect 669370 74897 669426 74953
rect 669494 74897 669550 74953
rect 669618 74897 669674 74953
rect 667882 74773 667938 74829
rect 668006 74773 668062 74829
rect 668130 74773 668186 74829
rect 668254 74773 668310 74829
rect 668378 74773 668434 74829
rect 668502 74773 668558 74829
rect 668626 74773 668682 74829
rect 668750 74773 668806 74829
rect 668874 74773 668930 74829
rect 668998 74773 669054 74829
rect 669122 74773 669178 74829
rect 669246 74773 669302 74829
rect 669370 74773 669426 74829
rect 669494 74773 669550 74829
rect 669618 74773 669674 74829
rect 667882 74649 667938 74705
rect 668006 74649 668062 74705
rect 668130 74649 668186 74705
rect 668254 74649 668310 74705
rect 668378 74649 668434 74705
rect 668502 74649 668558 74705
rect 668626 74649 668682 74705
rect 668750 74649 668806 74705
rect 668874 74649 668930 74705
rect 668998 74649 669054 74705
rect 669122 74649 669178 74705
rect 669246 74649 669302 74705
rect 669370 74649 669426 74705
rect 669494 74649 669550 74705
rect 669618 74649 669674 74705
rect 667882 74525 667938 74581
rect 668006 74525 668062 74581
rect 668130 74525 668186 74581
rect 668254 74525 668310 74581
rect 668378 74525 668434 74581
rect 668502 74525 668558 74581
rect 668626 74525 668682 74581
rect 668750 74525 668806 74581
rect 668874 74525 668930 74581
rect 668998 74525 669054 74581
rect 669122 74525 669178 74581
rect 669246 74525 669302 74581
rect 669370 74525 669426 74581
rect 669494 74525 669550 74581
rect 669618 74525 669674 74581
<< metal3 >>
rect 379272 941675 381172 941720
rect 379272 941655 379341 941675
rect 379397 941655 379483 941675
rect 379539 941655 379625 941675
rect 379681 941655 379767 941675
rect 379823 941655 379909 941675
rect 379965 941655 381172 941675
rect 379272 941599 379326 941655
rect 379397 941619 379450 941655
rect 379539 941619 379574 941655
rect 379681 941619 379698 941655
rect 379382 941599 379450 941619
rect 379506 941599 379574 941619
rect 379630 941599 379698 941619
rect 379754 941619 379767 941655
rect 379878 941619 379909 941655
rect 379754 941599 379822 941619
rect 379878 941599 379946 941619
rect 380002 941599 381172 941655
rect 379272 941533 381172 941599
rect 379272 941531 379341 941533
rect 379397 941531 379483 941533
rect 379539 941531 379625 941533
rect 379681 941531 379767 941533
rect 379823 941531 379909 941533
rect 379965 941531 381172 941533
rect 379272 941475 379326 941531
rect 379397 941477 379450 941531
rect 379539 941477 379574 941531
rect 379681 941477 379698 941531
rect 379382 941475 379450 941477
rect 379506 941475 379574 941477
rect 379630 941475 379698 941477
rect 379754 941477 379767 941531
rect 379878 941477 379909 941531
rect 379754 941475 379822 941477
rect 379878 941475 379946 941477
rect 380002 941475 381172 941531
rect 379272 941407 381172 941475
rect 379272 941351 379326 941407
rect 379382 941391 379450 941407
rect 379506 941391 379574 941407
rect 379630 941391 379698 941407
rect 379397 941351 379450 941391
rect 379539 941351 379574 941391
rect 379681 941351 379698 941391
rect 379754 941391 379822 941407
rect 379878 941391 379946 941407
rect 379754 941351 379767 941391
rect 379878 941351 379909 941391
rect 380002 941351 381172 941407
rect 379272 941335 379341 941351
rect 379397 941335 379483 941351
rect 379539 941335 379625 941351
rect 379681 941335 379767 941351
rect 379823 941335 379909 941351
rect 379965 941335 381172 941351
rect 379272 941283 381172 941335
rect 379272 941227 379326 941283
rect 379382 941249 379450 941283
rect 379506 941249 379574 941283
rect 379630 941249 379698 941283
rect 379397 941227 379450 941249
rect 379539 941227 379574 941249
rect 379681 941227 379698 941249
rect 379754 941249 379822 941283
rect 379878 941249 379946 941283
rect 379754 941227 379767 941249
rect 379878 941227 379909 941249
rect 380002 941227 381172 941283
rect 379272 941193 379341 941227
rect 379397 941193 379483 941227
rect 379539 941193 379625 941227
rect 379681 941193 379767 941227
rect 379823 941193 379909 941227
rect 379965 941193 381172 941227
rect 379272 941159 381172 941193
rect 379272 941103 379326 941159
rect 379382 941107 379450 941159
rect 379506 941107 379574 941159
rect 379630 941107 379698 941159
rect 379397 941103 379450 941107
rect 379539 941103 379574 941107
rect 379681 941103 379698 941107
rect 379754 941107 379822 941159
rect 379878 941107 379946 941159
rect 379754 941103 379767 941107
rect 379878 941103 379909 941107
rect 380002 941103 381172 941159
rect 379272 941051 379341 941103
rect 379397 941051 379483 941103
rect 379539 941051 379625 941103
rect 379681 941051 379767 941103
rect 379823 941051 379909 941103
rect 379965 941051 381172 941103
rect 379272 941035 381172 941051
rect 379272 940979 379326 941035
rect 379382 940979 379450 941035
rect 379506 940979 379574 941035
rect 379630 940979 379698 941035
rect 379754 940979 379822 941035
rect 379878 940979 379946 941035
rect 380002 940979 381172 941035
rect 379272 940965 381172 940979
rect 379272 940911 379341 940965
rect 379397 940911 379483 940965
rect 379539 940911 379625 940965
rect 379681 940911 379767 940965
rect 379823 940911 379909 940965
rect 379965 940911 381172 940965
rect 379272 940855 379326 940911
rect 379397 940909 379450 940911
rect 379539 940909 379574 940911
rect 379681 940909 379698 940911
rect 379382 940855 379450 940909
rect 379506 940855 379574 940909
rect 379630 940855 379698 940909
rect 379754 940909 379767 940911
rect 379878 940909 379909 940911
rect 379754 940855 379822 940909
rect 379878 940855 379946 940909
rect 380002 940855 381172 940911
rect 379272 940823 381172 940855
rect 379272 940787 379341 940823
rect 379397 940787 379483 940823
rect 379539 940787 379625 940823
rect 379681 940787 379767 940823
rect 379823 940787 379909 940823
rect 379965 940787 381172 940823
rect 379272 940731 379326 940787
rect 379397 940767 379450 940787
rect 379539 940767 379574 940787
rect 379681 940767 379698 940787
rect 379382 940731 379450 940767
rect 379506 940731 379574 940767
rect 379630 940731 379698 940767
rect 379754 940767 379767 940787
rect 379878 940767 379909 940787
rect 379754 940731 379822 940767
rect 379878 940731 379946 940767
rect 380002 940731 381172 940787
rect 379272 940681 381172 940731
rect 379272 940663 379341 940681
rect 379397 940663 379483 940681
rect 379539 940663 379625 940681
rect 379681 940663 379767 940681
rect 379823 940663 379909 940681
rect 379965 940663 381172 940681
rect 379272 940607 379326 940663
rect 379397 940625 379450 940663
rect 379539 940625 379574 940663
rect 379681 940625 379698 940663
rect 379382 940607 379450 940625
rect 379506 940607 379574 940625
rect 379630 940607 379698 940625
rect 379754 940625 379767 940663
rect 379878 940625 379909 940663
rect 379754 940607 379822 940625
rect 379878 940607 379946 940625
rect 380002 940607 381172 940663
rect 379272 940539 381172 940607
rect 379272 940483 379326 940539
rect 379397 940483 379450 940539
rect 379539 940483 379574 940539
rect 379681 940483 379698 940539
rect 379754 940483 379767 940539
rect 379878 940483 379909 940539
rect 380002 940483 381172 940539
rect 379272 940415 381172 940483
rect 379272 940359 379326 940415
rect 379382 940397 379450 940415
rect 379506 940397 379574 940415
rect 379630 940397 379698 940415
rect 379397 940359 379450 940397
rect 379539 940359 379574 940397
rect 379681 940359 379698 940397
rect 379754 940397 379822 940415
rect 379878 940397 379946 940415
rect 379754 940359 379767 940397
rect 379878 940359 379909 940397
rect 380002 940359 381172 940415
rect 379272 940341 379341 940359
rect 379397 940341 379483 940359
rect 379539 940341 379625 940359
rect 379681 940341 379767 940359
rect 379823 940341 379909 940359
rect 379965 940341 381172 940359
rect 379272 940291 381172 940341
rect 379272 940235 379326 940291
rect 379382 940255 379450 940291
rect 379506 940255 379574 940291
rect 379630 940255 379698 940291
rect 379397 940235 379450 940255
rect 379539 940235 379574 940255
rect 379681 940235 379698 940255
rect 379754 940255 379822 940291
rect 379878 940255 379946 940291
rect 379754 940235 379767 940255
rect 379878 940235 379909 940255
rect 380002 940235 381172 940291
rect 379272 940199 379341 940235
rect 379397 940199 379483 940235
rect 379539 940199 379625 940235
rect 379681 940199 379767 940235
rect 379823 940199 379909 940235
rect 379965 940199 381172 940235
rect 379272 940167 381172 940199
rect 379272 940111 379326 940167
rect 379382 940113 379450 940167
rect 379506 940113 379574 940167
rect 379630 940113 379698 940167
rect 379397 940111 379450 940113
rect 379539 940111 379574 940113
rect 379681 940111 379698 940113
rect 379754 940113 379822 940167
rect 379878 940113 379946 940167
rect 379754 940111 379767 940113
rect 379878 940111 379909 940113
rect 380002 940111 381172 940167
rect 379272 940057 379341 940111
rect 379397 940057 379483 940111
rect 379539 940057 379625 940111
rect 379681 940057 379767 940111
rect 379823 940057 379909 940111
rect 379965 940057 381172 940111
rect 379272 940043 381172 940057
rect 379272 939987 379326 940043
rect 379382 939987 379450 940043
rect 379506 939987 379574 940043
rect 379630 939987 379698 940043
rect 379754 939987 379822 940043
rect 379878 939987 379946 940043
rect 380002 939987 381172 940043
rect 379272 939971 381172 939987
rect 379272 939919 379341 939971
rect 379397 939919 379483 939971
rect 379539 939919 379625 939971
rect 379681 939919 379767 939971
rect 379823 939919 379909 939971
rect 379965 939919 381172 939971
rect 379272 939863 379326 939919
rect 379397 939915 379450 939919
rect 379539 939915 379574 939919
rect 379681 939915 379698 939919
rect 379382 939863 379450 939915
rect 379506 939863 379574 939915
rect 379630 939863 379698 939915
rect 379754 939915 379767 939919
rect 379878 939915 379909 939919
rect 379754 939863 379822 939915
rect 379878 939863 379946 939915
rect 380002 939863 381172 939919
rect 379272 939829 381172 939863
rect 379272 939773 379341 939829
rect 379397 939773 379483 939829
rect 379539 939773 379625 939829
rect 379681 939773 379767 939829
rect 379823 939773 379909 939829
rect 379965 939773 381172 939829
rect 379272 939720 381172 939773
rect 381752 941675 383802 941720
rect 381752 941619 381829 941675
rect 381885 941655 381971 941675
rect 382027 941655 382113 941675
rect 382169 941655 382255 941675
rect 382311 941655 382397 941675
rect 382453 941655 382539 941675
rect 382595 941655 382681 941675
rect 382737 941655 382823 941675
rect 382879 941655 382965 941675
rect 383021 941655 383107 941675
rect 383163 941655 383249 941675
rect 383305 941655 383391 941675
rect 383447 941655 383533 941675
rect 383589 941655 383675 941675
rect 383731 941655 383802 941675
rect 381752 941599 381832 941619
rect 381888 941599 381956 941655
rect 382027 941619 382080 941655
rect 382169 941619 382204 941655
rect 382311 941619 382328 941655
rect 382012 941599 382080 941619
rect 382136 941599 382204 941619
rect 382260 941599 382328 941619
rect 382384 941619 382397 941655
rect 382508 941619 382539 941655
rect 382632 941619 382681 941655
rect 382756 941619 382823 941655
rect 382384 941599 382452 941619
rect 382508 941599 382576 941619
rect 382632 941599 382700 941619
rect 382756 941599 382824 941619
rect 382880 941599 382948 941655
rect 383021 941619 383072 941655
rect 383163 941619 383196 941655
rect 383305 941619 383320 941655
rect 383004 941599 383072 941619
rect 383128 941599 383196 941619
rect 383252 941599 383320 941619
rect 383376 941619 383391 941655
rect 383500 941619 383533 941655
rect 383624 941619 383675 941655
rect 383376 941599 383444 941619
rect 383500 941599 383568 941619
rect 383624 941599 383692 941619
rect 383748 941599 383802 941655
rect 381752 941533 383802 941599
rect 381752 941477 381829 941533
rect 381885 941531 381971 941533
rect 382027 941531 382113 941533
rect 382169 941531 382255 941533
rect 382311 941531 382397 941533
rect 382453 941531 382539 941533
rect 382595 941531 382681 941533
rect 382737 941531 382823 941533
rect 382879 941531 382965 941533
rect 383021 941531 383107 941533
rect 383163 941531 383249 941533
rect 383305 941531 383391 941533
rect 383447 941531 383533 941533
rect 383589 941531 383675 941533
rect 383731 941531 383802 941533
rect 381752 941475 381832 941477
rect 381888 941475 381956 941531
rect 382027 941477 382080 941531
rect 382169 941477 382204 941531
rect 382311 941477 382328 941531
rect 382012 941475 382080 941477
rect 382136 941475 382204 941477
rect 382260 941475 382328 941477
rect 382384 941477 382397 941531
rect 382508 941477 382539 941531
rect 382632 941477 382681 941531
rect 382756 941477 382823 941531
rect 382384 941475 382452 941477
rect 382508 941475 382576 941477
rect 382632 941475 382700 941477
rect 382756 941475 382824 941477
rect 382880 941475 382948 941531
rect 383021 941477 383072 941531
rect 383163 941477 383196 941531
rect 383305 941477 383320 941531
rect 383004 941475 383072 941477
rect 383128 941475 383196 941477
rect 383252 941475 383320 941477
rect 383376 941477 383391 941531
rect 383500 941477 383533 941531
rect 383624 941477 383675 941531
rect 383376 941475 383444 941477
rect 383500 941475 383568 941477
rect 383624 941475 383692 941477
rect 383748 941475 383802 941531
rect 381752 941407 383802 941475
rect 381752 941391 381832 941407
rect 381752 941335 381829 941391
rect 381888 941351 381956 941407
rect 382012 941391 382080 941407
rect 382136 941391 382204 941407
rect 382260 941391 382328 941407
rect 382027 941351 382080 941391
rect 382169 941351 382204 941391
rect 382311 941351 382328 941391
rect 382384 941391 382452 941407
rect 382508 941391 382576 941407
rect 382632 941391 382700 941407
rect 382756 941391 382824 941407
rect 382384 941351 382397 941391
rect 382508 941351 382539 941391
rect 382632 941351 382681 941391
rect 382756 941351 382823 941391
rect 382880 941351 382948 941407
rect 383004 941391 383072 941407
rect 383128 941391 383196 941407
rect 383252 941391 383320 941407
rect 383021 941351 383072 941391
rect 383163 941351 383196 941391
rect 383305 941351 383320 941391
rect 383376 941391 383444 941407
rect 383500 941391 383568 941407
rect 383624 941391 383692 941407
rect 383376 941351 383391 941391
rect 383500 941351 383533 941391
rect 383624 941351 383675 941391
rect 383748 941351 383802 941407
rect 381885 941335 381971 941351
rect 382027 941335 382113 941351
rect 382169 941335 382255 941351
rect 382311 941335 382397 941351
rect 382453 941335 382539 941351
rect 382595 941335 382681 941351
rect 382737 941335 382823 941351
rect 382879 941335 382965 941351
rect 383021 941335 383107 941351
rect 383163 941335 383249 941351
rect 383305 941335 383391 941351
rect 383447 941335 383533 941351
rect 383589 941335 383675 941351
rect 383731 941335 383802 941351
rect 381752 941283 383802 941335
rect 381752 941249 381832 941283
rect 381752 941193 381829 941249
rect 381888 941227 381956 941283
rect 382012 941249 382080 941283
rect 382136 941249 382204 941283
rect 382260 941249 382328 941283
rect 382027 941227 382080 941249
rect 382169 941227 382204 941249
rect 382311 941227 382328 941249
rect 382384 941249 382452 941283
rect 382508 941249 382576 941283
rect 382632 941249 382700 941283
rect 382756 941249 382824 941283
rect 382384 941227 382397 941249
rect 382508 941227 382539 941249
rect 382632 941227 382681 941249
rect 382756 941227 382823 941249
rect 382880 941227 382948 941283
rect 383004 941249 383072 941283
rect 383128 941249 383196 941283
rect 383252 941249 383320 941283
rect 383021 941227 383072 941249
rect 383163 941227 383196 941249
rect 383305 941227 383320 941249
rect 383376 941249 383444 941283
rect 383500 941249 383568 941283
rect 383624 941249 383692 941283
rect 383376 941227 383391 941249
rect 383500 941227 383533 941249
rect 383624 941227 383675 941249
rect 383748 941227 383802 941283
rect 381885 941193 381971 941227
rect 382027 941193 382113 941227
rect 382169 941193 382255 941227
rect 382311 941193 382397 941227
rect 382453 941193 382539 941227
rect 382595 941193 382681 941227
rect 382737 941193 382823 941227
rect 382879 941193 382965 941227
rect 383021 941193 383107 941227
rect 383163 941193 383249 941227
rect 383305 941193 383391 941227
rect 383447 941193 383533 941227
rect 383589 941193 383675 941227
rect 383731 941193 383802 941227
rect 381752 941159 383802 941193
rect 381752 941107 381832 941159
rect 381752 941051 381829 941107
rect 381888 941103 381956 941159
rect 382012 941107 382080 941159
rect 382136 941107 382204 941159
rect 382260 941107 382328 941159
rect 382027 941103 382080 941107
rect 382169 941103 382204 941107
rect 382311 941103 382328 941107
rect 382384 941107 382452 941159
rect 382508 941107 382576 941159
rect 382632 941107 382700 941159
rect 382756 941107 382824 941159
rect 382384 941103 382397 941107
rect 382508 941103 382539 941107
rect 382632 941103 382681 941107
rect 382756 941103 382823 941107
rect 382880 941103 382948 941159
rect 383004 941107 383072 941159
rect 383128 941107 383196 941159
rect 383252 941107 383320 941159
rect 383021 941103 383072 941107
rect 383163 941103 383196 941107
rect 383305 941103 383320 941107
rect 383376 941107 383444 941159
rect 383500 941107 383568 941159
rect 383624 941107 383692 941159
rect 383376 941103 383391 941107
rect 383500 941103 383533 941107
rect 383624 941103 383675 941107
rect 383748 941103 383802 941159
rect 381885 941051 381971 941103
rect 382027 941051 382113 941103
rect 382169 941051 382255 941103
rect 382311 941051 382397 941103
rect 382453 941051 382539 941103
rect 382595 941051 382681 941103
rect 382737 941051 382823 941103
rect 382879 941051 382965 941103
rect 383021 941051 383107 941103
rect 383163 941051 383249 941103
rect 383305 941051 383391 941103
rect 383447 941051 383533 941103
rect 383589 941051 383675 941103
rect 383731 941051 383802 941103
rect 381752 941035 383802 941051
rect 381752 940979 381832 941035
rect 381888 940979 381956 941035
rect 382012 940979 382080 941035
rect 382136 940979 382204 941035
rect 382260 940979 382328 941035
rect 382384 940979 382452 941035
rect 382508 940979 382576 941035
rect 382632 940979 382700 941035
rect 382756 940979 382824 941035
rect 382880 940979 382948 941035
rect 383004 940979 383072 941035
rect 383128 940979 383196 941035
rect 383252 940979 383320 941035
rect 383376 940979 383444 941035
rect 383500 940979 383568 941035
rect 383624 940979 383692 941035
rect 383748 940979 383802 941035
rect 381752 940965 383802 940979
rect 381752 940909 381829 940965
rect 381885 940911 381971 940965
rect 382027 940911 382113 940965
rect 382169 940911 382255 940965
rect 382311 940911 382397 940965
rect 382453 940911 382539 940965
rect 382595 940911 382681 940965
rect 382737 940911 382823 940965
rect 382879 940911 382965 940965
rect 383021 940911 383107 940965
rect 383163 940911 383249 940965
rect 383305 940911 383391 940965
rect 383447 940911 383533 940965
rect 383589 940911 383675 940965
rect 383731 940911 383802 940965
rect 381752 940855 381832 940909
rect 381888 940855 381956 940911
rect 382027 940909 382080 940911
rect 382169 940909 382204 940911
rect 382311 940909 382328 940911
rect 382012 940855 382080 940909
rect 382136 940855 382204 940909
rect 382260 940855 382328 940909
rect 382384 940909 382397 940911
rect 382508 940909 382539 940911
rect 382632 940909 382681 940911
rect 382756 940909 382823 940911
rect 382384 940855 382452 940909
rect 382508 940855 382576 940909
rect 382632 940855 382700 940909
rect 382756 940855 382824 940909
rect 382880 940855 382948 940911
rect 383021 940909 383072 940911
rect 383163 940909 383196 940911
rect 383305 940909 383320 940911
rect 383004 940855 383072 940909
rect 383128 940855 383196 940909
rect 383252 940855 383320 940909
rect 383376 940909 383391 940911
rect 383500 940909 383533 940911
rect 383624 940909 383675 940911
rect 383376 940855 383444 940909
rect 383500 940855 383568 940909
rect 383624 940855 383692 940909
rect 383748 940855 383802 940911
rect 381752 940823 383802 940855
rect 381752 940767 381829 940823
rect 381885 940787 381971 940823
rect 382027 940787 382113 940823
rect 382169 940787 382255 940823
rect 382311 940787 382397 940823
rect 382453 940787 382539 940823
rect 382595 940787 382681 940823
rect 382737 940787 382823 940823
rect 382879 940787 382965 940823
rect 383021 940787 383107 940823
rect 383163 940787 383249 940823
rect 383305 940787 383391 940823
rect 383447 940787 383533 940823
rect 383589 940787 383675 940823
rect 383731 940787 383802 940823
rect 381752 940731 381832 940767
rect 381888 940731 381956 940787
rect 382027 940767 382080 940787
rect 382169 940767 382204 940787
rect 382311 940767 382328 940787
rect 382012 940731 382080 940767
rect 382136 940731 382204 940767
rect 382260 940731 382328 940767
rect 382384 940767 382397 940787
rect 382508 940767 382539 940787
rect 382632 940767 382681 940787
rect 382756 940767 382823 940787
rect 382384 940731 382452 940767
rect 382508 940731 382576 940767
rect 382632 940731 382700 940767
rect 382756 940731 382824 940767
rect 382880 940731 382948 940787
rect 383021 940767 383072 940787
rect 383163 940767 383196 940787
rect 383305 940767 383320 940787
rect 383004 940731 383072 940767
rect 383128 940731 383196 940767
rect 383252 940731 383320 940767
rect 383376 940767 383391 940787
rect 383500 940767 383533 940787
rect 383624 940767 383675 940787
rect 383376 940731 383444 940767
rect 383500 940731 383568 940767
rect 383624 940731 383692 940767
rect 383748 940731 383802 940787
rect 381752 940681 383802 940731
rect 381752 940625 381829 940681
rect 381885 940663 381971 940681
rect 382027 940663 382113 940681
rect 382169 940663 382255 940681
rect 382311 940663 382397 940681
rect 382453 940663 382539 940681
rect 382595 940663 382681 940681
rect 382737 940663 382823 940681
rect 382879 940663 382965 940681
rect 383021 940663 383107 940681
rect 383163 940663 383249 940681
rect 383305 940663 383391 940681
rect 383447 940663 383533 940681
rect 383589 940663 383675 940681
rect 383731 940663 383802 940681
rect 381752 940607 381832 940625
rect 381888 940607 381956 940663
rect 382027 940625 382080 940663
rect 382169 940625 382204 940663
rect 382311 940625 382328 940663
rect 382012 940607 382080 940625
rect 382136 940607 382204 940625
rect 382260 940607 382328 940625
rect 382384 940625 382397 940663
rect 382508 940625 382539 940663
rect 382632 940625 382681 940663
rect 382756 940625 382823 940663
rect 382384 940607 382452 940625
rect 382508 940607 382576 940625
rect 382632 940607 382700 940625
rect 382756 940607 382824 940625
rect 382880 940607 382948 940663
rect 383021 940625 383072 940663
rect 383163 940625 383196 940663
rect 383305 940625 383320 940663
rect 383004 940607 383072 940625
rect 383128 940607 383196 940625
rect 383252 940607 383320 940625
rect 383376 940625 383391 940663
rect 383500 940625 383533 940663
rect 383624 940625 383675 940663
rect 383376 940607 383444 940625
rect 383500 940607 383568 940625
rect 383624 940607 383692 940625
rect 383748 940607 383802 940663
rect 381752 940539 383802 940607
rect 381752 940483 381829 940539
rect 381888 940483 381956 940539
rect 382027 940483 382080 940539
rect 382169 940483 382204 940539
rect 382311 940483 382328 940539
rect 382384 940483 382397 940539
rect 382508 940483 382539 940539
rect 382632 940483 382681 940539
rect 382756 940483 382823 940539
rect 382880 940483 382948 940539
rect 383021 940483 383072 940539
rect 383163 940483 383196 940539
rect 383305 940483 383320 940539
rect 383376 940483 383391 940539
rect 383500 940483 383533 940539
rect 383624 940483 383675 940539
rect 383748 940483 383802 940539
rect 381752 940415 383802 940483
rect 381752 940397 381832 940415
rect 381752 940341 381829 940397
rect 381888 940359 381956 940415
rect 382012 940397 382080 940415
rect 382136 940397 382204 940415
rect 382260 940397 382328 940415
rect 382027 940359 382080 940397
rect 382169 940359 382204 940397
rect 382311 940359 382328 940397
rect 382384 940397 382452 940415
rect 382508 940397 382576 940415
rect 382632 940397 382700 940415
rect 382756 940397 382824 940415
rect 382384 940359 382397 940397
rect 382508 940359 382539 940397
rect 382632 940359 382681 940397
rect 382756 940359 382823 940397
rect 382880 940359 382948 940415
rect 383004 940397 383072 940415
rect 383128 940397 383196 940415
rect 383252 940397 383320 940415
rect 383021 940359 383072 940397
rect 383163 940359 383196 940397
rect 383305 940359 383320 940397
rect 383376 940397 383444 940415
rect 383500 940397 383568 940415
rect 383624 940397 383692 940415
rect 383376 940359 383391 940397
rect 383500 940359 383533 940397
rect 383624 940359 383675 940397
rect 383748 940359 383802 940415
rect 381885 940341 381971 940359
rect 382027 940341 382113 940359
rect 382169 940341 382255 940359
rect 382311 940341 382397 940359
rect 382453 940341 382539 940359
rect 382595 940341 382681 940359
rect 382737 940341 382823 940359
rect 382879 940341 382965 940359
rect 383021 940341 383107 940359
rect 383163 940341 383249 940359
rect 383305 940341 383391 940359
rect 383447 940341 383533 940359
rect 383589 940341 383675 940359
rect 383731 940341 383802 940359
rect 381752 940291 383802 940341
rect 381752 940255 381832 940291
rect 381752 940199 381829 940255
rect 381888 940235 381956 940291
rect 382012 940255 382080 940291
rect 382136 940255 382204 940291
rect 382260 940255 382328 940291
rect 382027 940235 382080 940255
rect 382169 940235 382204 940255
rect 382311 940235 382328 940255
rect 382384 940255 382452 940291
rect 382508 940255 382576 940291
rect 382632 940255 382700 940291
rect 382756 940255 382824 940291
rect 382384 940235 382397 940255
rect 382508 940235 382539 940255
rect 382632 940235 382681 940255
rect 382756 940235 382823 940255
rect 382880 940235 382948 940291
rect 383004 940255 383072 940291
rect 383128 940255 383196 940291
rect 383252 940255 383320 940291
rect 383021 940235 383072 940255
rect 383163 940235 383196 940255
rect 383305 940235 383320 940255
rect 383376 940255 383444 940291
rect 383500 940255 383568 940291
rect 383624 940255 383692 940291
rect 383376 940235 383391 940255
rect 383500 940235 383533 940255
rect 383624 940235 383675 940255
rect 383748 940235 383802 940291
rect 381885 940199 381971 940235
rect 382027 940199 382113 940235
rect 382169 940199 382255 940235
rect 382311 940199 382397 940235
rect 382453 940199 382539 940235
rect 382595 940199 382681 940235
rect 382737 940199 382823 940235
rect 382879 940199 382965 940235
rect 383021 940199 383107 940235
rect 383163 940199 383249 940235
rect 383305 940199 383391 940235
rect 383447 940199 383533 940235
rect 383589 940199 383675 940235
rect 383731 940199 383802 940235
rect 381752 940167 383802 940199
rect 381752 940113 381832 940167
rect 381752 940057 381829 940113
rect 381888 940111 381956 940167
rect 382012 940113 382080 940167
rect 382136 940113 382204 940167
rect 382260 940113 382328 940167
rect 382027 940111 382080 940113
rect 382169 940111 382204 940113
rect 382311 940111 382328 940113
rect 382384 940113 382452 940167
rect 382508 940113 382576 940167
rect 382632 940113 382700 940167
rect 382756 940113 382824 940167
rect 382384 940111 382397 940113
rect 382508 940111 382539 940113
rect 382632 940111 382681 940113
rect 382756 940111 382823 940113
rect 382880 940111 382948 940167
rect 383004 940113 383072 940167
rect 383128 940113 383196 940167
rect 383252 940113 383320 940167
rect 383021 940111 383072 940113
rect 383163 940111 383196 940113
rect 383305 940111 383320 940113
rect 383376 940113 383444 940167
rect 383500 940113 383568 940167
rect 383624 940113 383692 940167
rect 383376 940111 383391 940113
rect 383500 940111 383533 940113
rect 383624 940111 383675 940113
rect 383748 940111 383802 940167
rect 381885 940057 381971 940111
rect 382027 940057 382113 940111
rect 382169 940057 382255 940111
rect 382311 940057 382397 940111
rect 382453 940057 382539 940111
rect 382595 940057 382681 940111
rect 382737 940057 382823 940111
rect 382879 940057 382965 940111
rect 383021 940057 383107 940111
rect 383163 940057 383249 940111
rect 383305 940057 383391 940111
rect 383447 940057 383533 940111
rect 383589 940057 383675 940111
rect 383731 940057 383802 940111
rect 381752 940043 383802 940057
rect 381752 939987 381832 940043
rect 381888 939987 381956 940043
rect 382012 939987 382080 940043
rect 382136 939987 382204 940043
rect 382260 939987 382328 940043
rect 382384 939987 382452 940043
rect 382508 939987 382576 940043
rect 382632 939987 382700 940043
rect 382756 939987 382824 940043
rect 382880 939987 382948 940043
rect 383004 939987 383072 940043
rect 383128 939987 383196 940043
rect 383252 939987 383320 940043
rect 383376 939987 383444 940043
rect 383500 939987 383568 940043
rect 383624 939987 383692 940043
rect 383748 939987 383802 940043
rect 381752 939971 383802 939987
rect 381752 939915 381829 939971
rect 381885 939919 381971 939971
rect 382027 939919 382113 939971
rect 382169 939919 382255 939971
rect 382311 939919 382397 939971
rect 382453 939919 382539 939971
rect 382595 939919 382681 939971
rect 382737 939919 382823 939971
rect 382879 939919 382965 939971
rect 383021 939919 383107 939971
rect 383163 939919 383249 939971
rect 383305 939919 383391 939971
rect 383447 939919 383533 939971
rect 383589 939919 383675 939971
rect 383731 939919 383802 939971
rect 381752 939863 381832 939915
rect 381888 939863 381956 939919
rect 382027 939915 382080 939919
rect 382169 939915 382204 939919
rect 382311 939915 382328 939919
rect 382012 939863 382080 939915
rect 382136 939863 382204 939915
rect 382260 939863 382328 939915
rect 382384 939915 382397 939919
rect 382508 939915 382539 939919
rect 382632 939915 382681 939919
rect 382756 939915 382823 939919
rect 382384 939863 382452 939915
rect 382508 939863 382576 939915
rect 382632 939863 382700 939915
rect 382756 939863 382824 939915
rect 382880 939863 382948 939919
rect 383021 939915 383072 939919
rect 383163 939915 383196 939919
rect 383305 939915 383320 939919
rect 383004 939863 383072 939915
rect 383128 939863 383196 939915
rect 383252 939863 383320 939915
rect 383376 939915 383391 939919
rect 383500 939915 383533 939919
rect 383624 939915 383675 939919
rect 383376 939863 383444 939915
rect 383500 939863 383568 939915
rect 383624 939863 383692 939915
rect 383748 939863 383802 939919
rect 381752 939829 383802 939863
rect 381752 939773 381829 939829
rect 381885 939773 381971 939829
rect 382027 939773 382113 939829
rect 382169 939773 382255 939829
rect 382311 939773 382397 939829
rect 382453 939773 382539 939829
rect 382595 939773 382681 939829
rect 382737 939773 382823 939829
rect 382879 939773 382965 939829
rect 383021 939773 383107 939829
rect 383163 939773 383249 939829
rect 383305 939773 383391 939829
rect 383447 939773 383533 939829
rect 383589 939773 383675 939829
rect 383731 939773 383802 939829
rect 381752 939720 383802 939773
rect 384122 941675 386172 941720
rect 384122 941619 384199 941675
rect 384255 941655 384341 941675
rect 384397 941655 384483 941675
rect 384539 941655 384625 941675
rect 384681 941655 384767 941675
rect 384823 941655 384909 941675
rect 384965 941655 385051 941675
rect 385107 941655 385193 941675
rect 385249 941655 385335 941675
rect 385391 941655 385477 941675
rect 385533 941655 385619 941675
rect 385675 941655 385761 941675
rect 385817 941655 385903 941675
rect 385959 941655 386045 941675
rect 386101 941655 386172 941675
rect 384122 941599 384202 941619
rect 384258 941599 384326 941655
rect 384397 941619 384450 941655
rect 384539 941619 384574 941655
rect 384681 941619 384698 941655
rect 384382 941599 384450 941619
rect 384506 941599 384574 941619
rect 384630 941599 384698 941619
rect 384754 941619 384767 941655
rect 384878 941619 384909 941655
rect 385002 941619 385051 941655
rect 385126 941619 385193 941655
rect 384754 941599 384822 941619
rect 384878 941599 384946 941619
rect 385002 941599 385070 941619
rect 385126 941599 385194 941619
rect 385250 941599 385318 941655
rect 385391 941619 385442 941655
rect 385533 941619 385566 941655
rect 385675 941619 385690 941655
rect 385374 941599 385442 941619
rect 385498 941599 385566 941619
rect 385622 941599 385690 941619
rect 385746 941619 385761 941655
rect 385870 941619 385903 941655
rect 385994 941619 386045 941655
rect 385746 941599 385814 941619
rect 385870 941599 385938 941619
rect 385994 941599 386062 941619
rect 386118 941599 386172 941655
rect 384122 941533 386172 941599
rect 384122 941477 384199 941533
rect 384255 941531 384341 941533
rect 384397 941531 384483 941533
rect 384539 941531 384625 941533
rect 384681 941531 384767 941533
rect 384823 941531 384909 941533
rect 384965 941531 385051 941533
rect 385107 941531 385193 941533
rect 385249 941531 385335 941533
rect 385391 941531 385477 941533
rect 385533 941531 385619 941533
rect 385675 941531 385761 941533
rect 385817 941531 385903 941533
rect 385959 941531 386045 941533
rect 386101 941531 386172 941533
rect 384122 941475 384202 941477
rect 384258 941475 384326 941531
rect 384397 941477 384450 941531
rect 384539 941477 384574 941531
rect 384681 941477 384698 941531
rect 384382 941475 384450 941477
rect 384506 941475 384574 941477
rect 384630 941475 384698 941477
rect 384754 941477 384767 941531
rect 384878 941477 384909 941531
rect 385002 941477 385051 941531
rect 385126 941477 385193 941531
rect 384754 941475 384822 941477
rect 384878 941475 384946 941477
rect 385002 941475 385070 941477
rect 385126 941475 385194 941477
rect 385250 941475 385318 941531
rect 385391 941477 385442 941531
rect 385533 941477 385566 941531
rect 385675 941477 385690 941531
rect 385374 941475 385442 941477
rect 385498 941475 385566 941477
rect 385622 941475 385690 941477
rect 385746 941477 385761 941531
rect 385870 941477 385903 941531
rect 385994 941477 386045 941531
rect 385746 941475 385814 941477
rect 385870 941475 385938 941477
rect 385994 941475 386062 941477
rect 386118 941475 386172 941531
rect 384122 941407 386172 941475
rect 384122 941391 384202 941407
rect 384122 941335 384199 941391
rect 384258 941351 384326 941407
rect 384382 941391 384450 941407
rect 384506 941391 384574 941407
rect 384630 941391 384698 941407
rect 384397 941351 384450 941391
rect 384539 941351 384574 941391
rect 384681 941351 384698 941391
rect 384754 941391 384822 941407
rect 384878 941391 384946 941407
rect 385002 941391 385070 941407
rect 385126 941391 385194 941407
rect 384754 941351 384767 941391
rect 384878 941351 384909 941391
rect 385002 941351 385051 941391
rect 385126 941351 385193 941391
rect 385250 941351 385318 941407
rect 385374 941391 385442 941407
rect 385498 941391 385566 941407
rect 385622 941391 385690 941407
rect 385391 941351 385442 941391
rect 385533 941351 385566 941391
rect 385675 941351 385690 941391
rect 385746 941391 385814 941407
rect 385870 941391 385938 941407
rect 385994 941391 386062 941407
rect 385746 941351 385761 941391
rect 385870 941351 385903 941391
rect 385994 941351 386045 941391
rect 386118 941351 386172 941407
rect 384255 941335 384341 941351
rect 384397 941335 384483 941351
rect 384539 941335 384625 941351
rect 384681 941335 384767 941351
rect 384823 941335 384909 941351
rect 384965 941335 385051 941351
rect 385107 941335 385193 941351
rect 385249 941335 385335 941351
rect 385391 941335 385477 941351
rect 385533 941335 385619 941351
rect 385675 941335 385761 941351
rect 385817 941335 385903 941351
rect 385959 941335 386045 941351
rect 386101 941335 386172 941351
rect 384122 941283 386172 941335
rect 384122 941249 384202 941283
rect 384122 941193 384199 941249
rect 384258 941227 384326 941283
rect 384382 941249 384450 941283
rect 384506 941249 384574 941283
rect 384630 941249 384698 941283
rect 384397 941227 384450 941249
rect 384539 941227 384574 941249
rect 384681 941227 384698 941249
rect 384754 941249 384822 941283
rect 384878 941249 384946 941283
rect 385002 941249 385070 941283
rect 385126 941249 385194 941283
rect 384754 941227 384767 941249
rect 384878 941227 384909 941249
rect 385002 941227 385051 941249
rect 385126 941227 385193 941249
rect 385250 941227 385318 941283
rect 385374 941249 385442 941283
rect 385498 941249 385566 941283
rect 385622 941249 385690 941283
rect 385391 941227 385442 941249
rect 385533 941227 385566 941249
rect 385675 941227 385690 941249
rect 385746 941249 385814 941283
rect 385870 941249 385938 941283
rect 385994 941249 386062 941283
rect 385746 941227 385761 941249
rect 385870 941227 385903 941249
rect 385994 941227 386045 941249
rect 386118 941227 386172 941283
rect 384255 941193 384341 941227
rect 384397 941193 384483 941227
rect 384539 941193 384625 941227
rect 384681 941193 384767 941227
rect 384823 941193 384909 941227
rect 384965 941193 385051 941227
rect 385107 941193 385193 941227
rect 385249 941193 385335 941227
rect 385391 941193 385477 941227
rect 385533 941193 385619 941227
rect 385675 941193 385761 941227
rect 385817 941193 385903 941227
rect 385959 941193 386045 941227
rect 386101 941193 386172 941227
rect 384122 941159 386172 941193
rect 384122 941107 384202 941159
rect 384122 941051 384199 941107
rect 384258 941103 384326 941159
rect 384382 941107 384450 941159
rect 384506 941107 384574 941159
rect 384630 941107 384698 941159
rect 384397 941103 384450 941107
rect 384539 941103 384574 941107
rect 384681 941103 384698 941107
rect 384754 941107 384822 941159
rect 384878 941107 384946 941159
rect 385002 941107 385070 941159
rect 385126 941107 385194 941159
rect 384754 941103 384767 941107
rect 384878 941103 384909 941107
rect 385002 941103 385051 941107
rect 385126 941103 385193 941107
rect 385250 941103 385318 941159
rect 385374 941107 385442 941159
rect 385498 941107 385566 941159
rect 385622 941107 385690 941159
rect 385391 941103 385442 941107
rect 385533 941103 385566 941107
rect 385675 941103 385690 941107
rect 385746 941107 385814 941159
rect 385870 941107 385938 941159
rect 385994 941107 386062 941159
rect 385746 941103 385761 941107
rect 385870 941103 385903 941107
rect 385994 941103 386045 941107
rect 386118 941103 386172 941159
rect 384255 941051 384341 941103
rect 384397 941051 384483 941103
rect 384539 941051 384625 941103
rect 384681 941051 384767 941103
rect 384823 941051 384909 941103
rect 384965 941051 385051 941103
rect 385107 941051 385193 941103
rect 385249 941051 385335 941103
rect 385391 941051 385477 941103
rect 385533 941051 385619 941103
rect 385675 941051 385761 941103
rect 385817 941051 385903 941103
rect 385959 941051 386045 941103
rect 386101 941051 386172 941103
rect 384122 941035 386172 941051
rect 384122 940979 384202 941035
rect 384258 940979 384326 941035
rect 384382 940979 384450 941035
rect 384506 940979 384574 941035
rect 384630 940979 384698 941035
rect 384754 940979 384822 941035
rect 384878 940979 384946 941035
rect 385002 940979 385070 941035
rect 385126 940979 385194 941035
rect 385250 940979 385318 941035
rect 385374 940979 385442 941035
rect 385498 940979 385566 941035
rect 385622 940979 385690 941035
rect 385746 940979 385814 941035
rect 385870 940979 385938 941035
rect 385994 940979 386062 941035
rect 386118 940979 386172 941035
rect 384122 940965 386172 940979
rect 384122 940909 384199 940965
rect 384255 940911 384341 940965
rect 384397 940911 384483 940965
rect 384539 940911 384625 940965
rect 384681 940911 384767 940965
rect 384823 940911 384909 940965
rect 384965 940911 385051 940965
rect 385107 940911 385193 940965
rect 385249 940911 385335 940965
rect 385391 940911 385477 940965
rect 385533 940911 385619 940965
rect 385675 940911 385761 940965
rect 385817 940911 385903 940965
rect 385959 940911 386045 940965
rect 386101 940911 386172 940965
rect 384122 940855 384202 940909
rect 384258 940855 384326 940911
rect 384397 940909 384450 940911
rect 384539 940909 384574 940911
rect 384681 940909 384698 940911
rect 384382 940855 384450 940909
rect 384506 940855 384574 940909
rect 384630 940855 384698 940909
rect 384754 940909 384767 940911
rect 384878 940909 384909 940911
rect 385002 940909 385051 940911
rect 385126 940909 385193 940911
rect 384754 940855 384822 940909
rect 384878 940855 384946 940909
rect 385002 940855 385070 940909
rect 385126 940855 385194 940909
rect 385250 940855 385318 940911
rect 385391 940909 385442 940911
rect 385533 940909 385566 940911
rect 385675 940909 385690 940911
rect 385374 940855 385442 940909
rect 385498 940855 385566 940909
rect 385622 940855 385690 940909
rect 385746 940909 385761 940911
rect 385870 940909 385903 940911
rect 385994 940909 386045 940911
rect 385746 940855 385814 940909
rect 385870 940855 385938 940909
rect 385994 940855 386062 940909
rect 386118 940855 386172 940911
rect 384122 940823 386172 940855
rect 384122 940767 384199 940823
rect 384255 940787 384341 940823
rect 384397 940787 384483 940823
rect 384539 940787 384625 940823
rect 384681 940787 384767 940823
rect 384823 940787 384909 940823
rect 384965 940787 385051 940823
rect 385107 940787 385193 940823
rect 385249 940787 385335 940823
rect 385391 940787 385477 940823
rect 385533 940787 385619 940823
rect 385675 940787 385761 940823
rect 385817 940787 385903 940823
rect 385959 940787 386045 940823
rect 386101 940787 386172 940823
rect 384122 940731 384202 940767
rect 384258 940731 384326 940787
rect 384397 940767 384450 940787
rect 384539 940767 384574 940787
rect 384681 940767 384698 940787
rect 384382 940731 384450 940767
rect 384506 940731 384574 940767
rect 384630 940731 384698 940767
rect 384754 940767 384767 940787
rect 384878 940767 384909 940787
rect 385002 940767 385051 940787
rect 385126 940767 385193 940787
rect 384754 940731 384822 940767
rect 384878 940731 384946 940767
rect 385002 940731 385070 940767
rect 385126 940731 385194 940767
rect 385250 940731 385318 940787
rect 385391 940767 385442 940787
rect 385533 940767 385566 940787
rect 385675 940767 385690 940787
rect 385374 940731 385442 940767
rect 385498 940731 385566 940767
rect 385622 940731 385690 940767
rect 385746 940767 385761 940787
rect 385870 940767 385903 940787
rect 385994 940767 386045 940787
rect 385746 940731 385814 940767
rect 385870 940731 385938 940767
rect 385994 940731 386062 940767
rect 386118 940731 386172 940787
rect 384122 940681 386172 940731
rect 384122 940625 384199 940681
rect 384255 940663 384341 940681
rect 384397 940663 384483 940681
rect 384539 940663 384625 940681
rect 384681 940663 384767 940681
rect 384823 940663 384909 940681
rect 384965 940663 385051 940681
rect 385107 940663 385193 940681
rect 385249 940663 385335 940681
rect 385391 940663 385477 940681
rect 385533 940663 385619 940681
rect 385675 940663 385761 940681
rect 385817 940663 385903 940681
rect 385959 940663 386045 940681
rect 386101 940663 386172 940681
rect 384122 940607 384202 940625
rect 384258 940607 384326 940663
rect 384397 940625 384450 940663
rect 384539 940625 384574 940663
rect 384681 940625 384698 940663
rect 384382 940607 384450 940625
rect 384506 940607 384574 940625
rect 384630 940607 384698 940625
rect 384754 940625 384767 940663
rect 384878 940625 384909 940663
rect 385002 940625 385051 940663
rect 385126 940625 385193 940663
rect 384754 940607 384822 940625
rect 384878 940607 384946 940625
rect 385002 940607 385070 940625
rect 385126 940607 385194 940625
rect 385250 940607 385318 940663
rect 385391 940625 385442 940663
rect 385533 940625 385566 940663
rect 385675 940625 385690 940663
rect 385374 940607 385442 940625
rect 385498 940607 385566 940625
rect 385622 940607 385690 940625
rect 385746 940625 385761 940663
rect 385870 940625 385903 940663
rect 385994 940625 386045 940663
rect 385746 940607 385814 940625
rect 385870 940607 385938 940625
rect 385994 940607 386062 940625
rect 386118 940607 386172 940663
rect 384122 940539 386172 940607
rect 384122 940483 384199 940539
rect 384258 940483 384326 940539
rect 384397 940483 384450 940539
rect 384539 940483 384574 940539
rect 384681 940483 384698 940539
rect 384754 940483 384767 940539
rect 384878 940483 384909 940539
rect 385002 940483 385051 940539
rect 385126 940483 385193 940539
rect 385250 940483 385318 940539
rect 385391 940483 385442 940539
rect 385533 940483 385566 940539
rect 385675 940483 385690 940539
rect 385746 940483 385761 940539
rect 385870 940483 385903 940539
rect 385994 940483 386045 940539
rect 386118 940483 386172 940539
rect 384122 940415 386172 940483
rect 384122 940397 384202 940415
rect 384122 940341 384199 940397
rect 384258 940359 384326 940415
rect 384382 940397 384450 940415
rect 384506 940397 384574 940415
rect 384630 940397 384698 940415
rect 384397 940359 384450 940397
rect 384539 940359 384574 940397
rect 384681 940359 384698 940397
rect 384754 940397 384822 940415
rect 384878 940397 384946 940415
rect 385002 940397 385070 940415
rect 385126 940397 385194 940415
rect 384754 940359 384767 940397
rect 384878 940359 384909 940397
rect 385002 940359 385051 940397
rect 385126 940359 385193 940397
rect 385250 940359 385318 940415
rect 385374 940397 385442 940415
rect 385498 940397 385566 940415
rect 385622 940397 385690 940415
rect 385391 940359 385442 940397
rect 385533 940359 385566 940397
rect 385675 940359 385690 940397
rect 385746 940397 385814 940415
rect 385870 940397 385938 940415
rect 385994 940397 386062 940415
rect 385746 940359 385761 940397
rect 385870 940359 385903 940397
rect 385994 940359 386045 940397
rect 386118 940359 386172 940415
rect 384255 940341 384341 940359
rect 384397 940341 384483 940359
rect 384539 940341 384625 940359
rect 384681 940341 384767 940359
rect 384823 940341 384909 940359
rect 384965 940341 385051 940359
rect 385107 940341 385193 940359
rect 385249 940341 385335 940359
rect 385391 940341 385477 940359
rect 385533 940341 385619 940359
rect 385675 940341 385761 940359
rect 385817 940341 385903 940359
rect 385959 940341 386045 940359
rect 386101 940341 386172 940359
rect 384122 940291 386172 940341
rect 384122 940255 384202 940291
rect 384122 940199 384199 940255
rect 384258 940235 384326 940291
rect 384382 940255 384450 940291
rect 384506 940255 384574 940291
rect 384630 940255 384698 940291
rect 384397 940235 384450 940255
rect 384539 940235 384574 940255
rect 384681 940235 384698 940255
rect 384754 940255 384822 940291
rect 384878 940255 384946 940291
rect 385002 940255 385070 940291
rect 385126 940255 385194 940291
rect 384754 940235 384767 940255
rect 384878 940235 384909 940255
rect 385002 940235 385051 940255
rect 385126 940235 385193 940255
rect 385250 940235 385318 940291
rect 385374 940255 385442 940291
rect 385498 940255 385566 940291
rect 385622 940255 385690 940291
rect 385391 940235 385442 940255
rect 385533 940235 385566 940255
rect 385675 940235 385690 940255
rect 385746 940255 385814 940291
rect 385870 940255 385938 940291
rect 385994 940255 386062 940291
rect 385746 940235 385761 940255
rect 385870 940235 385903 940255
rect 385994 940235 386045 940255
rect 386118 940235 386172 940291
rect 384255 940199 384341 940235
rect 384397 940199 384483 940235
rect 384539 940199 384625 940235
rect 384681 940199 384767 940235
rect 384823 940199 384909 940235
rect 384965 940199 385051 940235
rect 385107 940199 385193 940235
rect 385249 940199 385335 940235
rect 385391 940199 385477 940235
rect 385533 940199 385619 940235
rect 385675 940199 385761 940235
rect 385817 940199 385903 940235
rect 385959 940199 386045 940235
rect 386101 940199 386172 940235
rect 384122 940167 386172 940199
rect 384122 940113 384202 940167
rect 384122 940057 384199 940113
rect 384258 940111 384326 940167
rect 384382 940113 384450 940167
rect 384506 940113 384574 940167
rect 384630 940113 384698 940167
rect 384397 940111 384450 940113
rect 384539 940111 384574 940113
rect 384681 940111 384698 940113
rect 384754 940113 384822 940167
rect 384878 940113 384946 940167
rect 385002 940113 385070 940167
rect 385126 940113 385194 940167
rect 384754 940111 384767 940113
rect 384878 940111 384909 940113
rect 385002 940111 385051 940113
rect 385126 940111 385193 940113
rect 385250 940111 385318 940167
rect 385374 940113 385442 940167
rect 385498 940113 385566 940167
rect 385622 940113 385690 940167
rect 385391 940111 385442 940113
rect 385533 940111 385566 940113
rect 385675 940111 385690 940113
rect 385746 940113 385814 940167
rect 385870 940113 385938 940167
rect 385994 940113 386062 940167
rect 385746 940111 385761 940113
rect 385870 940111 385903 940113
rect 385994 940111 386045 940113
rect 386118 940111 386172 940167
rect 384255 940057 384341 940111
rect 384397 940057 384483 940111
rect 384539 940057 384625 940111
rect 384681 940057 384767 940111
rect 384823 940057 384909 940111
rect 384965 940057 385051 940111
rect 385107 940057 385193 940111
rect 385249 940057 385335 940111
rect 385391 940057 385477 940111
rect 385533 940057 385619 940111
rect 385675 940057 385761 940111
rect 385817 940057 385903 940111
rect 385959 940057 386045 940111
rect 386101 940057 386172 940111
rect 384122 940043 386172 940057
rect 384122 939987 384202 940043
rect 384258 939987 384326 940043
rect 384382 939987 384450 940043
rect 384506 939987 384574 940043
rect 384630 939987 384698 940043
rect 384754 939987 384822 940043
rect 384878 939987 384946 940043
rect 385002 939987 385070 940043
rect 385126 939987 385194 940043
rect 385250 939987 385318 940043
rect 385374 939987 385442 940043
rect 385498 939987 385566 940043
rect 385622 939987 385690 940043
rect 385746 939987 385814 940043
rect 385870 939987 385938 940043
rect 385994 939987 386062 940043
rect 386118 939987 386172 940043
rect 384122 939971 386172 939987
rect 384122 939915 384199 939971
rect 384255 939919 384341 939971
rect 384397 939919 384483 939971
rect 384539 939919 384625 939971
rect 384681 939919 384767 939971
rect 384823 939919 384909 939971
rect 384965 939919 385051 939971
rect 385107 939919 385193 939971
rect 385249 939919 385335 939971
rect 385391 939919 385477 939971
rect 385533 939919 385619 939971
rect 385675 939919 385761 939971
rect 385817 939919 385903 939971
rect 385959 939919 386045 939971
rect 386101 939919 386172 939971
rect 384122 939863 384202 939915
rect 384258 939863 384326 939919
rect 384397 939915 384450 939919
rect 384539 939915 384574 939919
rect 384681 939915 384698 939919
rect 384382 939863 384450 939915
rect 384506 939863 384574 939915
rect 384630 939863 384698 939915
rect 384754 939915 384767 939919
rect 384878 939915 384909 939919
rect 385002 939915 385051 939919
rect 385126 939915 385193 939919
rect 384754 939863 384822 939915
rect 384878 939863 384946 939915
rect 385002 939863 385070 939915
rect 385126 939863 385194 939915
rect 385250 939863 385318 939919
rect 385391 939915 385442 939919
rect 385533 939915 385566 939919
rect 385675 939915 385690 939919
rect 385374 939863 385442 939915
rect 385498 939863 385566 939915
rect 385622 939863 385690 939915
rect 385746 939915 385761 939919
rect 385870 939915 385903 939919
rect 385994 939915 386045 939919
rect 385746 939863 385814 939915
rect 385870 939863 385938 939915
rect 385994 939863 386062 939915
rect 386118 939863 386172 939919
rect 384122 939829 386172 939863
rect 384122 939773 384199 939829
rect 384255 939773 384341 939829
rect 384397 939773 384483 939829
rect 384539 939773 384625 939829
rect 384681 939773 384767 939829
rect 384823 939773 384909 939829
rect 384965 939773 385051 939829
rect 385107 939773 385193 939829
rect 385249 939773 385335 939829
rect 385391 939773 385477 939829
rect 385533 939773 385619 939829
rect 385675 939773 385761 939829
rect 385817 939773 385903 939829
rect 385959 939773 386045 939829
rect 386101 939773 386172 939829
rect 384122 939720 386172 939773
rect 386828 941675 388878 941720
rect 386828 941619 386905 941675
rect 386961 941655 387047 941675
rect 387103 941655 387189 941675
rect 387245 941655 387331 941675
rect 387387 941655 387473 941675
rect 387529 941655 387615 941675
rect 387671 941655 387757 941675
rect 387813 941655 387899 941675
rect 387955 941655 388041 941675
rect 388097 941655 388183 941675
rect 388239 941655 388325 941675
rect 388381 941655 388467 941675
rect 388523 941655 388609 941675
rect 388665 941655 388751 941675
rect 388807 941655 388878 941675
rect 386828 941599 386908 941619
rect 386964 941599 387032 941655
rect 387103 941619 387156 941655
rect 387245 941619 387280 941655
rect 387387 941619 387404 941655
rect 387088 941599 387156 941619
rect 387212 941599 387280 941619
rect 387336 941599 387404 941619
rect 387460 941619 387473 941655
rect 387584 941619 387615 941655
rect 387708 941619 387757 941655
rect 387832 941619 387899 941655
rect 387460 941599 387528 941619
rect 387584 941599 387652 941619
rect 387708 941599 387776 941619
rect 387832 941599 387900 941619
rect 387956 941599 388024 941655
rect 388097 941619 388148 941655
rect 388239 941619 388272 941655
rect 388381 941619 388396 941655
rect 388080 941599 388148 941619
rect 388204 941599 388272 941619
rect 388328 941599 388396 941619
rect 388452 941619 388467 941655
rect 388576 941619 388609 941655
rect 388700 941619 388751 941655
rect 388452 941599 388520 941619
rect 388576 941599 388644 941619
rect 388700 941599 388768 941619
rect 388824 941599 388878 941655
rect 386828 941533 388878 941599
rect 386828 941477 386905 941533
rect 386961 941531 387047 941533
rect 387103 941531 387189 941533
rect 387245 941531 387331 941533
rect 387387 941531 387473 941533
rect 387529 941531 387615 941533
rect 387671 941531 387757 941533
rect 387813 941531 387899 941533
rect 387955 941531 388041 941533
rect 388097 941531 388183 941533
rect 388239 941531 388325 941533
rect 388381 941531 388467 941533
rect 388523 941531 388609 941533
rect 388665 941531 388751 941533
rect 388807 941531 388878 941533
rect 386828 941475 386908 941477
rect 386964 941475 387032 941531
rect 387103 941477 387156 941531
rect 387245 941477 387280 941531
rect 387387 941477 387404 941531
rect 387088 941475 387156 941477
rect 387212 941475 387280 941477
rect 387336 941475 387404 941477
rect 387460 941477 387473 941531
rect 387584 941477 387615 941531
rect 387708 941477 387757 941531
rect 387832 941477 387899 941531
rect 387460 941475 387528 941477
rect 387584 941475 387652 941477
rect 387708 941475 387776 941477
rect 387832 941475 387900 941477
rect 387956 941475 388024 941531
rect 388097 941477 388148 941531
rect 388239 941477 388272 941531
rect 388381 941477 388396 941531
rect 388080 941475 388148 941477
rect 388204 941475 388272 941477
rect 388328 941475 388396 941477
rect 388452 941477 388467 941531
rect 388576 941477 388609 941531
rect 388700 941477 388751 941531
rect 388452 941475 388520 941477
rect 388576 941475 388644 941477
rect 388700 941475 388768 941477
rect 388824 941475 388878 941531
rect 386828 941407 388878 941475
rect 386828 941391 386908 941407
rect 386828 941335 386905 941391
rect 386964 941351 387032 941407
rect 387088 941391 387156 941407
rect 387212 941391 387280 941407
rect 387336 941391 387404 941407
rect 387103 941351 387156 941391
rect 387245 941351 387280 941391
rect 387387 941351 387404 941391
rect 387460 941391 387528 941407
rect 387584 941391 387652 941407
rect 387708 941391 387776 941407
rect 387832 941391 387900 941407
rect 387460 941351 387473 941391
rect 387584 941351 387615 941391
rect 387708 941351 387757 941391
rect 387832 941351 387899 941391
rect 387956 941351 388024 941407
rect 388080 941391 388148 941407
rect 388204 941391 388272 941407
rect 388328 941391 388396 941407
rect 388097 941351 388148 941391
rect 388239 941351 388272 941391
rect 388381 941351 388396 941391
rect 388452 941391 388520 941407
rect 388576 941391 388644 941407
rect 388700 941391 388768 941407
rect 388452 941351 388467 941391
rect 388576 941351 388609 941391
rect 388700 941351 388751 941391
rect 388824 941351 388878 941407
rect 386961 941335 387047 941351
rect 387103 941335 387189 941351
rect 387245 941335 387331 941351
rect 387387 941335 387473 941351
rect 387529 941335 387615 941351
rect 387671 941335 387757 941351
rect 387813 941335 387899 941351
rect 387955 941335 388041 941351
rect 388097 941335 388183 941351
rect 388239 941335 388325 941351
rect 388381 941335 388467 941351
rect 388523 941335 388609 941351
rect 388665 941335 388751 941351
rect 388807 941335 388878 941351
rect 386828 941283 388878 941335
rect 386828 941249 386908 941283
rect 386828 941193 386905 941249
rect 386964 941227 387032 941283
rect 387088 941249 387156 941283
rect 387212 941249 387280 941283
rect 387336 941249 387404 941283
rect 387103 941227 387156 941249
rect 387245 941227 387280 941249
rect 387387 941227 387404 941249
rect 387460 941249 387528 941283
rect 387584 941249 387652 941283
rect 387708 941249 387776 941283
rect 387832 941249 387900 941283
rect 387460 941227 387473 941249
rect 387584 941227 387615 941249
rect 387708 941227 387757 941249
rect 387832 941227 387899 941249
rect 387956 941227 388024 941283
rect 388080 941249 388148 941283
rect 388204 941249 388272 941283
rect 388328 941249 388396 941283
rect 388097 941227 388148 941249
rect 388239 941227 388272 941249
rect 388381 941227 388396 941249
rect 388452 941249 388520 941283
rect 388576 941249 388644 941283
rect 388700 941249 388768 941283
rect 388452 941227 388467 941249
rect 388576 941227 388609 941249
rect 388700 941227 388751 941249
rect 388824 941227 388878 941283
rect 386961 941193 387047 941227
rect 387103 941193 387189 941227
rect 387245 941193 387331 941227
rect 387387 941193 387473 941227
rect 387529 941193 387615 941227
rect 387671 941193 387757 941227
rect 387813 941193 387899 941227
rect 387955 941193 388041 941227
rect 388097 941193 388183 941227
rect 388239 941193 388325 941227
rect 388381 941193 388467 941227
rect 388523 941193 388609 941227
rect 388665 941193 388751 941227
rect 388807 941193 388878 941227
rect 386828 941159 388878 941193
rect 386828 941107 386908 941159
rect 386828 941051 386905 941107
rect 386964 941103 387032 941159
rect 387088 941107 387156 941159
rect 387212 941107 387280 941159
rect 387336 941107 387404 941159
rect 387103 941103 387156 941107
rect 387245 941103 387280 941107
rect 387387 941103 387404 941107
rect 387460 941107 387528 941159
rect 387584 941107 387652 941159
rect 387708 941107 387776 941159
rect 387832 941107 387900 941159
rect 387460 941103 387473 941107
rect 387584 941103 387615 941107
rect 387708 941103 387757 941107
rect 387832 941103 387899 941107
rect 387956 941103 388024 941159
rect 388080 941107 388148 941159
rect 388204 941107 388272 941159
rect 388328 941107 388396 941159
rect 388097 941103 388148 941107
rect 388239 941103 388272 941107
rect 388381 941103 388396 941107
rect 388452 941107 388520 941159
rect 388576 941107 388644 941159
rect 388700 941107 388768 941159
rect 388452 941103 388467 941107
rect 388576 941103 388609 941107
rect 388700 941103 388751 941107
rect 388824 941103 388878 941159
rect 386961 941051 387047 941103
rect 387103 941051 387189 941103
rect 387245 941051 387331 941103
rect 387387 941051 387473 941103
rect 387529 941051 387615 941103
rect 387671 941051 387757 941103
rect 387813 941051 387899 941103
rect 387955 941051 388041 941103
rect 388097 941051 388183 941103
rect 388239 941051 388325 941103
rect 388381 941051 388467 941103
rect 388523 941051 388609 941103
rect 388665 941051 388751 941103
rect 388807 941051 388878 941103
rect 386828 941035 388878 941051
rect 386828 940979 386908 941035
rect 386964 940979 387032 941035
rect 387088 940979 387156 941035
rect 387212 940979 387280 941035
rect 387336 940979 387404 941035
rect 387460 940979 387528 941035
rect 387584 940979 387652 941035
rect 387708 940979 387776 941035
rect 387832 940979 387900 941035
rect 387956 940979 388024 941035
rect 388080 940979 388148 941035
rect 388204 940979 388272 941035
rect 388328 940979 388396 941035
rect 388452 940979 388520 941035
rect 388576 940979 388644 941035
rect 388700 940979 388768 941035
rect 388824 940979 388878 941035
rect 386828 940965 388878 940979
rect 386828 940909 386905 940965
rect 386961 940911 387047 940965
rect 387103 940911 387189 940965
rect 387245 940911 387331 940965
rect 387387 940911 387473 940965
rect 387529 940911 387615 940965
rect 387671 940911 387757 940965
rect 387813 940911 387899 940965
rect 387955 940911 388041 940965
rect 388097 940911 388183 940965
rect 388239 940911 388325 940965
rect 388381 940911 388467 940965
rect 388523 940911 388609 940965
rect 388665 940911 388751 940965
rect 388807 940911 388878 940965
rect 386828 940855 386908 940909
rect 386964 940855 387032 940911
rect 387103 940909 387156 940911
rect 387245 940909 387280 940911
rect 387387 940909 387404 940911
rect 387088 940855 387156 940909
rect 387212 940855 387280 940909
rect 387336 940855 387404 940909
rect 387460 940909 387473 940911
rect 387584 940909 387615 940911
rect 387708 940909 387757 940911
rect 387832 940909 387899 940911
rect 387460 940855 387528 940909
rect 387584 940855 387652 940909
rect 387708 940855 387776 940909
rect 387832 940855 387900 940909
rect 387956 940855 388024 940911
rect 388097 940909 388148 940911
rect 388239 940909 388272 940911
rect 388381 940909 388396 940911
rect 388080 940855 388148 940909
rect 388204 940855 388272 940909
rect 388328 940855 388396 940909
rect 388452 940909 388467 940911
rect 388576 940909 388609 940911
rect 388700 940909 388751 940911
rect 388452 940855 388520 940909
rect 388576 940855 388644 940909
rect 388700 940855 388768 940909
rect 388824 940855 388878 940911
rect 386828 940823 388878 940855
rect 386828 940767 386905 940823
rect 386961 940787 387047 940823
rect 387103 940787 387189 940823
rect 387245 940787 387331 940823
rect 387387 940787 387473 940823
rect 387529 940787 387615 940823
rect 387671 940787 387757 940823
rect 387813 940787 387899 940823
rect 387955 940787 388041 940823
rect 388097 940787 388183 940823
rect 388239 940787 388325 940823
rect 388381 940787 388467 940823
rect 388523 940787 388609 940823
rect 388665 940787 388751 940823
rect 388807 940787 388878 940823
rect 386828 940731 386908 940767
rect 386964 940731 387032 940787
rect 387103 940767 387156 940787
rect 387245 940767 387280 940787
rect 387387 940767 387404 940787
rect 387088 940731 387156 940767
rect 387212 940731 387280 940767
rect 387336 940731 387404 940767
rect 387460 940767 387473 940787
rect 387584 940767 387615 940787
rect 387708 940767 387757 940787
rect 387832 940767 387899 940787
rect 387460 940731 387528 940767
rect 387584 940731 387652 940767
rect 387708 940731 387776 940767
rect 387832 940731 387900 940767
rect 387956 940731 388024 940787
rect 388097 940767 388148 940787
rect 388239 940767 388272 940787
rect 388381 940767 388396 940787
rect 388080 940731 388148 940767
rect 388204 940731 388272 940767
rect 388328 940731 388396 940767
rect 388452 940767 388467 940787
rect 388576 940767 388609 940787
rect 388700 940767 388751 940787
rect 388452 940731 388520 940767
rect 388576 940731 388644 940767
rect 388700 940731 388768 940767
rect 388824 940731 388878 940787
rect 386828 940681 388878 940731
rect 386828 940625 386905 940681
rect 386961 940663 387047 940681
rect 387103 940663 387189 940681
rect 387245 940663 387331 940681
rect 387387 940663 387473 940681
rect 387529 940663 387615 940681
rect 387671 940663 387757 940681
rect 387813 940663 387899 940681
rect 387955 940663 388041 940681
rect 388097 940663 388183 940681
rect 388239 940663 388325 940681
rect 388381 940663 388467 940681
rect 388523 940663 388609 940681
rect 388665 940663 388751 940681
rect 388807 940663 388878 940681
rect 386828 940607 386908 940625
rect 386964 940607 387032 940663
rect 387103 940625 387156 940663
rect 387245 940625 387280 940663
rect 387387 940625 387404 940663
rect 387088 940607 387156 940625
rect 387212 940607 387280 940625
rect 387336 940607 387404 940625
rect 387460 940625 387473 940663
rect 387584 940625 387615 940663
rect 387708 940625 387757 940663
rect 387832 940625 387899 940663
rect 387460 940607 387528 940625
rect 387584 940607 387652 940625
rect 387708 940607 387776 940625
rect 387832 940607 387900 940625
rect 387956 940607 388024 940663
rect 388097 940625 388148 940663
rect 388239 940625 388272 940663
rect 388381 940625 388396 940663
rect 388080 940607 388148 940625
rect 388204 940607 388272 940625
rect 388328 940607 388396 940625
rect 388452 940625 388467 940663
rect 388576 940625 388609 940663
rect 388700 940625 388751 940663
rect 388452 940607 388520 940625
rect 388576 940607 388644 940625
rect 388700 940607 388768 940625
rect 388824 940607 388878 940663
rect 386828 940539 388878 940607
rect 386828 940483 386905 940539
rect 386964 940483 387032 940539
rect 387103 940483 387156 940539
rect 387245 940483 387280 940539
rect 387387 940483 387404 940539
rect 387460 940483 387473 940539
rect 387584 940483 387615 940539
rect 387708 940483 387757 940539
rect 387832 940483 387899 940539
rect 387956 940483 388024 940539
rect 388097 940483 388148 940539
rect 388239 940483 388272 940539
rect 388381 940483 388396 940539
rect 388452 940483 388467 940539
rect 388576 940483 388609 940539
rect 388700 940483 388751 940539
rect 388824 940483 388878 940539
rect 386828 940415 388878 940483
rect 386828 940397 386908 940415
rect 386828 940341 386905 940397
rect 386964 940359 387032 940415
rect 387088 940397 387156 940415
rect 387212 940397 387280 940415
rect 387336 940397 387404 940415
rect 387103 940359 387156 940397
rect 387245 940359 387280 940397
rect 387387 940359 387404 940397
rect 387460 940397 387528 940415
rect 387584 940397 387652 940415
rect 387708 940397 387776 940415
rect 387832 940397 387900 940415
rect 387460 940359 387473 940397
rect 387584 940359 387615 940397
rect 387708 940359 387757 940397
rect 387832 940359 387899 940397
rect 387956 940359 388024 940415
rect 388080 940397 388148 940415
rect 388204 940397 388272 940415
rect 388328 940397 388396 940415
rect 388097 940359 388148 940397
rect 388239 940359 388272 940397
rect 388381 940359 388396 940397
rect 388452 940397 388520 940415
rect 388576 940397 388644 940415
rect 388700 940397 388768 940415
rect 388452 940359 388467 940397
rect 388576 940359 388609 940397
rect 388700 940359 388751 940397
rect 388824 940359 388878 940415
rect 386961 940341 387047 940359
rect 387103 940341 387189 940359
rect 387245 940341 387331 940359
rect 387387 940341 387473 940359
rect 387529 940341 387615 940359
rect 387671 940341 387757 940359
rect 387813 940341 387899 940359
rect 387955 940341 388041 940359
rect 388097 940341 388183 940359
rect 388239 940341 388325 940359
rect 388381 940341 388467 940359
rect 388523 940341 388609 940359
rect 388665 940341 388751 940359
rect 388807 940341 388878 940359
rect 386828 940291 388878 940341
rect 386828 940255 386908 940291
rect 386828 940199 386905 940255
rect 386964 940235 387032 940291
rect 387088 940255 387156 940291
rect 387212 940255 387280 940291
rect 387336 940255 387404 940291
rect 387103 940235 387156 940255
rect 387245 940235 387280 940255
rect 387387 940235 387404 940255
rect 387460 940255 387528 940291
rect 387584 940255 387652 940291
rect 387708 940255 387776 940291
rect 387832 940255 387900 940291
rect 387460 940235 387473 940255
rect 387584 940235 387615 940255
rect 387708 940235 387757 940255
rect 387832 940235 387899 940255
rect 387956 940235 388024 940291
rect 388080 940255 388148 940291
rect 388204 940255 388272 940291
rect 388328 940255 388396 940291
rect 388097 940235 388148 940255
rect 388239 940235 388272 940255
rect 388381 940235 388396 940255
rect 388452 940255 388520 940291
rect 388576 940255 388644 940291
rect 388700 940255 388768 940291
rect 388452 940235 388467 940255
rect 388576 940235 388609 940255
rect 388700 940235 388751 940255
rect 388824 940235 388878 940291
rect 386961 940199 387047 940235
rect 387103 940199 387189 940235
rect 387245 940199 387331 940235
rect 387387 940199 387473 940235
rect 387529 940199 387615 940235
rect 387671 940199 387757 940235
rect 387813 940199 387899 940235
rect 387955 940199 388041 940235
rect 388097 940199 388183 940235
rect 388239 940199 388325 940235
rect 388381 940199 388467 940235
rect 388523 940199 388609 940235
rect 388665 940199 388751 940235
rect 388807 940199 388878 940235
rect 386828 940167 388878 940199
rect 386828 940113 386908 940167
rect 386828 940057 386905 940113
rect 386964 940111 387032 940167
rect 387088 940113 387156 940167
rect 387212 940113 387280 940167
rect 387336 940113 387404 940167
rect 387103 940111 387156 940113
rect 387245 940111 387280 940113
rect 387387 940111 387404 940113
rect 387460 940113 387528 940167
rect 387584 940113 387652 940167
rect 387708 940113 387776 940167
rect 387832 940113 387900 940167
rect 387460 940111 387473 940113
rect 387584 940111 387615 940113
rect 387708 940111 387757 940113
rect 387832 940111 387899 940113
rect 387956 940111 388024 940167
rect 388080 940113 388148 940167
rect 388204 940113 388272 940167
rect 388328 940113 388396 940167
rect 388097 940111 388148 940113
rect 388239 940111 388272 940113
rect 388381 940111 388396 940113
rect 388452 940113 388520 940167
rect 388576 940113 388644 940167
rect 388700 940113 388768 940167
rect 388452 940111 388467 940113
rect 388576 940111 388609 940113
rect 388700 940111 388751 940113
rect 388824 940111 388878 940167
rect 386961 940057 387047 940111
rect 387103 940057 387189 940111
rect 387245 940057 387331 940111
rect 387387 940057 387473 940111
rect 387529 940057 387615 940111
rect 387671 940057 387757 940111
rect 387813 940057 387899 940111
rect 387955 940057 388041 940111
rect 388097 940057 388183 940111
rect 388239 940057 388325 940111
rect 388381 940057 388467 940111
rect 388523 940057 388609 940111
rect 388665 940057 388751 940111
rect 388807 940057 388878 940111
rect 386828 940043 388878 940057
rect 386828 939987 386908 940043
rect 386964 939987 387032 940043
rect 387088 939987 387156 940043
rect 387212 939987 387280 940043
rect 387336 939987 387404 940043
rect 387460 939987 387528 940043
rect 387584 939987 387652 940043
rect 387708 939987 387776 940043
rect 387832 939987 387900 940043
rect 387956 939987 388024 940043
rect 388080 939987 388148 940043
rect 388204 939987 388272 940043
rect 388328 939987 388396 940043
rect 388452 939987 388520 940043
rect 388576 939987 388644 940043
rect 388700 939987 388768 940043
rect 388824 939987 388878 940043
rect 386828 939971 388878 939987
rect 386828 939915 386905 939971
rect 386961 939919 387047 939971
rect 387103 939919 387189 939971
rect 387245 939919 387331 939971
rect 387387 939919 387473 939971
rect 387529 939919 387615 939971
rect 387671 939919 387757 939971
rect 387813 939919 387899 939971
rect 387955 939919 388041 939971
rect 388097 939919 388183 939971
rect 388239 939919 388325 939971
rect 388381 939919 388467 939971
rect 388523 939919 388609 939971
rect 388665 939919 388751 939971
rect 388807 939919 388878 939971
rect 386828 939863 386908 939915
rect 386964 939863 387032 939919
rect 387103 939915 387156 939919
rect 387245 939915 387280 939919
rect 387387 939915 387404 939919
rect 387088 939863 387156 939915
rect 387212 939863 387280 939915
rect 387336 939863 387404 939915
rect 387460 939915 387473 939919
rect 387584 939915 387615 939919
rect 387708 939915 387757 939919
rect 387832 939915 387899 939919
rect 387460 939863 387528 939915
rect 387584 939863 387652 939915
rect 387708 939863 387776 939915
rect 387832 939863 387900 939915
rect 387956 939863 388024 939919
rect 388097 939915 388148 939919
rect 388239 939915 388272 939919
rect 388381 939915 388396 939919
rect 388080 939863 388148 939915
rect 388204 939863 388272 939915
rect 388328 939863 388396 939915
rect 388452 939915 388467 939919
rect 388576 939915 388609 939919
rect 388700 939915 388751 939919
rect 388452 939863 388520 939915
rect 388576 939863 388644 939915
rect 388700 939863 388768 939915
rect 388824 939863 388878 939919
rect 386828 939829 388878 939863
rect 386828 939773 386905 939829
rect 386961 939773 387047 939829
rect 387103 939773 387189 939829
rect 387245 939773 387331 939829
rect 387387 939773 387473 939829
rect 387529 939773 387615 939829
rect 387671 939773 387757 939829
rect 387813 939773 387899 939829
rect 387955 939773 388041 939829
rect 388097 939773 388183 939829
rect 388239 939773 388325 939829
rect 388381 939773 388467 939829
rect 388523 939773 388609 939829
rect 388665 939773 388751 939829
rect 388807 939773 388878 939829
rect 386828 939720 388878 939773
rect 389198 941675 391248 941720
rect 389198 941619 389275 941675
rect 389331 941655 389417 941675
rect 389473 941655 389559 941675
rect 389615 941655 389701 941675
rect 389757 941655 389843 941675
rect 389899 941655 389985 941675
rect 390041 941655 390127 941675
rect 390183 941655 390269 941675
rect 390325 941655 390411 941675
rect 390467 941655 390553 941675
rect 390609 941655 390695 941675
rect 390751 941655 390837 941675
rect 390893 941655 390979 941675
rect 391035 941655 391121 941675
rect 391177 941655 391248 941675
rect 389198 941599 389278 941619
rect 389334 941599 389402 941655
rect 389473 941619 389526 941655
rect 389615 941619 389650 941655
rect 389757 941619 389774 941655
rect 389458 941599 389526 941619
rect 389582 941599 389650 941619
rect 389706 941599 389774 941619
rect 389830 941619 389843 941655
rect 389954 941619 389985 941655
rect 390078 941619 390127 941655
rect 390202 941619 390269 941655
rect 389830 941599 389898 941619
rect 389954 941599 390022 941619
rect 390078 941599 390146 941619
rect 390202 941599 390270 941619
rect 390326 941599 390394 941655
rect 390467 941619 390518 941655
rect 390609 941619 390642 941655
rect 390751 941619 390766 941655
rect 390450 941599 390518 941619
rect 390574 941599 390642 941619
rect 390698 941599 390766 941619
rect 390822 941619 390837 941655
rect 390946 941619 390979 941655
rect 391070 941619 391121 941655
rect 390822 941599 390890 941619
rect 390946 941599 391014 941619
rect 391070 941599 391138 941619
rect 391194 941599 391248 941655
rect 389198 941533 391248 941599
rect 389198 941477 389275 941533
rect 389331 941531 389417 941533
rect 389473 941531 389559 941533
rect 389615 941531 389701 941533
rect 389757 941531 389843 941533
rect 389899 941531 389985 941533
rect 390041 941531 390127 941533
rect 390183 941531 390269 941533
rect 390325 941531 390411 941533
rect 390467 941531 390553 941533
rect 390609 941531 390695 941533
rect 390751 941531 390837 941533
rect 390893 941531 390979 941533
rect 391035 941531 391121 941533
rect 391177 941531 391248 941533
rect 389198 941475 389278 941477
rect 389334 941475 389402 941531
rect 389473 941477 389526 941531
rect 389615 941477 389650 941531
rect 389757 941477 389774 941531
rect 389458 941475 389526 941477
rect 389582 941475 389650 941477
rect 389706 941475 389774 941477
rect 389830 941477 389843 941531
rect 389954 941477 389985 941531
rect 390078 941477 390127 941531
rect 390202 941477 390269 941531
rect 389830 941475 389898 941477
rect 389954 941475 390022 941477
rect 390078 941475 390146 941477
rect 390202 941475 390270 941477
rect 390326 941475 390394 941531
rect 390467 941477 390518 941531
rect 390609 941477 390642 941531
rect 390751 941477 390766 941531
rect 390450 941475 390518 941477
rect 390574 941475 390642 941477
rect 390698 941475 390766 941477
rect 390822 941477 390837 941531
rect 390946 941477 390979 941531
rect 391070 941477 391121 941531
rect 390822 941475 390890 941477
rect 390946 941475 391014 941477
rect 391070 941475 391138 941477
rect 391194 941475 391248 941531
rect 389198 941407 391248 941475
rect 389198 941391 389278 941407
rect 389198 941335 389275 941391
rect 389334 941351 389402 941407
rect 389458 941391 389526 941407
rect 389582 941391 389650 941407
rect 389706 941391 389774 941407
rect 389473 941351 389526 941391
rect 389615 941351 389650 941391
rect 389757 941351 389774 941391
rect 389830 941391 389898 941407
rect 389954 941391 390022 941407
rect 390078 941391 390146 941407
rect 390202 941391 390270 941407
rect 389830 941351 389843 941391
rect 389954 941351 389985 941391
rect 390078 941351 390127 941391
rect 390202 941351 390269 941391
rect 390326 941351 390394 941407
rect 390450 941391 390518 941407
rect 390574 941391 390642 941407
rect 390698 941391 390766 941407
rect 390467 941351 390518 941391
rect 390609 941351 390642 941391
rect 390751 941351 390766 941391
rect 390822 941391 390890 941407
rect 390946 941391 391014 941407
rect 391070 941391 391138 941407
rect 390822 941351 390837 941391
rect 390946 941351 390979 941391
rect 391070 941351 391121 941391
rect 391194 941351 391248 941407
rect 389331 941335 389417 941351
rect 389473 941335 389559 941351
rect 389615 941335 389701 941351
rect 389757 941335 389843 941351
rect 389899 941335 389985 941351
rect 390041 941335 390127 941351
rect 390183 941335 390269 941351
rect 390325 941335 390411 941351
rect 390467 941335 390553 941351
rect 390609 941335 390695 941351
rect 390751 941335 390837 941351
rect 390893 941335 390979 941351
rect 391035 941335 391121 941351
rect 391177 941335 391248 941351
rect 389198 941283 391248 941335
rect 389198 941249 389278 941283
rect 389198 941193 389275 941249
rect 389334 941227 389402 941283
rect 389458 941249 389526 941283
rect 389582 941249 389650 941283
rect 389706 941249 389774 941283
rect 389473 941227 389526 941249
rect 389615 941227 389650 941249
rect 389757 941227 389774 941249
rect 389830 941249 389898 941283
rect 389954 941249 390022 941283
rect 390078 941249 390146 941283
rect 390202 941249 390270 941283
rect 389830 941227 389843 941249
rect 389954 941227 389985 941249
rect 390078 941227 390127 941249
rect 390202 941227 390269 941249
rect 390326 941227 390394 941283
rect 390450 941249 390518 941283
rect 390574 941249 390642 941283
rect 390698 941249 390766 941283
rect 390467 941227 390518 941249
rect 390609 941227 390642 941249
rect 390751 941227 390766 941249
rect 390822 941249 390890 941283
rect 390946 941249 391014 941283
rect 391070 941249 391138 941283
rect 390822 941227 390837 941249
rect 390946 941227 390979 941249
rect 391070 941227 391121 941249
rect 391194 941227 391248 941283
rect 389331 941193 389417 941227
rect 389473 941193 389559 941227
rect 389615 941193 389701 941227
rect 389757 941193 389843 941227
rect 389899 941193 389985 941227
rect 390041 941193 390127 941227
rect 390183 941193 390269 941227
rect 390325 941193 390411 941227
rect 390467 941193 390553 941227
rect 390609 941193 390695 941227
rect 390751 941193 390837 941227
rect 390893 941193 390979 941227
rect 391035 941193 391121 941227
rect 391177 941193 391248 941227
rect 389198 941159 391248 941193
rect 389198 941107 389278 941159
rect 389198 941051 389275 941107
rect 389334 941103 389402 941159
rect 389458 941107 389526 941159
rect 389582 941107 389650 941159
rect 389706 941107 389774 941159
rect 389473 941103 389526 941107
rect 389615 941103 389650 941107
rect 389757 941103 389774 941107
rect 389830 941107 389898 941159
rect 389954 941107 390022 941159
rect 390078 941107 390146 941159
rect 390202 941107 390270 941159
rect 389830 941103 389843 941107
rect 389954 941103 389985 941107
rect 390078 941103 390127 941107
rect 390202 941103 390269 941107
rect 390326 941103 390394 941159
rect 390450 941107 390518 941159
rect 390574 941107 390642 941159
rect 390698 941107 390766 941159
rect 390467 941103 390518 941107
rect 390609 941103 390642 941107
rect 390751 941103 390766 941107
rect 390822 941107 390890 941159
rect 390946 941107 391014 941159
rect 391070 941107 391138 941159
rect 390822 941103 390837 941107
rect 390946 941103 390979 941107
rect 391070 941103 391121 941107
rect 391194 941103 391248 941159
rect 389331 941051 389417 941103
rect 389473 941051 389559 941103
rect 389615 941051 389701 941103
rect 389757 941051 389843 941103
rect 389899 941051 389985 941103
rect 390041 941051 390127 941103
rect 390183 941051 390269 941103
rect 390325 941051 390411 941103
rect 390467 941051 390553 941103
rect 390609 941051 390695 941103
rect 390751 941051 390837 941103
rect 390893 941051 390979 941103
rect 391035 941051 391121 941103
rect 391177 941051 391248 941103
rect 389198 941035 391248 941051
rect 389198 940979 389278 941035
rect 389334 940979 389402 941035
rect 389458 940979 389526 941035
rect 389582 940979 389650 941035
rect 389706 940979 389774 941035
rect 389830 940979 389898 941035
rect 389954 940979 390022 941035
rect 390078 940979 390146 941035
rect 390202 940979 390270 941035
rect 390326 940979 390394 941035
rect 390450 940979 390518 941035
rect 390574 940979 390642 941035
rect 390698 940979 390766 941035
rect 390822 940979 390890 941035
rect 390946 940979 391014 941035
rect 391070 940979 391138 941035
rect 391194 940979 391248 941035
rect 389198 940965 391248 940979
rect 389198 940909 389275 940965
rect 389331 940911 389417 940965
rect 389473 940911 389559 940965
rect 389615 940911 389701 940965
rect 389757 940911 389843 940965
rect 389899 940911 389985 940965
rect 390041 940911 390127 940965
rect 390183 940911 390269 940965
rect 390325 940911 390411 940965
rect 390467 940911 390553 940965
rect 390609 940911 390695 940965
rect 390751 940911 390837 940965
rect 390893 940911 390979 940965
rect 391035 940911 391121 940965
rect 391177 940911 391248 940965
rect 389198 940855 389278 940909
rect 389334 940855 389402 940911
rect 389473 940909 389526 940911
rect 389615 940909 389650 940911
rect 389757 940909 389774 940911
rect 389458 940855 389526 940909
rect 389582 940855 389650 940909
rect 389706 940855 389774 940909
rect 389830 940909 389843 940911
rect 389954 940909 389985 940911
rect 390078 940909 390127 940911
rect 390202 940909 390269 940911
rect 389830 940855 389898 940909
rect 389954 940855 390022 940909
rect 390078 940855 390146 940909
rect 390202 940855 390270 940909
rect 390326 940855 390394 940911
rect 390467 940909 390518 940911
rect 390609 940909 390642 940911
rect 390751 940909 390766 940911
rect 390450 940855 390518 940909
rect 390574 940855 390642 940909
rect 390698 940855 390766 940909
rect 390822 940909 390837 940911
rect 390946 940909 390979 940911
rect 391070 940909 391121 940911
rect 390822 940855 390890 940909
rect 390946 940855 391014 940909
rect 391070 940855 391138 940909
rect 391194 940855 391248 940911
rect 389198 940823 391248 940855
rect 389198 940767 389275 940823
rect 389331 940787 389417 940823
rect 389473 940787 389559 940823
rect 389615 940787 389701 940823
rect 389757 940787 389843 940823
rect 389899 940787 389985 940823
rect 390041 940787 390127 940823
rect 390183 940787 390269 940823
rect 390325 940787 390411 940823
rect 390467 940787 390553 940823
rect 390609 940787 390695 940823
rect 390751 940787 390837 940823
rect 390893 940787 390979 940823
rect 391035 940787 391121 940823
rect 391177 940787 391248 940823
rect 389198 940731 389278 940767
rect 389334 940731 389402 940787
rect 389473 940767 389526 940787
rect 389615 940767 389650 940787
rect 389757 940767 389774 940787
rect 389458 940731 389526 940767
rect 389582 940731 389650 940767
rect 389706 940731 389774 940767
rect 389830 940767 389843 940787
rect 389954 940767 389985 940787
rect 390078 940767 390127 940787
rect 390202 940767 390269 940787
rect 389830 940731 389898 940767
rect 389954 940731 390022 940767
rect 390078 940731 390146 940767
rect 390202 940731 390270 940767
rect 390326 940731 390394 940787
rect 390467 940767 390518 940787
rect 390609 940767 390642 940787
rect 390751 940767 390766 940787
rect 390450 940731 390518 940767
rect 390574 940731 390642 940767
rect 390698 940731 390766 940767
rect 390822 940767 390837 940787
rect 390946 940767 390979 940787
rect 391070 940767 391121 940787
rect 390822 940731 390890 940767
rect 390946 940731 391014 940767
rect 391070 940731 391138 940767
rect 391194 940731 391248 940787
rect 389198 940681 391248 940731
rect 389198 940625 389275 940681
rect 389331 940663 389417 940681
rect 389473 940663 389559 940681
rect 389615 940663 389701 940681
rect 389757 940663 389843 940681
rect 389899 940663 389985 940681
rect 390041 940663 390127 940681
rect 390183 940663 390269 940681
rect 390325 940663 390411 940681
rect 390467 940663 390553 940681
rect 390609 940663 390695 940681
rect 390751 940663 390837 940681
rect 390893 940663 390979 940681
rect 391035 940663 391121 940681
rect 391177 940663 391248 940681
rect 389198 940607 389278 940625
rect 389334 940607 389402 940663
rect 389473 940625 389526 940663
rect 389615 940625 389650 940663
rect 389757 940625 389774 940663
rect 389458 940607 389526 940625
rect 389582 940607 389650 940625
rect 389706 940607 389774 940625
rect 389830 940625 389843 940663
rect 389954 940625 389985 940663
rect 390078 940625 390127 940663
rect 390202 940625 390269 940663
rect 389830 940607 389898 940625
rect 389954 940607 390022 940625
rect 390078 940607 390146 940625
rect 390202 940607 390270 940625
rect 390326 940607 390394 940663
rect 390467 940625 390518 940663
rect 390609 940625 390642 940663
rect 390751 940625 390766 940663
rect 390450 940607 390518 940625
rect 390574 940607 390642 940625
rect 390698 940607 390766 940625
rect 390822 940625 390837 940663
rect 390946 940625 390979 940663
rect 391070 940625 391121 940663
rect 390822 940607 390890 940625
rect 390946 940607 391014 940625
rect 391070 940607 391138 940625
rect 391194 940607 391248 940663
rect 389198 940539 391248 940607
rect 389198 940483 389275 940539
rect 389334 940483 389402 940539
rect 389473 940483 389526 940539
rect 389615 940483 389650 940539
rect 389757 940483 389774 940539
rect 389830 940483 389843 940539
rect 389954 940483 389985 940539
rect 390078 940483 390127 940539
rect 390202 940483 390269 940539
rect 390326 940483 390394 940539
rect 390467 940483 390518 940539
rect 390609 940483 390642 940539
rect 390751 940483 390766 940539
rect 390822 940483 390837 940539
rect 390946 940483 390979 940539
rect 391070 940483 391121 940539
rect 391194 940483 391248 940539
rect 389198 940415 391248 940483
rect 389198 940397 389278 940415
rect 389198 940341 389275 940397
rect 389334 940359 389402 940415
rect 389458 940397 389526 940415
rect 389582 940397 389650 940415
rect 389706 940397 389774 940415
rect 389473 940359 389526 940397
rect 389615 940359 389650 940397
rect 389757 940359 389774 940397
rect 389830 940397 389898 940415
rect 389954 940397 390022 940415
rect 390078 940397 390146 940415
rect 390202 940397 390270 940415
rect 389830 940359 389843 940397
rect 389954 940359 389985 940397
rect 390078 940359 390127 940397
rect 390202 940359 390269 940397
rect 390326 940359 390394 940415
rect 390450 940397 390518 940415
rect 390574 940397 390642 940415
rect 390698 940397 390766 940415
rect 390467 940359 390518 940397
rect 390609 940359 390642 940397
rect 390751 940359 390766 940397
rect 390822 940397 390890 940415
rect 390946 940397 391014 940415
rect 391070 940397 391138 940415
rect 390822 940359 390837 940397
rect 390946 940359 390979 940397
rect 391070 940359 391121 940397
rect 391194 940359 391248 940415
rect 389331 940341 389417 940359
rect 389473 940341 389559 940359
rect 389615 940341 389701 940359
rect 389757 940341 389843 940359
rect 389899 940341 389985 940359
rect 390041 940341 390127 940359
rect 390183 940341 390269 940359
rect 390325 940341 390411 940359
rect 390467 940341 390553 940359
rect 390609 940341 390695 940359
rect 390751 940341 390837 940359
rect 390893 940341 390979 940359
rect 391035 940341 391121 940359
rect 391177 940341 391248 940359
rect 389198 940291 391248 940341
rect 389198 940255 389278 940291
rect 389198 940199 389275 940255
rect 389334 940235 389402 940291
rect 389458 940255 389526 940291
rect 389582 940255 389650 940291
rect 389706 940255 389774 940291
rect 389473 940235 389526 940255
rect 389615 940235 389650 940255
rect 389757 940235 389774 940255
rect 389830 940255 389898 940291
rect 389954 940255 390022 940291
rect 390078 940255 390146 940291
rect 390202 940255 390270 940291
rect 389830 940235 389843 940255
rect 389954 940235 389985 940255
rect 390078 940235 390127 940255
rect 390202 940235 390269 940255
rect 390326 940235 390394 940291
rect 390450 940255 390518 940291
rect 390574 940255 390642 940291
rect 390698 940255 390766 940291
rect 390467 940235 390518 940255
rect 390609 940235 390642 940255
rect 390751 940235 390766 940255
rect 390822 940255 390890 940291
rect 390946 940255 391014 940291
rect 391070 940255 391138 940291
rect 390822 940235 390837 940255
rect 390946 940235 390979 940255
rect 391070 940235 391121 940255
rect 391194 940235 391248 940291
rect 389331 940199 389417 940235
rect 389473 940199 389559 940235
rect 389615 940199 389701 940235
rect 389757 940199 389843 940235
rect 389899 940199 389985 940235
rect 390041 940199 390127 940235
rect 390183 940199 390269 940235
rect 390325 940199 390411 940235
rect 390467 940199 390553 940235
rect 390609 940199 390695 940235
rect 390751 940199 390837 940235
rect 390893 940199 390979 940235
rect 391035 940199 391121 940235
rect 391177 940199 391248 940235
rect 389198 940167 391248 940199
rect 389198 940113 389278 940167
rect 389198 940057 389275 940113
rect 389334 940111 389402 940167
rect 389458 940113 389526 940167
rect 389582 940113 389650 940167
rect 389706 940113 389774 940167
rect 389473 940111 389526 940113
rect 389615 940111 389650 940113
rect 389757 940111 389774 940113
rect 389830 940113 389898 940167
rect 389954 940113 390022 940167
rect 390078 940113 390146 940167
rect 390202 940113 390270 940167
rect 389830 940111 389843 940113
rect 389954 940111 389985 940113
rect 390078 940111 390127 940113
rect 390202 940111 390269 940113
rect 390326 940111 390394 940167
rect 390450 940113 390518 940167
rect 390574 940113 390642 940167
rect 390698 940113 390766 940167
rect 390467 940111 390518 940113
rect 390609 940111 390642 940113
rect 390751 940111 390766 940113
rect 390822 940113 390890 940167
rect 390946 940113 391014 940167
rect 391070 940113 391138 940167
rect 390822 940111 390837 940113
rect 390946 940111 390979 940113
rect 391070 940111 391121 940113
rect 391194 940111 391248 940167
rect 389331 940057 389417 940111
rect 389473 940057 389559 940111
rect 389615 940057 389701 940111
rect 389757 940057 389843 940111
rect 389899 940057 389985 940111
rect 390041 940057 390127 940111
rect 390183 940057 390269 940111
rect 390325 940057 390411 940111
rect 390467 940057 390553 940111
rect 390609 940057 390695 940111
rect 390751 940057 390837 940111
rect 390893 940057 390979 940111
rect 391035 940057 391121 940111
rect 391177 940057 391248 940111
rect 389198 940043 391248 940057
rect 389198 939987 389278 940043
rect 389334 939987 389402 940043
rect 389458 939987 389526 940043
rect 389582 939987 389650 940043
rect 389706 939987 389774 940043
rect 389830 939987 389898 940043
rect 389954 939987 390022 940043
rect 390078 939987 390146 940043
rect 390202 939987 390270 940043
rect 390326 939987 390394 940043
rect 390450 939987 390518 940043
rect 390574 939987 390642 940043
rect 390698 939987 390766 940043
rect 390822 939987 390890 940043
rect 390946 939987 391014 940043
rect 391070 939987 391138 940043
rect 391194 939987 391248 940043
rect 389198 939971 391248 939987
rect 389198 939915 389275 939971
rect 389331 939919 389417 939971
rect 389473 939919 389559 939971
rect 389615 939919 389701 939971
rect 389757 939919 389843 939971
rect 389899 939919 389985 939971
rect 390041 939919 390127 939971
rect 390183 939919 390269 939971
rect 390325 939919 390411 939971
rect 390467 939919 390553 939971
rect 390609 939919 390695 939971
rect 390751 939919 390837 939971
rect 390893 939919 390979 939971
rect 391035 939919 391121 939971
rect 391177 939919 391248 939971
rect 389198 939863 389278 939915
rect 389334 939863 389402 939919
rect 389473 939915 389526 939919
rect 389615 939915 389650 939919
rect 389757 939915 389774 939919
rect 389458 939863 389526 939915
rect 389582 939863 389650 939915
rect 389706 939863 389774 939915
rect 389830 939915 389843 939919
rect 389954 939915 389985 939919
rect 390078 939915 390127 939919
rect 390202 939915 390269 939919
rect 389830 939863 389898 939915
rect 389954 939863 390022 939915
rect 390078 939863 390146 939915
rect 390202 939863 390270 939915
rect 390326 939863 390394 939919
rect 390467 939915 390518 939919
rect 390609 939915 390642 939919
rect 390751 939915 390766 939919
rect 390450 939863 390518 939915
rect 390574 939863 390642 939915
rect 390698 939863 390766 939915
rect 390822 939915 390837 939919
rect 390946 939915 390979 939919
rect 391070 939915 391121 939919
rect 390822 939863 390890 939915
rect 390946 939863 391014 939915
rect 391070 939863 391138 939915
rect 391194 939863 391248 939919
rect 389198 939829 391248 939863
rect 389198 939773 389275 939829
rect 389331 939773 389417 939829
rect 389473 939773 389559 939829
rect 389615 939773 389701 939829
rect 389757 939773 389843 939829
rect 389899 939773 389985 939829
rect 390041 939773 390127 939829
rect 390183 939773 390269 939829
rect 390325 939773 390411 939829
rect 390467 939773 390553 939829
rect 390609 939773 390695 939829
rect 390751 939773 390837 939829
rect 390893 939773 390979 939829
rect 391035 939773 391121 939829
rect 391177 939773 391248 939829
rect 389198 939720 391248 939773
rect 391828 941675 393728 941720
rect 391828 941655 391897 941675
rect 391953 941655 392039 941675
rect 392095 941655 392181 941675
rect 392237 941655 392323 941675
rect 392379 941655 392465 941675
rect 392521 941655 392607 941675
rect 392663 941655 392749 941675
rect 392805 941655 392891 941675
rect 392947 941655 393033 941675
rect 393089 941655 393175 941675
rect 393231 941655 393317 941675
rect 393373 941655 393459 941675
rect 393515 941655 393601 941675
rect 393657 941655 393728 941675
rect 391828 941599 391882 941655
rect 391953 941619 392006 941655
rect 392095 941619 392130 941655
rect 392237 941619 392254 941655
rect 391938 941599 392006 941619
rect 392062 941599 392130 941619
rect 392186 941599 392254 941619
rect 392310 941619 392323 941655
rect 392434 941619 392465 941655
rect 392558 941619 392607 941655
rect 392682 941619 392749 941655
rect 392310 941599 392378 941619
rect 392434 941599 392502 941619
rect 392558 941599 392626 941619
rect 392682 941599 392750 941619
rect 392806 941599 392874 941655
rect 392947 941619 392998 941655
rect 393089 941619 393122 941655
rect 393231 941619 393246 941655
rect 392930 941599 392998 941619
rect 393054 941599 393122 941619
rect 393178 941599 393246 941619
rect 393302 941619 393317 941655
rect 393426 941619 393459 941655
rect 393550 941619 393601 941655
rect 393302 941599 393370 941619
rect 393426 941599 393494 941619
rect 393550 941599 393618 941619
rect 393674 941599 393728 941655
rect 391828 941533 393728 941599
rect 391828 941531 391897 941533
rect 391953 941531 392039 941533
rect 392095 941531 392181 941533
rect 392237 941531 392323 941533
rect 392379 941531 392465 941533
rect 392521 941531 392607 941533
rect 392663 941531 392749 941533
rect 392805 941531 392891 941533
rect 392947 941531 393033 941533
rect 393089 941531 393175 941533
rect 393231 941531 393317 941533
rect 393373 941531 393459 941533
rect 393515 941531 393601 941533
rect 393657 941531 393728 941533
rect 391828 941475 391882 941531
rect 391953 941477 392006 941531
rect 392095 941477 392130 941531
rect 392237 941477 392254 941531
rect 391938 941475 392006 941477
rect 392062 941475 392130 941477
rect 392186 941475 392254 941477
rect 392310 941477 392323 941531
rect 392434 941477 392465 941531
rect 392558 941477 392607 941531
rect 392682 941477 392749 941531
rect 392310 941475 392378 941477
rect 392434 941475 392502 941477
rect 392558 941475 392626 941477
rect 392682 941475 392750 941477
rect 392806 941475 392874 941531
rect 392947 941477 392998 941531
rect 393089 941477 393122 941531
rect 393231 941477 393246 941531
rect 392930 941475 392998 941477
rect 393054 941475 393122 941477
rect 393178 941475 393246 941477
rect 393302 941477 393317 941531
rect 393426 941477 393459 941531
rect 393550 941477 393601 941531
rect 393302 941475 393370 941477
rect 393426 941475 393494 941477
rect 393550 941475 393618 941477
rect 393674 941475 393728 941531
rect 391828 941407 393728 941475
rect 391828 941351 391882 941407
rect 391938 941391 392006 941407
rect 392062 941391 392130 941407
rect 392186 941391 392254 941407
rect 391953 941351 392006 941391
rect 392095 941351 392130 941391
rect 392237 941351 392254 941391
rect 392310 941391 392378 941407
rect 392434 941391 392502 941407
rect 392558 941391 392626 941407
rect 392682 941391 392750 941407
rect 392310 941351 392323 941391
rect 392434 941351 392465 941391
rect 392558 941351 392607 941391
rect 392682 941351 392749 941391
rect 392806 941351 392874 941407
rect 392930 941391 392998 941407
rect 393054 941391 393122 941407
rect 393178 941391 393246 941407
rect 392947 941351 392998 941391
rect 393089 941351 393122 941391
rect 393231 941351 393246 941391
rect 393302 941391 393370 941407
rect 393426 941391 393494 941407
rect 393550 941391 393618 941407
rect 393302 941351 393317 941391
rect 393426 941351 393459 941391
rect 393550 941351 393601 941391
rect 393674 941351 393728 941407
rect 391828 941335 391897 941351
rect 391953 941335 392039 941351
rect 392095 941335 392181 941351
rect 392237 941335 392323 941351
rect 392379 941335 392465 941351
rect 392521 941335 392607 941351
rect 392663 941335 392749 941351
rect 392805 941335 392891 941351
rect 392947 941335 393033 941351
rect 393089 941335 393175 941351
rect 393231 941335 393317 941351
rect 393373 941335 393459 941351
rect 393515 941335 393601 941351
rect 393657 941335 393728 941351
rect 391828 941283 393728 941335
rect 391828 941227 391882 941283
rect 391938 941249 392006 941283
rect 392062 941249 392130 941283
rect 392186 941249 392254 941283
rect 391953 941227 392006 941249
rect 392095 941227 392130 941249
rect 392237 941227 392254 941249
rect 392310 941249 392378 941283
rect 392434 941249 392502 941283
rect 392558 941249 392626 941283
rect 392682 941249 392750 941283
rect 392310 941227 392323 941249
rect 392434 941227 392465 941249
rect 392558 941227 392607 941249
rect 392682 941227 392749 941249
rect 392806 941227 392874 941283
rect 392930 941249 392998 941283
rect 393054 941249 393122 941283
rect 393178 941249 393246 941283
rect 392947 941227 392998 941249
rect 393089 941227 393122 941249
rect 393231 941227 393246 941249
rect 393302 941249 393370 941283
rect 393426 941249 393494 941283
rect 393550 941249 393618 941283
rect 393302 941227 393317 941249
rect 393426 941227 393459 941249
rect 393550 941227 393601 941249
rect 393674 941227 393728 941283
rect 391828 941193 391897 941227
rect 391953 941193 392039 941227
rect 392095 941193 392181 941227
rect 392237 941193 392323 941227
rect 392379 941193 392465 941227
rect 392521 941193 392607 941227
rect 392663 941193 392749 941227
rect 392805 941193 392891 941227
rect 392947 941193 393033 941227
rect 393089 941193 393175 941227
rect 393231 941193 393317 941227
rect 393373 941193 393459 941227
rect 393515 941193 393601 941227
rect 393657 941193 393728 941227
rect 391828 941159 393728 941193
rect 391828 941103 391882 941159
rect 391938 941107 392006 941159
rect 392062 941107 392130 941159
rect 392186 941107 392254 941159
rect 391953 941103 392006 941107
rect 392095 941103 392130 941107
rect 392237 941103 392254 941107
rect 392310 941107 392378 941159
rect 392434 941107 392502 941159
rect 392558 941107 392626 941159
rect 392682 941107 392750 941159
rect 392310 941103 392323 941107
rect 392434 941103 392465 941107
rect 392558 941103 392607 941107
rect 392682 941103 392749 941107
rect 392806 941103 392874 941159
rect 392930 941107 392998 941159
rect 393054 941107 393122 941159
rect 393178 941107 393246 941159
rect 392947 941103 392998 941107
rect 393089 941103 393122 941107
rect 393231 941103 393246 941107
rect 393302 941107 393370 941159
rect 393426 941107 393494 941159
rect 393550 941107 393618 941159
rect 393302 941103 393317 941107
rect 393426 941103 393459 941107
rect 393550 941103 393601 941107
rect 393674 941103 393728 941159
rect 391828 941051 391897 941103
rect 391953 941051 392039 941103
rect 392095 941051 392181 941103
rect 392237 941051 392323 941103
rect 392379 941051 392465 941103
rect 392521 941051 392607 941103
rect 392663 941051 392749 941103
rect 392805 941051 392891 941103
rect 392947 941051 393033 941103
rect 393089 941051 393175 941103
rect 393231 941051 393317 941103
rect 393373 941051 393459 941103
rect 393515 941051 393601 941103
rect 393657 941051 393728 941103
rect 391828 941035 393728 941051
rect 391828 940979 391882 941035
rect 391938 940979 392006 941035
rect 392062 940979 392130 941035
rect 392186 940979 392254 941035
rect 392310 940979 392378 941035
rect 392434 940979 392502 941035
rect 392558 940979 392626 941035
rect 392682 940979 392750 941035
rect 392806 940979 392874 941035
rect 392930 940979 392998 941035
rect 393054 940979 393122 941035
rect 393178 940979 393246 941035
rect 393302 940979 393370 941035
rect 393426 940979 393494 941035
rect 393550 940979 393618 941035
rect 393674 940979 393728 941035
rect 391828 940965 393728 940979
rect 391828 940911 391897 940965
rect 391953 940911 392039 940965
rect 392095 940911 392181 940965
rect 392237 940911 392323 940965
rect 392379 940911 392465 940965
rect 392521 940911 392607 940965
rect 392663 940911 392749 940965
rect 392805 940911 392891 940965
rect 392947 940911 393033 940965
rect 393089 940911 393175 940965
rect 393231 940911 393317 940965
rect 393373 940911 393459 940965
rect 393515 940911 393601 940965
rect 393657 940911 393728 940965
rect 391828 940855 391882 940911
rect 391953 940909 392006 940911
rect 392095 940909 392130 940911
rect 392237 940909 392254 940911
rect 391938 940855 392006 940909
rect 392062 940855 392130 940909
rect 392186 940855 392254 940909
rect 392310 940909 392323 940911
rect 392434 940909 392465 940911
rect 392558 940909 392607 940911
rect 392682 940909 392749 940911
rect 392310 940855 392378 940909
rect 392434 940855 392502 940909
rect 392558 940855 392626 940909
rect 392682 940855 392750 940909
rect 392806 940855 392874 940911
rect 392947 940909 392998 940911
rect 393089 940909 393122 940911
rect 393231 940909 393246 940911
rect 392930 940855 392998 940909
rect 393054 940855 393122 940909
rect 393178 940855 393246 940909
rect 393302 940909 393317 940911
rect 393426 940909 393459 940911
rect 393550 940909 393601 940911
rect 393302 940855 393370 940909
rect 393426 940855 393494 940909
rect 393550 940855 393618 940909
rect 393674 940855 393728 940911
rect 391828 940823 393728 940855
rect 391828 940787 391897 940823
rect 391953 940787 392039 940823
rect 392095 940787 392181 940823
rect 392237 940787 392323 940823
rect 392379 940787 392465 940823
rect 392521 940787 392607 940823
rect 392663 940787 392749 940823
rect 392805 940787 392891 940823
rect 392947 940787 393033 940823
rect 393089 940787 393175 940823
rect 393231 940787 393317 940823
rect 393373 940787 393459 940823
rect 393515 940787 393601 940823
rect 393657 940787 393728 940823
rect 391828 940731 391882 940787
rect 391953 940767 392006 940787
rect 392095 940767 392130 940787
rect 392237 940767 392254 940787
rect 391938 940731 392006 940767
rect 392062 940731 392130 940767
rect 392186 940731 392254 940767
rect 392310 940767 392323 940787
rect 392434 940767 392465 940787
rect 392558 940767 392607 940787
rect 392682 940767 392749 940787
rect 392310 940731 392378 940767
rect 392434 940731 392502 940767
rect 392558 940731 392626 940767
rect 392682 940731 392750 940767
rect 392806 940731 392874 940787
rect 392947 940767 392998 940787
rect 393089 940767 393122 940787
rect 393231 940767 393246 940787
rect 392930 940731 392998 940767
rect 393054 940731 393122 940767
rect 393178 940731 393246 940767
rect 393302 940767 393317 940787
rect 393426 940767 393459 940787
rect 393550 940767 393601 940787
rect 393302 940731 393370 940767
rect 393426 940731 393494 940767
rect 393550 940731 393618 940767
rect 393674 940731 393728 940787
rect 391828 940681 393728 940731
rect 391828 940663 391897 940681
rect 391953 940663 392039 940681
rect 392095 940663 392181 940681
rect 392237 940663 392323 940681
rect 392379 940663 392465 940681
rect 392521 940663 392607 940681
rect 392663 940663 392749 940681
rect 392805 940663 392891 940681
rect 392947 940663 393033 940681
rect 393089 940663 393175 940681
rect 393231 940663 393317 940681
rect 393373 940663 393459 940681
rect 393515 940663 393601 940681
rect 393657 940663 393728 940681
rect 391828 940607 391882 940663
rect 391953 940625 392006 940663
rect 392095 940625 392130 940663
rect 392237 940625 392254 940663
rect 391938 940607 392006 940625
rect 392062 940607 392130 940625
rect 392186 940607 392254 940625
rect 392310 940625 392323 940663
rect 392434 940625 392465 940663
rect 392558 940625 392607 940663
rect 392682 940625 392749 940663
rect 392310 940607 392378 940625
rect 392434 940607 392502 940625
rect 392558 940607 392626 940625
rect 392682 940607 392750 940625
rect 392806 940607 392874 940663
rect 392947 940625 392998 940663
rect 393089 940625 393122 940663
rect 393231 940625 393246 940663
rect 392930 940607 392998 940625
rect 393054 940607 393122 940625
rect 393178 940607 393246 940625
rect 393302 940625 393317 940663
rect 393426 940625 393459 940663
rect 393550 940625 393601 940663
rect 393302 940607 393370 940625
rect 393426 940607 393494 940625
rect 393550 940607 393618 940625
rect 393674 940607 393728 940663
rect 391828 940539 393728 940607
rect 391828 940483 391882 940539
rect 391953 940483 392006 940539
rect 392095 940483 392130 940539
rect 392237 940483 392254 940539
rect 392310 940483 392323 940539
rect 392434 940483 392465 940539
rect 392558 940483 392607 940539
rect 392682 940483 392749 940539
rect 392806 940483 392874 940539
rect 392947 940483 392998 940539
rect 393089 940483 393122 940539
rect 393231 940483 393246 940539
rect 393302 940483 393317 940539
rect 393426 940483 393459 940539
rect 393550 940483 393601 940539
rect 393674 940483 393728 940539
rect 391828 940415 393728 940483
rect 391828 940359 391882 940415
rect 391938 940397 392006 940415
rect 392062 940397 392130 940415
rect 392186 940397 392254 940415
rect 391953 940359 392006 940397
rect 392095 940359 392130 940397
rect 392237 940359 392254 940397
rect 392310 940397 392378 940415
rect 392434 940397 392502 940415
rect 392558 940397 392626 940415
rect 392682 940397 392750 940415
rect 392310 940359 392323 940397
rect 392434 940359 392465 940397
rect 392558 940359 392607 940397
rect 392682 940359 392749 940397
rect 392806 940359 392874 940415
rect 392930 940397 392998 940415
rect 393054 940397 393122 940415
rect 393178 940397 393246 940415
rect 392947 940359 392998 940397
rect 393089 940359 393122 940397
rect 393231 940359 393246 940397
rect 393302 940397 393370 940415
rect 393426 940397 393494 940415
rect 393550 940397 393618 940415
rect 393302 940359 393317 940397
rect 393426 940359 393459 940397
rect 393550 940359 393601 940397
rect 393674 940359 393728 940415
rect 391828 940341 391897 940359
rect 391953 940341 392039 940359
rect 392095 940341 392181 940359
rect 392237 940341 392323 940359
rect 392379 940341 392465 940359
rect 392521 940341 392607 940359
rect 392663 940341 392749 940359
rect 392805 940341 392891 940359
rect 392947 940341 393033 940359
rect 393089 940341 393175 940359
rect 393231 940341 393317 940359
rect 393373 940341 393459 940359
rect 393515 940341 393601 940359
rect 393657 940341 393728 940359
rect 391828 940291 393728 940341
rect 391828 940235 391882 940291
rect 391938 940255 392006 940291
rect 392062 940255 392130 940291
rect 392186 940255 392254 940291
rect 391953 940235 392006 940255
rect 392095 940235 392130 940255
rect 392237 940235 392254 940255
rect 392310 940255 392378 940291
rect 392434 940255 392502 940291
rect 392558 940255 392626 940291
rect 392682 940255 392750 940291
rect 392310 940235 392323 940255
rect 392434 940235 392465 940255
rect 392558 940235 392607 940255
rect 392682 940235 392749 940255
rect 392806 940235 392874 940291
rect 392930 940255 392998 940291
rect 393054 940255 393122 940291
rect 393178 940255 393246 940291
rect 392947 940235 392998 940255
rect 393089 940235 393122 940255
rect 393231 940235 393246 940255
rect 393302 940255 393370 940291
rect 393426 940255 393494 940291
rect 393550 940255 393618 940291
rect 393302 940235 393317 940255
rect 393426 940235 393459 940255
rect 393550 940235 393601 940255
rect 393674 940235 393728 940291
rect 391828 940199 391897 940235
rect 391953 940199 392039 940235
rect 392095 940199 392181 940235
rect 392237 940199 392323 940235
rect 392379 940199 392465 940235
rect 392521 940199 392607 940235
rect 392663 940199 392749 940235
rect 392805 940199 392891 940235
rect 392947 940199 393033 940235
rect 393089 940199 393175 940235
rect 393231 940199 393317 940235
rect 393373 940199 393459 940235
rect 393515 940199 393601 940235
rect 393657 940199 393728 940235
rect 391828 940167 393728 940199
rect 391828 940111 391882 940167
rect 391938 940113 392006 940167
rect 392062 940113 392130 940167
rect 392186 940113 392254 940167
rect 391953 940111 392006 940113
rect 392095 940111 392130 940113
rect 392237 940111 392254 940113
rect 392310 940113 392378 940167
rect 392434 940113 392502 940167
rect 392558 940113 392626 940167
rect 392682 940113 392750 940167
rect 392310 940111 392323 940113
rect 392434 940111 392465 940113
rect 392558 940111 392607 940113
rect 392682 940111 392749 940113
rect 392806 940111 392874 940167
rect 392930 940113 392998 940167
rect 393054 940113 393122 940167
rect 393178 940113 393246 940167
rect 392947 940111 392998 940113
rect 393089 940111 393122 940113
rect 393231 940111 393246 940113
rect 393302 940113 393370 940167
rect 393426 940113 393494 940167
rect 393550 940113 393618 940167
rect 393302 940111 393317 940113
rect 393426 940111 393459 940113
rect 393550 940111 393601 940113
rect 393674 940111 393728 940167
rect 391828 940057 391897 940111
rect 391953 940057 392039 940111
rect 392095 940057 392181 940111
rect 392237 940057 392323 940111
rect 392379 940057 392465 940111
rect 392521 940057 392607 940111
rect 392663 940057 392749 940111
rect 392805 940057 392891 940111
rect 392947 940057 393033 940111
rect 393089 940057 393175 940111
rect 393231 940057 393317 940111
rect 393373 940057 393459 940111
rect 393515 940057 393601 940111
rect 393657 940057 393728 940111
rect 391828 940043 393728 940057
rect 391828 939987 391882 940043
rect 391938 939987 392006 940043
rect 392062 939987 392130 940043
rect 392186 939987 392254 940043
rect 392310 939987 392378 940043
rect 392434 939987 392502 940043
rect 392558 939987 392626 940043
rect 392682 939987 392750 940043
rect 392806 939987 392874 940043
rect 392930 939987 392998 940043
rect 393054 939987 393122 940043
rect 393178 939987 393246 940043
rect 393302 939987 393370 940043
rect 393426 939987 393494 940043
rect 393550 939987 393618 940043
rect 393674 939987 393728 940043
rect 391828 939971 393728 939987
rect 391828 939919 391897 939971
rect 391953 939919 392039 939971
rect 392095 939919 392181 939971
rect 392237 939919 392323 939971
rect 392379 939919 392465 939971
rect 392521 939919 392607 939971
rect 392663 939919 392749 939971
rect 392805 939919 392891 939971
rect 392947 939919 393033 939971
rect 393089 939919 393175 939971
rect 393231 939919 393317 939971
rect 393373 939919 393459 939971
rect 393515 939919 393601 939971
rect 393657 939919 393728 939971
rect 391828 939863 391882 939919
rect 391953 939915 392006 939919
rect 392095 939915 392130 939919
rect 392237 939915 392254 939919
rect 391938 939863 392006 939915
rect 392062 939863 392130 939915
rect 392186 939863 392254 939915
rect 392310 939915 392323 939919
rect 392434 939915 392465 939919
rect 392558 939915 392607 939919
rect 392682 939915 392749 939919
rect 392310 939863 392378 939915
rect 392434 939863 392502 939915
rect 392558 939863 392626 939915
rect 392682 939863 392750 939915
rect 392806 939863 392874 939919
rect 392947 939915 392998 939919
rect 393089 939915 393122 939919
rect 393231 939915 393246 939919
rect 392930 939863 392998 939915
rect 393054 939863 393122 939915
rect 393178 939863 393246 939915
rect 393302 939915 393317 939919
rect 393426 939915 393459 939919
rect 393550 939915 393601 939919
rect 393302 939863 393370 939915
rect 393426 939863 393494 939915
rect 393550 939863 393618 939915
rect 393674 939863 393728 939919
rect 391828 939829 393728 939863
rect 391828 939773 391897 939829
rect 391953 939773 392039 939829
rect 392095 939773 392181 939829
rect 392237 939773 392323 939829
rect 392379 939773 392465 939829
rect 392521 939773 392607 939829
rect 392663 939773 392749 939829
rect 392805 939773 392891 939829
rect 392947 939773 393033 939829
rect 393089 939773 393175 939829
rect 393231 939773 393317 939829
rect 393373 939773 393459 939829
rect 393515 939773 393601 939829
rect 393657 939773 393728 939829
rect 391828 939720 393728 939773
rect 599272 941675 601172 941720
rect 599272 941655 599341 941675
rect 599397 941655 599483 941675
rect 599539 941655 599625 941675
rect 599681 941655 599767 941675
rect 599823 941655 599909 941675
rect 599965 941655 600051 941675
rect 600107 941655 600193 941675
rect 600249 941655 600335 941675
rect 600391 941655 600477 941675
rect 600533 941655 600619 941675
rect 600675 941655 600761 941675
rect 600817 941655 600903 941675
rect 600959 941655 601045 941675
rect 601101 941655 601172 941675
rect 599272 941599 599326 941655
rect 599397 941619 599450 941655
rect 599539 941619 599574 941655
rect 599681 941619 599698 941655
rect 599382 941599 599450 941619
rect 599506 941599 599574 941619
rect 599630 941599 599698 941619
rect 599754 941619 599767 941655
rect 599878 941619 599909 941655
rect 600002 941619 600051 941655
rect 600126 941619 600193 941655
rect 599754 941599 599822 941619
rect 599878 941599 599946 941619
rect 600002 941599 600070 941619
rect 600126 941599 600194 941619
rect 600250 941599 600318 941655
rect 600391 941619 600442 941655
rect 600533 941619 600566 941655
rect 600675 941619 600690 941655
rect 600374 941599 600442 941619
rect 600498 941599 600566 941619
rect 600622 941599 600690 941619
rect 600746 941619 600761 941655
rect 600870 941619 600903 941655
rect 600994 941619 601045 941655
rect 600746 941599 600814 941619
rect 600870 941599 600938 941619
rect 600994 941599 601062 941619
rect 601118 941599 601172 941655
rect 599272 941533 601172 941599
rect 599272 941531 599341 941533
rect 599397 941531 599483 941533
rect 599539 941531 599625 941533
rect 599681 941531 599767 941533
rect 599823 941531 599909 941533
rect 599965 941531 600051 941533
rect 600107 941531 600193 941533
rect 600249 941531 600335 941533
rect 600391 941531 600477 941533
rect 600533 941531 600619 941533
rect 600675 941531 600761 941533
rect 600817 941531 600903 941533
rect 600959 941531 601045 941533
rect 601101 941531 601172 941533
rect 599272 941475 599326 941531
rect 599397 941477 599450 941531
rect 599539 941477 599574 941531
rect 599681 941477 599698 941531
rect 599382 941475 599450 941477
rect 599506 941475 599574 941477
rect 599630 941475 599698 941477
rect 599754 941477 599767 941531
rect 599878 941477 599909 941531
rect 600002 941477 600051 941531
rect 600126 941477 600193 941531
rect 599754 941475 599822 941477
rect 599878 941475 599946 941477
rect 600002 941475 600070 941477
rect 600126 941475 600194 941477
rect 600250 941475 600318 941531
rect 600391 941477 600442 941531
rect 600533 941477 600566 941531
rect 600675 941477 600690 941531
rect 600374 941475 600442 941477
rect 600498 941475 600566 941477
rect 600622 941475 600690 941477
rect 600746 941477 600761 941531
rect 600870 941477 600903 941531
rect 600994 941477 601045 941531
rect 600746 941475 600814 941477
rect 600870 941475 600938 941477
rect 600994 941475 601062 941477
rect 601118 941475 601172 941531
rect 599272 941407 601172 941475
rect 599272 941351 599326 941407
rect 599382 941391 599450 941407
rect 599506 941391 599574 941407
rect 599630 941391 599698 941407
rect 599397 941351 599450 941391
rect 599539 941351 599574 941391
rect 599681 941351 599698 941391
rect 599754 941391 599822 941407
rect 599878 941391 599946 941407
rect 600002 941391 600070 941407
rect 600126 941391 600194 941407
rect 599754 941351 599767 941391
rect 599878 941351 599909 941391
rect 600002 941351 600051 941391
rect 600126 941351 600193 941391
rect 600250 941351 600318 941407
rect 600374 941391 600442 941407
rect 600498 941391 600566 941407
rect 600622 941391 600690 941407
rect 600391 941351 600442 941391
rect 600533 941351 600566 941391
rect 600675 941351 600690 941391
rect 600746 941391 600814 941407
rect 600870 941391 600938 941407
rect 600994 941391 601062 941407
rect 600746 941351 600761 941391
rect 600870 941351 600903 941391
rect 600994 941351 601045 941391
rect 601118 941351 601172 941407
rect 599272 941335 599341 941351
rect 599397 941335 599483 941351
rect 599539 941335 599625 941351
rect 599681 941335 599767 941351
rect 599823 941335 599909 941351
rect 599965 941335 600051 941351
rect 600107 941335 600193 941351
rect 600249 941335 600335 941351
rect 600391 941335 600477 941351
rect 600533 941335 600619 941351
rect 600675 941335 600761 941351
rect 600817 941335 600903 941351
rect 600959 941335 601045 941351
rect 601101 941335 601172 941351
rect 599272 941283 601172 941335
rect 599272 941227 599326 941283
rect 599382 941249 599450 941283
rect 599506 941249 599574 941283
rect 599630 941249 599698 941283
rect 599397 941227 599450 941249
rect 599539 941227 599574 941249
rect 599681 941227 599698 941249
rect 599754 941249 599822 941283
rect 599878 941249 599946 941283
rect 600002 941249 600070 941283
rect 600126 941249 600194 941283
rect 599754 941227 599767 941249
rect 599878 941227 599909 941249
rect 600002 941227 600051 941249
rect 600126 941227 600193 941249
rect 600250 941227 600318 941283
rect 600374 941249 600442 941283
rect 600498 941249 600566 941283
rect 600622 941249 600690 941283
rect 600391 941227 600442 941249
rect 600533 941227 600566 941249
rect 600675 941227 600690 941249
rect 600746 941249 600814 941283
rect 600870 941249 600938 941283
rect 600994 941249 601062 941283
rect 600746 941227 600761 941249
rect 600870 941227 600903 941249
rect 600994 941227 601045 941249
rect 601118 941227 601172 941283
rect 599272 941193 599341 941227
rect 599397 941193 599483 941227
rect 599539 941193 599625 941227
rect 599681 941193 599767 941227
rect 599823 941193 599909 941227
rect 599965 941193 600051 941227
rect 600107 941193 600193 941227
rect 600249 941193 600335 941227
rect 600391 941193 600477 941227
rect 600533 941193 600619 941227
rect 600675 941193 600761 941227
rect 600817 941193 600903 941227
rect 600959 941193 601045 941227
rect 601101 941193 601172 941227
rect 599272 941159 601172 941193
rect 599272 941103 599326 941159
rect 599382 941107 599450 941159
rect 599506 941107 599574 941159
rect 599630 941107 599698 941159
rect 599397 941103 599450 941107
rect 599539 941103 599574 941107
rect 599681 941103 599698 941107
rect 599754 941107 599822 941159
rect 599878 941107 599946 941159
rect 600002 941107 600070 941159
rect 600126 941107 600194 941159
rect 599754 941103 599767 941107
rect 599878 941103 599909 941107
rect 600002 941103 600051 941107
rect 600126 941103 600193 941107
rect 600250 941103 600318 941159
rect 600374 941107 600442 941159
rect 600498 941107 600566 941159
rect 600622 941107 600690 941159
rect 600391 941103 600442 941107
rect 600533 941103 600566 941107
rect 600675 941103 600690 941107
rect 600746 941107 600814 941159
rect 600870 941107 600938 941159
rect 600994 941107 601062 941159
rect 600746 941103 600761 941107
rect 600870 941103 600903 941107
rect 600994 941103 601045 941107
rect 601118 941103 601172 941159
rect 599272 941051 599341 941103
rect 599397 941051 599483 941103
rect 599539 941051 599625 941103
rect 599681 941051 599767 941103
rect 599823 941051 599909 941103
rect 599965 941051 600051 941103
rect 600107 941051 600193 941103
rect 600249 941051 600335 941103
rect 600391 941051 600477 941103
rect 600533 941051 600619 941103
rect 600675 941051 600761 941103
rect 600817 941051 600903 941103
rect 600959 941051 601045 941103
rect 601101 941051 601172 941103
rect 599272 941035 601172 941051
rect 599272 940979 599326 941035
rect 599382 940979 599450 941035
rect 599506 940979 599574 941035
rect 599630 940979 599698 941035
rect 599754 940979 599822 941035
rect 599878 940979 599946 941035
rect 600002 940979 600070 941035
rect 600126 940979 600194 941035
rect 600250 940979 600318 941035
rect 600374 940979 600442 941035
rect 600498 940979 600566 941035
rect 600622 940979 600690 941035
rect 600746 940979 600814 941035
rect 600870 940979 600938 941035
rect 600994 940979 601062 941035
rect 601118 940979 601172 941035
rect 599272 940965 601172 940979
rect 599272 940911 599341 940965
rect 599397 940911 599483 940965
rect 599539 940911 599625 940965
rect 599681 940911 599767 940965
rect 599823 940911 599909 940965
rect 599965 940911 600051 940965
rect 600107 940911 600193 940965
rect 600249 940911 600335 940965
rect 600391 940911 600477 940965
rect 600533 940911 600619 940965
rect 600675 940911 600761 940965
rect 600817 940911 600903 940965
rect 600959 940911 601045 940965
rect 601101 940911 601172 940965
rect 599272 940855 599326 940911
rect 599397 940909 599450 940911
rect 599539 940909 599574 940911
rect 599681 940909 599698 940911
rect 599382 940855 599450 940909
rect 599506 940855 599574 940909
rect 599630 940855 599698 940909
rect 599754 940909 599767 940911
rect 599878 940909 599909 940911
rect 600002 940909 600051 940911
rect 600126 940909 600193 940911
rect 599754 940855 599822 940909
rect 599878 940855 599946 940909
rect 600002 940855 600070 940909
rect 600126 940855 600194 940909
rect 600250 940855 600318 940911
rect 600391 940909 600442 940911
rect 600533 940909 600566 940911
rect 600675 940909 600690 940911
rect 600374 940855 600442 940909
rect 600498 940855 600566 940909
rect 600622 940855 600690 940909
rect 600746 940909 600761 940911
rect 600870 940909 600903 940911
rect 600994 940909 601045 940911
rect 600746 940855 600814 940909
rect 600870 940855 600938 940909
rect 600994 940855 601062 940909
rect 601118 940855 601172 940911
rect 599272 940823 601172 940855
rect 599272 940787 599341 940823
rect 599397 940787 599483 940823
rect 599539 940787 599625 940823
rect 599681 940787 599767 940823
rect 599823 940787 599909 940823
rect 599965 940787 600051 940823
rect 600107 940787 600193 940823
rect 600249 940787 600335 940823
rect 600391 940787 600477 940823
rect 600533 940787 600619 940823
rect 600675 940787 600761 940823
rect 600817 940787 600903 940823
rect 600959 940787 601045 940823
rect 601101 940787 601172 940823
rect 599272 940731 599326 940787
rect 599397 940767 599450 940787
rect 599539 940767 599574 940787
rect 599681 940767 599698 940787
rect 599382 940731 599450 940767
rect 599506 940731 599574 940767
rect 599630 940731 599698 940767
rect 599754 940767 599767 940787
rect 599878 940767 599909 940787
rect 600002 940767 600051 940787
rect 600126 940767 600193 940787
rect 599754 940731 599822 940767
rect 599878 940731 599946 940767
rect 600002 940731 600070 940767
rect 600126 940731 600194 940767
rect 600250 940731 600318 940787
rect 600391 940767 600442 940787
rect 600533 940767 600566 940787
rect 600675 940767 600690 940787
rect 600374 940731 600442 940767
rect 600498 940731 600566 940767
rect 600622 940731 600690 940767
rect 600746 940767 600761 940787
rect 600870 940767 600903 940787
rect 600994 940767 601045 940787
rect 600746 940731 600814 940767
rect 600870 940731 600938 940767
rect 600994 940731 601062 940767
rect 601118 940731 601172 940787
rect 599272 940681 601172 940731
rect 599272 940663 599341 940681
rect 599397 940663 599483 940681
rect 599539 940663 599625 940681
rect 599681 940663 599767 940681
rect 599823 940663 599909 940681
rect 599965 940663 600051 940681
rect 600107 940663 600193 940681
rect 600249 940663 600335 940681
rect 600391 940663 600477 940681
rect 600533 940663 600619 940681
rect 600675 940663 600761 940681
rect 600817 940663 600903 940681
rect 600959 940663 601045 940681
rect 601101 940663 601172 940681
rect 599272 940607 599326 940663
rect 599397 940625 599450 940663
rect 599539 940625 599574 940663
rect 599681 940625 599698 940663
rect 599382 940607 599450 940625
rect 599506 940607 599574 940625
rect 599630 940607 599698 940625
rect 599754 940625 599767 940663
rect 599878 940625 599909 940663
rect 600002 940625 600051 940663
rect 600126 940625 600193 940663
rect 599754 940607 599822 940625
rect 599878 940607 599946 940625
rect 600002 940607 600070 940625
rect 600126 940607 600194 940625
rect 600250 940607 600318 940663
rect 600391 940625 600442 940663
rect 600533 940625 600566 940663
rect 600675 940625 600690 940663
rect 600374 940607 600442 940625
rect 600498 940607 600566 940625
rect 600622 940607 600690 940625
rect 600746 940625 600761 940663
rect 600870 940625 600903 940663
rect 600994 940625 601045 940663
rect 600746 940607 600814 940625
rect 600870 940607 600938 940625
rect 600994 940607 601062 940625
rect 601118 940607 601172 940663
rect 599272 940539 601172 940607
rect 599272 940483 599326 940539
rect 599397 940483 599450 940539
rect 599539 940483 599574 940539
rect 599681 940483 599698 940539
rect 599754 940483 599767 940539
rect 599878 940483 599909 940539
rect 600002 940483 600051 940539
rect 600126 940483 600193 940539
rect 600250 940483 600318 940539
rect 600391 940483 600442 940539
rect 600533 940483 600566 940539
rect 600675 940483 600690 940539
rect 600746 940483 600761 940539
rect 600870 940483 600903 940539
rect 600994 940483 601045 940539
rect 601118 940483 601172 940539
rect 599272 940415 601172 940483
rect 599272 940359 599326 940415
rect 599382 940397 599450 940415
rect 599506 940397 599574 940415
rect 599630 940397 599698 940415
rect 599397 940359 599450 940397
rect 599539 940359 599574 940397
rect 599681 940359 599698 940397
rect 599754 940397 599822 940415
rect 599878 940397 599946 940415
rect 600002 940397 600070 940415
rect 600126 940397 600194 940415
rect 599754 940359 599767 940397
rect 599878 940359 599909 940397
rect 600002 940359 600051 940397
rect 600126 940359 600193 940397
rect 600250 940359 600318 940415
rect 600374 940397 600442 940415
rect 600498 940397 600566 940415
rect 600622 940397 600690 940415
rect 600391 940359 600442 940397
rect 600533 940359 600566 940397
rect 600675 940359 600690 940397
rect 600746 940397 600814 940415
rect 600870 940397 600938 940415
rect 600994 940397 601062 940415
rect 600746 940359 600761 940397
rect 600870 940359 600903 940397
rect 600994 940359 601045 940397
rect 601118 940359 601172 940415
rect 599272 940341 599341 940359
rect 599397 940341 599483 940359
rect 599539 940341 599625 940359
rect 599681 940341 599767 940359
rect 599823 940341 599909 940359
rect 599965 940341 600051 940359
rect 600107 940341 600193 940359
rect 600249 940341 600335 940359
rect 600391 940341 600477 940359
rect 600533 940341 600619 940359
rect 600675 940341 600761 940359
rect 600817 940341 600903 940359
rect 600959 940341 601045 940359
rect 601101 940341 601172 940359
rect 599272 940291 601172 940341
rect 599272 940235 599326 940291
rect 599382 940255 599450 940291
rect 599506 940255 599574 940291
rect 599630 940255 599698 940291
rect 599397 940235 599450 940255
rect 599539 940235 599574 940255
rect 599681 940235 599698 940255
rect 599754 940255 599822 940291
rect 599878 940255 599946 940291
rect 600002 940255 600070 940291
rect 600126 940255 600194 940291
rect 599754 940235 599767 940255
rect 599878 940235 599909 940255
rect 600002 940235 600051 940255
rect 600126 940235 600193 940255
rect 600250 940235 600318 940291
rect 600374 940255 600442 940291
rect 600498 940255 600566 940291
rect 600622 940255 600690 940291
rect 600391 940235 600442 940255
rect 600533 940235 600566 940255
rect 600675 940235 600690 940255
rect 600746 940255 600814 940291
rect 600870 940255 600938 940291
rect 600994 940255 601062 940291
rect 600746 940235 600761 940255
rect 600870 940235 600903 940255
rect 600994 940235 601045 940255
rect 601118 940235 601172 940291
rect 599272 940199 599341 940235
rect 599397 940199 599483 940235
rect 599539 940199 599625 940235
rect 599681 940199 599767 940235
rect 599823 940199 599909 940235
rect 599965 940199 600051 940235
rect 600107 940199 600193 940235
rect 600249 940199 600335 940235
rect 600391 940199 600477 940235
rect 600533 940199 600619 940235
rect 600675 940199 600761 940235
rect 600817 940199 600903 940235
rect 600959 940199 601045 940235
rect 601101 940199 601172 940235
rect 599272 940167 601172 940199
rect 599272 940111 599326 940167
rect 599382 940113 599450 940167
rect 599506 940113 599574 940167
rect 599630 940113 599698 940167
rect 599397 940111 599450 940113
rect 599539 940111 599574 940113
rect 599681 940111 599698 940113
rect 599754 940113 599822 940167
rect 599878 940113 599946 940167
rect 600002 940113 600070 940167
rect 600126 940113 600194 940167
rect 599754 940111 599767 940113
rect 599878 940111 599909 940113
rect 600002 940111 600051 940113
rect 600126 940111 600193 940113
rect 600250 940111 600318 940167
rect 600374 940113 600442 940167
rect 600498 940113 600566 940167
rect 600622 940113 600690 940167
rect 600391 940111 600442 940113
rect 600533 940111 600566 940113
rect 600675 940111 600690 940113
rect 600746 940113 600814 940167
rect 600870 940113 600938 940167
rect 600994 940113 601062 940167
rect 600746 940111 600761 940113
rect 600870 940111 600903 940113
rect 600994 940111 601045 940113
rect 601118 940111 601172 940167
rect 599272 940057 599341 940111
rect 599397 940057 599483 940111
rect 599539 940057 599625 940111
rect 599681 940057 599767 940111
rect 599823 940057 599909 940111
rect 599965 940057 600051 940111
rect 600107 940057 600193 940111
rect 600249 940057 600335 940111
rect 600391 940057 600477 940111
rect 600533 940057 600619 940111
rect 600675 940057 600761 940111
rect 600817 940057 600903 940111
rect 600959 940057 601045 940111
rect 601101 940057 601172 940111
rect 599272 940043 601172 940057
rect 599272 939987 599326 940043
rect 599382 939987 599450 940043
rect 599506 939987 599574 940043
rect 599630 939987 599698 940043
rect 599754 939987 599822 940043
rect 599878 939987 599946 940043
rect 600002 939987 600070 940043
rect 600126 939987 600194 940043
rect 600250 939987 600318 940043
rect 600374 939987 600442 940043
rect 600498 939987 600566 940043
rect 600622 939987 600690 940043
rect 600746 939987 600814 940043
rect 600870 939987 600938 940043
rect 600994 939987 601062 940043
rect 601118 939987 601172 940043
rect 599272 939971 601172 939987
rect 599272 939919 599341 939971
rect 599397 939919 599483 939971
rect 599539 939919 599625 939971
rect 599681 939919 599767 939971
rect 599823 939919 599909 939971
rect 599965 939919 600051 939971
rect 600107 939919 600193 939971
rect 600249 939919 600335 939971
rect 600391 939919 600477 939971
rect 600533 939919 600619 939971
rect 600675 939919 600761 939971
rect 600817 939919 600903 939971
rect 600959 939919 601045 939971
rect 601101 939919 601172 939971
rect 599272 939863 599326 939919
rect 599397 939915 599450 939919
rect 599539 939915 599574 939919
rect 599681 939915 599698 939919
rect 599382 939863 599450 939915
rect 599506 939863 599574 939915
rect 599630 939863 599698 939915
rect 599754 939915 599767 939919
rect 599878 939915 599909 939919
rect 600002 939915 600051 939919
rect 600126 939915 600193 939919
rect 599754 939863 599822 939915
rect 599878 939863 599946 939915
rect 600002 939863 600070 939915
rect 600126 939863 600194 939915
rect 600250 939863 600318 939919
rect 600391 939915 600442 939919
rect 600533 939915 600566 939919
rect 600675 939915 600690 939919
rect 600374 939863 600442 939915
rect 600498 939863 600566 939915
rect 600622 939863 600690 939915
rect 600746 939915 600761 939919
rect 600870 939915 600903 939919
rect 600994 939915 601045 939919
rect 600746 939863 600814 939915
rect 600870 939863 600938 939915
rect 600994 939863 601062 939915
rect 601118 939863 601172 939919
rect 599272 939829 601172 939863
rect 599272 939773 599341 939829
rect 599397 939773 599483 939829
rect 599539 939773 599625 939829
rect 599681 939773 599767 939829
rect 599823 939773 599909 939829
rect 599965 939773 600051 939829
rect 600107 939773 600193 939829
rect 600249 939773 600335 939829
rect 600391 939773 600477 939829
rect 600533 939773 600619 939829
rect 600675 939773 600761 939829
rect 600817 939773 600903 939829
rect 600959 939773 601045 939829
rect 601101 939773 601172 939829
rect 599272 939720 601172 939773
rect 601752 941675 603802 941720
rect 601752 941619 601829 941675
rect 601885 941655 601971 941675
rect 602027 941655 602113 941675
rect 602169 941655 602255 941675
rect 602311 941655 602397 941675
rect 602453 941655 602539 941675
rect 602595 941655 602681 941675
rect 602737 941655 602823 941675
rect 602879 941655 602965 941675
rect 603021 941655 603107 941675
rect 603163 941655 603249 941675
rect 603305 941655 603391 941675
rect 603447 941655 603533 941675
rect 603589 941655 603675 941675
rect 603731 941655 603802 941675
rect 601752 941599 601832 941619
rect 601888 941599 601956 941655
rect 602027 941619 602080 941655
rect 602169 941619 602204 941655
rect 602311 941619 602328 941655
rect 602012 941599 602080 941619
rect 602136 941599 602204 941619
rect 602260 941599 602328 941619
rect 602384 941619 602397 941655
rect 602508 941619 602539 941655
rect 602632 941619 602681 941655
rect 602756 941619 602823 941655
rect 602384 941599 602452 941619
rect 602508 941599 602576 941619
rect 602632 941599 602700 941619
rect 602756 941599 602824 941619
rect 602880 941599 602948 941655
rect 603021 941619 603072 941655
rect 603163 941619 603196 941655
rect 603305 941619 603320 941655
rect 603004 941599 603072 941619
rect 603128 941599 603196 941619
rect 603252 941599 603320 941619
rect 603376 941619 603391 941655
rect 603500 941619 603533 941655
rect 603624 941619 603675 941655
rect 603376 941599 603444 941619
rect 603500 941599 603568 941619
rect 603624 941599 603692 941619
rect 603748 941599 603802 941655
rect 601752 941533 603802 941599
rect 601752 941477 601829 941533
rect 601885 941531 601971 941533
rect 602027 941531 602113 941533
rect 602169 941531 602255 941533
rect 602311 941531 602397 941533
rect 602453 941531 602539 941533
rect 602595 941531 602681 941533
rect 602737 941531 602823 941533
rect 602879 941531 602965 941533
rect 603021 941531 603107 941533
rect 603163 941531 603249 941533
rect 603305 941531 603391 941533
rect 603447 941531 603533 941533
rect 603589 941531 603675 941533
rect 603731 941531 603802 941533
rect 601752 941475 601832 941477
rect 601888 941475 601956 941531
rect 602027 941477 602080 941531
rect 602169 941477 602204 941531
rect 602311 941477 602328 941531
rect 602012 941475 602080 941477
rect 602136 941475 602204 941477
rect 602260 941475 602328 941477
rect 602384 941477 602397 941531
rect 602508 941477 602539 941531
rect 602632 941477 602681 941531
rect 602756 941477 602823 941531
rect 602384 941475 602452 941477
rect 602508 941475 602576 941477
rect 602632 941475 602700 941477
rect 602756 941475 602824 941477
rect 602880 941475 602948 941531
rect 603021 941477 603072 941531
rect 603163 941477 603196 941531
rect 603305 941477 603320 941531
rect 603004 941475 603072 941477
rect 603128 941475 603196 941477
rect 603252 941475 603320 941477
rect 603376 941477 603391 941531
rect 603500 941477 603533 941531
rect 603624 941477 603675 941531
rect 603376 941475 603444 941477
rect 603500 941475 603568 941477
rect 603624 941475 603692 941477
rect 603748 941475 603802 941531
rect 601752 941407 603802 941475
rect 601752 941391 601832 941407
rect 601752 941335 601829 941391
rect 601888 941351 601956 941407
rect 602012 941391 602080 941407
rect 602136 941391 602204 941407
rect 602260 941391 602328 941407
rect 602027 941351 602080 941391
rect 602169 941351 602204 941391
rect 602311 941351 602328 941391
rect 602384 941391 602452 941407
rect 602508 941391 602576 941407
rect 602632 941391 602700 941407
rect 602756 941391 602824 941407
rect 602384 941351 602397 941391
rect 602508 941351 602539 941391
rect 602632 941351 602681 941391
rect 602756 941351 602823 941391
rect 602880 941351 602948 941407
rect 603004 941391 603072 941407
rect 603128 941391 603196 941407
rect 603252 941391 603320 941407
rect 603021 941351 603072 941391
rect 603163 941351 603196 941391
rect 603305 941351 603320 941391
rect 603376 941391 603444 941407
rect 603500 941391 603568 941407
rect 603624 941391 603692 941407
rect 603376 941351 603391 941391
rect 603500 941351 603533 941391
rect 603624 941351 603675 941391
rect 603748 941351 603802 941407
rect 601885 941335 601971 941351
rect 602027 941335 602113 941351
rect 602169 941335 602255 941351
rect 602311 941335 602397 941351
rect 602453 941335 602539 941351
rect 602595 941335 602681 941351
rect 602737 941335 602823 941351
rect 602879 941335 602965 941351
rect 603021 941335 603107 941351
rect 603163 941335 603249 941351
rect 603305 941335 603391 941351
rect 603447 941335 603533 941351
rect 603589 941335 603675 941351
rect 603731 941335 603802 941351
rect 601752 941283 603802 941335
rect 601752 941249 601832 941283
rect 601752 941193 601829 941249
rect 601888 941227 601956 941283
rect 602012 941249 602080 941283
rect 602136 941249 602204 941283
rect 602260 941249 602328 941283
rect 602027 941227 602080 941249
rect 602169 941227 602204 941249
rect 602311 941227 602328 941249
rect 602384 941249 602452 941283
rect 602508 941249 602576 941283
rect 602632 941249 602700 941283
rect 602756 941249 602824 941283
rect 602384 941227 602397 941249
rect 602508 941227 602539 941249
rect 602632 941227 602681 941249
rect 602756 941227 602823 941249
rect 602880 941227 602948 941283
rect 603004 941249 603072 941283
rect 603128 941249 603196 941283
rect 603252 941249 603320 941283
rect 603021 941227 603072 941249
rect 603163 941227 603196 941249
rect 603305 941227 603320 941249
rect 603376 941249 603444 941283
rect 603500 941249 603568 941283
rect 603624 941249 603692 941283
rect 603376 941227 603391 941249
rect 603500 941227 603533 941249
rect 603624 941227 603675 941249
rect 603748 941227 603802 941283
rect 601885 941193 601971 941227
rect 602027 941193 602113 941227
rect 602169 941193 602255 941227
rect 602311 941193 602397 941227
rect 602453 941193 602539 941227
rect 602595 941193 602681 941227
rect 602737 941193 602823 941227
rect 602879 941193 602965 941227
rect 603021 941193 603107 941227
rect 603163 941193 603249 941227
rect 603305 941193 603391 941227
rect 603447 941193 603533 941227
rect 603589 941193 603675 941227
rect 603731 941193 603802 941227
rect 601752 941159 603802 941193
rect 601752 941107 601832 941159
rect 601752 941051 601829 941107
rect 601888 941103 601956 941159
rect 602012 941107 602080 941159
rect 602136 941107 602204 941159
rect 602260 941107 602328 941159
rect 602027 941103 602080 941107
rect 602169 941103 602204 941107
rect 602311 941103 602328 941107
rect 602384 941107 602452 941159
rect 602508 941107 602576 941159
rect 602632 941107 602700 941159
rect 602756 941107 602824 941159
rect 602384 941103 602397 941107
rect 602508 941103 602539 941107
rect 602632 941103 602681 941107
rect 602756 941103 602823 941107
rect 602880 941103 602948 941159
rect 603004 941107 603072 941159
rect 603128 941107 603196 941159
rect 603252 941107 603320 941159
rect 603021 941103 603072 941107
rect 603163 941103 603196 941107
rect 603305 941103 603320 941107
rect 603376 941107 603444 941159
rect 603500 941107 603568 941159
rect 603624 941107 603692 941159
rect 603376 941103 603391 941107
rect 603500 941103 603533 941107
rect 603624 941103 603675 941107
rect 603748 941103 603802 941159
rect 601885 941051 601971 941103
rect 602027 941051 602113 941103
rect 602169 941051 602255 941103
rect 602311 941051 602397 941103
rect 602453 941051 602539 941103
rect 602595 941051 602681 941103
rect 602737 941051 602823 941103
rect 602879 941051 602965 941103
rect 603021 941051 603107 941103
rect 603163 941051 603249 941103
rect 603305 941051 603391 941103
rect 603447 941051 603533 941103
rect 603589 941051 603675 941103
rect 603731 941051 603802 941103
rect 601752 941035 603802 941051
rect 601752 940979 601832 941035
rect 601888 940979 601956 941035
rect 602012 940979 602080 941035
rect 602136 940979 602204 941035
rect 602260 940979 602328 941035
rect 602384 940979 602452 941035
rect 602508 940979 602576 941035
rect 602632 940979 602700 941035
rect 602756 940979 602824 941035
rect 602880 940979 602948 941035
rect 603004 940979 603072 941035
rect 603128 940979 603196 941035
rect 603252 940979 603320 941035
rect 603376 940979 603444 941035
rect 603500 940979 603568 941035
rect 603624 940979 603692 941035
rect 603748 940979 603802 941035
rect 601752 940965 603802 940979
rect 601752 940909 601829 940965
rect 601885 940911 601971 940965
rect 602027 940911 602113 940965
rect 602169 940911 602255 940965
rect 602311 940911 602397 940965
rect 602453 940911 602539 940965
rect 602595 940911 602681 940965
rect 602737 940911 602823 940965
rect 602879 940911 602965 940965
rect 603021 940911 603107 940965
rect 603163 940911 603249 940965
rect 603305 940911 603391 940965
rect 603447 940911 603533 940965
rect 603589 940911 603675 940965
rect 603731 940911 603802 940965
rect 601752 940855 601832 940909
rect 601888 940855 601956 940911
rect 602027 940909 602080 940911
rect 602169 940909 602204 940911
rect 602311 940909 602328 940911
rect 602012 940855 602080 940909
rect 602136 940855 602204 940909
rect 602260 940855 602328 940909
rect 602384 940909 602397 940911
rect 602508 940909 602539 940911
rect 602632 940909 602681 940911
rect 602756 940909 602823 940911
rect 602384 940855 602452 940909
rect 602508 940855 602576 940909
rect 602632 940855 602700 940909
rect 602756 940855 602824 940909
rect 602880 940855 602948 940911
rect 603021 940909 603072 940911
rect 603163 940909 603196 940911
rect 603305 940909 603320 940911
rect 603004 940855 603072 940909
rect 603128 940855 603196 940909
rect 603252 940855 603320 940909
rect 603376 940909 603391 940911
rect 603500 940909 603533 940911
rect 603624 940909 603675 940911
rect 603376 940855 603444 940909
rect 603500 940855 603568 940909
rect 603624 940855 603692 940909
rect 603748 940855 603802 940911
rect 601752 940823 603802 940855
rect 601752 940767 601829 940823
rect 601885 940787 601971 940823
rect 602027 940787 602113 940823
rect 602169 940787 602255 940823
rect 602311 940787 602397 940823
rect 602453 940787 602539 940823
rect 602595 940787 602681 940823
rect 602737 940787 602823 940823
rect 602879 940787 602965 940823
rect 603021 940787 603107 940823
rect 603163 940787 603249 940823
rect 603305 940787 603391 940823
rect 603447 940787 603533 940823
rect 603589 940787 603675 940823
rect 603731 940787 603802 940823
rect 601752 940731 601832 940767
rect 601888 940731 601956 940787
rect 602027 940767 602080 940787
rect 602169 940767 602204 940787
rect 602311 940767 602328 940787
rect 602012 940731 602080 940767
rect 602136 940731 602204 940767
rect 602260 940731 602328 940767
rect 602384 940767 602397 940787
rect 602508 940767 602539 940787
rect 602632 940767 602681 940787
rect 602756 940767 602823 940787
rect 602384 940731 602452 940767
rect 602508 940731 602576 940767
rect 602632 940731 602700 940767
rect 602756 940731 602824 940767
rect 602880 940731 602948 940787
rect 603021 940767 603072 940787
rect 603163 940767 603196 940787
rect 603305 940767 603320 940787
rect 603004 940731 603072 940767
rect 603128 940731 603196 940767
rect 603252 940731 603320 940767
rect 603376 940767 603391 940787
rect 603500 940767 603533 940787
rect 603624 940767 603675 940787
rect 603376 940731 603444 940767
rect 603500 940731 603568 940767
rect 603624 940731 603692 940767
rect 603748 940731 603802 940787
rect 601752 940681 603802 940731
rect 601752 940625 601829 940681
rect 601885 940663 601971 940681
rect 602027 940663 602113 940681
rect 602169 940663 602255 940681
rect 602311 940663 602397 940681
rect 602453 940663 602539 940681
rect 602595 940663 602681 940681
rect 602737 940663 602823 940681
rect 602879 940663 602965 940681
rect 603021 940663 603107 940681
rect 603163 940663 603249 940681
rect 603305 940663 603391 940681
rect 603447 940663 603533 940681
rect 603589 940663 603675 940681
rect 603731 940663 603802 940681
rect 601752 940607 601832 940625
rect 601888 940607 601956 940663
rect 602027 940625 602080 940663
rect 602169 940625 602204 940663
rect 602311 940625 602328 940663
rect 602012 940607 602080 940625
rect 602136 940607 602204 940625
rect 602260 940607 602328 940625
rect 602384 940625 602397 940663
rect 602508 940625 602539 940663
rect 602632 940625 602681 940663
rect 602756 940625 602823 940663
rect 602384 940607 602452 940625
rect 602508 940607 602576 940625
rect 602632 940607 602700 940625
rect 602756 940607 602824 940625
rect 602880 940607 602948 940663
rect 603021 940625 603072 940663
rect 603163 940625 603196 940663
rect 603305 940625 603320 940663
rect 603004 940607 603072 940625
rect 603128 940607 603196 940625
rect 603252 940607 603320 940625
rect 603376 940625 603391 940663
rect 603500 940625 603533 940663
rect 603624 940625 603675 940663
rect 603376 940607 603444 940625
rect 603500 940607 603568 940625
rect 603624 940607 603692 940625
rect 603748 940607 603802 940663
rect 601752 940539 603802 940607
rect 601752 940483 601829 940539
rect 601888 940483 601956 940539
rect 602027 940483 602080 940539
rect 602169 940483 602204 940539
rect 602311 940483 602328 940539
rect 602384 940483 602397 940539
rect 602508 940483 602539 940539
rect 602632 940483 602681 940539
rect 602756 940483 602823 940539
rect 602880 940483 602948 940539
rect 603021 940483 603072 940539
rect 603163 940483 603196 940539
rect 603305 940483 603320 940539
rect 603376 940483 603391 940539
rect 603500 940483 603533 940539
rect 603624 940483 603675 940539
rect 603748 940483 603802 940539
rect 601752 940415 603802 940483
rect 601752 940397 601832 940415
rect 601752 940341 601829 940397
rect 601888 940359 601956 940415
rect 602012 940397 602080 940415
rect 602136 940397 602204 940415
rect 602260 940397 602328 940415
rect 602027 940359 602080 940397
rect 602169 940359 602204 940397
rect 602311 940359 602328 940397
rect 602384 940397 602452 940415
rect 602508 940397 602576 940415
rect 602632 940397 602700 940415
rect 602756 940397 602824 940415
rect 602384 940359 602397 940397
rect 602508 940359 602539 940397
rect 602632 940359 602681 940397
rect 602756 940359 602823 940397
rect 602880 940359 602948 940415
rect 603004 940397 603072 940415
rect 603128 940397 603196 940415
rect 603252 940397 603320 940415
rect 603021 940359 603072 940397
rect 603163 940359 603196 940397
rect 603305 940359 603320 940397
rect 603376 940397 603444 940415
rect 603500 940397 603568 940415
rect 603624 940397 603692 940415
rect 603376 940359 603391 940397
rect 603500 940359 603533 940397
rect 603624 940359 603675 940397
rect 603748 940359 603802 940415
rect 601885 940341 601971 940359
rect 602027 940341 602113 940359
rect 602169 940341 602255 940359
rect 602311 940341 602397 940359
rect 602453 940341 602539 940359
rect 602595 940341 602681 940359
rect 602737 940341 602823 940359
rect 602879 940341 602965 940359
rect 603021 940341 603107 940359
rect 603163 940341 603249 940359
rect 603305 940341 603391 940359
rect 603447 940341 603533 940359
rect 603589 940341 603675 940359
rect 603731 940341 603802 940359
rect 601752 940291 603802 940341
rect 601752 940255 601832 940291
rect 601752 940199 601829 940255
rect 601888 940235 601956 940291
rect 602012 940255 602080 940291
rect 602136 940255 602204 940291
rect 602260 940255 602328 940291
rect 602027 940235 602080 940255
rect 602169 940235 602204 940255
rect 602311 940235 602328 940255
rect 602384 940255 602452 940291
rect 602508 940255 602576 940291
rect 602632 940255 602700 940291
rect 602756 940255 602824 940291
rect 602384 940235 602397 940255
rect 602508 940235 602539 940255
rect 602632 940235 602681 940255
rect 602756 940235 602823 940255
rect 602880 940235 602948 940291
rect 603004 940255 603072 940291
rect 603128 940255 603196 940291
rect 603252 940255 603320 940291
rect 603021 940235 603072 940255
rect 603163 940235 603196 940255
rect 603305 940235 603320 940255
rect 603376 940255 603444 940291
rect 603500 940255 603568 940291
rect 603624 940255 603692 940291
rect 603376 940235 603391 940255
rect 603500 940235 603533 940255
rect 603624 940235 603675 940255
rect 603748 940235 603802 940291
rect 601885 940199 601971 940235
rect 602027 940199 602113 940235
rect 602169 940199 602255 940235
rect 602311 940199 602397 940235
rect 602453 940199 602539 940235
rect 602595 940199 602681 940235
rect 602737 940199 602823 940235
rect 602879 940199 602965 940235
rect 603021 940199 603107 940235
rect 603163 940199 603249 940235
rect 603305 940199 603391 940235
rect 603447 940199 603533 940235
rect 603589 940199 603675 940235
rect 603731 940199 603802 940235
rect 601752 940167 603802 940199
rect 601752 940113 601832 940167
rect 601752 940057 601829 940113
rect 601888 940111 601956 940167
rect 602012 940113 602080 940167
rect 602136 940113 602204 940167
rect 602260 940113 602328 940167
rect 602027 940111 602080 940113
rect 602169 940111 602204 940113
rect 602311 940111 602328 940113
rect 602384 940113 602452 940167
rect 602508 940113 602576 940167
rect 602632 940113 602700 940167
rect 602756 940113 602824 940167
rect 602384 940111 602397 940113
rect 602508 940111 602539 940113
rect 602632 940111 602681 940113
rect 602756 940111 602823 940113
rect 602880 940111 602948 940167
rect 603004 940113 603072 940167
rect 603128 940113 603196 940167
rect 603252 940113 603320 940167
rect 603021 940111 603072 940113
rect 603163 940111 603196 940113
rect 603305 940111 603320 940113
rect 603376 940113 603444 940167
rect 603500 940113 603568 940167
rect 603624 940113 603692 940167
rect 603376 940111 603391 940113
rect 603500 940111 603533 940113
rect 603624 940111 603675 940113
rect 603748 940111 603802 940167
rect 601885 940057 601971 940111
rect 602027 940057 602113 940111
rect 602169 940057 602255 940111
rect 602311 940057 602397 940111
rect 602453 940057 602539 940111
rect 602595 940057 602681 940111
rect 602737 940057 602823 940111
rect 602879 940057 602965 940111
rect 603021 940057 603107 940111
rect 603163 940057 603249 940111
rect 603305 940057 603391 940111
rect 603447 940057 603533 940111
rect 603589 940057 603675 940111
rect 603731 940057 603802 940111
rect 601752 940043 603802 940057
rect 601752 939987 601832 940043
rect 601888 939987 601956 940043
rect 602012 939987 602080 940043
rect 602136 939987 602204 940043
rect 602260 939987 602328 940043
rect 602384 939987 602452 940043
rect 602508 939987 602576 940043
rect 602632 939987 602700 940043
rect 602756 939987 602824 940043
rect 602880 939987 602948 940043
rect 603004 939987 603072 940043
rect 603128 939987 603196 940043
rect 603252 939987 603320 940043
rect 603376 939987 603444 940043
rect 603500 939987 603568 940043
rect 603624 939987 603692 940043
rect 603748 939987 603802 940043
rect 601752 939971 603802 939987
rect 601752 939915 601829 939971
rect 601885 939919 601971 939971
rect 602027 939919 602113 939971
rect 602169 939919 602255 939971
rect 602311 939919 602397 939971
rect 602453 939919 602539 939971
rect 602595 939919 602681 939971
rect 602737 939919 602823 939971
rect 602879 939919 602965 939971
rect 603021 939919 603107 939971
rect 603163 939919 603249 939971
rect 603305 939919 603391 939971
rect 603447 939919 603533 939971
rect 603589 939919 603675 939971
rect 603731 939919 603802 939971
rect 601752 939863 601832 939915
rect 601888 939863 601956 939919
rect 602027 939915 602080 939919
rect 602169 939915 602204 939919
rect 602311 939915 602328 939919
rect 602012 939863 602080 939915
rect 602136 939863 602204 939915
rect 602260 939863 602328 939915
rect 602384 939915 602397 939919
rect 602508 939915 602539 939919
rect 602632 939915 602681 939919
rect 602756 939915 602823 939919
rect 602384 939863 602452 939915
rect 602508 939863 602576 939915
rect 602632 939863 602700 939915
rect 602756 939863 602824 939915
rect 602880 939863 602948 939919
rect 603021 939915 603072 939919
rect 603163 939915 603196 939919
rect 603305 939915 603320 939919
rect 603004 939863 603072 939915
rect 603128 939863 603196 939915
rect 603252 939863 603320 939915
rect 603376 939915 603391 939919
rect 603500 939915 603533 939919
rect 603624 939915 603675 939919
rect 603376 939863 603444 939915
rect 603500 939863 603568 939915
rect 603624 939863 603692 939915
rect 603748 939863 603802 939919
rect 601752 939829 603802 939863
rect 601752 939773 601829 939829
rect 601885 939773 601971 939829
rect 602027 939773 602113 939829
rect 602169 939773 602255 939829
rect 602311 939773 602397 939829
rect 602453 939773 602539 939829
rect 602595 939773 602681 939829
rect 602737 939773 602823 939829
rect 602879 939773 602965 939829
rect 603021 939773 603107 939829
rect 603163 939773 603249 939829
rect 603305 939773 603391 939829
rect 603447 939773 603533 939829
rect 603589 939773 603675 939829
rect 603731 939773 603802 939829
rect 601752 939720 603802 939773
rect 604122 941675 606172 941720
rect 604122 941619 605051 941675
rect 605107 941655 605193 941675
rect 605249 941655 605335 941675
rect 605391 941655 605477 941675
rect 605533 941655 605619 941675
rect 605675 941655 605761 941675
rect 605817 941655 605903 941675
rect 605959 941655 606045 941675
rect 606101 941655 606172 941675
rect 605126 941619 605193 941655
rect 604122 941599 605070 941619
rect 605126 941599 605194 941619
rect 605250 941599 605318 941655
rect 605391 941619 605442 941655
rect 605533 941619 605566 941655
rect 605675 941619 605690 941655
rect 605374 941599 605442 941619
rect 605498 941599 605566 941619
rect 605622 941599 605690 941619
rect 605746 941619 605761 941655
rect 605870 941619 605903 941655
rect 605994 941619 606045 941655
rect 605746 941599 605814 941619
rect 605870 941599 605938 941619
rect 605994 941599 606062 941619
rect 606118 941599 606172 941655
rect 604122 941533 606172 941599
rect 604122 941477 605051 941533
rect 605107 941531 605193 941533
rect 605249 941531 605335 941533
rect 605391 941531 605477 941533
rect 605533 941531 605619 941533
rect 605675 941531 605761 941533
rect 605817 941531 605903 941533
rect 605959 941531 606045 941533
rect 606101 941531 606172 941533
rect 605126 941477 605193 941531
rect 604122 941475 605070 941477
rect 605126 941475 605194 941477
rect 605250 941475 605318 941531
rect 605391 941477 605442 941531
rect 605533 941477 605566 941531
rect 605675 941477 605690 941531
rect 605374 941475 605442 941477
rect 605498 941475 605566 941477
rect 605622 941475 605690 941477
rect 605746 941477 605761 941531
rect 605870 941477 605903 941531
rect 605994 941477 606045 941531
rect 605746 941475 605814 941477
rect 605870 941475 605938 941477
rect 605994 941475 606062 941477
rect 606118 941475 606172 941531
rect 604122 941407 606172 941475
rect 604122 941391 605070 941407
rect 605126 941391 605194 941407
rect 604122 941335 605051 941391
rect 605126 941351 605193 941391
rect 605250 941351 605318 941407
rect 605374 941391 605442 941407
rect 605498 941391 605566 941407
rect 605622 941391 605690 941407
rect 605391 941351 605442 941391
rect 605533 941351 605566 941391
rect 605675 941351 605690 941391
rect 605746 941391 605814 941407
rect 605870 941391 605938 941407
rect 605994 941391 606062 941407
rect 605746 941351 605761 941391
rect 605870 941351 605903 941391
rect 605994 941351 606045 941391
rect 606118 941351 606172 941407
rect 605107 941335 605193 941351
rect 605249 941335 605335 941351
rect 605391 941335 605477 941351
rect 605533 941335 605619 941351
rect 605675 941335 605761 941351
rect 605817 941335 605903 941351
rect 605959 941335 606045 941351
rect 606101 941335 606172 941351
rect 604122 941283 606172 941335
rect 604122 941249 605070 941283
rect 605126 941249 605194 941283
rect 604122 941193 605051 941249
rect 605126 941227 605193 941249
rect 605250 941227 605318 941283
rect 605374 941249 605442 941283
rect 605498 941249 605566 941283
rect 605622 941249 605690 941283
rect 605391 941227 605442 941249
rect 605533 941227 605566 941249
rect 605675 941227 605690 941249
rect 605746 941249 605814 941283
rect 605870 941249 605938 941283
rect 605994 941249 606062 941283
rect 605746 941227 605761 941249
rect 605870 941227 605903 941249
rect 605994 941227 606045 941249
rect 606118 941227 606172 941283
rect 605107 941193 605193 941227
rect 605249 941193 605335 941227
rect 605391 941193 605477 941227
rect 605533 941193 605619 941227
rect 605675 941193 605761 941227
rect 605817 941193 605903 941227
rect 605959 941193 606045 941227
rect 606101 941193 606172 941227
rect 604122 941159 606172 941193
rect 604122 941107 605070 941159
rect 605126 941107 605194 941159
rect 604122 941051 605051 941107
rect 605126 941103 605193 941107
rect 605250 941103 605318 941159
rect 605374 941107 605442 941159
rect 605498 941107 605566 941159
rect 605622 941107 605690 941159
rect 605391 941103 605442 941107
rect 605533 941103 605566 941107
rect 605675 941103 605690 941107
rect 605746 941107 605814 941159
rect 605870 941107 605938 941159
rect 605994 941107 606062 941159
rect 605746 941103 605761 941107
rect 605870 941103 605903 941107
rect 605994 941103 606045 941107
rect 606118 941103 606172 941159
rect 605107 941051 605193 941103
rect 605249 941051 605335 941103
rect 605391 941051 605477 941103
rect 605533 941051 605619 941103
rect 605675 941051 605761 941103
rect 605817 941051 605903 941103
rect 605959 941051 606045 941103
rect 606101 941051 606172 941103
rect 604122 941035 606172 941051
rect 604122 940979 605070 941035
rect 605126 940979 605194 941035
rect 605250 940979 605318 941035
rect 605374 940979 605442 941035
rect 605498 940979 605566 941035
rect 605622 940979 605690 941035
rect 605746 940979 605814 941035
rect 605870 940979 605938 941035
rect 605994 940979 606062 941035
rect 606118 940979 606172 941035
rect 604122 940965 606172 940979
rect 604122 940909 605051 940965
rect 605107 940911 605193 940965
rect 605249 940911 605335 940965
rect 605391 940911 605477 940965
rect 605533 940911 605619 940965
rect 605675 940911 605761 940965
rect 605817 940911 605903 940965
rect 605959 940911 606045 940965
rect 606101 940911 606172 940965
rect 605126 940909 605193 940911
rect 604122 940855 605070 940909
rect 605126 940855 605194 940909
rect 605250 940855 605318 940911
rect 605391 940909 605442 940911
rect 605533 940909 605566 940911
rect 605675 940909 605690 940911
rect 605374 940855 605442 940909
rect 605498 940855 605566 940909
rect 605622 940855 605690 940909
rect 605746 940909 605761 940911
rect 605870 940909 605903 940911
rect 605994 940909 606045 940911
rect 605746 940855 605814 940909
rect 605870 940855 605938 940909
rect 605994 940855 606062 940909
rect 606118 940855 606172 940911
rect 604122 940823 606172 940855
rect 604122 940767 605051 940823
rect 605107 940787 605193 940823
rect 605249 940787 605335 940823
rect 605391 940787 605477 940823
rect 605533 940787 605619 940823
rect 605675 940787 605761 940823
rect 605817 940787 605903 940823
rect 605959 940787 606045 940823
rect 606101 940787 606172 940823
rect 605126 940767 605193 940787
rect 604122 940731 605070 940767
rect 605126 940731 605194 940767
rect 605250 940731 605318 940787
rect 605391 940767 605442 940787
rect 605533 940767 605566 940787
rect 605675 940767 605690 940787
rect 605374 940731 605442 940767
rect 605498 940731 605566 940767
rect 605622 940731 605690 940767
rect 605746 940767 605761 940787
rect 605870 940767 605903 940787
rect 605994 940767 606045 940787
rect 605746 940731 605814 940767
rect 605870 940731 605938 940767
rect 605994 940731 606062 940767
rect 606118 940731 606172 940787
rect 604122 940681 606172 940731
rect 604122 940625 605051 940681
rect 605107 940663 605193 940681
rect 605249 940663 605335 940681
rect 605391 940663 605477 940681
rect 605533 940663 605619 940681
rect 605675 940663 605761 940681
rect 605817 940663 605903 940681
rect 605959 940663 606045 940681
rect 606101 940663 606172 940681
rect 605126 940625 605193 940663
rect 604122 940607 605070 940625
rect 605126 940607 605194 940625
rect 605250 940607 605318 940663
rect 605391 940625 605442 940663
rect 605533 940625 605566 940663
rect 605675 940625 605690 940663
rect 605374 940607 605442 940625
rect 605498 940607 605566 940625
rect 605622 940607 605690 940625
rect 605746 940625 605761 940663
rect 605870 940625 605903 940663
rect 605994 940625 606045 940663
rect 605746 940607 605814 940625
rect 605870 940607 605938 940625
rect 605994 940607 606062 940625
rect 606118 940607 606172 940663
rect 604122 940539 606172 940607
rect 604122 940483 605051 940539
rect 605126 940483 605193 940539
rect 605250 940483 605318 940539
rect 605391 940483 605442 940539
rect 605533 940483 605566 940539
rect 605675 940483 605690 940539
rect 605746 940483 605761 940539
rect 605870 940483 605903 940539
rect 605994 940483 606045 940539
rect 606118 940483 606172 940539
rect 604122 940415 606172 940483
rect 604122 940397 605070 940415
rect 605126 940397 605194 940415
rect 604122 940341 605051 940397
rect 605126 940359 605193 940397
rect 605250 940359 605318 940415
rect 605374 940397 605442 940415
rect 605498 940397 605566 940415
rect 605622 940397 605690 940415
rect 605391 940359 605442 940397
rect 605533 940359 605566 940397
rect 605675 940359 605690 940397
rect 605746 940397 605814 940415
rect 605870 940397 605938 940415
rect 605994 940397 606062 940415
rect 605746 940359 605761 940397
rect 605870 940359 605903 940397
rect 605994 940359 606045 940397
rect 606118 940359 606172 940415
rect 605107 940341 605193 940359
rect 605249 940341 605335 940359
rect 605391 940341 605477 940359
rect 605533 940341 605619 940359
rect 605675 940341 605761 940359
rect 605817 940341 605903 940359
rect 605959 940341 606045 940359
rect 606101 940341 606172 940359
rect 604122 940291 606172 940341
rect 604122 940255 605070 940291
rect 605126 940255 605194 940291
rect 604122 940199 605051 940255
rect 605126 940235 605193 940255
rect 605250 940235 605318 940291
rect 605374 940255 605442 940291
rect 605498 940255 605566 940291
rect 605622 940255 605690 940291
rect 605391 940235 605442 940255
rect 605533 940235 605566 940255
rect 605675 940235 605690 940255
rect 605746 940255 605814 940291
rect 605870 940255 605938 940291
rect 605994 940255 606062 940291
rect 605746 940235 605761 940255
rect 605870 940235 605903 940255
rect 605994 940235 606045 940255
rect 606118 940235 606172 940291
rect 605107 940199 605193 940235
rect 605249 940199 605335 940235
rect 605391 940199 605477 940235
rect 605533 940199 605619 940235
rect 605675 940199 605761 940235
rect 605817 940199 605903 940235
rect 605959 940199 606045 940235
rect 606101 940199 606172 940235
rect 604122 940167 606172 940199
rect 604122 940113 605070 940167
rect 605126 940113 605194 940167
rect 604122 940057 605051 940113
rect 605126 940111 605193 940113
rect 605250 940111 605318 940167
rect 605374 940113 605442 940167
rect 605498 940113 605566 940167
rect 605622 940113 605690 940167
rect 605391 940111 605442 940113
rect 605533 940111 605566 940113
rect 605675 940111 605690 940113
rect 605746 940113 605814 940167
rect 605870 940113 605938 940167
rect 605994 940113 606062 940167
rect 605746 940111 605761 940113
rect 605870 940111 605903 940113
rect 605994 940111 606045 940113
rect 606118 940111 606172 940167
rect 605107 940057 605193 940111
rect 605249 940057 605335 940111
rect 605391 940057 605477 940111
rect 605533 940057 605619 940111
rect 605675 940057 605761 940111
rect 605817 940057 605903 940111
rect 605959 940057 606045 940111
rect 606101 940057 606172 940111
rect 604122 940043 606172 940057
rect 604122 939987 605070 940043
rect 605126 939987 605194 940043
rect 605250 939987 605318 940043
rect 605374 939987 605442 940043
rect 605498 939987 605566 940043
rect 605622 939987 605690 940043
rect 605746 939987 605814 940043
rect 605870 939987 605938 940043
rect 605994 939987 606062 940043
rect 606118 939987 606172 940043
rect 604122 939971 606172 939987
rect 604122 939915 605051 939971
rect 605107 939919 605193 939971
rect 605249 939919 605335 939971
rect 605391 939919 605477 939971
rect 605533 939919 605619 939971
rect 605675 939919 605761 939971
rect 605817 939919 605903 939971
rect 605959 939919 606045 939971
rect 606101 939919 606172 939971
rect 605126 939915 605193 939919
rect 604122 939863 605070 939915
rect 605126 939863 605194 939915
rect 605250 939863 605318 939919
rect 605391 939915 605442 939919
rect 605533 939915 605566 939919
rect 605675 939915 605690 939919
rect 605374 939863 605442 939915
rect 605498 939863 605566 939915
rect 605622 939863 605690 939915
rect 605746 939915 605761 939919
rect 605870 939915 605903 939919
rect 605994 939915 606045 939919
rect 605746 939863 605814 939915
rect 605870 939863 605938 939915
rect 605994 939863 606062 939915
rect 606118 939863 606172 939919
rect 604122 939829 606172 939863
rect 604122 939773 605051 939829
rect 605107 939773 605193 939829
rect 605249 939773 605335 939829
rect 605391 939773 605477 939829
rect 605533 939773 605619 939829
rect 605675 939773 605761 939829
rect 605817 939773 605903 939829
rect 605959 939773 606045 939829
rect 606101 939773 606172 939829
rect 604122 939720 606172 939773
rect 606828 941675 608878 941720
rect 606828 941619 606905 941675
rect 606961 941655 607047 941675
rect 607103 941655 607189 941675
rect 607245 941655 607331 941675
rect 607387 941655 607473 941675
rect 607529 941655 607615 941675
rect 607671 941655 607757 941675
rect 607813 941655 607899 941675
rect 607955 941655 608041 941675
rect 608097 941655 608183 941675
rect 608239 941655 608325 941675
rect 608381 941655 608467 941675
rect 608523 941655 608609 941675
rect 608665 941655 608751 941675
rect 608807 941655 608878 941675
rect 606828 941599 606908 941619
rect 606964 941599 607032 941655
rect 607103 941619 607156 941655
rect 607245 941619 607280 941655
rect 607387 941619 607404 941655
rect 607088 941599 607156 941619
rect 607212 941599 607280 941619
rect 607336 941599 607404 941619
rect 607460 941619 607473 941655
rect 607584 941619 607615 941655
rect 607708 941619 607757 941655
rect 607832 941619 607899 941655
rect 607460 941599 607528 941619
rect 607584 941599 607652 941619
rect 607708 941599 607776 941619
rect 607832 941599 607900 941619
rect 607956 941599 608024 941655
rect 608097 941619 608148 941655
rect 608239 941619 608272 941655
rect 608381 941619 608396 941655
rect 608080 941599 608148 941619
rect 608204 941599 608272 941619
rect 608328 941599 608396 941619
rect 608452 941619 608467 941655
rect 608576 941619 608609 941655
rect 608700 941619 608751 941655
rect 608452 941599 608520 941619
rect 608576 941599 608644 941619
rect 608700 941599 608768 941619
rect 608824 941599 608878 941655
rect 606828 941533 608878 941599
rect 606828 941477 606905 941533
rect 606961 941531 607047 941533
rect 607103 941531 607189 941533
rect 607245 941531 607331 941533
rect 607387 941531 607473 941533
rect 607529 941531 607615 941533
rect 607671 941531 607757 941533
rect 607813 941531 607899 941533
rect 607955 941531 608041 941533
rect 608097 941531 608183 941533
rect 608239 941531 608325 941533
rect 608381 941531 608467 941533
rect 608523 941531 608609 941533
rect 608665 941531 608751 941533
rect 608807 941531 608878 941533
rect 606828 941475 606908 941477
rect 606964 941475 607032 941531
rect 607103 941477 607156 941531
rect 607245 941477 607280 941531
rect 607387 941477 607404 941531
rect 607088 941475 607156 941477
rect 607212 941475 607280 941477
rect 607336 941475 607404 941477
rect 607460 941477 607473 941531
rect 607584 941477 607615 941531
rect 607708 941477 607757 941531
rect 607832 941477 607899 941531
rect 607460 941475 607528 941477
rect 607584 941475 607652 941477
rect 607708 941475 607776 941477
rect 607832 941475 607900 941477
rect 607956 941475 608024 941531
rect 608097 941477 608148 941531
rect 608239 941477 608272 941531
rect 608381 941477 608396 941531
rect 608080 941475 608148 941477
rect 608204 941475 608272 941477
rect 608328 941475 608396 941477
rect 608452 941477 608467 941531
rect 608576 941477 608609 941531
rect 608700 941477 608751 941531
rect 608452 941475 608520 941477
rect 608576 941475 608644 941477
rect 608700 941475 608768 941477
rect 608824 941475 608878 941531
rect 606828 941407 608878 941475
rect 606828 941391 606908 941407
rect 606828 941335 606905 941391
rect 606964 941351 607032 941407
rect 607088 941391 607156 941407
rect 607212 941391 607280 941407
rect 607336 941391 607404 941407
rect 607103 941351 607156 941391
rect 607245 941351 607280 941391
rect 607387 941351 607404 941391
rect 607460 941391 607528 941407
rect 607584 941391 607652 941407
rect 607708 941391 607776 941407
rect 607832 941391 607900 941407
rect 607460 941351 607473 941391
rect 607584 941351 607615 941391
rect 607708 941351 607757 941391
rect 607832 941351 607899 941391
rect 607956 941351 608024 941407
rect 608080 941391 608148 941407
rect 608204 941391 608272 941407
rect 608328 941391 608396 941407
rect 608097 941351 608148 941391
rect 608239 941351 608272 941391
rect 608381 941351 608396 941391
rect 608452 941391 608520 941407
rect 608576 941391 608644 941407
rect 608700 941391 608768 941407
rect 608452 941351 608467 941391
rect 608576 941351 608609 941391
rect 608700 941351 608751 941391
rect 608824 941351 608878 941407
rect 606961 941335 607047 941351
rect 607103 941335 607189 941351
rect 607245 941335 607331 941351
rect 607387 941335 607473 941351
rect 607529 941335 607615 941351
rect 607671 941335 607757 941351
rect 607813 941335 607899 941351
rect 607955 941335 608041 941351
rect 608097 941335 608183 941351
rect 608239 941335 608325 941351
rect 608381 941335 608467 941351
rect 608523 941335 608609 941351
rect 608665 941335 608751 941351
rect 608807 941335 608878 941351
rect 606828 941283 608878 941335
rect 606828 941249 606908 941283
rect 606828 941193 606905 941249
rect 606964 941227 607032 941283
rect 607088 941249 607156 941283
rect 607212 941249 607280 941283
rect 607336 941249 607404 941283
rect 607103 941227 607156 941249
rect 607245 941227 607280 941249
rect 607387 941227 607404 941249
rect 607460 941249 607528 941283
rect 607584 941249 607652 941283
rect 607708 941249 607776 941283
rect 607832 941249 607900 941283
rect 607460 941227 607473 941249
rect 607584 941227 607615 941249
rect 607708 941227 607757 941249
rect 607832 941227 607899 941249
rect 607956 941227 608024 941283
rect 608080 941249 608148 941283
rect 608204 941249 608272 941283
rect 608328 941249 608396 941283
rect 608097 941227 608148 941249
rect 608239 941227 608272 941249
rect 608381 941227 608396 941249
rect 608452 941249 608520 941283
rect 608576 941249 608644 941283
rect 608700 941249 608768 941283
rect 608452 941227 608467 941249
rect 608576 941227 608609 941249
rect 608700 941227 608751 941249
rect 608824 941227 608878 941283
rect 606961 941193 607047 941227
rect 607103 941193 607189 941227
rect 607245 941193 607331 941227
rect 607387 941193 607473 941227
rect 607529 941193 607615 941227
rect 607671 941193 607757 941227
rect 607813 941193 607899 941227
rect 607955 941193 608041 941227
rect 608097 941193 608183 941227
rect 608239 941193 608325 941227
rect 608381 941193 608467 941227
rect 608523 941193 608609 941227
rect 608665 941193 608751 941227
rect 608807 941193 608878 941227
rect 606828 941159 608878 941193
rect 606828 941107 606908 941159
rect 606828 941051 606905 941107
rect 606964 941103 607032 941159
rect 607088 941107 607156 941159
rect 607212 941107 607280 941159
rect 607336 941107 607404 941159
rect 607103 941103 607156 941107
rect 607245 941103 607280 941107
rect 607387 941103 607404 941107
rect 607460 941107 607528 941159
rect 607584 941107 607652 941159
rect 607708 941107 607776 941159
rect 607832 941107 607900 941159
rect 607460 941103 607473 941107
rect 607584 941103 607615 941107
rect 607708 941103 607757 941107
rect 607832 941103 607899 941107
rect 607956 941103 608024 941159
rect 608080 941107 608148 941159
rect 608204 941107 608272 941159
rect 608328 941107 608396 941159
rect 608097 941103 608148 941107
rect 608239 941103 608272 941107
rect 608381 941103 608396 941107
rect 608452 941107 608520 941159
rect 608576 941107 608644 941159
rect 608700 941107 608768 941159
rect 608452 941103 608467 941107
rect 608576 941103 608609 941107
rect 608700 941103 608751 941107
rect 608824 941103 608878 941159
rect 606961 941051 607047 941103
rect 607103 941051 607189 941103
rect 607245 941051 607331 941103
rect 607387 941051 607473 941103
rect 607529 941051 607615 941103
rect 607671 941051 607757 941103
rect 607813 941051 607899 941103
rect 607955 941051 608041 941103
rect 608097 941051 608183 941103
rect 608239 941051 608325 941103
rect 608381 941051 608467 941103
rect 608523 941051 608609 941103
rect 608665 941051 608751 941103
rect 608807 941051 608878 941103
rect 606828 941035 608878 941051
rect 606828 940979 606908 941035
rect 606964 940979 607032 941035
rect 607088 940979 607156 941035
rect 607212 940979 607280 941035
rect 607336 940979 607404 941035
rect 607460 940979 607528 941035
rect 607584 940979 607652 941035
rect 607708 940979 607776 941035
rect 607832 940979 607900 941035
rect 607956 940979 608024 941035
rect 608080 940979 608148 941035
rect 608204 940979 608272 941035
rect 608328 940979 608396 941035
rect 608452 940979 608520 941035
rect 608576 940979 608644 941035
rect 608700 940979 608768 941035
rect 608824 940979 608878 941035
rect 606828 940965 608878 940979
rect 606828 940909 606905 940965
rect 606961 940911 607047 940965
rect 607103 940911 607189 940965
rect 607245 940911 607331 940965
rect 607387 940911 607473 940965
rect 607529 940911 607615 940965
rect 607671 940911 607757 940965
rect 607813 940911 607899 940965
rect 607955 940911 608041 940965
rect 608097 940911 608183 940965
rect 608239 940911 608325 940965
rect 608381 940911 608467 940965
rect 608523 940911 608609 940965
rect 608665 940911 608751 940965
rect 608807 940911 608878 940965
rect 606828 940855 606908 940909
rect 606964 940855 607032 940911
rect 607103 940909 607156 940911
rect 607245 940909 607280 940911
rect 607387 940909 607404 940911
rect 607088 940855 607156 940909
rect 607212 940855 607280 940909
rect 607336 940855 607404 940909
rect 607460 940909 607473 940911
rect 607584 940909 607615 940911
rect 607708 940909 607757 940911
rect 607832 940909 607899 940911
rect 607460 940855 607528 940909
rect 607584 940855 607652 940909
rect 607708 940855 607776 940909
rect 607832 940855 607900 940909
rect 607956 940855 608024 940911
rect 608097 940909 608148 940911
rect 608239 940909 608272 940911
rect 608381 940909 608396 940911
rect 608080 940855 608148 940909
rect 608204 940855 608272 940909
rect 608328 940855 608396 940909
rect 608452 940909 608467 940911
rect 608576 940909 608609 940911
rect 608700 940909 608751 940911
rect 608452 940855 608520 940909
rect 608576 940855 608644 940909
rect 608700 940855 608768 940909
rect 608824 940855 608878 940911
rect 606828 940823 608878 940855
rect 606828 940767 606905 940823
rect 606961 940787 607047 940823
rect 607103 940787 607189 940823
rect 607245 940787 607331 940823
rect 607387 940787 607473 940823
rect 607529 940787 607615 940823
rect 607671 940787 607757 940823
rect 607813 940787 607899 940823
rect 607955 940787 608041 940823
rect 608097 940787 608183 940823
rect 608239 940787 608325 940823
rect 608381 940787 608467 940823
rect 608523 940787 608609 940823
rect 608665 940787 608751 940823
rect 608807 940787 608878 940823
rect 606828 940731 606908 940767
rect 606964 940731 607032 940787
rect 607103 940767 607156 940787
rect 607245 940767 607280 940787
rect 607387 940767 607404 940787
rect 607088 940731 607156 940767
rect 607212 940731 607280 940767
rect 607336 940731 607404 940767
rect 607460 940767 607473 940787
rect 607584 940767 607615 940787
rect 607708 940767 607757 940787
rect 607832 940767 607899 940787
rect 607460 940731 607528 940767
rect 607584 940731 607652 940767
rect 607708 940731 607776 940767
rect 607832 940731 607900 940767
rect 607956 940731 608024 940787
rect 608097 940767 608148 940787
rect 608239 940767 608272 940787
rect 608381 940767 608396 940787
rect 608080 940731 608148 940767
rect 608204 940731 608272 940767
rect 608328 940731 608396 940767
rect 608452 940767 608467 940787
rect 608576 940767 608609 940787
rect 608700 940767 608751 940787
rect 608452 940731 608520 940767
rect 608576 940731 608644 940767
rect 608700 940731 608768 940767
rect 608824 940731 608878 940787
rect 606828 940681 608878 940731
rect 606828 940625 606905 940681
rect 606961 940663 607047 940681
rect 607103 940663 607189 940681
rect 607245 940663 607331 940681
rect 607387 940663 607473 940681
rect 607529 940663 607615 940681
rect 607671 940663 607757 940681
rect 607813 940663 607899 940681
rect 607955 940663 608041 940681
rect 608097 940663 608183 940681
rect 608239 940663 608325 940681
rect 608381 940663 608467 940681
rect 608523 940663 608609 940681
rect 608665 940663 608751 940681
rect 608807 940663 608878 940681
rect 606828 940607 606908 940625
rect 606964 940607 607032 940663
rect 607103 940625 607156 940663
rect 607245 940625 607280 940663
rect 607387 940625 607404 940663
rect 607088 940607 607156 940625
rect 607212 940607 607280 940625
rect 607336 940607 607404 940625
rect 607460 940625 607473 940663
rect 607584 940625 607615 940663
rect 607708 940625 607757 940663
rect 607832 940625 607899 940663
rect 607460 940607 607528 940625
rect 607584 940607 607652 940625
rect 607708 940607 607776 940625
rect 607832 940607 607900 940625
rect 607956 940607 608024 940663
rect 608097 940625 608148 940663
rect 608239 940625 608272 940663
rect 608381 940625 608396 940663
rect 608080 940607 608148 940625
rect 608204 940607 608272 940625
rect 608328 940607 608396 940625
rect 608452 940625 608467 940663
rect 608576 940625 608609 940663
rect 608700 940625 608751 940663
rect 608452 940607 608520 940625
rect 608576 940607 608644 940625
rect 608700 940607 608768 940625
rect 608824 940607 608878 940663
rect 606828 940539 608878 940607
rect 606828 940483 606905 940539
rect 606964 940483 607032 940539
rect 607103 940483 607156 940539
rect 607245 940483 607280 940539
rect 607387 940483 607404 940539
rect 607460 940483 607473 940539
rect 607584 940483 607615 940539
rect 607708 940483 607757 940539
rect 607832 940483 607899 940539
rect 607956 940483 608024 940539
rect 608097 940483 608148 940539
rect 608239 940483 608272 940539
rect 608381 940483 608396 940539
rect 608452 940483 608467 940539
rect 608576 940483 608609 940539
rect 608700 940483 608751 940539
rect 608824 940483 608878 940539
rect 606828 940415 608878 940483
rect 606828 940397 606908 940415
rect 606828 940341 606905 940397
rect 606964 940359 607032 940415
rect 607088 940397 607156 940415
rect 607212 940397 607280 940415
rect 607336 940397 607404 940415
rect 607103 940359 607156 940397
rect 607245 940359 607280 940397
rect 607387 940359 607404 940397
rect 607460 940397 607528 940415
rect 607584 940397 607652 940415
rect 607708 940397 607776 940415
rect 607832 940397 607900 940415
rect 607460 940359 607473 940397
rect 607584 940359 607615 940397
rect 607708 940359 607757 940397
rect 607832 940359 607899 940397
rect 607956 940359 608024 940415
rect 608080 940397 608148 940415
rect 608204 940397 608272 940415
rect 608328 940397 608396 940415
rect 608097 940359 608148 940397
rect 608239 940359 608272 940397
rect 608381 940359 608396 940397
rect 608452 940397 608520 940415
rect 608576 940397 608644 940415
rect 608700 940397 608768 940415
rect 608452 940359 608467 940397
rect 608576 940359 608609 940397
rect 608700 940359 608751 940397
rect 608824 940359 608878 940415
rect 606961 940341 607047 940359
rect 607103 940341 607189 940359
rect 607245 940341 607331 940359
rect 607387 940341 607473 940359
rect 607529 940341 607615 940359
rect 607671 940341 607757 940359
rect 607813 940341 607899 940359
rect 607955 940341 608041 940359
rect 608097 940341 608183 940359
rect 608239 940341 608325 940359
rect 608381 940341 608467 940359
rect 608523 940341 608609 940359
rect 608665 940341 608751 940359
rect 608807 940341 608878 940359
rect 606828 940291 608878 940341
rect 606828 940255 606908 940291
rect 606828 940199 606905 940255
rect 606964 940235 607032 940291
rect 607088 940255 607156 940291
rect 607212 940255 607280 940291
rect 607336 940255 607404 940291
rect 607103 940235 607156 940255
rect 607245 940235 607280 940255
rect 607387 940235 607404 940255
rect 607460 940255 607528 940291
rect 607584 940255 607652 940291
rect 607708 940255 607776 940291
rect 607832 940255 607900 940291
rect 607460 940235 607473 940255
rect 607584 940235 607615 940255
rect 607708 940235 607757 940255
rect 607832 940235 607899 940255
rect 607956 940235 608024 940291
rect 608080 940255 608148 940291
rect 608204 940255 608272 940291
rect 608328 940255 608396 940291
rect 608097 940235 608148 940255
rect 608239 940235 608272 940255
rect 608381 940235 608396 940255
rect 608452 940255 608520 940291
rect 608576 940255 608644 940291
rect 608700 940255 608768 940291
rect 608452 940235 608467 940255
rect 608576 940235 608609 940255
rect 608700 940235 608751 940255
rect 608824 940235 608878 940291
rect 606961 940199 607047 940235
rect 607103 940199 607189 940235
rect 607245 940199 607331 940235
rect 607387 940199 607473 940235
rect 607529 940199 607615 940235
rect 607671 940199 607757 940235
rect 607813 940199 607899 940235
rect 607955 940199 608041 940235
rect 608097 940199 608183 940235
rect 608239 940199 608325 940235
rect 608381 940199 608467 940235
rect 608523 940199 608609 940235
rect 608665 940199 608751 940235
rect 608807 940199 608878 940235
rect 606828 940167 608878 940199
rect 606828 940113 606908 940167
rect 606828 940057 606905 940113
rect 606964 940111 607032 940167
rect 607088 940113 607156 940167
rect 607212 940113 607280 940167
rect 607336 940113 607404 940167
rect 607103 940111 607156 940113
rect 607245 940111 607280 940113
rect 607387 940111 607404 940113
rect 607460 940113 607528 940167
rect 607584 940113 607652 940167
rect 607708 940113 607776 940167
rect 607832 940113 607900 940167
rect 607460 940111 607473 940113
rect 607584 940111 607615 940113
rect 607708 940111 607757 940113
rect 607832 940111 607899 940113
rect 607956 940111 608024 940167
rect 608080 940113 608148 940167
rect 608204 940113 608272 940167
rect 608328 940113 608396 940167
rect 608097 940111 608148 940113
rect 608239 940111 608272 940113
rect 608381 940111 608396 940113
rect 608452 940113 608520 940167
rect 608576 940113 608644 940167
rect 608700 940113 608768 940167
rect 608452 940111 608467 940113
rect 608576 940111 608609 940113
rect 608700 940111 608751 940113
rect 608824 940111 608878 940167
rect 606961 940057 607047 940111
rect 607103 940057 607189 940111
rect 607245 940057 607331 940111
rect 607387 940057 607473 940111
rect 607529 940057 607615 940111
rect 607671 940057 607757 940111
rect 607813 940057 607899 940111
rect 607955 940057 608041 940111
rect 608097 940057 608183 940111
rect 608239 940057 608325 940111
rect 608381 940057 608467 940111
rect 608523 940057 608609 940111
rect 608665 940057 608751 940111
rect 608807 940057 608878 940111
rect 606828 940043 608878 940057
rect 606828 939987 606908 940043
rect 606964 939987 607032 940043
rect 607088 939987 607156 940043
rect 607212 939987 607280 940043
rect 607336 939987 607404 940043
rect 607460 939987 607528 940043
rect 607584 939987 607652 940043
rect 607708 939987 607776 940043
rect 607832 939987 607900 940043
rect 607956 939987 608024 940043
rect 608080 939987 608148 940043
rect 608204 939987 608272 940043
rect 608328 939987 608396 940043
rect 608452 939987 608520 940043
rect 608576 939987 608644 940043
rect 608700 939987 608768 940043
rect 608824 939987 608878 940043
rect 606828 939971 608878 939987
rect 606828 939915 606905 939971
rect 606961 939919 607047 939971
rect 607103 939919 607189 939971
rect 607245 939919 607331 939971
rect 607387 939919 607473 939971
rect 607529 939919 607615 939971
rect 607671 939919 607757 939971
rect 607813 939919 607899 939971
rect 607955 939919 608041 939971
rect 608097 939919 608183 939971
rect 608239 939919 608325 939971
rect 608381 939919 608467 939971
rect 608523 939919 608609 939971
rect 608665 939919 608751 939971
rect 608807 939919 608878 939971
rect 606828 939863 606908 939915
rect 606964 939863 607032 939919
rect 607103 939915 607156 939919
rect 607245 939915 607280 939919
rect 607387 939915 607404 939919
rect 607088 939863 607156 939915
rect 607212 939863 607280 939915
rect 607336 939863 607404 939915
rect 607460 939915 607473 939919
rect 607584 939915 607615 939919
rect 607708 939915 607757 939919
rect 607832 939915 607899 939919
rect 607460 939863 607528 939915
rect 607584 939863 607652 939915
rect 607708 939863 607776 939915
rect 607832 939863 607900 939915
rect 607956 939863 608024 939919
rect 608097 939915 608148 939919
rect 608239 939915 608272 939919
rect 608381 939915 608396 939919
rect 608080 939863 608148 939915
rect 608204 939863 608272 939915
rect 608328 939863 608396 939915
rect 608452 939915 608467 939919
rect 608576 939915 608609 939919
rect 608700 939915 608751 939919
rect 608452 939863 608520 939915
rect 608576 939863 608644 939915
rect 608700 939863 608768 939915
rect 608824 939863 608878 939919
rect 606828 939829 608878 939863
rect 606828 939773 606905 939829
rect 606961 939773 607047 939829
rect 607103 939773 607189 939829
rect 607245 939773 607331 939829
rect 607387 939773 607473 939829
rect 607529 939773 607615 939829
rect 607671 939773 607757 939829
rect 607813 939773 607899 939829
rect 607955 939773 608041 939829
rect 608097 939773 608183 939829
rect 608239 939773 608325 939829
rect 608381 939773 608467 939829
rect 608523 939773 608609 939829
rect 608665 939773 608751 939829
rect 608807 939773 608878 939829
rect 606828 939720 608878 939773
rect 609198 941675 611248 941720
rect 609198 941619 609275 941675
rect 609331 941655 609417 941675
rect 609473 941655 609559 941675
rect 609615 941655 609701 941675
rect 609757 941655 609843 941675
rect 609899 941655 609985 941675
rect 610041 941655 610127 941675
rect 610183 941655 610269 941675
rect 610325 941655 610411 941675
rect 610467 941655 610553 941675
rect 610609 941655 610695 941675
rect 610751 941655 610837 941675
rect 610893 941655 610979 941675
rect 611035 941655 611121 941675
rect 611177 941655 611248 941675
rect 609198 941599 609278 941619
rect 609334 941599 609402 941655
rect 609473 941619 609526 941655
rect 609615 941619 609650 941655
rect 609757 941619 609774 941655
rect 609458 941599 609526 941619
rect 609582 941599 609650 941619
rect 609706 941599 609774 941619
rect 609830 941619 609843 941655
rect 609954 941619 609985 941655
rect 610078 941619 610127 941655
rect 610202 941619 610269 941655
rect 609830 941599 609898 941619
rect 609954 941599 610022 941619
rect 610078 941599 610146 941619
rect 610202 941599 610270 941619
rect 610326 941599 610394 941655
rect 610467 941619 610518 941655
rect 610609 941619 610642 941655
rect 610751 941619 610766 941655
rect 610450 941599 610518 941619
rect 610574 941599 610642 941619
rect 610698 941599 610766 941619
rect 610822 941619 610837 941655
rect 610946 941619 610979 941655
rect 611070 941619 611121 941655
rect 610822 941599 610890 941619
rect 610946 941599 611014 941619
rect 611070 941599 611138 941619
rect 611194 941599 611248 941655
rect 609198 941533 611248 941599
rect 609198 941477 609275 941533
rect 609331 941531 609417 941533
rect 609473 941531 609559 941533
rect 609615 941531 609701 941533
rect 609757 941531 609843 941533
rect 609899 941531 609985 941533
rect 610041 941531 610127 941533
rect 610183 941531 610269 941533
rect 610325 941531 610411 941533
rect 610467 941531 610553 941533
rect 610609 941531 610695 941533
rect 610751 941531 610837 941533
rect 610893 941531 610979 941533
rect 611035 941531 611121 941533
rect 611177 941531 611248 941533
rect 609198 941475 609278 941477
rect 609334 941475 609402 941531
rect 609473 941477 609526 941531
rect 609615 941477 609650 941531
rect 609757 941477 609774 941531
rect 609458 941475 609526 941477
rect 609582 941475 609650 941477
rect 609706 941475 609774 941477
rect 609830 941477 609843 941531
rect 609954 941477 609985 941531
rect 610078 941477 610127 941531
rect 610202 941477 610269 941531
rect 609830 941475 609898 941477
rect 609954 941475 610022 941477
rect 610078 941475 610146 941477
rect 610202 941475 610270 941477
rect 610326 941475 610394 941531
rect 610467 941477 610518 941531
rect 610609 941477 610642 941531
rect 610751 941477 610766 941531
rect 610450 941475 610518 941477
rect 610574 941475 610642 941477
rect 610698 941475 610766 941477
rect 610822 941477 610837 941531
rect 610946 941477 610979 941531
rect 611070 941477 611121 941531
rect 610822 941475 610890 941477
rect 610946 941475 611014 941477
rect 611070 941475 611138 941477
rect 611194 941475 611248 941531
rect 609198 941407 611248 941475
rect 609198 941391 609278 941407
rect 609198 941335 609275 941391
rect 609334 941351 609402 941407
rect 609458 941391 609526 941407
rect 609582 941391 609650 941407
rect 609706 941391 609774 941407
rect 609473 941351 609526 941391
rect 609615 941351 609650 941391
rect 609757 941351 609774 941391
rect 609830 941391 609898 941407
rect 609954 941391 610022 941407
rect 610078 941391 610146 941407
rect 610202 941391 610270 941407
rect 609830 941351 609843 941391
rect 609954 941351 609985 941391
rect 610078 941351 610127 941391
rect 610202 941351 610269 941391
rect 610326 941351 610394 941407
rect 610450 941391 610518 941407
rect 610574 941391 610642 941407
rect 610698 941391 610766 941407
rect 610467 941351 610518 941391
rect 610609 941351 610642 941391
rect 610751 941351 610766 941391
rect 610822 941391 610890 941407
rect 610946 941391 611014 941407
rect 611070 941391 611138 941407
rect 610822 941351 610837 941391
rect 610946 941351 610979 941391
rect 611070 941351 611121 941391
rect 611194 941351 611248 941407
rect 609331 941335 609417 941351
rect 609473 941335 609559 941351
rect 609615 941335 609701 941351
rect 609757 941335 609843 941351
rect 609899 941335 609985 941351
rect 610041 941335 610127 941351
rect 610183 941335 610269 941351
rect 610325 941335 610411 941351
rect 610467 941335 610553 941351
rect 610609 941335 610695 941351
rect 610751 941335 610837 941351
rect 610893 941335 610979 941351
rect 611035 941335 611121 941351
rect 611177 941335 611248 941351
rect 609198 941283 611248 941335
rect 609198 941249 609278 941283
rect 609198 941193 609275 941249
rect 609334 941227 609402 941283
rect 609458 941249 609526 941283
rect 609582 941249 609650 941283
rect 609706 941249 609774 941283
rect 609473 941227 609526 941249
rect 609615 941227 609650 941249
rect 609757 941227 609774 941249
rect 609830 941249 609898 941283
rect 609954 941249 610022 941283
rect 610078 941249 610146 941283
rect 610202 941249 610270 941283
rect 609830 941227 609843 941249
rect 609954 941227 609985 941249
rect 610078 941227 610127 941249
rect 610202 941227 610269 941249
rect 610326 941227 610394 941283
rect 610450 941249 610518 941283
rect 610574 941249 610642 941283
rect 610698 941249 610766 941283
rect 610467 941227 610518 941249
rect 610609 941227 610642 941249
rect 610751 941227 610766 941249
rect 610822 941249 610890 941283
rect 610946 941249 611014 941283
rect 611070 941249 611138 941283
rect 610822 941227 610837 941249
rect 610946 941227 610979 941249
rect 611070 941227 611121 941249
rect 611194 941227 611248 941283
rect 609331 941193 609417 941227
rect 609473 941193 609559 941227
rect 609615 941193 609701 941227
rect 609757 941193 609843 941227
rect 609899 941193 609985 941227
rect 610041 941193 610127 941227
rect 610183 941193 610269 941227
rect 610325 941193 610411 941227
rect 610467 941193 610553 941227
rect 610609 941193 610695 941227
rect 610751 941193 610837 941227
rect 610893 941193 610979 941227
rect 611035 941193 611121 941227
rect 611177 941193 611248 941227
rect 609198 941159 611248 941193
rect 609198 941107 609278 941159
rect 609198 941051 609275 941107
rect 609334 941103 609402 941159
rect 609458 941107 609526 941159
rect 609582 941107 609650 941159
rect 609706 941107 609774 941159
rect 609473 941103 609526 941107
rect 609615 941103 609650 941107
rect 609757 941103 609774 941107
rect 609830 941107 609898 941159
rect 609954 941107 610022 941159
rect 610078 941107 610146 941159
rect 610202 941107 610270 941159
rect 609830 941103 609843 941107
rect 609954 941103 609985 941107
rect 610078 941103 610127 941107
rect 610202 941103 610269 941107
rect 610326 941103 610394 941159
rect 610450 941107 610518 941159
rect 610574 941107 610642 941159
rect 610698 941107 610766 941159
rect 610467 941103 610518 941107
rect 610609 941103 610642 941107
rect 610751 941103 610766 941107
rect 610822 941107 610890 941159
rect 610946 941107 611014 941159
rect 611070 941107 611138 941159
rect 610822 941103 610837 941107
rect 610946 941103 610979 941107
rect 611070 941103 611121 941107
rect 611194 941103 611248 941159
rect 609331 941051 609417 941103
rect 609473 941051 609559 941103
rect 609615 941051 609701 941103
rect 609757 941051 609843 941103
rect 609899 941051 609985 941103
rect 610041 941051 610127 941103
rect 610183 941051 610269 941103
rect 610325 941051 610411 941103
rect 610467 941051 610553 941103
rect 610609 941051 610695 941103
rect 610751 941051 610837 941103
rect 610893 941051 610979 941103
rect 611035 941051 611121 941103
rect 611177 941051 611248 941103
rect 609198 941035 611248 941051
rect 609198 940979 609278 941035
rect 609334 940979 609402 941035
rect 609458 940979 609526 941035
rect 609582 940979 609650 941035
rect 609706 940979 609774 941035
rect 609830 940979 609898 941035
rect 609954 940979 610022 941035
rect 610078 940979 610146 941035
rect 610202 940979 610270 941035
rect 610326 940979 610394 941035
rect 610450 940979 610518 941035
rect 610574 940979 610642 941035
rect 610698 940979 610766 941035
rect 610822 940979 610890 941035
rect 610946 940979 611014 941035
rect 611070 940979 611138 941035
rect 611194 940979 611248 941035
rect 609198 940965 611248 940979
rect 609198 940909 609275 940965
rect 609331 940911 609417 940965
rect 609473 940911 609559 940965
rect 609615 940911 609701 940965
rect 609757 940911 609843 940965
rect 609899 940911 609985 940965
rect 610041 940911 610127 940965
rect 610183 940911 610269 940965
rect 610325 940911 610411 940965
rect 610467 940911 610553 940965
rect 610609 940911 610695 940965
rect 610751 940911 610837 940965
rect 610893 940911 610979 940965
rect 611035 940911 611121 940965
rect 611177 940911 611248 940965
rect 609198 940855 609278 940909
rect 609334 940855 609402 940911
rect 609473 940909 609526 940911
rect 609615 940909 609650 940911
rect 609757 940909 609774 940911
rect 609458 940855 609526 940909
rect 609582 940855 609650 940909
rect 609706 940855 609774 940909
rect 609830 940909 609843 940911
rect 609954 940909 609985 940911
rect 610078 940909 610127 940911
rect 610202 940909 610269 940911
rect 609830 940855 609898 940909
rect 609954 940855 610022 940909
rect 610078 940855 610146 940909
rect 610202 940855 610270 940909
rect 610326 940855 610394 940911
rect 610467 940909 610518 940911
rect 610609 940909 610642 940911
rect 610751 940909 610766 940911
rect 610450 940855 610518 940909
rect 610574 940855 610642 940909
rect 610698 940855 610766 940909
rect 610822 940909 610837 940911
rect 610946 940909 610979 940911
rect 611070 940909 611121 940911
rect 610822 940855 610890 940909
rect 610946 940855 611014 940909
rect 611070 940855 611138 940909
rect 611194 940855 611248 940911
rect 609198 940823 611248 940855
rect 609198 940767 609275 940823
rect 609331 940787 609417 940823
rect 609473 940787 609559 940823
rect 609615 940787 609701 940823
rect 609757 940787 609843 940823
rect 609899 940787 609985 940823
rect 610041 940787 610127 940823
rect 610183 940787 610269 940823
rect 610325 940787 610411 940823
rect 610467 940787 610553 940823
rect 610609 940787 610695 940823
rect 610751 940787 610837 940823
rect 610893 940787 610979 940823
rect 611035 940787 611121 940823
rect 611177 940787 611248 940823
rect 609198 940731 609278 940767
rect 609334 940731 609402 940787
rect 609473 940767 609526 940787
rect 609615 940767 609650 940787
rect 609757 940767 609774 940787
rect 609458 940731 609526 940767
rect 609582 940731 609650 940767
rect 609706 940731 609774 940767
rect 609830 940767 609843 940787
rect 609954 940767 609985 940787
rect 610078 940767 610127 940787
rect 610202 940767 610269 940787
rect 609830 940731 609898 940767
rect 609954 940731 610022 940767
rect 610078 940731 610146 940767
rect 610202 940731 610270 940767
rect 610326 940731 610394 940787
rect 610467 940767 610518 940787
rect 610609 940767 610642 940787
rect 610751 940767 610766 940787
rect 610450 940731 610518 940767
rect 610574 940731 610642 940767
rect 610698 940731 610766 940767
rect 610822 940767 610837 940787
rect 610946 940767 610979 940787
rect 611070 940767 611121 940787
rect 610822 940731 610890 940767
rect 610946 940731 611014 940767
rect 611070 940731 611138 940767
rect 611194 940731 611248 940787
rect 609198 940681 611248 940731
rect 609198 940625 609275 940681
rect 609331 940663 609417 940681
rect 609473 940663 609559 940681
rect 609615 940663 609701 940681
rect 609757 940663 609843 940681
rect 609899 940663 609985 940681
rect 610041 940663 610127 940681
rect 610183 940663 610269 940681
rect 610325 940663 610411 940681
rect 610467 940663 610553 940681
rect 610609 940663 610695 940681
rect 610751 940663 610837 940681
rect 610893 940663 610979 940681
rect 611035 940663 611121 940681
rect 611177 940663 611248 940681
rect 609198 940607 609278 940625
rect 609334 940607 609402 940663
rect 609473 940625 609526 940663
rect 609615 940625 609650 940663
rect 609757 940625 609774 940663
rect 609458 940607 609526 940625
rect 609582 940607 609650 940625
rect 609706 940607 609774 940625
rect 609830 940625 609843 940663
rect 609954 940625 609985 940663
rect 610078 940625 610127 940663
rect 610202 940625 610269 940663
rect 609830 940607 609898 940625
rect 609954 940607 610022 940625
rect 610078 940607 610146 940625
rect 610202 940607 610270 940625
rect 610326 940607 610394 940663
rect 610467 940625 610518 940663
rect 610609 940625 610642 940663
rect 610751 940625 610766 940663
rect 610450 940607 610518 940625
rect 610574 940607 610642 940625
rect 610698 940607 610766 940625
rect 610822 940625 610837 940663
rect 610946 940625 610979 940663
rect 611070 940625 611121 940663
rect 610822 940607 610890 940625
rect 610946 940607 611014 940625
rect 611070 940607 611138 940625
rect 611194 940607 611248 940663
rect 609198 940539 611248 940607
rect 609198 940483 609275 940539
rect 609334 940483 609402 940539
rect 609473 940483 609526 940539
rect 609615 940483 609650 940539
rect 609757 940483 609774 940539
rect 609830 940483 609843 940539
rect 609954 940483 609985 940539
rect 610078 940483 610127 940539
rect 610202 940483 610269 940539
rect 610326 940483 610394 940539
rect 610467 940483 610518 940539
rect 610609 940483 610642 940539
rect 610751 940483 610766 940539
rect 610822 940483 610837 940539
rect 610946 940483 610979 940539
rect 611070 940483 611121 940539
rect 611194 940483 611248 940539
rect 609198 940415 611248 940483
rect 609198 940397 609278 940415
rect 609198 940341 609275 940397
rect 609334 940359 609402 940415
rect 609458 940397 609526 940415
rect 609582 940397 609650 940415
rect 609706 940397 609774 940415
rect 609473 940359 609526 940397
rect 609615 940359 609650 940397
rect 609757 940359 609774 940397
rect 609830 940397 609898 940415
rect 609954 940397 610022 940415
rect 610078 940397 610146 940415
rect 610202 940397 610270 940415
rect 609830 940359 609843 940397
rect 609954 940359 609985 940397
rect 610078 940359 610127 940397
rect 610202 940359 610269 940397
rect 610326 940359 610394 940415
rect 610450 940397 610518 940415
rect 610574 940397 610642 940415
rect 610698 940397 610766 940415
rect 610467 940359 610518 940397
rect 610609 940359 610642 940397
rect 610751 940359 610766 940397
rect 610822 940397 610890 940415
rect 610946 940397 611014 940415
rect 611070 940397 611138 940415
rect 610822 940359 610837 940397
rect 610946 940359 610979 940397
rect 611070 940359 611121 940397
rect 611194 940359 611248 940415
rect 609331 940341 609417 940359
rect 609473 940341 609559 940359
rect 609615 940341 609701 940359
rect 609757 940341 609843 940359
rect 609899 940341 609985 940359
rect 610041 940341 610127 940359
rect 610183 940341 610269 940359
rect 610325 940341 610411 940359
rect 610467 940341 610553 940359
rect 610609 940341 610695 940359
rect 610751 940341 610837 940359
rect 610893 940341 610979 940359
rect 611035 940341 611121 940359
rect 611177 940341 611248 940359
rect 609198 940291 611248 940341
rect 609198 940255 609278 940291
rect 609198 940199 609275 940255
rect 609334 940235 609402 940291
rect 609458 940255 609526 940291
rect 609582 940255 609650 940291
rect 609706 940255 609774 940291
rect 609473 940235 609526 940255
rect 609615 940235 609650 940255
rect 609757 940235 609774 940255
rect 609830 940255 609898 940291
rect 609954 940255 610022 940291
rect 610078 940255 610146 940291
rect 610202 940255 610270 940291
rect 609830 940235 609843 940255
rect 609954 940235 609985 940255
rect 610078 940235 610127 940255
rect 610202 940235 610269 940255
rect 610326 940235 610394 940291
rect 610450 940255 610518 940291
rect 610574 940255 610642 940291
rect 610698 940255 610766 940291
rect 610467 940235 610518 940255
rect 610609 940235 610642 940255
rect 610751 940235 610766 940255
rect 610822 940255 610890 940291
rect 610946 940255 611014 940291
rect 611070 940255 611138 940291
rect 610822 940235 610837 940255
rect 610946 940235 610979 940255
rect 611070 940235 611121 940255
rect 611194 940235 611248 940291
rect 609331 940199 609417 940235
rect 609473 940199 609559 940235
rect 609615 940199 609701 940235
rect 609757 940199 609843 940235
rect 609899 940199 609985 940235
rect 610041 940199 610127 940235
rect 610183 940199 610269 940235
rect 610325 940199 610411 940235
rect 610467 940199 610553 940235
rect 610609 940199 610695 940235
rect 610751 940199 610837 940235
rect 610893 940199 610979 940235
rect 611035 940199 611121 940235
rect 611177 940199 611248 940235
rect 609198 940167 611248 940199
rect 609198 940113 609278 940167
rect 609198 940057 609275 940113
rect 609334 940111 609402 940167
rect 609458 940113 609526 940167
rect 609582 940113 609650 940167
rect 609706 940113 609774 940167
rect 609473 940111 609526 940113
rect 609615 940111 609650 940113
rect 609757 940111 609774 940113
rect 609830 940113 609898 940167
rect 609954 940113 610022 940167
rect 610078 940113 610146 940167
rect 610202 940113 610270 940167
rect 609830 940111 609843 940113
rect 609954 940111 609985 940113
rect 610078 940111 610127 940113
rect 610202 940111 610269 940113
rect 610326 940111 610394 940167
rect 610450 940113 610518 940167
rect 610574 940113 610642 940167
rect 610698 940113 610766 940167
rect 610467 940111 610518 940113
rect 610609 940111 610642 940113
rect 610751 940111 610766 940113
rect 610822 940113 610890 940167
rect 610946 940113 611014 940167
rect 611070 940113 611138 940167
rect 610822 940111 610837 940113
rect 610946 940111 610979 940113
rect 611070 940111 611121 940113
rect 611194 940111 611248 940167
rect 609331 940057 609417 940111
rect 609473 940057 609559 940111
rect 609615 940057 609701 940111
rect 609757 940057 609843 940111
rect 609899 940057 609985 940111
rect 610041 940057 610127 940111
rect 610183 940057 610269 940111
rect 610325 940057 610411 940111
rect 610467 940057 610553 940111
rect 610609 940057 610695 940111
rect 610751 940057 610837 940111
rect 610893 940057 610979 940111
rect 611035 940057 611121 940111
rect 611177 940057 611248 940111
rect 609198 940043 611248 940057
rect 609198 939987 609278 940043
rect 609334 939987 609402 940043
rect 609458 939987 609526 940043
rect 609582 939987 609650 940043
rect 609706 939987 609774 940043
rect 609830 939987 609898 940043
rect 609954 939987 610022 940043
rect 610078 939987 610146 940043
rect 610202 939987 610270 940043
rect 610326 939987 610394 940043
rect 610450 939987 610518 940043
rect 610574 939987 610642 940043
rect 610698 939987 610766 940043
rect 610822 939987 610890 940043
rect 610946 939987 611014 940043
rect 611070 939987 611138 940043
rect 611194 939987 611248 940043
rect 609198 939971 611248 939987
rect 609198 939915 609275 939971
rect 609331 939919 609417 939971
rect 609473 939919 609559 939971
rect 609615 939919 609701 939971
rect 609757 939919 609843 939971
rect 609899 939919 609985 939971
rect 610041 939919 610127 939971
rect 610183 939919 610269 939971
rect 610325 939919 610411 939971
rect 610467 939919 610553 939971
rect 610609 939919 610695 939971
rect 610751 939919 610837 939971
rect 610893 939919 610979 939971
rect 611035 939919 611121 939971
rect 611177 939919 611248 939971
rect 609198 939863 609278 939915
rect 609334 939863 609402 939919
rect 609473 939915 609526 939919
rect 609615 939915 609650 939919
rect 609757 939915 609774 939919
rect 609458 939863 609526 939915
rect 609582 939863 609650 939915
rect 609706 939863 609774 939915
rect 609830 939915 609843 939919
rect 609954 939915 609985 939919
rect 610078 939915 610127 939919
rect 610202 939915 610269 939919
rect 609830 939863 609898 939915
rect 609954 939863 610022 939915
rect 610078 939863 610146 939915
rect 610202 939863 610270 939915
rect 610326 939863 610394 939919
rect 610467 939915 610518 939919
rect 610609 939915 610642 939919
rect 610751 939915 610766 939919
rect 610450 939863 610518 939915
rect 610574 939863 610642 939915
rect 610698 939863 610766 939915
rect 610822 939915 610837 939919
rect 610946 939915 610979 939919
rect 611070 939915 611121 939919
rect 610822 939863 610890 939915
rect 610946 939863 611014 939915
rect 611070 939863 611138 939915
rect 611194 939863 611248 939919
rect 609198 939829 611248 939863
rect 609198 939773 609275 939829
rect 609331 939773 609417 939829
rect 609473 939773 609559 939829
rect 609615 939773 609701 939829
rect 609757 939773 609843 939829
rect 609899 939773 609985 939829
rect 610041 939773 610127 939829
rect 610183 939773 610269 939829
rect 610325 939773 610411 939829
rect 610467 939773 610553 939829
rect 610609 939773 610695 939829
rect 610751 939773 610837 939829
rect 610893 939773 610979 939829
rect 611035 939773 611121 939829
rect 611177 939773 611248 939829
rect 609198 939720 611248 939773
rect 611828 941675 613728 941720
rect 611828 941655 611897 941675
rect 611953 941655 612039 941675
rect 612095 941655 612181 941675
rect 612237 941655 612323 941675
rect 612379 941655 612465 941675
rect 612521 941655 612607 941675
rect 612663 941655 612749 941675
rect 612805 941655 612891 941675
rect 612947 941655 613033 941675
rect 613089 941655 613175 941675
rect 613231 941655 613317 941675
rect 613373 941655 613459 941675
rect 613515 941655 613601 941675
rect 613657 941655 613728 941675
rect 611828 941599 611882 941655
rect 611953 941619 612006 941655
rect 612095 941619 612130 941655
rect 612237 941619 612254 941655
rect 611938 941599 612006 941619
rect 612062 941599 612130 941619
rect 612186 941599 612254 941619
rect 612310 941619 612323 941655
rect 612434 941619 612465 941655
rect 612558 941619 612607 941655
rect 612682 941619 612749 941655
rect 612310 941599 612378 941619
rect 612434 941599 612502 941619
rect 612558 941599 612626 941619
rect 612682 941599 612750 941619
rect 612806 941599 612874 941655
rect 612947 941619 612998 941655
rect 613089 941619 613122 941655
rect 613231 941619 613246 941655
rect 612930 941599 612998 941619
rect 613054 941599 613122 941619
rect 613178 941599 613246 941619
rect 613302 941619 613317 941655
rect 613426 941619 613459 941655
rect 613550 941619 613601 941655
rect 613302 941599 613370 941619
rect 613426 941599 613494 941619
rect 613550 941599 613618 941619
rect 613674 941599 613728 941655
rect 611828 941533 613728 941599
rect 611828 941531 611897 941533
rect 611953 941531 612039 941533
rect 612095 941531 612181 941533
rect 612237 941531 612323 941533
rect 612379 941531 612465 941533
rect 612521 941531 612607 941533
rect 612663 941531 612749 941533
rect 612805 941531 612891 941533
rect 612947 941531 613033 941533
rect 613089 941531 613175 941533
rect 613231 941531 613317 941533
rect 613373 941531 613459 941533
rect 613515 941531 613601 941533
rect 613657 941531 613728 941533
rect 611828 941475 611882 941531
rect 611953 941477 612006 941531
rect 612095 941477 612130 941531
rect 612237 941477 612254 941531
rect 611938 941475 612006 941477
rect 612062 941475 612130 941477
rect 612186 941475 612254 941477
rect 612310 941477 612323 941531
rect 612434 941477 612465 941531
rect 612558 941477 612607 941531
rect 612682 941477 612749 941531
rect 612310 941475 612378 941477
rect 612434 941475 612502 941477
rect 612558 941475 612626 941477
rect 612682 941475 612750 941477
rect 612806 941475 612874 941531
rect 612947 941477 612998 941531
rect 613089 941477 613122 941531
rect 613231 941477 613246 941531
rect 612930 941475 612998 941477
rect 613054 941475 613122 941477
rect 613178 941475 613246 941477
rect 613302 941477 613317 941531
rect 613426 941477 613459 941531
rect 613550 941477 613601 941531
rect 613302 941475 613370 941477
rect 613426 941475 613494 941477
rect 613550 941475 613618 941477
rect 613674 941475 613728 941531
rect 611828 941407 613728 941475
rect 611828 941351 611882 941407
rect 611938 941391 612006 941407
rect 612062 941391 612130 941407
rect 612186 941391 612254 941407
rect 611953 941351 612006 941391
rect 612095 941351 612130 941391
rect 612237 941351 612254 941391
rect 612310 941391 612378 941407
rect 612434 941391 612502 941407
rect 612558 941391 612626 941407
rect 612682 941391 612750 941407
rect 612310 941351 612323 941391
rect 612434 941351 612465 941391
rect 612558 941351 612607 941391
rect 612682 941351 612749 941391
rect 612806 941351 612874 941407
rect 612930 941391 612998 941407
rect 613054 941391 613122 941407
rect 613178 941391 613246 941407
rect 612947 941351 612998 941391
rect 613089 941351 613122 941391
rect 613231 941351 613246 941391
rect 613302 941391 613370 941407
rect 613426 941391 613494 941407
rect 613550 941391 613618 941407
rect 613302 941351 613317 941391
rect 613426 941351 613459 941391
rect 613550 941351 613601 941391
rect 613674 941351 613728 941407
rect 611828 941335 611897 941351
rect 611953 941335 612039 941351
rect 612095 941335 612181 941351
rect 612237 941335 612323 941351
rect 612379 941335 612465 941351
rect 612521 941335 612607 941351
rect 612663 941335 612749 941351
rect 612805 941335 612891 941351
rect 612947 941335 613033 941351
rect 613089 941335 613175 941351
rect 613231 941335 613317 941351
rect 613373 941335 613459 941351
rect 613515 941335 613601 941351
rect 613657 941335 613728 941351
rect 611828 941283 613728 941335
rect 611828 941227 611882 941283
rect 611938 941249 612006 941283
rect 612062 941249 612130 941283
rect 612186 941249 612254 941283
rect 611953 941227 612006 941249
rect 612095 941227 612130 941249
rect 612237 941227 612254 941249
rect 612310 941249 612378 941283
rect 612434 941249 612502 941283
rect 612558 941249 612626 941283
rect 612682 941249 612750 941283
rect 612310 941227 612323 941249
rect 612434 941227 612465 941249
rect 612558 941227 612607 941249
rect 612682 941227 612749 941249
rect 612806 941227 612874 941283
rect 612930 941249 612998 941283
rect 613054 941249 613122 941283
rect 613178 941249 613246 941283
rect 612947 941227 612998 941249
rect 613089 941227 613122 941249
rect 613231 941227 613246 941249
rect 613302 941249 613370 941283
rect 613426 941249 613494 941283
rect 613550 941249 613618 941283
rect 613302 941227 613317 941249
rect 613426 941227 613459 941249
rect 613550 941227 613601 941249
rect 613674 941227 613728 941283
rect 611828 941193 611897 941227
rect 611953 941193 612039 941227
rect 612095 941193 612181 941227
rect 612237 941193 612323 941227
rect 612379 941193 612465 941227
rect 612521 941193 612607 941227
rect 612663 941193 612749 941227
rect 612805 941193 612891 941227
rect 612947 941193 613033 941227
rect 613089 941193 613175 941227
rect 613231 941193 613317 941227
rect 613373 941193 613459 941227
rect 613515 941193 613601 941227
rect 613657 941193 613728 941227
rect 611828 941159 613728 941193
rect 611828 941103 611882 941159
rect 611938 941107 612006 941159
rect 612062 941107 612130 941159
rect 612186 941107 612254 941159
rect 611953 941103 612006 941107
rect 612095 941103 612130 941107
rect 612237 941103 612254 941107
rect 612310 941107 612378 941159
rect 612434 941107 612502 941159
rect 612558 941107 612626 941159
rect 612682 941107 612750 941159
rect 612310 941103 612323 941107
rect 612434 941103 612465 941107
rect 612558 941103 612607 941107
rect 612682 941103 612749 941107
rect 612806 941103 612874 941159
rect 612930 941107 612998 941159
rect 613054 941107 613122 941159
rect 613178 941107 613246 941159
rect 612947 941103 612998 941107
rect 613089 941103 613122 941107
rect 613231 941103 613246 941107
rect 613302 941107 613370 941159
rect 613426 941107 613494 941159
rect 613550 941107 613618 941159
rect 613302 941103 613317 941107
rect 613426 941103 613459 941107
rect 613550 941103 613601 941107
rect 613674 941103 613728 941159
rect 611828 941051 611897 941103
rect 611953 941051 612039 941103
rect 612095 941051 612181 941103
rect 612237 941051 612323 941103
rect 612379 941051 612465 941103
rect 612521 941051 612607 941103
rect 612663 941051 612749 941103
rect 612805 941051 612891 941103
rect 612947 941051 613033 941103
rect 613089 941051 613175 941103
rect 613231 941051 613317 941103
rect 613373 941051 613459 941103
rect 613515 941051 613601 941103
rect 613657 941051 613728 941103
rect 611828 941035 613728 941051
rect 611828 940979 611882 941035
rect 611938 940979 612006 941035
rect 612062 940979 612130 941035
rect 612186 940979 612254 941035
rect 612310 940979 612378 941035
rect 612434 940979 612502 941035
rect 612558 940979 612626 941035
rect 612682 940979 612750 941035
rect 612806 940979 612874 941035
rect 612930 940979 612998 941035
rect 613054 940979 613122 941035
rect 613178 940979 613246 941035
rect 613302 940979 613370 941035
rect 613426 940979 613494 941035
rect 613550 940979 613618 941035
rect 613674 940979 613728 941035
rect 611828 940965 613728 940979
rect 611828 940911 611897 940965
rect 611953 940911 612039 940965
rect 612095 940911 612181 940965
rect 612237 940911 612323 940965
rect 612379 940911 612465 940965
rect 612521 940911 612607 940965
rect 612663 940911 612749 940965
rect 612805 940911 612891 940965
rect 612947 940911 613033 940965
rect 613089 940911 613175 940965
rect 613231 940911 613317 940965
rect 613373 940911 613459 940965
rect 613515 940911 613601 940965
rect 613657 940911 613728 940965
rect 611828 940855 611882 940911
rect 611953 940909 612006 940911
rect 612095 940909 612130 940911
rect 612237 940909 612254 940911
rect 611938 940855 612006 940909
rect 612062 940855 612130 940909
rect 612186 940855 612254 940909
rect 612310 940909 612323 940911
rect 612434 940909 612465 940911
rect 612558 940909 612607 940911
rect 612682 940909 612749 940911
rect 612310 940855 612378 940909
rect 612434 940855 612502 940909
rect 612558 940855 612626 940909
rect 612682 940855 612750 940909
rect 612806 940855 612874 940911
rect 612947 940909 612998 940911
rect 613089 940909 613122 940911
rect 613231 940909 613246 940911
rect 612930 940855 612998 940909
rect 613054 940855 613122 940909
rect 613178 940855 613246 940909
rect 613302 940909 613317 940911
rect 613426 940909 613459 940911
rect 613550 940909 613601 940911
rect 613302 940855 613370 940909
rect 613426 940855 613494 940909
rect 613550 940855 613618 940909
rect 613674 940855 613728 940911
rect 611828 940823 613728 940855
rect 611828 940787 611897 940823
rect 611953 940787 612039 940823
rect 612095 940787 612181 940823
rect 612237 940787 612323 940823
rect 612379 940787 612465 940823
rect 612521 940787 612607 940823
rect 612663 940787 612749 940823
rect 612805 940787 612891 940823
rect 612947 940787 613033 940823
rect 613089 940787 613175 940823
rect 613231 940787 613317 940823
rect 613373 940787 613459 940823
rect 613515 940787 613601 940823
rect 613657 940787 613728 940823
rect 611828 940731 611882 940787
rect 611953 940767 612006 940787
rect 612095 940767 612130 940787
rect 612237 940767 612254 940787
rect 611938 940731 612006 940767
rect 612062 940731 612130 940767
rect 612186 940731 612254 940767
rect 612310 940767 612323 940787
rect 612434 940767 612465 940787
rect 612558 940767 612607 940787
rect 612682 940767 612749 940787
rect 612310 940731 612378 940767
rect 612434 940731 612502 940767
rect 612558 940731 612626 940767
rect 612682 940731 612750 940767
rect 612806 940731 612874 940787
rect 612947 940767 612998 940787
rect 613089 940767 613122 940787
rect 613231 940767 613246 940787
rect 612930 940731 612998 940767
rect 613054 940731 613122 940767
rect 613178 940731 613246 940767
rect 613302 940767 613317 940787
rect 613426 940767 613459 940787
rect 613550 940767 613601 940787
rect 613302 940731 613370 940767
rect 613426 940731 613494 940767
rect 613550 940731 613618 940767
rect 613674 940731 613728 940787
rect 611828 940681 613728 940731
rect 611828 940663 611897 940681
rect 611953 940663 612039 940681
rect 612095 940663 612181 940681
rect 612237 940663 612323 940681
rect 612379 940663 612465 940681
rect 612521 940663 612607 940681
rect 612663 940663 612749 940681
rect 612805 940663 612891 940681
rect 612947 940663 613033 940681
rect 613089 940663 613175 940681
rect 613231 940663 613317 940681
rect 613373 940663 613459 940681
rect 613515 940663 613601 940681
rect 613657 940663 613728 940681
rect 611828 940607 611882 940663
rect 611953 940625 612006 940663
rect 612095 940625 612130 940663
rect 612237 940625 612254 940663
rect 611938 940607 612006 940625
rect 612062 940607 612130 940625
rect 612186 940607 612254 940625
rect 612310 940625 612323 940663
rect 612434 940625 612465 940663
rect 612558 940625 612607 940663
rect 612682 940625 612749 940663
rect 612310 940607 612378 940625
rect 612434 940607 612502 940625
rect 612558 940607 612626 940625
rect 612682 940607 612750 940625
rect 612806 940607 612874 940663
rect 612947 940625 612998 940663
rect 613089 940625 613122 940663
rect 613231 940625 613246 940663
rect 612930 940607 612998 940625
rect 613054 940607 613122 940625
rect 613178 940607 613246 940625
rect 613302 940625 613317 940663
rect 613426 940625 613459 940663
rect 613550 940625 613601 940663
rect 613302 940607 613370 940625
rect 613426 940607 613494 940625
rect 613550 940607 613618 940625
rect 613674 940607 613728 940663
rect 611828 940539 613728 940607
rect 611828 940483 611882 940539
rect 611953 940483 612006 940539
rect 612095 940483 612130 940539
rect 612237 940483 612254 940539
rect 612310 940483 612323 940539
rect 612434 940483 612465 940539
rect 612558 940483 612607 940539
rect 612682 940483 612749 940539
rect 612806 940483 612874 940539
rect 612947 940483 612998 940539
rect 613089 940483 613122 940539
rect 613231 940483 613246 940539
rect 613302 940483 613317 940539
rect 613426 940483 613459 940539
rect 613550 940483 613601 940539
rect 613674 940483 613728 940539
rect 611828 940415 613728 940483
rect 611828 940359 611882 940415
rect 611938 940397 612006 940415
rect 612062 940397 612130 940415
rect 612186 940397 612254 940415
rect 611953 940359 612006 940397
rect 612095 940359 612130 940397
rect 612237 940359 612254 940397
rect 612310 940397 612378 940415
rect 612434 940397 612502 940415
rect 612558 940397 612626 940415
rect 612682 940397 612750 940415
rect 612310 940359 612323 940397
rect 612434 940359 612465 940397
rect 612558 940359 612607 940397
rect 612682 940359 612749 940397
rect 612806 940359 612874 940415
rect 612930 940397 612998 940415
rect 613054 940397 613122 940415
rect 613178 940397 613246 940415
rect 612947 940359 612998 940397
rect 613089 940359 613122 940397
rect 613231 940359 613246 940397
rect 613302 940397 613370 940415
rect 613426 940397 613494 940415
rect 613550 940397 613618 940415
rect 613302 940359 613317 940397
rect 613426 940359 613459 940397
rect 613550 940359 613601 940397
rect 613674 940359 613728 940415
rect 611828 940341 611897 940359
rect 611953 940341 612039 940359
rect 612095 940341 612181 940359
rect 612237 940341 612323 940359
rect 612379 940341 612465 940359
rect 612521 940341 612607 940359
rect 612663 940341 612749 940359
rect 612805 940341 612891 940359
rect 612947 940341 613033 940359
rect 613089 940341 613175 940359
rect 613231 940341 613317 940359
rect 613373 940341 613459 940359
rect 613515 940341 613601 940359
rect 613657 940341 613728 940359
rect 611828 940291 613728 940341
rect 611828 940235 611882 940291
rect 611938 940255 612006 940291
rect 612062 940255 612130 940291
rect 612186 940255 612254 940291
rect 611953 940235 612006 940255
rect 612095 940235 612130 940255
rect 612237 940235 612254 940255
rect 612310 940255 612378 940291
rect 612434 940255 612502 940291
rect 612558 940255 612626 940291
rect 612682 940255 612750 940291
rect 612310 940235 612323 940255
rect 612434 940235 612465 940255
rect 612558 940235 612607 940255
rect 612682 940235 612749 940255
rect 612806 940235 612874 940291
rect 612930 940255 612998 940291
rect 613054 940255 613122 940291
rect 613178 940255 613246 940291
rect 612947 940235 612998 940255
rect 613089 940235 613122 940255
rect 613231 940235 613246 940255
rect 613302 940255 613370 940291
rect 613426 940255 613494 940291
rect 613550 940255 613618 940291
rect 613302 940235 613317 940255
rect 613426 940235 613459 940255
rect 613550 940235 613601 940255
rect 613674 940235 613728 940291
rect 611828 940199 611897 940235
rect 611953 940199 612039 940235
rect 612095 940199 612181 940235
rect 612237 940199 612323 940235
rect 612379 940199 612465 940235
rect 612521 940199 612607 940235
rect 612663 940199 612749 940235
rect 612805 940199 612891 940235
rect 612947 940199 613033 940235
rect 613089 940199 613175 940235
rect 613231 940199 613317 940235
rect 613373 940199 613459 940235
rect 613515 940199 613601 940235
rect 613657 940199 613728 940235
rect 611828 940167 613728 940199
rect 611828 940111 611882 940167
rect 611938 940113 612006 940167
rect 612062 940113 612130 940167
rect 612186 940113 612254 940167
rect 611953 940111 612006 940113
rect 612095 940111 612130 940113
rect 612237 940111 612254 940113
rect 612310 940113 612378 940167
rect 612434 940113 612502 940167
rect 612558 940113 612626 940167
rect 612682 940113 612750 940167
rect 612310 940111 612323 940113
rect 612434 940111 612465 940113
rect 612558 940111 612607 940113
rect 612682 940111 612749 940113
rect 612806 940111 612874 940167
rect 612930 940113 612998 940167
rect 613054 940113 613122 940167
rect 613178 940113 613246 940167
rect 612947 940111 612998 940113
rect 613089 940111 613122 940113
rect 613231 940111 613246 940113
rect 613302 940113 613370 940167
rect 613426 940113 613494 940167
rect 613550 940113 613618 940167
rect 613302 940111 613317 940113
rect 613426 940111 613459 940113
rect 613550 940111 613601 940113
rect 613674 940111 613728 940167
rect 611828 940057 611897 940111
rect 611953 940057 612039 940111
rect 612095 940057 612181 940111
rect 612237 940057 612323 940111
rect 612379 940057 612465 940111
rect 612521 940057 612607 940111
rect 612663 940057 612749 940111
rect 612805 940057 612891 940111
rect 612947 940057 613033 940111
rect 613089 940057 613175 940111
rect 613231 940057 613317 940111
rect 613373 940057 613459 940111
rect 613515 940057 613601 940111
rect 613657 940057 613728 940111
rect 611828 940043 613728 940057
rect 611828 939987 611882 940043
rect 611938 939987 612006 940043
rect 612062 939987 612130 940043
rect 612186 939987 612254 940043
rect 612310 939987 612378 940043
rect 612434 939987 612502 940043
rect 612558 939987 612626 940043
rect 612682 939987 612750 940043
rect 612806 939987 612874 940043
rect 612930 939987 612998 940043
rect 613054 939987 613122 940043
rect 613178 939987 613246 940043
rect 613302 939987 613370 940043
rect 613426 939987 613494 940043
rect 613550 939987 613618 940043
rect 613674 939987 613728 940043
rect 611828 939971 613728 939987
rect 611828 939919 611897 939971
rect 611953 939919 612039 939971
rect 612095 939919 612181 939971
rect 612237 939919 612323 939971
rect 612379 939919 612465 939971
rect 612521 939919 612607 939971
rect 612663 939919 612749 939971
rect 612805 939919 612891 939971
rect 612947 939919 613033 939971
rect 613089 939919 613175 939971
rect 613231 939919 613317 939971
rect 613373 939919 613459 939971
rect 613515 939919 613601 939971
rect 613657 939919 613728 939971
rect 611828 939863 611882 939919
rect 611953 939915 612006 939919
rect 612095 939915 612130 939919
rect 612237 939915 612254 939919
rect 611938 939863 612006 939915
rect 612062 939863 612130 939915
rect 612186 939863 612254 939915
rect 612310 939915 612323 939919
rect 612434 939915 612465 939919
rect 612558 939915 612607 939919
rect 612682 939915 612749 939919
rect 612310 939863 612378 939915
rect 612434 939863 612502 939915
rect 612558 939863 612626 939915
rect 612682 939863 612750 939915
rect 612806 939863 612874 939919
rect 612947 939915 612998 939919
rect 613089 939915 613122 939919
rect 613231 939915 613246 939919
rect 612930 939863 612998 939915
rect 613054 939863 613122 939915
rect 613178 939863 613246 939915
rect 613302 939915 613317 939919
rect 613426 939915 613459 939919
rect 613550 939915 613601 939919
rect 613302 939863 613370 939915
rect 613426 939863 613494 939915
rect 613550 939863 613618 939915
rect 613674 939863 613728 939919
rect 611828 939829 613728 939863
rect 611828 939773 611897 939829
rect 611953 939773 612039 939829
rect 612095 939773 612181 939829
rect 612237 939773 612323 939829
rect 612379 939773 612465 939829
rect 612521 939773 612607 939829
rect 612663 939773 612749 939829
rect 612805 939773 612891 939829
rect 612947 939773 613033 939829
rect 613089 939773 613175 939829
rect 613231 939773 613317 939829
rect 613373 939773 613459 939829
rect 613515 939773 613601 939829
rect 613657 939773 613728 939829
rect 611828 939720 613728 939773
rect 70000 878661 75816 878728
rect 70000 878605 70047 878661
rect 70103 878605 70171 878661
rect 70227 878605 70295 878661
rect 70351 878605 70419 878661
rect 70475 878650 75816 878661
rect 70475 878605 73866 878650
rect 70000 878594 73866 878605
rect 73922 878594 74008 878650
rect 74064 878594 74150 878650
rect 74206 878594 74292 878650
rect 74348 878594 74434 878650
rect 74490 878594 74576 878650
rect 74632 878594 74718 878650
rect 74774 878594 74860 878650
rect 74916 878594 75002 878650
rect 75058 878594 75144 878650
rect 75200 878594 75286 878650
rect 75342 878594 75428 878650
rect 75484 878594 75570 878650
rect 75626 878594 75712 878650
rect 75768 878594 75816 878650
rect 70000 878537 75816 878594
rect 70000 878481 70047 878537
rect 70103 878481 70171 878537
rect 70227 878481 70295 878537
rect 70351 878481 70419 878537
rect 70475 878508 75816 878537
rect 70475 878481 73866 878508
rect 70000 878452 73866 878481
rect 73922 878452 74008 878508
rect 74064 878452 74150 878508
rect 74206 878452 74292 878508
rect 74348 878452 74434 878508
rect 74490 878452 74576 878508
rect 74632 878452 74718 878508
rect 74774 878452 74860 878508
rect 74916 878452 75002 878508
rect 75058 878452 75144 878508
rect 75200 878452 75286 878508
rect 75342 878452 75428 878508
rect 75484 878452 75570 878508
rect 75626 878452 75712 878508
rect 75768 878452 75816 878508
rect 70000 878413 75816 878452
rect 70000 878357 70047 878413
rect 70103 878357 70171 878413
rect 70227 878357 70295 878413
rect 70351 878357 70419 878413
rect 70475 878366 75816 878413
rect 70475 878357 73866 878366
rect 70000 878310 73866 878357
rect 73922 878310 74008 878366
rect 74064 878310 74150 878366
rect 74206 878310 74292 878366
rect 74348 878310 74434 878366
rect 74490 878310 74576 878366
rect 74632 878310 74718 878366
rect 74774 878310 74860 878366
rect 74916 878310 75002 878366
rect 75058 878310 75144 878366
rect 75200 878310 75286 878366
rect 75342 878310 75428 878366
rect 75484 878310 75570 878366
rect 75626 878310 75712 878366
rect 75768 878310 75816 878366
rect 70000 878289 75816 878310
rect 70000 878233 70047 878289
rect 70103 878233 70171 878289
rect 70227 878233 70295 878289
rect 70351 878233 70419 878289
rect 70475 878233 75816 878289
rect 70000 878224 75816 878233
rect 70000 878168 73866 878224
rect 73922 878168 74008 878224
rect 74064 878168 74150 878224
rect 74206 878168 74292 878224
rect 74348 878168 74434 878224
rect 74490 878168 74576 878224
rect 74632 878168 74718 878224
rect 74774 878168 74860 878224
rect 74916 878168 75002 878224
rect 75058 878168 75144 878224
rect 75200 878168 75286 878224
rect 75342 878168 75428 878224
rect 75484 878168 75570 878224
rect 75626 878168 75712 878224
rect 75768 878168 75816 878224
rect 70000 878165 75816 878168
rect 70000 878109 70047 878165
rect 70103 878109 70171 878165
rect 70227 878109 70295 878165
rect 70351 878109 70419 878165
rect 70475 878109 75816 878165
rect 70000 878082 75816 878109
rect 70000 878041 73866 878082
rect 70000 877985 70047 878041
rect 70103 877985 70171 878041
rect 70227 877985 70295 878041
rect 70351 877985 70419 878041
rect 70475 878026 73866 878041
rect 73922 878026 74008 878082
rect 74064 878026 74150 878082
rect 74206 878026 74292 878082
rect 74348 878026 74434 878082
rect 74490 878026 74576 878082
rect 74632 878026 74718 878082
rect 74774 878026 74860 878082
rect 74916 878026 75002 878082
rect 75058 878026 75144 878082
rect 75200 878026 75286 878082
rect 75342 878026 75428 878082
rect 75484 878026 75570 878082
rect 75626 878026 75712 878082
rect 75768 878026 75816 878082
rect 70475 877985 75816 878026
rect 70000 877940 75816 877985
rect 70000 877917 73866 877940
rect 70000 877861 70047 877917
rect 70103 877861 70171 877917
rect 70227 877861 70295 877917
rect 70351 877861 70419 877917
rect 70475 877884 73866 877917
rect 73922 877884 74008 877940
rect 74064 877884 74150 877940
rect 74206 877884 74292 877940
rect 74348 877884 74434 877940
rect 74490 877884 74576 877940
rect 74632 877884 74718 877940
rect 74774 877884 74860 877940
rect 74916 877884 75002 877940
rect 75058 877884 75144 877940
rect 75200 877884 75286 877940
rect 75342 877884 75428 877940
rect 75484 877884 75570 877940
rect 75626 877884 75712 877940
rect 75768 877884 75816 877940
rect 70475 877861 75816 877884
rect 70000 877798 75816 877861
rect 70000 877793 73866 877798
rect 70000 877737 70047 877793
rect 70103 877737 70171 877793
rect 70227 877737 70295 877793
rect 70351 877737 70419 877793
rect 70475 877742 73866 877793
rect 73922 877742 74008 877798
rect 74064 877742 74150 877798
rect 74206 877742 74292 877798
rect 74348 877742 74434 877798
rect 74490 877742 74576 877798
rect 74632 877742 74718 877798
rect 74774 877742 74860 877798
rect 74916 877742 75002 877798
rect 75058 877742 75144 877798
rect 75200 877742 75286 877798
rect 75342 877742 75428 877798
rect 75484 877742 75570 877798
rect 75626 877742 75712 877798
rect 75768 877742 75816 877798
rect 70475 877737 75816 877742
rect 70000 877669 75816 877737
rect 70000 877613 70047 877669
rect 70103 877613 70171 877669
rect 70227 877613 70295 877669
rect 70351 877613 70419 877669
rect 70475 877656 75816 877669
rect 70475 877613 73866 877656
rect 70000 877600 73866 877613
rect 73922 877600 74008 877656
rect 74064 877600 74150 877656
rect 74206 877600 74292 877656
rect 74348 877600 74434 877656
rect 74490 877600 74576 877656
rect 74632 877600 74718 877656
rect 74774 877600 74860 877656
rect 74916 877600 75002 877656
rect 75058 877600 75144 877656
rect 75200 877600 75286 877656
rect 75342 877600 75428 877656
rect 75484 877600 75570 877656
rect 75626 877600 75712 877656
rect 75768 877600 75816 877656
rect 70000 877545 75816 877600
rect 70000 877489 70047 877545
rect 70103 877489 70171 877545
rect 70227 877489 70295 877545
rect 70351 877489 70419 877545
rect 70475 877514 75816 877545
rect 70475 877489 73866 877514
rect 70000 877458 73866 877489
rect 73922 877458 74008 877514
rect 74064 877458 74150 877514
rect 74206 877458 74292 877514
rect 74348 877458 74434 877514
rect 74490 877458 74576 877514
rect 74632 877458 74718 877514
rect 74774 877458 74860 877514
rect 74916 877458 75002 877514
rect 75058 877458 75144 877514
rect 75200 877458 75286 877514
rect 75342 877458 75428 877514
rect 75484 877458 75570 877514
rect 75626 877458 75712 877514
rect 75768 877458 75816 877514
rect 70000 877421 75816 877458
rect 70000 877365 70047 877421
rect 70103 877365 70171 877421
rect 70227 877365 70295 877421
rect 70351 877365 70419 877421
rect 70475 877372 75816 877421
rect 70475 877365 73866 877372
rect 70000 877316 73866 877365
rect 73922 877316 74008 877372
rect 74064 877316 74150 877372
rect 74206 877316 74292 877372
rect 74348 877316 74434 877372
rect 74490 877316 74576 877372
rect 74632 877316 74718 877372
rect 74774 877316 74860 877372
rect 74916 877316 75002 877372
rect 75058 877316 75144 877372
rect 75200 877316 75286 877372
rect 75342 877316 75428 877372
rect 75484 877316 75570 877372
rect 75626 877316 75712 877372
rect 75768 877316 75816 877372
rect 70000 877297 75816 877316
rect 70000 877241 70047 877297
rect 70103 877241 70171 877297
rect 70227 877241 70295 877297
rect 70351 877241 70419 877297
rect 70475 877241 75816 877297
rect 70000 877230 75816 877241
rect 70000 877174 73866 877230
rect 73922 877174 74008 877230
rect 74064 877174 74150 877230
rect 74206 877174 74292 877230
rect 74348 877174 74434 877230
rect 74490 877174 74576 877230
rect 74632 877174 74718 877230
rect 74774 877174 74860 877230
rect 74916 877174 75002 877230
rect 75058 877174 75144 877230
rect 75200 877174 75286 877230
rect 75342 877174 75428 877230
rect 75484 877174 75570 877230
rect 75626 877174 75712 877230
rect 75768 877174 75816 877230
rect 70000 877173 75816 877174
rect 70000 877117 70047 877173
rect 70103 877117 70171 877173
rect 70227 877117 70295 877173
rect 70351 877117 70419 877173
rect 70475 877117 75816 877173
rect 70000 877088 75816 877117
rect 70000 877049 73866 877088
rect 70000 876993 70047 877049
rect 70103 876993 70171 877049
rect 70227 876993 70295 877049
rect 70351 876993 70419 877049
rect 70475 877032 73866 877049
rect 73922 877032 74008 877088
rect 74064 877032 74150 877088
rect 74206 877032 74292 877088
rect 74348 877032 74434 877088
rect 74490 877032 74576 877088
rect 74632 877032 74718 877088
rect 74774 877032 74860 877088
rect 74916 877032 75002 877088
rect 75058 877032 75144 877088
rect 75200 877032 75286 877088
rect 75342 877032 75428 877088
rect 75484 877032 75570 877088
rect 75626 877032 75712 877088
rect 75768 877032 75816 877088
rect 70475 876993 75816 877032
rect 70000 876946 75816 876993
rect 70000 876925 73866 876946
rect 70000 876869 70047 876925
rect 70103 876869 70171 876925
rect 70227 876869 70295 876925
rect 70351 876869 70419 876925
rect 70475 876890 73866 876925
rect 73922 876890 74008 876946
rect 74064 876890 74150 876946
rect 74206 876890 74292 876946
rect 74348 876890 74434 876946
rect 74490 876890 74576 876946
rect 74632 876890 74718 876946
rect 74774 876890 74860 876946
rect 74916 876890 75002 876946
rect 75058 876890 75144 876946
rect 75200 876890 75286 876946
rect 75342 876890 75428 876946
rect 75484 876890 75570 876946
rect 75626 876890 75712 876946
rect 75768 876890 75816 876946
rect 70475 876869 75816 876890
rect 70000 876828 75816 876869
rect 699992 877687 706000 877728
rect 699992 877666 705525 877687
rect 699992 877610 700040 877666
rect 700096 877610 700182 877666
rect 700238 877610 700324 877666
rect 700380 877610 700466 877666
rect 700522 877610 700608 877666
rect 700664 877610 700750 877666
rect 700806 877610 700892 877666
rect 700948 877610 701034 877666
rect 701090 877610 701176 877666
rect 701232 877610 701318 877666
rect 701374 877610 701460 877666
rect 701516 877610 701602 877666
rect 701658 877610 701744 877666
rect 701800 877610 701886 877666
rect 701942 877631 705525 877666
rect 705581 877631 705649 877687
rect 705705 877631 705773 877687
rect 705829 877631 705897 877687
rect 705953 877631 706000 877687
rect 701942 877610 706000 877631
rect 699992 877563 706000 877610
rect 699992 877524 705525 877563
rect 699992 877468 700040 877524
rect 700096 877468 700182 877524
rect 700238 877468 700324 877524
rect 700380 877468 700466 877524
rect 700522 877468 700608 877524
rect 700664 877468 700750 877524
rect 700806 877468 700892 877524
rect 700948 877468 701034 877524
rect 701090 877468 701176 877524
rect 701232 877468 701318 877524
rect 701374 877468 701460 877524
rect 701516 877468 701602 877524
rect 701658 877468 701744 877524
rect 701800 877468 701886 877524
rect 701942 877507 705525 877524
rect 705581 877507 705649 877563
rect 705705 877507 705773 877563
rect 705829 877507 705897 877563
rect 705953 877507 706000 877563
rect 701942 877468 706000 877507
rect 699992 877439 706000 877468
rect 699992 877383 705525 877439
rect 705581 877383 705649 877439
rect 705705 877383 705773 877439
rect 705829 877383 705897 877439
rect 705953 877383 706000 877439
rect 699992 877382 706000 877383
rect 699992 877326 700040 877382
rect 700096 877326 700182 877382
rect 700238 877326 700324 877382
rect 700380 877326 700466 877382
rect 700522 877326 700608 877382
rect 700664 877326 700750 877382
rect 700806 877326 700892 877382
rect 700948 877326 701034 877382
rect 701090 877326 701176 877382
rect 701232 877326 701318 877382
rect 701374 877326 701460 877382
rect 701516 877326 701602 877382
rect 701658 877326 701744 877382
rect 701800 877326 701886 877382
rect 701942 877326 706000 877382
rect 699992 877315 706000 877326
rect 699992 877259 705525 877315
rect 705581 877259 705649 877315
rect 705705 877259 705773 877315
rect 705829 877259 705897 877315
rect 705953 877259 706000 877315
rect 699992 877240 706000 877259
rect 699992 877184 700040 877240
rect 700096 877184 700182 877240
rect 700238 877184 700324 877240
rect 700380 877184 700466 877240
rect 700522 877184 700608 877240
rect 700664 877184 700750 877240
rect 700806 877184 700892 877240
rect 700948 877184 701034 877240
rect 701090 877184 701176 877240
rect 701232 877184 701318 877240
rect 701374 877184 701460 877240
rect 701516 877184 701602 877240
rect 701658 877184 701744 877240
rect 701800 877184 701886 877240
rect 701942 877191 706000 877240
rect 701942 877184 705525 877191
rect 699992 877135 705525 877184
rect 705581 877135 705649 877191
rect 705705 877135 705773 877191
rect 705829 877135 705897 877191
rect 705953 877135 706000 877191
rect 699992 877098 706000 877135
rect 699992 877042 700040 877098
rect 700096 877042 700182 877098
rect 700238 877042 700324 877098
rect 700380 877042 700466 877098
rect 700522 877042 700608 877098
rect 700664 877042 700750 877098
rect 700806 877042 700892 877098
rect 700948 877042 701034 877098
rect 701090 877042 701176 877098
rect 701232 877042 701318 877098
rect 701374 877042 701460 877098
rect 701516 877042 701602 877098
rect 701658 877042 701744 877098
rect 701800 877042 701886 877098
rect 701942 877067 706000 877098
rect 701942 877042 705525 877067
rect 699992 877011 705525 877042
rect 705581 877011 705649 877067
rect 705705 877011 705773 877067
rect 705829 877011 705897 877067
rect 705953 877011 706000 877067
rect 699992 876956 706000 877011
rect 699992 876900 700040 876956
rect 700096 876900 700182 876956
rect 700238 876900 700324 876956
rect 700380 876900 700466 876956
rect 700522 876900 700608 876956
rect 700664 876900 700750 876956
rect 700806 876900 700892 876956
rect 700948 876900 701034 876956
rect 701090 876900 701176 876956
rect 701232 876900 701318 876956
rect 701374 876900 701460 876956
rect 701516 876900 701602 876956
rect 701658 876900 701744 876956
rect 701800 876900 701886 876956
rect 701942 876943 706000 876956
rect 701942 876900 705525 876943
rect 699992 876887 705525 876900
rect 705581 876887 705649 876943
rect 705705 876887 705773 876943
rect 705829 876887 705897 876943
rect 705953 876887 706000 876943
rect 699992 876819 706000 876887
rect 699992 876814 705525 876819
rect 699992 876758 700040 876814
rect 700096 876758 700182 876814
rect 700238 876758 700324 876814
rect 700380 876758 700466 876814
rect 700522 876758 700608 876814
rect 700664 876758 700750 876814
rect 700806 876758 700892 876814
rect 700948 876758 701034 876814
rect 701090 876758 701176 876814
rect 701232 876758 701318 876814
rect 701374 876758 701460 876814
rect 701516 876758 701602 876814
rect 701658 876758 701744 876814
rect 701800 876758 701886 876814
rect 701942 876763 705525 876814
rect 705581 876763 705649 876819
rect 705705 876763 705773 876819
rect 705829 876763 705897 876819
rect 705953 876763 706000 876819
rect 701942 876758 706000 876763
rect 699992 876695 706000 876758
rect 699992 876672 705525 876695
rect 699992 876616 700040 876672
rect 700096 876616 700182 876672
rect 700238 876616 700324 876672
rect 700380 876616 700466 876672
rect 700522 876616 700608 876672
rect 700664 876616 700750 876672
rect 700806 876616 700892 876672
rect 700948 876616 701034 876672
rect 701090 876616 701176 876672
rect 701232 876616 701318 876672
rect 701374 876616 701460 876672
rect 701516 876616 701602 876672
rect 701658 876616 701744 876672
rect 701800 876616 701886 876672
rect 701942 876639 705525 876672
rect 705581 876639 705649 876695
rect 705705 876639 705773 876695
rect 705829 876639 705897 876695
rect 705953 876639 706000 876695
rect 701942 876616 706000 876639
rect 699992 876571 706000 876616
rect 699992 876530 705525 876571
rect 699992 876474 700040 876530
rect 700096 876474 700182 876530
rect 700238 876474 700324 876530
rect 700380 876474 700466 876530
rect 700522 876474 700608 876530
rect 700664 876474 700750 876530
rect 700806 876474 700892 876530
rect 700948 876474 701034 876530
rect 701090 876474 701176 876530
rect 701232 876474 701318 876530
rect 701374 876474 701460 876530
rect 701516 876474 701602 876530
rect 701658 876474 701744 876530
rect 701800 876474 701886 876530
rect 701942 876515 705525 876530
rect 705581 876515 705649 876571
rect 705705 876515 705773 876571
rect 705829 876515 705897 876571
rect 705953 876515 706000 876571
rect 701942 876474 706000 876515
rect 699992 876447 706000 876474
rect 699992 876391 705525 876447
rect 705581 876391 705649 876447
rect 705705 876391 705773 876447
rect 705829 876391 705897 876447
rect 705953 876391 706000 876447
rect 699992 876388 706000 876391
rect 699992 876332 700040 876388
rect 700096 876332 700182 876388
rect 700238 876332 700324 876388
rect 700380 876332 700466 876388
rect 700522 876332 700608 876388
rect 700664 876332 700750 876388
rect 700806 876332 700892 876388
rect 700948 876332 701034 876388
rect 701090 876332 701176 876388
rect 701232 876332 701318 876388
rect 701374 876332 701460 876388
rect 701516 876332 701602 876388
rect 701658 876332 701744 876388
rect 701800 876332 701886 876388
rect 701942 876332 706000 876388
rect 699992 876323 706000 876332
rect 699992 876267 705525 876323
rect 705581 876267 705649 876323
rect 705705 876267 705773 876323
rect 705829 876267 705897 876323
rect 705953 876267 706000 876323
rect 70000 876181 75816 876248
rect 70000 876125 70047 876181
rect 70103 876125 70171 876181
rect 70227 876125 70295 876181
rect 70351 876125 70419 876181
rect 70475 876169 75816 876181
rect 70475 876125 73855 876169
rect 70000 876113 73855 876125
rect 73911 876113 73997 876169
rect 74053 876113 74139 876169
rect 74195 876113 74281 876169
rect 74337 876113 74423 876169
rect 74479 876113 74565 876169
rect 74621 876113 74707 876169
rect 74763 876113 74849 876169
rect 74905 876113 74991 876169
rect 75047 876113 75133 876169
rect 75189 876113 75275 876169
rect 75331 876113 75417 876169
rect 75473 876113 75559 876169
rect 75615 876113 75701 876169
rect 75757 876113 75816 876169
rect 70000 876057 75816 876113
rect 70000 876001 70047 876057
rect 70103 876001 70171 876057
rect 70227 876001 70295 876057
rect 70351 876001 70419 876057
rect 70475 876027 75816 876057
rect 70475 876001 73855 876027
rect 70000 875971 73855 876001
rect 73911 875971 73997 876027
rect 74053 875971 74139 876027
rect 74195 875971 74281 876027
rect 74337 875971 74423 876027
rect 74479 875971 74565 876027
rect 74621 875971 74707 876027
rect 74763 875971 74849 876027
rect 74905 875971 74991 876027
rect 75047 875971 75133 876027
rect 75189 875971 75275 876027
rect 75331 875971 75417 876027
rect 75473 875971 75559 876027
rect 75615 875971 75701 876027
rect 75757 875971 75816 876027
rect 70000 875933 75816 875971
rect 70000 875877 70047 875933
rect 70103 875877 70171 875933
rect 70227 875877 70295 875933
rect 70351 875877 70419 875933
rect 70475 875885 75816 875933
rect 70475 875877 73855 875885
rect 70000 875829 73855 875877
rect 73911 875829 73997 875885
rect 74053 875829 74139 875885
rect 74195 875829 74281 875885
rect 74337 875829 74423 875885
rect 74479 875829 74565 875885
rect 74621 875829 74707 875885
rect 74763 875829 74849 875885
rect 74905 875829 74991 875885
rect 75047 875829 75133 875885
rect 75189 875829 75275 875885
rect 75331 875829 75417 875885
rect 75473 875829 75559 875885
rect 75615 875829 75701 875885
rect 75757 875829 75816 875885
rect 70000 875809 75816 875829
rect 699992 876246 706000 876267
rect 699992 876190 700040 876246
rect 700096 876190 700182 876246
rect 700238 876190 700324 876246
rect 700380 876190 700466 876246
rect 700522 876190 700608 876246
rect 700664 876190 700750 876246
rect 700806 876190 700892 876246
rect 700948 876190 701034 876246
rect 701090 876190 701176 876246
rect 701232 876190 701318 876246
rect 701374 876190 701460 876246
rect 701516 876190 701602 876246
rect 701658 876190 701744 876246
rect 701800 876190 701886 876246
rect 701942 876199 706000 876246
rect 701942 876190 705525 876199
rect 699992 876143 705525 876190
rect 705581 876143 705649 876199
rect 705705 876143 705773 876199
rect 705829 876143 705897 876199
rect 705953 876143 706000 876199
rect 699992 876104 706000 876143
rect 699992 876048 700040 876104
rect 700096 876048 700182 876104
rect 700238 876048 700324 876104
rect 700380 876048 700466 876104
rect 700522 876048 700608 876104
rect 700664 876048 700750 876104
rect 700806 876048 700892 876104
rect 700948 876048 701034 876104
rect 701090 876048 701176 876104
rect 701232 876048 701318 876104
rect 701374 876048 701460 876104
rect 701516 876048 701602 876104
rect 701658 876048 701744 876104
rect 701800 876048 701886 876104
rect 701942 876075 706000 876104
rect 701942 876048 705525 876075
rect 699992 876019 705525 876048
rect 705581 876019 705649 876075
rect 705705 876019 705773 876075
rect 705829 876019 705897 876075
rect 705953 876019 706000 876075
rect 699992 875962 706000 876019
rect 699992 875906 700040 875962
rect 700096 875906 700182 875962
rect 700238 875906 700324 875962
rect 700380 875906 700466 875962
rect 700522 875906 700608 875962
rect 700664 875906 700750 875962
rect 700806 875906 700892 875962
rect 700948 875906 701034 875962
rect 701090 875906 701176 875962
rect 701232 875906 701318 875962
rect 701374 875906 701460 875962
rect 701516 875906 701602 875962
rect 701658 875906 701744 875962
rect 701800 875906 701886 875962
rect 701942 875951 706000 875962
rect 701942 875906 705525 875951
rect 699992 875895 705525 875906
rect 705581 875895 705649 875951
rect 705705 875895 705773 875951
rect 705829 875895 705897 875951
rect 705953 875895 706000 875951
rect 699992 875828 706000 875895
rect 70000 875753 70047 875809
rect 70103 875753 70171 875809
rect 70227 875753 70295 875809
rect 70351 875753 70419 875809
rect 70475 875753 75816 875809
rect 70000 875743 75816 875753
rect 70000 875687 73855 875743
rect 73911 875687 73997 875743
rect 74053 875687 74139 875743
rect 74195 875687 74281 875743
rect 74337 875687 74423 875743
rect 74479 875687 74565 875743
rect 74621 875687 74707 875743
rect 74763 875687 74849 875743
rect 74905 875687 74991 875743
rect 75047 875687 75133 875743
rect 75189 875687 75275 875743
rect 75331 875687 75417 875743
rect 75473 875687 75559 875743
rect 75615 875687 75701 875743
rect 75757 875687 75816 875743
rect 70000 875685 75816 875687
rect 70000 875629 70047 875685
rect 70103 875629 70171 875685
rect 70227 875629 70295 875685
rect 70351 875629 70419 875685
rect 70475 875629 75816 875685
rect 70000 875601 75816 875629
rect 70000 875561 73855 875601
rect 70000 875505 70047 875561
rect 70103 875505 70171 875561
rect 70227 875505 70295 875561
rect 70351 875505 70419 875561
rect 70475 875545 73855 875561
rect 73911 875545 73997 875601
rect 74053 875545 74139 875601
rect 74195 875545 74281 875601
rect 74337 875545 74423 875601
rect 74479 875545 74565 875601
rect 74621 875545 74707 875601
rect 74763 875545 74849 875601
rect 74905 875545 74991 875601
rect 75047 875545 75133 875601
rect 75189 875545 75275 875601
rect 75331 875545 75417 875601
rect 75473 875545 75559 875601
rect 75615 875545 75701 875601
rect 75757 875545 75816 875601
rect 70475 875505 75816 875545
rect 70000 875459 75816 875505
rect 70000 875437 73855 875459
rect 70000 875381 70047 875437
rect 70103 875381 70171 875437
rect 70227 875381 70295 875437
rect 70351 875381 70419 875437
rect 70475 875403 73855 875437
rect 73911 875403 73997 875459
rect 74053 875403 74139 875459
rect 74195 875403 74281 875459
rect 74337 875403 74423 875459
rect 74479 875403 74565 875459
rect 74621 875403 74707 875459
rect 74763 875403 74849 875459
rect 74905 875403 74991 875459
rect 75047 875403 75133 875459
rect 75189 875403 75275 875459
rect 75331 875403 75417 875459
rect 75473 875403 75559 875459
rect 75615 875403 75701 875459
rect 75757 875403 75816 875459
rect 70475 875381 75816 875403
rect 70000 875317 75816 875381
rect 70000 875313 73855 875317
rect 70000 875257 70047 875313
rect 70103 875257 70171 875313
rect 70227 875257 70295 875313
rect 70351 875257 70419 875313
rect 70475 875261 73855 875313
rect 73911 875261 73997 875317
rect 74053 875261 74139 875317
rect 74195 875261 74281 875317
rect 74337 875261 74423 875317
rect 74479 875261 74565 875317
rect 74621 875261 74707 875317
rect 74763 875261 74849 875317
rect 74905 875261 74991 875317
rect 75047 875261 75133 875317
rect 75189 875261 75275 875317
rect 75331 875261 75417 875317
rect 75473 875261 75559 875317
rect 75615 875261 75701 875317
rect 75757 875261 75816 875317
rect 70475 875257 75816 875261
rect 70000 875189 75816 875257
rect 70000 875133 70047 875189
rect 70103 875133 70171 875189
rect 70227 875133 70295 875189
rect 70351 875133 70419 875189
rect 70475 875175 75816 875189
rect 70475 875133 73855 875175
rect 70000 875119 73855 875133
rect 73911 875119 73997 875175
rect 74053 875119 74139 875175
rect 74195 875119 74281 875175
rect 74337 875119 74423 875175
rect 74479 875119 74565 875175
rect 74621 875119 74707 875175
rect 74763 875119 74849 875175
rect 74905 875119 74991 875175
rect 75047 875119 75133 875175
rect 75189 875119 75275 875175
rect 75331 875119 75417 875175
rect 75473 875119 75559 875175
rect 75615 875119 75701 875175
rect 75757 875119 75816 875175
rect 70000 875065 75816 875119
rect 70000 875009 70047 875065
rect 70103 875009 70171 875065
rect 70227 875009 70295 875065
rect 70351 875009 70419 875065
rect 70475 875033 75816 875065
rect 70475 875009 73855 875033
rect 70000 874977 73855 875009
rect 73911 874977 73997 875033
rect 74053 874977 74139 875033
rect 74195 874977 74281 875033
rect 74337 874977 74423 875033
rect 74479 874977 74565 875033
rect 74621 874977 74707 875033
rect 74763 874977 74849 875033
rect 74905 874977 74991 875033
rect 75047 874977 75133 875033
rect 75189 874977 75275 875033
rect 75331 874977 75417 875033
rect 75473 874977 75559 875033
rect 75615 874977 75701 875033
rect 75757 874977 75816 875033
rect 70000 874941 75816 874977
rect 70000 874885 70047 874941
rect 70103 874885 70171 874941
rect 70227 874885 70295 874941
rect 70351 874885 70419 874941
rect 70475 874891 75816 874941
rect 70475 874885 73855 874891
rect 70000 874835 73855 874885
rect 73911 874835 73997 874891
rect 74053 874835 74139 874891
rect 74195 874835 74281 874891
rect 74337 874835 74423 874891
rect 74479 874835 74565 874891
rect 74621 874835 74707 874891
rect 74763 874835 74849 874891
rect 74905 874835 74991 874891
rect 75047 874835 75133 874891
rect 75189 874835 75275 874891
rect 75331 874835 75417 874891
rect 75473 874835 75559 874891
rect 75615 874835 75701 874891
rect 75757 874835 75816 874891
rect 70000 874817 75816 874835
rect 70000 874761 70047 874817
rect 70103 874761 70171 874817
rect 70227 874761 70295 874817
rect 70351 874761 70419 874817
rect 70475 874761 75816 874817
rect 70000 874749 75816 874761
rect 70000 874693 73855 874749
rect 73911 874693 73997 874749
rect 74053 874693 74139 874749
rect 74195 874693 74281 874749
rect 74337 874693 74423 874749
rect 74479 874693 74565 874749
rect 74621 874693 74707 874749
rect 74763 874693 74849 874749
rect 74905 874693 74991 874749
rect 75047 874693 75133 874749
rect 75189 874693 75275 874749
rect 75331 874693 75417 874749
rect 75473 874693 75559 874749
rect 75615 874693 75701 874749
rect 75757 874693 75816 874749
rect 70000 874637 70047 874693
rect 70103 874637 70171 874693
rect 70227 874637 70295 874693
rect 70351 874637 70419 874693
rect 70475 874637 75816 874693
rect 70000 874607 75816 874637
rect 70000 874569 73855 874607
rect 70000 874513 70047 874569
rect 70103 874513 70171 874569
rect 70227 874513 70295 874569
rect 70351 874513 70419 874569
rect 70475 874551 73855 874569
rect 73911 874551 73997 874607
rect 74053 874551 74139 874607
rect 74195 874551 74281 874607
rect 74337 874551 74423 874607
rect 74479 874551 74565 874607
rect 74621 874551 74707 874607
rect 74763 874551 74849 874607
rect 74905 874551 74991 874607
rect 75047 874551 75133 874607
rect 75189 874551 75275 874607
rect 75331 874551 75417 874607
rect 75473 874551 75559 874607
rect 75615 874551 75701 874607
rect 75757 874551 75816 874607
rect 70475 874513 75816 874551
rect 70000 874465 75816 874513
rect 70000 874445 73855 874465
rect 70000 874389 70047 874445
rect 70103 874389 70171 874445
rect 70227 874389 70295 874445
rect 70351 874389 70419 874445
rect 70475 874409 73855 874445
rect 73911 874409 73997 874465
rect 74053 874409 74139 874465
rect 74195 874409 74281 874465
rect 74337 874409 74423 874465
rect 74479 874409 74565 874465
rect 74621 874409 74707 874465
rect 74763 874409 74849 874465
rect 74905 874409 74991 874465
rect 75047 874409 75133 874465
rect 75189 874409 75275 874465
rect 75331 874409 75417 874465
rect 75473 874409 75559 874465
rect 75615 874409 75701 874465
rect 75757 874409 75816 874465
rect 70475 874389 75816 874409
rect 70000 874323 75816 874389
rect 70000 874321 73855 874323
rect 70000 874265 70047 874321
rect 70103 874265 70171 874321
rect 70227 874265 70295 874321
rect 70351 874265 70419 874321
rect 70475 874267 73855 874321
rect 73911 874267 73997 874323
rect 74053 874267 74139 874323
rect 74195 874267 74281 874323
rect 74337 874267 74423 874323
rect 74479 874267 74565 874323
rect 74621 874267 74707 874323
rect 74763 874267 74849 874323
rect 74905 874267 74991 874323
rect 75047 874267 75133 874323
rect 75189 874267 75275 874323
rect 75331 874267 75417 874323
rect 75473 874267 75559 874323
rect 75615 874267 75701 874323
rect 75757 874267 75816 874323
rect 70475 874265 75816 874267
rect 70000 874198 75816 874265
rect 699992 875181 706000 875248
rect 699992 875179 705525 875181
rect 699992 875123 700051 875179
rect 700107 875123 700193 875179
rect 700249 875123 700335 875179
rect 700391 875123 700477 875179
rect 700533 875123 700619 875179
rect 700675 875123 700761 875179
rect 700817 875123 700903 875179
rect 700959 875123 701045 875179
rect 701101 875123 701187 875179
rect 701243 875123 701329 875179
rect 701385 875123 701471 875179
rect 701527 875123 701613 875179
rect 701669 875123 701755 875179
rect 701811 875123 701897 875179
rect 701953 875125 705525 875179
rect 705581 875125 705649 875181
rect 705705 875125 705773 875181
rect 705829 875125 705897 875181
rect 705953 875125 706000 875181
rect 701953 875123 706000 875125
rect 699992 875057 706000 875123
rect 699992 875037 705525 875057
rect 699992 874981 700051 875037
rect 700107 874981 700193 875037
rect 700249 874981 700335 875037
rect 700391 874981 700477 875037
rect 700533 874981 700619 875037
rect 700675 874981 700761 875037
rect 700817 874981 700903 875037
rect 700959 874981 701045 875037
rect 701101 874981 701187 875037
rect 701243 874981 701329 875037
rect 701385 874981 701471 875037
rect 701527 874981 701613 875037
rect 701669 874981 701755 875037
rect 701811 874981 701897 875037
rect 701953 875001 705525 875037
rect 705581 875001 705649 875057
rect 705705 875001 705773 875057
rect 705829 875001 705897 875057
rect 705953 875001 706000 875057
rect 701953 874981 706000 875001
rect 699992 874933 706000 874981
rect 699992 874895 705525 874933
rect 699992 874839 700051 874895
rect 700107 874839 700193 874895
rect 700249 874839 700335 874895
rect 700391 874839 700477 874895
rect 700533 874839 700619 874895
rect 700675 874839 700761 874895
rect 700817 874839 700903 874895
rect 700959 874839 701045 874895
rect 701101 874839 701187 874895
rect 701243 874839 701329 874895
rect 701385 874839 701471 874895
rect 701527 874839 701613 874895
rect 701669 874839 701755 874895
rect 701811 874839 701897 874895
rect 701953 874877 705525 874895
rect 705581 874877 705649 874933
rect 705705 874877 705773 874933
rect 705829 874877 705897 874933
rect 705953 874877 706000 874933
rect 701953 874839 706000 874877
rect 699992 874809 706000 874839
rect 699992 874753 705525 874809
rect 705581 874753 705649 874809
rect 705705 874753 705773 874809
rect 705829 874753 705897 874809
rect 705953 874753 706000 874809
rect 699992 874697 700051 874753
rect 700107 874697 700193 874753
rect 700249 874697 700335 874753
rect 700391 874697 700477 874753
rect 700533 874697 700619 874753
rect 700675 874697 700761 874753
rect 700817 874697 700903 874753
rect 700959 874697 701045 874753
rect 701101 874697 701187 874753
rect 701243 874697 701329 874753
rect 701385 874697 701471 874753
rect 701527 874697 701613 874753
rect 701669 874697 701755 874753
rect 701811 874697 701897 874753
rect 701953 874697 706000 874753
rect 699992 874685 706000 874697
rect 699992 874629 705525 874685
rect 705581 874629 705649 874685
rect 705705 874629 705773 874685
rect 705829 874629 705897 874685
rect 705953 874629 706000 874685
rect 699992 874611 706000 874629
rect 699992 874555 700051 874611
rect 700107 874555 700193 874611
rect 700249 874555 700335 874611
rect 700391 874555 700477 874611
rect 700533 874555 700619 874611
rect 700675 874555 700761 874611
rect 700817 874555 700903 874611
rect 700959 874555 701045 874611
rect 701101 874555 701187 874611
rect 701243 874555 701329 874611
rect 701385 874555 701471 874611
rect 701527 874555 701613 874611
rect 701669 874555 701755 874611
rect 701811 874555 701897 874611
rect 701953 874561 706000 874611
rect 701953 874555 705525 874561
rect 699992 874505 705525 874555
rect 705581 874505 705649 874561
rect 705705 874505 705773 874561
rect 705829 874505 705897 874561
rect 705953 874505 706000 874561
rect 699992 874469 706000 874505
rect 699992 874413 700051 874469
rect 700107 874413 700193 874469
rect 700249 874413 700335 874469
rect 700391 874413 700477 874469
rect 700533 874413 700619 874469
rect 700675 874413 700761 874469
rect 700817 874413 700903 874469
rect 700959 874413 701045 874469
rect 701101 874413 701187 874469
rect 701243 874413 701329 874469
rect 701385 874413 701471 874469
rect 701527 874413 701613 874469
rect 701669 874413 701755 874469
rect 701811 874413 701897 874469
rect 701953 874437 706000 874469
rect 701953 874413 705525 874437
rect 699992 874381 705525 874413
rect 705581 874381 705649 874437
rect 705705 874381 705773 874437
rect 705829 874381 705897 874437
rect 705953 874381 706000 874437
rect 699992 874327 706000 874381
rect 699992 874271 700051 874327
rect 700107 874271 700193 874327
rect 700249 874271 700335 874327
rect 700391 874271 700477 874327
rect 700533 874271 700619 874327
rect 700675 874271 700761 874327
rect 700817 874271 700903 874327
rect 700959 874271 701045 874327
rect 701101 874271 701187 874327
rect 701243 874271 701329 874327
rect 701385 874271 701471 874327
rect 701527 874271 701613 874327
rect 701669 874271 701755 874327
rect 701811 874271 701897 874327
rect 701953 874313 706000 874327
rect 701953 874271 705525 874313
rect 699992 874257 705525 874271
rect 705581 874257 705649 874313
rect 705705 874257 705773 874313
rect 705829 874257 705897 874313
rect 705953 874257 706000 874313
rect 699992 874189 706000 874257
rect 699992 874185 705525 874189
rect 699992 874129 700051 874185
rect 700107 874129 700193 874185
rect 700249 874129 700335 874185
rect 700391 874129 700477 874185
rect 700533 874129 700619 874185
rect 700675 874129 700761 874185
rect 700817 874129 700903 874185
rect 700959 874129 701045 874185
rect 701101 874129 701187 874185
rect 701243 874129 701329 874185
rect 701385 874129 701471 874185
rect 701527 874129 701613 874185
rect 701669 874129 701755 874185
rect 701811 874129 701897 874185
rect 701953 874133 705525 874185
rect 705581 874133 705649 874189
rect 705705 874133 705773 874189
rect 705829 874133 705897 874189
rect 705953 874133 706000 874189
rect 701953 874129 706000 874133
rect 699992 874065 706000 874129
rect 699992 874043 705525 874065
rect 699992 873987 700051 874043
rect 700107 873987 700193 874043
rect 700249 873987 700335 874043
rect 700391 873987 700477 874043
rect 700533 873987 700619 874043
rect 700675 873987 700761 874043
rect 700817 873987 700903 874043
rect 700959 873987 701045 874043
rect 701101 873987 701187 874043
rect 701243 873987 701329 874043
rect 701385 873987 701471 874043
rect 701527 873987 701613 874043
rect 701669 873987 701755 874043
rect 701811 873987 701897 874043
rect 701953 874009 705525 874043
rect 705581 874009 705649 874065
rect 705705 874009 705773 874065
rect 705829 874009 705897 874065
rect 705953 874009 706000 874065
rect 701953 873987 706000 874009
rect 699992 873941 706000 873987
rect 699992 873901 705525 873941
rect 70000 873811 75816 873878
rect 70000 873755 70047 873811
rect 70103 873755 70171 873811
rect 70227 873755 70295 873811
rect 70351 873755 70419 873811
rect 70475 873799 75816 873811
rect 70475 873755 73855 873799
rect 70000 873743 73855 873755
rect 73911 873743 73997 873799
rect 74053 873743 74139 873799
rect 74195 873743 74281 873799
rect 74337 873743 74423 873799
rect 74479 873743 74565 873799
rect 74621 873743 74707 873799
rect 74763 873743 74849 873799
rect 74905 873743 74991 873799
rect 75047 873743 75133 873799
rect 75189 873743 75275 873799
rect 75331 873743 75417 873799
rect 75473 873743 75559 873799
rect 75615 873743 75701 873799
rect 75757 873743 75816 873799
rect 70000 873687 75816 873743
rect 70000 873631 70047 873687
rect 70103 873631 70171 873687
rect 70227 873631 70295 873687
rect 70351 873631 70419 873687
rect 70475 873657 75816 873687
rect 70475 873631 73855 873657
rect 70000 873601 73855 873631
rect 73911 873601 73997 873657
rect 74053 873601 74139 873657
rect 74195 873601 74281 873657
rect 74337 873601 74423 873657
rect 74479 873601 74565 873657
rect 74621 873601 74707 873657
rect 74763 873601 74849 873657
rect 74905 873601 74991 873657
rect 75047 873601 75133 873657
rect 75189 873601 75275 873657
rect 75331 873601 75417 873657
rect 75473 873601 75559 873657
rect 75615 873601 75701 873657
rect 75757 873601 75816 873657
rect 70000 873563 75816 873601
rect 70000 873507 70047 873563
rect 70103 873507 70171 873563
rect 70227 873507 70295 873563
rect 70351 873507 70419 873563
rect 70475 873515 75816 873563
rect 70475 873507 73855 873515
rect 70000 873459 73855 873507
rect 73911 873459 73997 873515
rect 74053 873459 74139 873515
rect 74195 873459 74281 873515
rect 74337 873459 74423 873515
rect 74479 873459 74565 873515
rect 74621 873459 74707 873515
rect 74763 873459 74849 873515
rect 74905 873459 74991 873515
rect 75047 873459 75133 873515
rect 75189 873459 75275 873515
rect 75331 873459 75417 873515
rect 75473 873459 75559 873515
rect 75615 873459 75701 873515
rect 75757 873459 75816 873515
rect 70000 873439 75816 873459
rect 70000 873383 70047 873439
rect 70103 873383 70171 873439
rect 70227 873383 70295 873439
rect 70351 873383 70419 873439
rect 70475 873383 75816 873439
rect 70000 873373 75816 873383
rect 70000 873317 73855 873373
rect 73911 873317 73997 873373
rect 74053 873317 74139 873373
rect 74195 873317 74281 873373
rect 74337 873317 74423 873373
rect 74479 873317 74565 873373
rect 74621 873317 74707 873373
rect 74763 873317 74849 873373
rect 74905 873317 74991 873373
rect 75047 873317 75133 873373
rect 75189 873317 75275 873373
rect 75331 873317 75417 873373
rect 75473 873317 75559 873373
rect 75615 873317 75701 873373
rect 75757 873317 75816 873373
rect 70000 873315 75816 873317
rect 70000 873259 70047 873315
rect 70103 873259 70171 873315
rect 70227 873259 70295 873315
rect 70351 873259 70419 873315
rect 70475 873259 75816 873315
rect 70000 873231 75816 873259
rect 70000 873191 73855 873231
rect 70000 873135 70047 873191
rect 70103 873135 70171 873191
rect 70227 873135 70295 873191
rect 70351 873135 70419 873191
rect 70475 873175 73855 873191
rect 73911 873175 73997 873231
rect 74053 873175 74139 873231
rect 74195 873175 74281 873231
rect 74337 873175 74423 873231
rect 74479 873175 74565 873231
rect 74621 873175 74707 873231
rect 74763 873175 74849 873231
rect 74905 873175 74991 873231
rect 75047 873175 75133 873231
rect 75189 873175 75275 873231
rect 75331 873175 75417 873231
rect 75473 873175 75559 873231
rect 75615 873175 75701 873231
rect 75757 873175 75816 873231
rect 699992 873845 700051 873901
rect 700107 873845 700193 873901
rect 700249 873845 700335 873901
rect 700391 873845 700477 873901
rect 700533 873845 700619 873901
rect 700675 873845 700761 873901
rect 700817 873845 700903 873901
rect 700959 873845 701045 873901
rect 701101 873845 701187 873901
rect 701243 873845 701329 873901
rect 701385 873845 701471 873901
rect 701527 873845 701613 873901
rect 701669 873845 701755 873901
rect 701811 873845 701897 873901
rect 701953 873885 705525 873901
rect 705581 873885 705649 873941
rect 705705 873885 705773 873941
rect 705829 873885 705897 873941
rect 705953 873885 706000 873941
rect 701953 873845 706000 873885
rect 699992 873817 706000 873845
rect 699992 873761 705525 873817
rect 705581 873761 705649 873817
rect 705705 873761 705773 873817
rect 705829 873761 705897 873817
rect 705953 873761 706000 873817
rect 699992 873759 706000 873761
rect 699992 873703 700051 873759
rect 700107 873703 700193 873759
rect 700249 873703 700335 873759
rect 700391 873703 700477 873759
rect 700533 873703 700619 873759
rect 700675 873703 700761 873759
rect 700817 873703 700903 873759
rect 700959 873703 701045 873759
rect 701101 873703 701187 873759
rect 701243 873703 701329 873759
rect 701385 873703 701471 873759
rect 701527 873703 701613 873759
rect 701669 873703 701755 873759
rect 701811 873703 701897 873759
rect 701953 873703 706000 873759
rect 699992 873693 706000 873703
rect 699992 873637 705525 873693
rect 705581 873637 705649 873693
rect 705705 873637 705773 873693
rect 705829 873637 705897 873693
rect 705953 873637 706000 873693
rect 699992 873617 706000 873637
rect 699992 873561 700051 873617
rect 700107 873561 700193 873617
rect 700249 873561 700335 873617
rect 700391 873561 700477 873617
rect 700533 873561 700619 873617
rect 700675 873561 700761 873617
rect 700817 873561 700903 873617
rect 700959 873561 701045 873617
rect 701101 873561 701187 873617
rect 701243 873561 701329 873617
rect 701385 873561 701471 873617
rect 701527 873561 701613 873617
rect 701669 873561 701755 873617
rect 701811 873561 701897 873617
rect 701953 873569 706000 873617
rect 701953 873561 705525 873569
rect 699992 873513 705525 873561
rect 705581 873513 705649 873569
rect 705705 873513 705773 873569
rect 705829 873513 705897 873569
rect 705953 873513 706000 873569
rect 699992 873475 706000 873513
rect 699992 873419 700051 873475
rect 700107 873419 700193 873475
rect 700249 873419 700335 873475
rect 700391 873419 700477 873475
rect 700533 873419 700619 873475
rect 700675 873419 700761 873475
rect 700817 873419 700903 873475
rect 700959 873419 701045 873475
rect 701101 873419 701187 873475
rect 701243 873419 701329 873475
rect 701385 873419 701471 873475
rect 701527 873419 701613 873475
rect 701669 873419 701755 873475
rect 701811 873419 701897 873475
rect 701953 873445 706000 873475
rect 701953 873419 705525 873445
rect 699992 873389 705525 873419
rect 705581 873389 705649 873445
rect 705705 873389 705773 873445
rect 705829 873389 705897 873445
rect 705953 873389 706000 873445
rect 699992 873333 706000 873389
rect 699992 873277 700051 873333
rect 700107 873277 700193 873333
rect 700249 873277 700335 873333
rect 700391 873277 700477 873333
rect 700533 873277 700619 873333
rect 700675 873277 700761 873333
rect 700817 873277 700903 873333
rect 700959 873277 701045 873333
rect 701101 873277 701187 873333
rect 701243 873277 701329 873333
rect 701385 873277 701471 873333
rect 701527 873277 701613 873333
rect 701669 873277 701755 873333
rect 701811 873277 701897 873333
rect 701953 873321 706000 873333
rect 701953 873277 705525 873321
rect 699992 873265 705525 873277
rect 705581 873265 705649 873321
rect 705705 873265 705773 873321
rect 705829 873265 705897 873321
rect 705953 873265 706000 873321
rect 699992 873198 706000 873265
rect 70475 873135 75816 873175
rect 70000 873089 75816 873135
rect 70000 873067 73855 873089
rect 70000 873011 70047 873067
rect 70103 873011 70171 873067
rect 70227 873011 70295 873067
rect 70351 873011 70419 873067
rect 70475 873033 73855 873067
rect 73911 873033 73997 873089
rect 74053 873033 74139 873089
rect 74195 873033 74281 873089
rect 74337 873033 74423 873089
rect 74479 873033 74565 873089
rect 74621 873033 74707 873089
rect 74763 873033 74849 873089
rect 74905 873033 74991 873089
rect 75047 873033 75133 873089
rect 75189 873033 75275 873089
rect 75331 873033 75417 873089
rect 75473 873033 75559 873089
rect 75615 873033 75701 873089
rect 75757 873033 75816 873089
rect 70475 873011 75816 873033
rect 70000 872947 75816 873011
rect 70000 872943 73855 872947
rect 70000 872887 70047 872943
rect 70103 872887 70171 872943
rect 70227 872887 70295 872943
rect 70351 872887 70419 872943
rect 70475 872891 73855 872943
rect 73911 872891 73997 872947
rect 74053 872891 74139 872947
rect 74195 872891 74281 872947
rect 74337 872891 74423 872947
rect 74479 872891 74565 872947
rect 74621 872891 74707 872947
rect 74763 872891 74849 872947
rect 74905 872891 74991 872947
rect 75047 872891 75133 872947
rect 75189 872891 75275 872947
rect 75331 872891 75417 872947
rect 75473 872891 75559 872947
rect 75615 872891 75701 872947
rect 75757 872891 75816 872947
rect 70475 872887 75816 872891
rect 70000 872819 75816 872887
rect 70000 872763 70047 872819
rect 70103 872763 70171 872819
rect 70227 872763 70295 872819
rect 70351 872763 70419 872819
rect 70475 872805 75816 872819
rect 70475 872763 73855 872805
rect 70000 872749 73855 872763
rect 73911 872749 73997 872805
rect 74053 872749 74139 872805
rect 74195 872749 74281 872805
rect 74337 872749 74423 872805
rect 74479 872749 74565 872805
rect 74621 872749 74707 872805
rect 74763 872749 74849 872805
rect 74905 872749 74991 872805
rect 75047 872749 75133 872805
rect 75189 872749 75275 872805
rect 75331 872749 75417 872805
rect 75473 872749 75559 872805
rect 75615 872749 75701 872805
rect 75757 872749 75816 872805
rect 70000 872695 75816 872749
rect 70000 872639 70047 872695
rect 70103 872639 70171 872695
rect 70227 872639 70295 872695
rect 70351 872639 70419 872695
rect 70475 872663 75816 872695
rect 70475 872639 73855 872663
rect 70000 872607 73855 872639
rect 73911 872607 73997 872663
rect 74053 872607 74139 872663
rect 74195 872607 74281 872663
rect 74337 872607 74423 872663
rect 74479 872607 74565 872663
rect 74621 872607 74707 872663
rect 74763 872607 74849 872663
rect 74905 872607 74991 872663
rect 75047 872607 75133 872663
rect 75189 872607 75275 872663
rect 75331 872607 75417 872663
rect 75473 872607 75559 872663
rect 75615 872607 75701 872663
rect 75757 872607 75816 872663
rect 70000 872571 75816 872607
rect 70000 872515 70047 872571
rect 70103 872515 70171 872571
rect 70227 872515 70295 872571
rect 70351 872515 70419 872571
rect 70475 872521 75816 872571
rect 70475 872515 73855 872521
rect 70000 872465 73855 872515
rect 73911 872465 73997 872521
rect 74053 872465 74139 872521
rect 74195 872465 74281 872521
rect 74337 872465 74423 872521
rect 74479 872465 74565 872521
rect 74621 872465 74707 872521
rect 74763 872465 74849 872521
rect 74905 872465 74991 872521
rect 75047 872465 75133 872521
rect 75189 872465 75275 872521
rect 75331 872465 75417 872521
rect 75473 872465 75559 872521
rect 75615 872465 75701 872521
rect 75757 872465 75816 872521
rect 70000 872447 75816 872465
rect 70000 872391 70047 872447
rect 70103 872391 70171 872447
rect 70227 872391 70295 872447
rect 70351 872391 70419 872447
rect 70475 872391 75816 872447
rect 70000 872379 75816 872391
rect 70000 872323 73855 872379
rect 73911 872323 73997 872379
rect 74053 872323 74139 872379
rect 74195 872323 74281 872379
rect 74337 872323 74423 872379
rect 74479 872323 74565 872379
rect 74621 872323 74707 872379
rect 74763 872323 74849 872379
rect 74905 872323 74991 872379
rect 75047 872323 75133 872379
rect 75189 872323 75275 872379
rect 75331 872323 75417 872379
rect 75473 872323 75559 872379
rect 75615 872323 75701 872379
rect 75757 872323 75816 872379
rect 70000 872267 70047 872323
rect 70103 872267 70171 872323
rect 70227 872267 70295 872323
rect 70351 872267 70419 872323
rect 70475 872267 75816 872323
rect 70000 872237 75816 872267
rect 70000 872199 73855 872237
rect 70000 872143 70047 872199
rect 70103 872143 70171 872199
rect 70227 872143 70295 872199
rect 70351 872143 70419 872199
rect 70475 872181 73855 872199
rect 73911 872181 73997 872237
rect 74053 872181 74139 872237
rect 74195 872181 74281 872237
rect 74337 872181 74423 872237
rect 74479 872181 74565 872237
rect 74621 872181 74707 872237
rect 74763 872181 74849 872237
rect 74905 872181 74991 872237
rect 75047 872181 75133 872237
rect 75189 872181 75275 872237
rect 75331 872181 75417 872237
rect 75473 872181 75559 872237
rect 75615 872181 75701 872237
rect 75757 872181 75816 872237
rect 70475 872143 75816 872181
rect 70000 872095 75816 872143
rect 70000 872075 73855 872095
rect 70000 872019 70047 872075
rect 70103 872019 70171 872075
rect 70227 872019 70295 872075
rect 70351 872019 70419 872075
rect 70475 872039 73855 872075
rect 73911 872039 73997 872095
rect 74053 872039 74139 872095
rect 74195 872039 74281 872095
rect 74337 872039 74423 872095
rect 74479 872039 74565 872095
rect 74621 872039 74707 872095
rect 74763 872039 74849 872095
rect 74905 872039 74991 872095
rect 75047 872039 75133 872095
rect 75189 872039 75275 872095
rect 75331 872039 75417 872095
rect 75473 872039 75559 872095
rect 75615 872039 75701 872095
rect 75757 872039 75816 872095
rect 70475 872019 75816 872039
rect 70000 871953 75816 872019
rect 70000 871951 73855 871953
rect 70000 871895 70047 871951
rect 70103 871895 70171 871951
rect 70227 871895 70295 871951
rect 70351 871895 70419 871951
rect 70475 871897 73855 871951
rect 73911 871897 73997 871953
rect 74053 871897 74139 871953
rect 74195 871897 74281 871953
rect 74337 871897 74423 871953
rect 74479 871897 74565 871953
rect 74621 871897 74707 871953
rect 74763 871897 74849 871953
rect 74905 871897 74991 871953
rect 75047 871897 75133 871953
rect 75189 871897 75275 871953
rect 75331 871897 75417 871953
rect 75473 871897 75559 871953
rect 75615 871897 75701 871953
rect 75757 871897 75816 871953
rect 70475 871895 75816 871897
rect 70000 871828 75816 871895
rect 699992 872811 706000 872878
rect 699992 872809 705525 872811
rect 699992 872753 700051 872809
rect 700107 872753 700193 872809
rect 700249 872753 700335 872809
rect 700391 872753 700477 872809
rect 700533 872753 700619 872809
rect 700675 872753 700761 872809
rect 700817 872753 700903 872809
rect 700959 872753 701045 872809
rect 701101 872753 701187 872809
rect 701243 872753 701329 872809
rect 701385 872753 701471 872809
rect 701527 872753 701613 872809
rect 701669 872753 701755 872809
rect 701811 872753 701897 872809
rect 701953 872755 705525 872809
rect 705581 872755 705649 872811
rect 705705 872755 705773 872811
rect 705829 872755 705897 872811
rect 705953 872755 706000 872811
rect 701953 872753 706000 872755
rect 699992 872687 706000 872753
rect 699992 872667 705525 872687
rect 699992 872611 700051 872667
rect 700107 872611 700193 872667
rect 700249 872611 700335 872667
rect 700391 872611 700477 872667
rect 700533 872611 700619 872667
rect 700675 872611 700761 872667
rect 700817 872611 700903 872667
rect 700959 872611 701045 872667
rect 701101 872611 701187 872667
rect 701243 872611 701329 872667
rect 701385 872611 701471 872667
rect 701527 872611 701613 872667
rect 701669 872611 701755 872667
rect 701811 872611 701897 872667
rect 701953 872631 705525 872667
rect 705581 872631 705649 872687
rect 705705 872631 705773 872687
rect 705829 872631 705897 872687
rect 705953 872631 706000 872687
rect 701953 872611 706000 872631
rect 699992 872563 706000 872611
rect 699992 872525 705525 872563
rect 699992 872469 700051 872525
rect 700107 872469 700193 872525
rect 700249 872469 700335 872525
rect 700391 872469 700477 872525
rect 700533 872469 700619 872525
rect 700675 872469 700761 872525
rect 700817 872469 700903 872525
rect 700959 872469 701045 872525
rect 701101 872469 701187 872525
rect 701243 872469 701329 872525
rect 701385 872469 701471 872525
rect 701527 872469 701613 872525
rect 701669 872469 701755 872525
rect 701811 872469 701897 872525
rect 701953 872507 705525 872525
rect 705581 872507 705649 872563
rect 705705 872507 705773 872563
rect 705829 872507 705897 872563
rect 705953 872507 706000 872563
rect 701953 872469 706000 872507
rect 699992 872439 706000 872469
rect 699992 872383 705525 872439
rect 705581 872383 705649 872439
rect 705705 872383 705773 872439
rect 705829 872383 705897 872439
rect 705953 872383 706000 872439
rect 699992 872327 700051 872383
rect 700107 872327 700193 872383
rect 700249 872327 700335 872383
rect 700391 872327 700477 872383
rect 700533 872327 700619 872383
rect 700675 872327 700761 872383
rect 700817 872327 700903 872383
rect 700959 872327 701045 872383
rect 701101 872327 701187 872383
rect 701243 872327 701329 872383
rect 701385 872327 701471 872383
rect 701527 872327 701613 872383
rect 701669 872327 701755 872383
rect 701811 872327 701897 872383
rect 701953 872327 706000 872383
rect 699992 872315 706000 872327
rect 699992 872259 705525 872315
rect 705581 872259 705649 872315
rect 705705 872259 705773 872315
rect 705829 872259 705897 872315
rect 705953 872259 706000 872315
rect 699992 872241 706000 872259
rect 699992 872185 700051 872241
rect 700107 872185 700193 872241
rect 700249 872185 700335 872241
rect 700391 872185 700477 872241
rect 700533 872185 700619 872241
rect 700675 872185 700761 872241
rect 700817 872185 700903 872241
rect 700959 872185 701045 872241
rect 701101 872185 701187 872241
rect 701243 872185 701329 872241
rect 701385 872185 701471 872241
rect 701527 872185 701613 872241
rect 701669 872185 701755 872241
rect 701811 872185 701897 872241
rect 701953 872191 706000 872241
rect 701953 872185 705525 872191
rect 699992 872135 705525 872185
rect 705581 872135 705649 872191
rect 705705 872135 705773 872191
rect 705829 872135 705897 872191
rect 705953 872135 706000 872191
rect 699992 872099 706000 872135
rect 699992 872043 700051 872099
rect 700107 872043 700193 872099
rect 700249 872043 700335 872099
rect 700391 872043 700477 872099
rect 700533 872043 700619 872099
rect 700675 872043 700761 872099
rect 700817 872043 700903 872099
rect 700959 872043 701045 872099
rect 701101 872043 701187 872099
rect 701243 872043 701329 872099
rect 701385 872043 701471 872099
rect 701527 872043 701613 872099
rect 701669 872043 701755 872099
rect 701811 872043 701897 872099
rect 701953 872067 706000 872099
rect 701953 872043 705525 872067
rect 699992 872011 705525 872043
rect 705581 872011 705649 872067
rect 705705 872011 705773 872067
rect 705829 872011 705897 872067
rect 705953 872011 706000 872067
rect 699992 871957 706000 872011
rect 699992 871901 700051 871957
rect 700107 871901 700193 871957
rect 700249 871901 700335 871957
rect 700391 871901 700477 871957
rect 700533 871901 700619 871957
rect 700675 871901 700761 871957
rect 700817 871901 700903 871957
rect 700959 871901 701045 871957
rect 701101 871901 701187 871957
rect 701243 871901 701329 871957
rect 701385 871901 701471 871957
rect 701527 871901 701613 871957
rect 701669 871901 701755 871957
rect 701811 871901 701897 871957
rect 701953 871943 706000 871957
rect 701953 871901 705525 871943
rect 699992 871887 705525 871901
rect 705581 871887 705649 871943
rect 705705 871887 705773 871943
rect 705829 871887 705897 871943
rect 705953 871887 706000 871943
rect 699992 871819 706000 871887
rect 699992 871815 705525 871819
rect 699992 871759 700051 871815
rect 700107 871759 700193 871815
rect 700249 871759 700335 871815
rect 700391 871759 700477 871815
rect 700533 871759 700619 871815
rect 700675 871759 700761 871815
rect 700817 871759 700903 871815
rect 700959 871759 701045 871815
rect 701101 871759 701187 871815
rect 701243 871759 701329 871815
rect 701385 871759 701471 871815
rect 701527 871759 701613 871815
rect 701669 871759 701755 871815
rect 701811 871759 701897 871815
rect 701953 871763 705525 871815
rect 705581 871763 705649 871819
rect 705705 871763 705773 871819
rect 705829 871763 705897 871819
rect 705953 871763 706000 871819
rect 701953 871759 706000 871763
rect 699992 871695 706000 871759
rect 699992 871673 705525 871695
rect 699992 871617 700051 871673
rect 700107 871617 700193 871673
rect 700249 871617 700335 871673
rect 700391 871617 700477 871673
rect 700533 871617 700619 871673
rect 700675 871617 700761 871673
rect 700817 871617 700903 871673
rect 700959 871617 701045 871673
rect 701101 871617 701187 871673
rect 701243 871617 701329 871673
rect 701385 871617 701471 871673
rect 701527 871617 701613 871673
rect 701669 871617 701755 871673
rect 701811 871617 701897 871673
rect 701953 871639 705525 871673
rect 705581 871639 705649 871695
rect 705705 871639 705773 871695
rect 705829 871639 705897 871695
rect 705953 871639 706000 871695
rect 701953 871617 706000 871639
rect 699992 871571 706000 871617
rect 699992 871531 705525 871571
rect 699992 871475 700051 871531
rect 700107 871475 700193 871531
rect 700249 871475 700335 871531
rect 700391 871475 700477 871531
rect 700533 871475 700619 871531
rect 700675 871475 700761 871531
rect 700817 871475 700903 871531
rect 700959 871475 701045 871531
rect 701101 871475 701187 871531
rect 701243 871475 701329 871531
rect 701385 871475 701471 871531
rect 701527 871475 701613 871531
rect 701669 871475 701755 871531
rect 701811 871475 701897 871531
rect 701953 871515 705525 871531
rect 705581 871515 705649 871571
rect 705705 871515 705773 871571
rect 705829 871515 705897 871571
rect 705953 871515 706000 871571
rect 701953 871475 706000 871515
rect 699992 871447 706000 871475
rect 699992 871391 705525 871447
rect 705581 871391 705649 871447
rect 705705 871391 705773 871447
rect 705829 871391 705897 871447
rect 705953 871391 706000 871447
rect 699992 871389 706000 871391
rect 699992 871333 700051 871389
rect 700107 871333 700193 871389
rect 700249 871333 700335 871389
rect 700391 871333 700477 871389
rect 700533 871333 700619 871389
rect 700675 871333 700761 871389
rect 700817 871333 700903 871389
rect 700959 871333 701045 871389
rect 701101 871333 701187 871389
rect 701243 871333 701329 871389
rect 701385 871333 701471 871389
rect 701527 871333 701613 871389
rect 701669 871333 701755 871389
rect 701811 871333 701897 871389
rect 701953 871333 706000 871389
rect 699992 871323 706000 871333
rect 699992 871267 705525 871323
rect 705581 871267 705649 871323
rect 705705 871267 705773 871323
rect 705829 871267 705897 871323
rect 705953 871267 706000 871323
rect 699992 871247 706000 871267
rect 699992 871191 700051 871247
rect 700107 871191 700193 871247
rect 700249 871191 700335 871247
rect 700391 871191 700477 871247
rect 700533 871191 700619 871247
rect 700675 871191 700761 871247
rect 700817 871191 700903 871247
rect 700959 871191 701045 871247
rect 701101 871191 701187 871247
rect 701243 871191 701329 871247
rect 701385 871191 701471 871247
rect 701527 871191 701613 871247
rect 701669 871191 701755 871247
rect 701811 871191 701897 871247
rect 701953 871199 706000 871247
rect 701953 871191 705525 871199
rect 70000 871105 75816 871172
rect 70000 871049 70047 871105
rect 70103 871049 70171 871105
rect 70227 871049 70295 871105
rect 70351 871049 70419 871105
rect 70475 871093 75816 871105
rect 70475 871049 73855 871093
rect 70000 871037 73855 871049
rect 73911 871037 73997 871093
rect 74053 871037 74139 871093
rect 74195 871037 74281 871093
rect 74337 871037 74423 871093
rect 74479 871037 74565 871093
rect 74621 871037 74707 871093
rect 74763 871037 74849 871093
rect 74905 871037 74991 871093
rect 75047 871037 75133 871093
rect 75189 871037 75275 871093
rect 75331 871037 75417 871093
rect 75473 871037 75559 871093
rect 75615 871037 75701 871093
rect 75757 871037 75816 871093
rect 70000 870981 75816 871037
rect 70000 870925 70047 870981
rect 70103 870925 70171 870981
rect 70227 870925 70295 870981
rect 70351 870925 70419 870981
rect 70475 870951 75816 870981
rect 70475 870925 73855 870951
rect 70000 870895 73855 870925
rect 73911 870895 73997 870951
rect 74053 870895 74139 870951
rect 74195 870895 74281 870951
rect 74337 870895 74423 870951
rect 74479 870895 74565 870951
rect 74621 870895 74707 870951
rect 74763 870895 74849 870951
rect 74905 870895 74991 870951
rect 75047 870895 75133 870951
rect 75189 870895 75275 870951
rect 75331 870895 75417 870951
rect 75473 870895 75559 870951
rect 75615 870895 75701 870951
rect 75757 870895 75816 870951
rect 70000 870857 75816 870895
rect 70000 870801 70047 870857
rect 70103 870801 70171 870857
rect 70227 870801 70295 870857
rect 70351 870801 70419 870857
rect 70475 870809 75816 870857
rect 699992 871143 705525 871191
rect 705581 871143 705649 871199
rect 705705 871143 705773 871199
rect 705829 871143 705897 871199
rect 705953 871143 706000 871199
rect 699992 871105 706000 871143
rect 699992 871049 700051 871105
rect 700107 871049 700193 871105
rect 700249 871049 700335 871105
rect 700391 871049 700477 871105
rect 700533 871049 700619 871105
rect 700675 871049 700761 871105
rect 700817 871049 700903 871105
rect 700959 871049 701045 871105
rect 701101 871049 701187 871105
rect 701243 871049 701329 871105
rect 701385 871049 701471 871105
rect 701527 871049 701613 871105
rect 701669 871049 701755 871105
rect 701811 871049 701897 871105
rect 701953 871075 706000 871105
rect 701953 871049 705525 871075
rect 699992 871019 705525 871049
rect 705581 871019 705649 871075
rect 705705 871019 705773 871075
rect 705829 871019 705897 871075
rect 705953 871019 706000 871075
rect 699992 870963 706000 871019
rect 699992 870907 700051 870963
rect 700107 870907 700193 870963
rect 700249 870907 700335 870963
rect 700391 870907 700477 870963
rect 700533 870907 700619 870963
rect 700675 870907 700761 870963
rect 700817 870907 700903 870963
rect 700959 870907 701045 870963
rect 701101 870907 701187 870963
rect 701243 870907 701329 870963
rect 701385 870907 701471 870963
rect 701527 870907 701613 870963
rect 701669 870907 701755 870963
rect 701811 870907 701897 870963
rect 701953 870951 706000 870963
rect 701953 870907 705525 870951
rect 699992 870895 705525 870907
rect 705581 870895 705649 870951
rect 705705 870895 705773 870951
rect 705829 870895 705897 870951
rect 705953 870895 706000 870951
rect 699992 870828 706000 870895
rect 70475 870801 73855 870809
rect 70000 870753 73855 870801
rect 73911 870753 73997 870809
rect 74053 870753 74139 870809
rect 74195 870753 74281 870809
rect 74337 870753 74423 870809
rect 74479 870753 74565 870809
rect 74621 870753 74707 870809
rect 74763 870753 74849 870809
rect 74905 870753 74991 870809
rect 75047 870753 75133 870809
rect 75189 870753 75275 870809
rect 75331 870753 75417 870809
rect 75473 870753 75559 870809
rect 75615 870753 75701 870809
rect 75757 870753 75816 870809
rect 70000 870733 75816 870753
rect 70000 870677 70047 870733
rect 70103 870677 70171 870733
rect 70227 870677 70295 870733
rect 70351 870677 70419 870733
rect 70475 870677 75816 870733
rect 70000 870667 75816 870677
rect 70000 870611 73855 870667
rect 73911 870611 73997 870667
rect 74053 870611 74139 870667
rect 74195 870611 74281 870667
rect 74337 870611 74423 870667
rect 74479 870611 74565 870667
rect 74621 870611 74707 870667
rect 74763 870611 74849 870667
rect 74905 870611 74991 870667
rect 75047 870611 75133 870667
rect 75189 870611 75275 870667
rect 75331 870611 75417 870667
rect 75473 870611 75559 870667
rect 75615 870611 75701 870667
rect 75757 870611 75816 870667
rect 70000 870609 75816 870611
rect 70000 870553 70047 870609
rect 70103 870553 70171 870609
rect 70227 870553 70295 870609
rect 70351 870553 70419 870609
rect 70475 870553 75816 870609
rect 70000 870525 75816 870553
rect 70000 870485 73855 870525
rect 70000 870429 70047 870485
rect 70103 870429 70171 870485
rect 70227 870429 70295 870485
rect 70351 870429 70419 870485
rect 70475 870469 73855 870485
rect 73911 870469 73997 870525
rect 74053 870469 74139 870525
rect 74195 870469 74281 870525
rect 74337 870469 74423 870525
rect 74479 870469 74565 870525
rect 74621 870469 74707 870525
rect 74763 870469 74849 870525
rect 74905 870469 74991 870525
rect 75047 870469 75133 870525
rect 75189 870469 75275 870525
rect 75331 870469 75417 870525
rect 75473 870469 75559 870525
rect 75615 870469 75701 870525
rect 75757 870469 75816 870525
rect 70475 870429 75816 870469
rect 70000 870383 75816 870429
rect 70000 870361 73855 870383
rect 70000 870305 70047 870361
rect 70103 870305 70171 870361
rect 70227 870305 70295 870361
rect 70351 870305 70419 870361
rect 70475 870327 73855 870361
rect 73911 870327 73997 870383
rect 74053 870327 74139 870383
rect 74195 870327 74281 870383
rect 74337 870327 74423 870383
rect 74479 870327 74565 870383
rect 74621 870327 74707 870383
rect 74763 870327 74849 870383
rect 74905 870327 74991 870383
rect 75047 870327 75133 870383
rect 75189 870327 75275 870383
rect 75331 870327 75417 870383
rect 75473 870327 75559 870383
rect 75615 870327 75701 870383
rect 75757 870327 75816 870383
rect 70475 870305 75816 870327
rect 70000 870241 75816 870305
rect 70000 870237 73855 870241
rect 70000 870181 70047 870237
rect 70103 870181 70171 870237
rect 70227 870181 70295 870237
rect 70351 870181 70419 870237
rect 70475 870185 73855 870237
rect 73911 870185 73997 870241
rect 74053 870185 74139 870241
rect 74195 870185 74281 870241
rect 74337 870185 74423 870241
rect 74479 870185 74565 870241
rect 74621 870185 74707 870241
rect 74763 870185 74849 870241
rect 74905 870185 74991 870241
rect 75047 870185 75133 870241
rect 75189 870185 75275 870241
rect 75331 870185 75417 870241
rect 75473 870185 75559 870241
rect 75615 870185 75701 870241
rect 75757 870185 75816 870241
rect 70475 870181 75816 870185
rect 70000 870113 75816 870181
rect 70000 870057 70047 870113
rect 70103 870057 70171 870113
rect 70227 870057 70295 870113
rect 70351 870057 70419 870113
rect 70475 870099 75816 870113
rect 70475 870057 73855 870099
rect 70000 870043 73855 870057
rect 73911 870043 73997 870099
rect 74053 870043 74139 870099
rect 74195 870043 74281 870099
rect 74337 870043 74423 870099
rect 74479 870043 74565 870099
rect 74621 870043 74707 870099
rect 74763 870043 74849 870099
rect 74905 870043 74991 870099
rect 75047 870043 75133 870099
rect 75189 870043 75275 870099
rect 75331 870043 75417 870099
rect 75473 870043 75559 870099
rect 75615 870043 75701 870099
rect 75757 870043 75816 870099
rect 70000 869989 75816 870043
rect 70000 869933 70047 869989
rect 70103 869933 70171 869989
rect 70227 869933 70295 869989
rect 70351 869933 70419 869989
rect 70475 869957 75816 869989
rect 70475 869933 73855 869957
rect 70000 869901 73855 869933
rect 73911 869901 73997 869957
rect 74053 869901 74139 869957
rect 74195 869901 74281 869957
rect 74337 869901 74423 869957
rect 74479 869901 74565 869957
rect 74621 869901 74707 869957
rect 74763 869901 74849 869957
rect 74905 869901 74991 869957
rect 75047 869901 75133 869957
rect 75189 869901 75275 869957
rect 75331 869901 75417 869957
rect 75473 869901 75559 869957
rect 75615 869901 75701 869957
rect 75757 869901 75816 869957
rect 70000 869865 75816 869901
rect 70000 869809 70047 869865
rect 70103 869809 70171 869865
rect 70227 869809 70295 869865
rect 70351 869809 70419 869865
rect 70475 869815 75816 869865
rect 70475 869809 73855 869815
rect 70000 869759 73855 869809
rect 73911 869759 73997 869815
rect 74053 869759 74139 869815
rect 74195 869759 74281 869815
rect 74337 869759 74423 869815
rect 74479 869759 74565 869815
rect 74621 869759 74707 869815
rect 74763 869759 74849 869815
rect 74905 869759 74991 869815
rect 75047 869759 75133 869815
rect 75189 869759 75275 869815
rect 75331 869759 75417 869815
rect 75473 869759 75559 869815
rect 75615 869759 75701 869815
rect 75757 869759 75816 869815
rect 70000 869741 75816 869759
rect 70000 869685 70047 869741
rect 70103 869685 70171 869741
rect 70227 869685 70295 869741
rect 70351 869685 70419 869741
rect 70475 869685 75816 869741
rect 70000 869673 75816 869685
rect 70000 869617 73855 869673
rect 73911 869617 73997 869673
rect 74053 869617 74139 869673
rect 74195 869617 74281 869673
rect 74337 869617 74423 869673
rect 74479 869617 74565 869673
rect 74621 869617 74707 869673
rect 74763 869617 74849 869673
rect 74905 869617 74991 869673
rect 75047 869617 75133 869673
rect 75189 869617 75275 869673
rect 75331 869617 75417 869673
rect 75473 869617 75559 869673
rect 75615 869617 75701 869673
rect 75757 869617 75816 869673
rect 70000 869561 70047 869617
rect 70103 869561 70171 869617
rect 70227 869561 70295 869617
rect 70351 869561 70419 869617
rect 70475 869561 75816 869617
rect 70000 869531 75816 869561
rect 70000 869493 73855 869531
rect 70000 869437 70047 869493
rect 70103 869437 70171 869493
rect 70227 869437 70295 869493
rect 70351 869437 70419 869493
rect 70475 869475 73855 869493
rect 73911 869475 73997 869531
rect 74053 869475 74139 869531
rect 74195 869475 74281 869531
rect 74337 869475 74423 869531
rect 74479 869475 74565 869531
rect 74621 869475 74707 869531
rect 74763 869475 74849 869531
rect 74905 869475 74991 869531
rect 75047 869475 75133 869531
rect 75189 869475 75275 869531
rect 75331 869475 75417 869531
rect 75473 869475 75559 869531
rect 75615 869475 75701 869531
rect 75757 869475 75816 869531
rect 70475 869437 75816 869475
rect 70000 869389 75816 869437
rect 70000 869369 73855 869389
rect 70000 869313 70047 869369
rect 70103 869313 70171 869369
rect 70227 869313 70295 869369
rect 70351 869313 70419 869369
rect 70475 869333 73855 869369
rect 73911 869333 73997 869389
rect 74053 869333 74139 869389
rect 74195 869333 74281 869389
rect 74337 869333 74423 869389
rect 74479 869333 74565 869389
rect 74621 869333 74707 869389
rect 74763 869333 74849 869389
rect 74905 869333 74991 869389
rect 75047 869333 75133 869389
rect 75189 869333 75275 869389
rect 75331 869333 75417 869389
rect 75473 869333 75559 869389
rect 75615 869333 75701 869389
rect 75757 869333 75816 869389
rect 70475 869313 75816 869333
rect 70000 869247 75816 869313
rect 70000 869245 73855 869247
rect 70000 869189 70047 869245
rect 70103 869189 70171 869245
rect 70227 869189 70295 869245
rect 70351 869189 70419 869245
rect 70475 869191 73855 869245
rect 73911 869191 73997 869247
rect 74053 869191 74139 869247
rect 74195 869191 74281 869247
rect 74337 869191 74423 869247
rect 74479 869191 74565 869247
rect 74621 869191 74707 869247
rect 74763 869191 74849 869247
rect 74905 869191 74991 869247
rect 75047 869191 75133 869247
rect 75189 869191 75275 869247
rect 75331 869191 75417 869247
rect 75473 869191 75559 869247
rect 75615 869191 75701 869247
rect 75757 869191 75816 869247
rect 70475 869189 75816 869191
rect 70000 869122 75816 869189
rect 699992 870105 706000 870172
rect 699992 870103 705525 870105
rect 699992 870047 700051 870103
rect 700107 870047 700193 870103
rect 700249 870047 700335 870103
rect 700391 870047 700477 870103
rect 700533 870047 700619 870103
rect 700675 870047 700761 870103
rect 700817 870047 700903 870103
rect 700959 870047 701045 870103
rect 701101 870047 701187 870103
rect 701243 870047 701329 870103
rect 701385 870047 701471 870103
rect 701527 870047 701613 870103
rect 701669 870047 701755 870103
rect 701811 870047 701897 870103
rect 701953 870049 705525 870103
rect 705581 870049 705649 870105
rect 705705 870049 705773 870105
rect 705829 870049 705897 870105
rect 705953 870049 706000 870105
rect 701953 870047 706000 870049
rect 699992 869981 706000 870047
rect 699992 869961 705525 869981
rect 699992 869905 700051 869961
rect 700107 869905 700193 869961
rect 700249 869905 700335 869961
rect 700391 869905 700477 869961
rect 700533 869905 700619 869961
rect 700675 869905 700761 869961
rect 700817 869905 700903 869961
rect 700959 869905 701045 869961
rect 701101 869905 701187 869961
rect 701243 869905 701329 869961
rect 701385 869905 701471 869961
rect 701527 869905 701613 869961
rect 701669 869905 701755 869961
rect 701811 869905 701897 869961
rect 701953 869925 705525 869961
rect 705581 869925 705649 869981
rect 705705 869925 705773 869981
rect 705829 869925 705897 869981
rect 705953 869925 706000 869981
rect 701953 869905 706000 869925
rect 699992 869857 706000 869905
rect 699992 869819 705525 869857
rect 699992 869763 700051 869819
rect 700107 869763 700193 869819
rect 700249 869763 700335 869819
rect 700391 869763 700477 869819
rect 700533 869763 700619 869819
rect 700675 869763 700761 869819
rect 700817 869763 700903 869819
rect 700959 869763 701045 869819
rect 701101 869763 701187 869819
rect 701243 869763 701329 869819
rect 701385 869763 701471 869819
rect 701527 869763 701613 869819
rect 701669 869763 701755 869819
rect 701811 869763 701897 869819
rect 701953 869801 705525 869819
rect 705581 869801 705649 869857
rect 705705 869801 705773 869857
rect 705829 869801 705897 869857
rect 705953 869801 706000 869857
rect 701953 869763 706000 869801
rect 699992 869733 706000 869763
rect 699992 869677 705525 869733
rect 705581 869677 705649 869733
rect 705705 869677 705773 869733
rect 705829 869677 705897 869733
rect 705953 869677 706000 869733
rect 699992 869621 700051 869677
rect 700107 869621 700193 869677
rect 700249 869621 700335 869677
rect 700391 869621 700477 869677
rect 700533 869621 700619 869677
rect 700675 869621 700761 869677
rect 700817 869621 700903 869677
rect 700959 869621 701045 869677
rect 701101 869621 701187 869677
rect 701243 869621 701329 869677
rect 701385 869621 701471 869677
rect 701527 869621 701613 869677
rect 701669 869621 701755 869677
rect 701811 869621 701897 869677
rect 701953 869621 706000 869677
rect 699992 869609 706000 869621
rect 699992 869553 705525 869609
rect 705581 869553 705649 869609
rect 705705 869553 705773 869609
rect 705829 869553 705897 869609
rect 705953 869553 706000 869609
rect 699992 869535 706000 869553
rect 699992 869479 700051 869535
rect 700107 869479 700193 869535
rect 700249 869479 700335 869535
rect 700391 869479 700477 869535
rect 700533 869479 700619 869535
rect 700675 869479 700761 869535
rect 700817 869479 700903 869535
rect 700959 869479 701045 869535
rect 701101 869479 701187 869535
rect 701243 869479 701329 869535
rect 701385 869479 701471 869535
rect 701527 869479 701613 869535
rect 701669 869479 701755 869535
rect 701811 869479 701897 869535
rect 701953 869485 706000 869535
rect 701953 869479 705525 869485
rect 699992 869429 705525 869479
rect 705581 869429 705649 869485
rect 705705 869429 705773 869485
rect 705829 869429 705897 869485
rect 705953 869429 706000 869485
rect 699992 869393 706000 869429
rect 699992 869337 700051 869393
rect 700107 869337 700193 869393
rect 700249 869337 700335 869393
rect 700391 869337 700477 869393
rect 700533 869337 700619 869393
rect 700675 869337 700761 869393
rect 700817 869337 700903 869393
rect 700959 869337 701045 869393
rect 701101 869337 701187 869393
rect 701243 869337 701329 869393
rect 701385 869337 701471 869393
rect 701527 869337 701613 869393
rect 701669 869337 701755 869393
rect 701811 869337 701897 869393
rect 701953 869361 706000 869393
rect 701953 869337 705525 869361
rect 699992 869305 705525 869337
rect 705581 869305 705649 869361
rect 705705 869305 705773 869361
rect 705829 869305 705897 869361
rect 705953 869305 706000 869361
rect 699992 869251 706000 869305
rect 699992 869195 700051 869251
rect 700107 869195 700193 869251
rect 700249 869195 700335 869251
rect 700391 869195 700477 869251
rect 700533 869195 700619 869251
rect 700675 869195 700761 869251
rect 700817 869195 700903 869251
rect 700959 869195 701045 869251
rect 701101 869195 701187 869251
rect 701243 869195 701329 869251
rect 701385 869195 701471 869251
rect 701527 869195 701613 869251
rect 701669 869195 701755 869251
rect 701811 869195 701897 869251
rect 701953 869237 706000 869251
rect 701953 869195 705525 869237
rect 699992 869181 705525 869195
rect 705581 869181 705649 869237
rect 705705 869181 705773 869237
rect 705829 869181 705897 869237
rect 705953 869181 706000 869237
rect 699992 869113 706000 869181
rect 699992 869109 705525 869113
rect 699992 869053 700051 869109
rect 700107 869053 700193 869109
rect 700249 869053 700335 869109
rect 700391 869053 700477 869109
rect 700533 869053 700619 869109
rect 700675 869053 700761 869109
rect 700817 869053 700903 869109
rect 700959 869053 701045 869109
rect 701101 869053 701187 869109
rect 701243 869053 701329 869109
rect 701385 869053 701471 869109
rect 701527 869053 701613 869109
rect 701669 869053 701755 869109
rect 701811 869053 701897 869109
rect 701953 869057 705525 869109
rect 705581 869057 705649 869113
rect 705705 869057 705773 869113
rect 705829 869057 705897 869113
rect 705953 869057 706000 869113
rect 701953 869053 706000 869057
rect 699992 868989 706000 869053
rect 699992 868967 705525 868989
rect 699992 868911 700051 868967
rect 700107 868911 700193 868967
rect 700249 868911 700335 868967
rect 700391 868911 700477 868967
rect 700533 868911 700619 868967
rect 700675 868911 700761 868967
rect 700817 868911 700903 868967
rect 700959 868911 701045 868967
rect 701101 868911 701187 868967
rect 701243 868911 701329 868967
rect 701385 868911 701471 868967
rect 701527 868911 701613 868967
rect 701669 868911 701755 868967
rect 701811 868911 701897 868967
rect 701953 868933 705525 868967
rect 705581 868933 705649 868989
rect 705705 868933 705773 868989
rect 705829 868933 705897 868989
rect 705953 868933 706000 868989
rect 701953 868911 706000 868933
rect 699992 868865 706000 868911
rect 699992 868825 705525 868865
rect 70000 868735 75816 868802
rect 70000 868679 70047 868735
rect 70103 868679 70171 868735
rect 70227 868679 70295 868735
rect 70351 868679 70419 868735
rect 70475 868723 75816 868735
rect 70475 868679 73855 868723
rect 70000 868667 73855 868679
rect 73911 868667 73997 868723
rect 74053 868667 74139 868723
rect 74195 868667 74281 868723
rect 74337 868667 74423 868723
rect 74479 868667 74565 868723
rect 74621 868667 74707 868723
rect 74763 868667 74849 868723
rect 74905 868667 74991 868723
rect 75047 868667 75133 868723
rect 75189 868667 75275 868723
rect 75331 868667 75417 868723
rect 75473 868667 75559 868723
rect 75615 868667 75701 868723
rect 75757 868667 75816 868723
rect 70000 868611 75816 868667
rect 70000 868555 70047 868611
rect 70103 868555 70171 868611
rect 70227 868555 70295 868611
rect 70351 868555 70419 868611
rect 70475 868581 75816 868611
rect 70475 868555 73855 868581
rect 70000 868525 73855 868555
rect 73911 868525 73997 868581
rect 74053 868525 74139 868581
rect 74195 868525 74281 868581
rect 74337 868525 74423 868581
rect 74479 868525 74565 868581
rect 74621 868525 74707 868581
rect 74763 868525 74849 868581
rect 74905 868525 74991 868581
rect 75047 868525 75133 868581
rect 75189 868525 75275 868581
rect 75331 868525 75417 868581
rect 75473 868525 75559 868581
rect 75615 868525 75701 868581
rect 75757 868525 75816 868581
rect 70000 868487 75816 868525
rect 70000 868431 70047 868487
rect 70103 868431 70171 868487
rect 70227 868431 70295 868487
rect 70351 868431 70419 868487
rect 70475 868439 75816 868487
rect 70475 868431 73855 868439
rect 70000 868383 73855 868431
rect 73911 868383 73997 868439
rect 74053 868383 74139 868439
rect 74195 868383 74281 868439
rect 74337 868383 74423 868439
rect 74479 868383 74565 868439
rect 74621 868383 74707 868439
rect 74763 868383 74849 868439
rect 74905 868383 74991 868439
rect 75047 868383 75133 868439
rect 75189 868383 75275 868439
rect 75331 868383 75417 868439
rect 75473 868383 75559 868439
rect 75615 868383 75701 868439
rect 75757 868383 75816 868439
rect 70000 868363 75816 868383
rect 70000 868307 70047 868363
rect 70103 868307 70171 868363
rect 70227 868307 70295 868363
rect 70351 868307 70419 868363
rect 70475 868307 75816 868363
rect 70000 868297 75816 868307
rect 70000 868241 73855 868297
rect 73911 868241 73997 868297
rect 74053 868241 74139 868297
rect 74195 868241 74281 868297
rect 74337 868241 74423 868297
rect 74479 868241 74565 868297
rect 74621 868241 74707 868297
rect 74763 868241 74849 868297
rect 74905 868241 74991 868297
rect 75047 868241 75133 868297
rect 75189 868241 75275 868297
rect 75331 868241 75417 868297
rect 75473 868241 75559 868297
rect 75615 868241 75701 868297
rect 75757 868241 75816 868297
rect 70000 868239 75816 868241
rect 70000 868183 70047 868239
rect 70103 868183 70171 868239
rect 70227 868183 70295 868239
rect 70351 868183 70419 868239
rect 70475 868183 75816 868239
rect 70000 868155 75816 868183
rect 70000 868115 73855 868155
rect 70000 868059 70047 868115
rect 70103 868059 70171 868115
rect 70227 868059 70295 868115
rect 70351 868059 70419 868115
rect 70475 868099 73855 868115
rect 73911 868099 73997 868155
rect 74053 868099 74139 868155
rect 74195 868099 74281 868155
rect 74337 868099 74423 868155
rect 74479 868099 74565 868155
rect 74621 868099 74707 868155
rect 74763 868099 74849 868155
rect 74905 868099 74991 868155
rect 75047 868099 75133 868155
rect 75189 868099 75275 868155
rect 75331 868099 75417 868155
rect 75473 868099 75559 868155
rect 75615 868099 75701 868155
rect 75757 868099 75816 868155
rect 699992 868769 700051 868825
rect 700107 868769 700193 868825
rect 700249 868769 700335 868825
rect 700391 868769 700477 868825
rect 700533 868769 700619 868825
rect 700675 868769 700761 868825
rect 700817 868769 700903 868825
rect 700959 868769 701045 868825
rect 701101 868769 701187 868825
rect 701243 868769 701329 868825
rect 701385 868769 701471 868825
rect 701527 868769 701613 868825
rect 701669 868769 701755 868825
rect 701811 868769 701897 868825
rect 701953 868809 705525 868825
rect 705581 868809 705649 868865
rect 705705 868809 705773 868865
rect 705829 868809 705897 868865
rect 705953 868809 706000 868865
rect 701953 868769 706000 868809
rect 699992 868741 706000 868769
rect 699992 868685 705525 868741
rect 705581 868685 705649 868741
rect 705705 868685 705773 868741
rect 705829 868685 705897 868741
rect 705953 868685 706000 868741
rect 699992 868683 706000 868685
rect 699992 868627 700051 868683
rect 700107 868627 700193 868683
rect 700249 868627 700335 868683
rect 700391 868627 700477 868683
rect 700533 868627 700619 868683
rect 700675 868627 700761 868683
rect 700817 868627 700903 868683
rect 700959 868627 701045 868683
rect 701101 868627 701187 868683
rect 701243 868627 701329 868683
rect 701385 868627 701471 868683
rect 701527 868627 701613 868683
rect 701669 868627 701755 868683
rect 701811 868627 701897 868683
rect 701953 868627 706000 868683
rect 699992 868617 706000 868627
rect 699992 868561 705525 868617
rect 705581 868561 705649 868617
rect 705705 868561 705773 868617
rect 705829 868561 705897 868617
rect 705953 868561 706000 868617
rect 699992 868541 706000 868561
rect 699992 868485 700051 868541
rect 700107 868485 700193 868541
rect 700249 868485 700335 868541
rect 700391 868485 700477 868541
rect 700533 868485 700619 868541
rect 700675 868485 700761 868541
rect 700817 868485 700903 868541
rect 700959 868485 701045 868541
rect 701101 868485 701187 868541
rect 701243 868485 701329 868541
rect 701385 868485 701471 868541
rect 701527 868485 701613 868541
rect 701669 868485 701755 868541
rect 701811 868485 701897 868541
rect 701953 868493 706000 868541
rect 701953 868485 705525 868493
rect 699992 868437 705525 868485
rect 705581 868437 705649 868493
rect 705705 868437 705773 868493
rect 705829 868437 705897 868493
rect 705953 868437 706000 868493
rect 699992 868399 706000 868437
rect 699992 868343 700051 868399
rect 700107 868343 700193 868399
rect 700249 868343 700335 868399
rect 700391 868343 700477 868399
rect 700533 868343 700619 868399
rect 700675 868343 700761 868399
rect 700817 868343 700903 868399
rect 700959 868343 701045 868399
rect 701101 868343 701187 868399
rect 701243 868343 701329 868399
rect 701385 868343 701471 868399
rect 701527 868343 701613 868399
rect 701669 868343 701755 868399
rect 701811 868343 701897 868399
rect 701953 868369 706000 868399
rect 701953 868343 705525 868369
rect 699992 868313 705525 868343
rect 705581 868313 705649 868369
rect 705705 868313 705773 868369
rect 705829 868313 705897 868369
rect 705953 868313 706000 868369
rect 699992 868257 706000 868313
rect 699992 868201 700051 868257
rect 700107 868201 700193 868257
rect 700249 868201 700335 868257
rect 700391 868201 700477 868257
rect 700533 868201 700619 868257
rect 700675 868201 700761 868257
rect 700817 868201 700903 868257
rect 700959 868201 701045 868257
rect 701101 868201 701187 868257
rect 701243 868201 701329 868257
rect 701385 868201 701471 868257
rect 701527 868201 701613 868257
rect 701669 868201 701755 868257
rect 701811 868201 701897 868257
rect 701953 868245 706000 868257
rect 701953 868201 705525 868245
rect 699992 868189 705525 868201
rect 705581 868189 705649 868245
rect 705705 868189 705773 868245
rect 705829 868189 705897 868245
rect 705953 868189 706000 868245
rect 699992 868122 706000 868189
rect 70475 868059 75816 868099
rect 70000 868013 75816 868059
rect 70000 867991 73855 868013
rect 70000 867935 70047 867991
rect 70103 867935 70171 867991
rect 70227 867935 70295 867991
rect 70351 867935 70419 867991
rect 70475 867957 73855 867991
rect 73911 867957 73997 868013
rect 74053 867957 74139 868013
rect 74195 867957 74281 868013
rect 74337 867957 74423 868013
rect 74479 867957 74565 868013
rect 74621 867957 74707 868013
rect 74763 867957 74849 868013
rect 74905 867957 74991 868013
rect 75047 867957 75133 868013
rect 75189 867957 75275 868013
rect 75331 867957 75417 868013
rect 75473 867957 75559 868013
rect 75615 867957 75701 868013
rect 75757 867957 75816 868013
rect 70475 867935 75816 867957
rect 70000 867871 75816 867935
rect 70000 867867 73855 867871
rect 70000 867811 70047 867867
rect 70103 867811 70171 867867
rect 70227 867811 70295 867867
rect 70351 867811 70419 867867
rect 70475 867815 73855 867867
rect 73911 867815 73997 867871
rect 74053 867815 74139 867871
rect 74195 867815 74281 867871
rect 74337 867815 74423 867871
rect 74479 867815 74565 867871
rect 74621 867815 74707 867871
rect 74763 867815 74849 867871
rect 74905 867815 74991 867871
rect 75047 867815 75133 867871
rect 75189 867815 75275 867871
rect 75331 867815 75417 867871
rect 75473 867815 75559 867871
rect 75615 867815 75701 867871
rect 75757 867815 75816 867871
rect 70475 867811 75816 867815
rect 70000 867743 75816 867811
rect 70000 867687 70047 867743
rect 70103 867687 70171 867743
rect 70227 867687 70295 867743
rect 70351 867687 70419 867743
rect 70475 867729 75816 867743
rect 70475 867687 73855 867729
rect 70000 867673 73855 867687
rect 73911 867673 73997 867729
rect 74053 867673 74139 867729
rect 74195 867673 74281 867729
rect 74337 867673 74423 867729
rect 74479 867673 74565 867729
rect 74621 867673 74707 867729
rect 74763 867673 74849 867729
rect 74905 867673 74991 867729
rect 75047 867673 75133 867729
rect 75189 867673 75275 867729
rect 75331 867673 75417 867729
rect 75473 867673 75559 867729
rect 75615 867673 75701 867729
rect 75757 867673 75816 867729
rect 70000 867619 75816 867673
rect 70000 867563 70047 867619
rect 70103 867563 70171 867619
rect 70227 867563 70295 867619
rect 70351 867563 70419 867619
rect 70475 867587 75816 867619
rect 70475 867563 73855 867587
rect 70000 867531 73855 867563
rect 73911 867531 73997 867587
rect 74053 867531 74139 867587
rect 74195 867531 74281 867587
rect 74337 867531 74423 867587
rect 74479 867531 74565 867587
rect 74621 867531 74707 867587
rect 74763 867531 74849 867587
rect 74905 867531 74991 867587
rect 75047 867531 75133 867587
rect 75189 867531 75275 867587
rect 75331 867531 75417 867587
rect 75473 867531 75559 867587
rect 75615 867531 75701 867587
rect 75757 867531 75816 867587
rect 70000 867495 75816 867531
rect 70000 867439 70047 867495
rect 70103 867439 70171 867495
rect 70227 867439 70295 867495
rect 70351 867439 70419 867495
rect 70475 867445 75816 867495
rect 70475 867439 73855 867445
rect 70000 867389 73855 867439
rect 73911 867389 73997 867445
rect 74053 867389 74139 867445
rect 74195 867389 74281 867445
rect 74337 867389 74423 867445
rect 74479 867389 74565 867445
rect 74621 867389 74707 867445
rect 74763 867389 74849 867445
rect 74905 867389 74991 867445
rect 75047 867389 75133 867445
rect 75189 867389 75275 867445
rect 75331 867389 75417 867445
rect 75473 867389 75559 867445
rect 75615 867389 75701 867445
rect 75757 867389 75816 867445
rect 70000 867371 75816 867389
rect 70000 867315 70047 867371
rect 70103 867315 70171 867371
rect 70227 867315 70295 867371
rect 70351 867315 70419 867371
rect 70475 867315 75816 867371
rect 70000 867303 75816 867315
rect 70000 867247 73855 867303
rect 73911 867247 73997 867303
rect 74053 867247 74139 867303
rect 74195 867247 74281 867303
rect 74337 867247 74423 867303
rect 74479 867247 74565 867303
rect 74621 867247 74707 867303
rect 74763 867247 74849 867303
rect 74905 867247 74991 867303
rect 75047 867247 75133 867303
rect 75189 867247 75275 867303
rect 75331 867247 75417 867303
rect 75473 867247 75559 867303
rect 75615 867247 75701 867303
rect 75757 867247 75816 867303
rect 70000 867191 70047 867247
rect 70103 867191 70171 867247
rect 70227 867191 70295 867247
rect 70351 867191 70419 867247
rect 70475 867191 75816 867247
rect 70000 867161 75816 867191
rect 70000 867123 73855 867161
rect 70000 867067 70047 867123
rect 70103 867067 70171 867123
rect 70227 867067 70295 867123
rect 70351 867067 70419 867123
rect 70475 867105 73855 867123
rect 73911 867105 73997 867161
rect 74053 867105 74139 867161
rect 74195 867105 74281 867161
rect 74337 867105 74423 867161
rect 74479 867105 74565 867161
rect 74621 867105 74707 867161
rect 74763 867105 74849 867161
rect 74905 867105 74991 867161
rect 75047 867105 75133 867161
rect 75189 867105 75275 867161
rect 75331 867105 75417 867161
rect 75473 867105 75559 867161
rect 75615 867105 75701 867161
rect 75757 867105 75816 867161
rect 70475 867067 75816 867105
rect 70000 867019 75816 867067
rect 70000 866999 73855 867019
rect 70000 866943 70047 866999
rect 70103 866943 70171 866999
rect 70227 866943 70295 866999
rect 70351 866943 70419 866999
rect 70475 866963 73855 866999
rect 73911 866963 73997 867019
rect 74053 866963 74139 867019
rect 74195 866963 74281 867019
rect 74337 866963 74423 867019
rect 74479 866963 74565 867019
rect 74621 866963 74707 867019
rect 74763 866963 74849 867019
rect 74905 866963 74991 867019
rect 75047 866963 75133 867019
rect 75189 866963 75275 867019
rect 75331 866963 75417 867019
rect 75473 866963 75559 867019
rect 75615 866963 75701 867019
rect 75757 866963 75816 867019
rect 70475 866943 75816 866963
rect 70000 866877 75816 866943
rect 70000 866875 73855 866877
rect 70000 866819 70047 866875
rect 70103 866819 70171 866875
rect 70227 866819 70295 866875
rect 70351 866819 70419 866875
rect 70475 866821 73855 866875
rect 73911 866821 73997 866877
rect 74053 866821 74139 866877
rect 74195 866821 74281 866877
rect 74337 866821 74423 866877
rect 74479 866821 74565 866877
rect 74621 866821 74707 866877
rect 74763 866821 74849 866877
rect 74905 866821 74991 866877
rect 75047 866821 75133 866877
rect 75189 866821 75275 866877
rect 75331 866821 75417 866877
rect 75473 866821 75559 866877
rect 75615 866821 75701 866877
rect 75757 866821 75816 866877
rect 70475 866819 75816 866821
rect 70000 866752 75816 866819
rect 699992 867735 706000 867802
rect 699992 867733 705525 867735
rect 699992 867677 700051 867733
rect 700107 867677 700193 867733
rect 700249 867677 700335 867733
rect 700391 867677 700477 867733
rect 700533 867677 700619 867733
rect 700675 867677 700761 867733
rect 700817 867677 700903 867733
rect 700959 867677 701045 867733
rect 701101 867677 701187 867733
rect 701243 867677 701329 867733
rect 701385 867677 701471 867733
rect 701527 867677 701613 867733
rect 701669 867677 701755 867733
rect 701811 867677 701897 867733
rect 701953 867679 705525 867733
rect 705581 867679 705649 867735
rect 705705 867679 705773 867735
rect 705829 867679 705897 867735
rect 705953 867679 706000 867735
rect 701953 867677 706000 867679
rect 699992 867611 706000 867677
rect 699992 867591 705525 867611
rect 699992 867535 700051 867591
rect 700107 867535 700193 867591
rect 700249 867535 700335 867591
rect 700391 867535 700477 867591
rect 700533 867535 700619 867591
rect 700675 867535 700761 867591
rect 700817 867535 700903 867591
rect 700959 867535 701045 867591
rect 701101 867535 701187 867591
rect 701243 867535 701329 867591
rect 701385 867535 701471 867591
rect 701527 867535 701613 867591
rect 701669 867535 701755 867591
rect 701811 867535 701897 867591
rect 701953 867555 705525 867591
rect 705581 867555 705649 867611
rect 705705 867555 705773 867611
rect 705829 867555 705897 867611
rect 705953 867555 706000 867611
rect 701953 867535 706000 867555
rect 699992 867487 706000 867535
rect 699992 867449 705525 867487
rect 699992 867393 700051 867449
rect 700107 867393 700193 867449
rect 700249 867393 700335 867449
rect 700391 867393 700477 867449
rect 700533 867393 700619 867449
rect 700675 867393 700761 867449
rect 700817 867393 700903 867449
rect 700959 867393 701045 867449
rect 701101 867393 701187 867449
rect 701243 867393 701329 867449
rect 701385 867393 701471 867449
rect 701527 867393 701613 867449
rect 701669 867393 701755 867449
rect 701811 867393 701897 867449
rect 701953 867431 705525 867449
rect 705581 867431 705649 867487
rect 705705 867431 705773 867487
rect 705829 867431 705897 867487
rect 705953 867431 706000 867487
rect 701953 867393 706000 867431
rect 699992 867363 706000 867393
rect 699992 867307 705525 867363
rect 705581 867307 705649 867363
rect 705705 867307 705773 867363
rect 705829 867307 705897 867363
rect 705953 867307 706000 867363
rect 699992 867251 700051 867307
rect 700107 867251 700193 867307
rect 700249 867251 700335 867307
rect 700391 867251 700477 867307
rect 700533 867251 700619 867307
rect 700675 867251 700761 867307
rect 700817 867251 700903 867307
rect 700959 867251 701045 867307
rect 701101 867251 701187 867307
rect 701243 867251 701329 867307
rect 701385 867251 701471 867307
rect 701527 867251 701613 867307
rect 701669 867251 701755 867307
rect 701811 867251 701897 867307
rect 701953 867251 706000 867307
rect 699992 867239 706000 867251
rect 699992 867183 705525 867239
rect 705581 867183 705649 867239
rect 705705 867183 705773 867239
rect 705829 867183 705897 867239
rect 705953 867183 706000 867239
rect 699992 867165 706000 867183
rect 699992 867109 700051 867165
rect 700107 867109 700193 867165
rect 700249 867109 700335 867165
rect 700391 867109 700477 867165
rect 700533 867109 700619 867165
rect 700675 867109 700761 867165
rect 700817 867109 700903 867165
rect 700959 867109 701045 867165
rect 701101 867109 701187 867165
rect 701243 867109 701329 867165
rect 701385 867109 701471 867165
rect 701527 867109 701613 867165
rect 701669 867109 701755 867165
rect 701811 867109 701897 867165
rect 701953 867115 706000 867165
rect 701953 867109 705525 867115
rect 699992 867059 705525 867109
rect 705581 867059 705649 867115
rect 705705 867059 705773 867115
rect 705829 867059 705897 867115
rect 705953 867059 706000 867115
rect 699992 867023 706000 867059
rect 699992 866967 700051 867023
rect 700107 866967 700193 867023
rect 700249 866967 700335 867023
rect 700391 866967 700477 867023
rect 700533 866967 700619 867023
rect 700675 866967 700761 867023
rect 700817 866967 700903 867023
rect 700959 866967 701045 867023
rect 701101 866967 701187 867023
rect 701243 866967 701329 867023
rect 701385 866967 701471 867023
rect 701527 866967 701613 867023
rect 701669 866967 701755 867023
rect 701811 866967 701897 867023
rect 701953 866991 706000 867023
rect 701953 866967 705525 866991
rect 699992 866935 705525 866967
rect 705581 866935 705649 866991
rect 705705 866935 705773 866991
rect 705829 866935 705897 866991
rect 705953 866935 706000 866991
rect 699992 866881 706000 866935
rect 699992 866825 700051 866881
rect 700107 866825 700193 866881
rect 700249 866825 700335 866881
rect 700391 866825 700477 866881
rect 700533 866825 700619 866881
rect 700675 866825 700761 866881
rect 700817 866825 700903 866881
rect 700959 866825 701045 866881
rect 701101 866825 701187 866881
rect 701243 866825 701329 866881
rect 701385 866825 701471 866881
rect 701527 866825 701613 866881
rect 701669 866825 701755 866881
rect 701811 866825 701897 866881
rect 701953 866867 706000 866881
rect 701953 866825 705525 866867
rect 699992 866811 705525 866825
rect 705581 866811 705649 866867
rect 705705 866811 705773 866867
rect 705829 866811 705897 866867
rect 705953 866811 706000 866867
rect 699992 866743 706000 866811
rect 699992 866739 705525 866743
rect 699992 866683 700051 866739
rect 700107 866683 700193 866739
rect 700249 866683 700335 866739
rect 700391 866683 700477 866739
rect 700533 866683 700619 866739
rect 700675 866683 700761 866739
rect 700817 866683 700903 866739
rect 700959 866683 701045 866739
rect 701101 866683 701187 866739
rect 701243 866683 701329 866739
rect 701385 866683 701471 866739
rect 701527 866683 701613 866739
rect 701669 866683 701755 866739
rect 701811 866683 701897 866739
rect 701953 866687 705525 866739
rect 705581 866687 705649 866743
rect 705705 866687 705773 866743
rect 705829 866687 705897 866743
rect 705953 866687 706000 866743
rect 701953 866683 706000 866687
rect 699992 866619 706000 866683
rect 699992 866597 705525 866619
rect 699992 866541 700051 866597
rect 700107 866541 700193 866597
rect 700249 866541 700335 866597
rect 700391 866541 700477 866597
rect 700533 866541 700619 866597
rect 700675 866541 700761 866597
rect 700817 866541 700903 866597
rect 700959 866541 701045 866597
rect 701101 866541 701187 866597
rect 701243 866541 701329 866597
rect 701385 866541 701471 866597
rect 701527 866541 701613 866597
rect 701669 866541 701755 866597
rect 701811 866541 701897 866597
rect 701953 866563 705525 866597
rect 705581 866563 705649 866619
rect 705705 866563 705773 866619
rect 705829 866563 705897 866619
rect 705953 866563 706000 866619
rect 701953 866541 706000 866563
rect 699992 866495 706000 866541
rect 699992 866455 705525 866495
rect 699992 866399 700051 866455
rect 700107 866399 700193 866455
rect 700249 866399 700335 866455
rect 700391 866399 700477 866455
rect 700533 866399 700619 866455
rect 700675 866399 700761 866455
rect 700817 866399 700903 866455
rect 700959 866399 701045 866455
rect 701101 866399 701187 866455
rect 701243 866399 701329 866455
rect 701385 866399 701471 866455
rect 701527 866399 701613 866455
rect 701669 866399 701755 866455
rect 701811 866399 701897 866455
rect 701953 866439 705525 866455
rect 705581 866439 705649 866495
rect 705705 866439 705773 866495
rect 705829 866439 705897 866495
rect 705953 866439 706000 866495
rect 701953 866399 706000 866439
rect 699992 866371 706000 866399
rect 699992 866315 705525 866371
rect 705581 866315 705649 866371
rect 705705 866315 705773 866371
rect 705829 866315 705897 866371
rect 705953 866315 706000 866371
rect 699992 866313 706000 866315
rect 699992 866257 700051 866313
rect 700107 866257 700193 866313
rect 700249 866257 700335 866313
rect 700391 866257 700477 866313
rect 700533 866257 700619 866313
rect 700675 866257 700761 866313
rect 700817 866257 700903 866313
rect 700959 866257 701045 866313
rect 701101 866257 701187 866313
rect 701243 866257 701329 866313
rect 701385 866257 701471 866313
rect 701527 866257 701613 866313
rect 701669 866257 701755 866313
rect 701811 866257 701897 866313
rect 701953 866257 706000 866313
rect 699992 866247 706000 866257
rect 699992 866191 705525 866247
rect 705581 866191 705649 866247
rect 705705 866191 705773 866247
rect 705829 866191 705897 866247
rect 705953 866191 706000 866247
rect 70000 866105 75816 866172
rect 70000 866049 70047 866105
rect 70103 866049 70171 866105
rect 70227 866049 70295 866105
rect 70351 866049 70419 866105
rect 70475 866094 75816 866105
rect 70475 866049 73866 866094
rect 70000 866038 73866 866049
rect 73922 866038 74008 866094
rect 74064 866038 74150 866094
rect 74206 866038 74292 866094
rect 74348 866038 74434 866094
rect 74490 866038 74576 866094
rect 74632 866038 74718 866094
rect 74774 866038 74860 866094
rect 74916 866038 75002 866094
rect 75058 866038 75144 866094
rect 75200 866038 75286 866094
rect 75342 866038 75428 866094
rect 75484 866038 75570 866094
rect 75626 866038 75712 866094
rect 75768 866038 75816 866094
rect 70000 865981 75816 866038
rect 70000 865925 70047 865981
rect 70103 865925 70171 865981
rect 70227 865925 70295 865981
rect 70351 865925 70419 865981
rect 70475 865952 75816 865981
rect 70475 865925 73866 865952
rect 70000 865896 73866 865925
rect 73922 865896 74008 865952
rect 74064 865896 74150 865952
rect 74206 865896 74292 865952
rect 74348 865896 74434 865952
rect 74490 865896 74576 865952
rect 74632 865896 74718 865952
rect 74774 865896 74860 865952
rect 74916 865896 75002 865952
rect 75058 865896 75144 865952
rect 75200 865896 75286 865952
rect 75342 865896 75428 865952
rect 75484 865896 75570 865952
rect 75626 865896 75712 865952
rect 75768 865896 75816 865952
rect 70000 865857 75816 865896
rect 70000 865801 70047 865857
rect 70103 865801 70171 865857
rect 70227 865801 70295 865857
rect 70351 865801 70419 865857
rect 70475 865810 75816 865857
rect 70475 865801 73866 865810
rect 70000 865754 73866 865801
rect 73922 865754 74008 865810
rect 74064 865754 74150 865810
rect 74206 865754 74292 865810
rect 74348 865754 74434 865810
rect 74490 865754 74576 865810
rect 74632 865754 74718 865810
rect 74774 865754 74860 865810
rect 74916 865754 75002 865810
rect 75058 865754 75144 865810
rect 75200 865754 75286 865810
rect 75342 865754 75428 865810
rect 75484 865754 75570 865810
rect 75626 865754 75712 865810
rect 75768 865754 75816 865810
rect 70000 865733 75816 865754
rect 699992 866171 706000 866191
rect 699992 866115 700051 866171
rect 700107 866115 700193 866171
rect 700249 866115 700335 866171
rect 700391 866115 700477 866171
rect 700533 866115 700619 866171
rect 700675 866115 700761 866171
rect 700817 866115 700903 866171
rect 700959 866115 701045 866171
rect 701101 866115 701187 866171
rect 701243 866115 701329 866171
rect 701385 866115 701471 866171
rect 701527 866115 701613 866171
rect 701669 866115 701755 866171
rect 701811 866115 701897 866171
rect 701953 866123 706000 866171
rect 701953 866115 705525 866123
rect 699992 866067 705525 866115
rect 705581 866067 705649 866123
rect 705705 866067 705773 866123
rect 705829 866067 705897 866123
rect 705953 866067 706000 866123
rect 699992 866029 706000 866067
rect 699992 865973 700051 866029
rect 700107 865973 700193 866029
rect 700249 865973 700335 866029
rect 700391 865973 700477 866029
rect 700533 865973 700619 866029
rect 700675 865973 700761 866029
rect 700817 865973 700903 866029
rect 700959 865973 701045 866029
rect 701101 865973 701187 866029
rect 701243 865973 701329 866029
rect 701385 865973 701471 866029
rect 701527 865973 701613 866029
rect 701669 865973 701755 866029
rect 701811 865973 701897 866029
rect 701953 865999 706000 866029
rect 701953 865973 705525 865999
rect 699992 865943 705525 865973
rect 705581 865943 705649 865999
rect 705705 865943 705773 865999
rect 705829 865943 705897 865999
rect 705953 865943 706000 865999
rect 699992 865887 706000 865943
rect 699992 865831 700051 865887
rect 700107 865831 700193 865887
rect 700249 865831 700335 865887
rect 700391 865831 700477 865887
rect 700533 865831 700619 865887
rect 700675 865831 700761 865887
rect 700817 865831 700903 865887
rect 700959 865831 701045 865887
rect 701101 865831 701187 865887
rect 701243 865831 701329 865887
rect 701385 865831 701471 865887
rect 701527 865831 701613 865887
rect 701669 865831 701755 865887
rect 701811 865831 701897 865887
rect 701953 865875 706000 865887
rect 701953 865831 705525 865875
rect 699992 865819 705525 865831
rect 705581 865819 705649 865875
rect 705705 865819 705773 865875
rect 705829 865819 705897 865875
rect 705953 865819 706000 865875
rect 699992 865752 706000 865819
rect 70000 865677 70047 865733
rect 70103 865677 70171 865733
rect 70227 865677 70295 865733
rect 70351 865677 70419 865733
rect 70475 865677 75816 865733
rect 70000 865668 75816 865677
rect 70000 865612 73866 865668
rect 73922 865612 74008 865668
rect 74064 865612 74150 865668
rect 74206 865612 74292 865668
rect 74348 865612 74434 865668
rect 74490 865612 74576 865668
rect 74632 865612 74718 865668
rect 74774 865612 74860 865668
rect 74916 865612 75002 865668
rect 75058 865612 75144 865668
rect 75200 865612 75286 865668
rect 75342 865612 75428 865668
rect 75484 865612 75570 865668
rect 75626 865612 75712 865668
rect 75768 865612 75816 865668
rect 70000 865609 75816 865612
rect 70000 865553 70047 865609
rect 70103 865553 70171 865609
rect 70227 865553 70295 865609
rect 70351 865553 70419 865609
rect 70475 865553 75816 865609
rect 70000 865526 75816 865553
rect 70000 865485 73866 865526
rect 70000 865429 70047 865485
rect 70103 865429 70171 865485
rect 70227 865429 70295 865485
rect 70351 865429 70419 865485
rect 70475 865470 73866 865485
rect 73922 865470 74008 865526
rect 74064 865470 74150 865526
rect 74206 865470 74292 865526
rect 74348 865470 74434 865526
rect 74490 865470 74576 865526
rect 74632 865470 74718 865526
rect 74774 865470 74860 865526
rect 74916 865470 75002 865526
rect 75058 865470 75144 865526
rect 75200 865470 75286 865526
rect 75342 865470 75428 865526
rect 75484 865470 75570 865526
rect 75626 865470 75712 865526
rect 75768 865470 75816 865526
rect 70475 865429 75816 865470
rect 70000 865384 75816 865429
rect 70000 865361 73866 865384
rect 70000 865305 70047 865361
rect 70103 865305 70171 865361
rect 70227 865305 70295 865361
rect 70351 865305 70419 865361
rect 70475 865328 73866 865361
rect 73922 865328 74008 865384
rect 74064 865328 74150 865384
rect 74206 865328 74292 865384
rect 74348 865328 74434 865384
rect 74490 865328 74576 865384
rect 74632 865328 74718 865384
rect 74774 865328 74860 865384
rect 74916 865328 75002 865384
rect 75058 865328 75144 865384
rect 75200 865328 75286 865384
rect 75342 865328 75428 865384
rect 75484 865328 75570 865384
rect 75626 865328 75712 865384
rect 75768 865328 75816 865384
rect 70475 865305 75816 865328
rect 70000 865242 75816 865305
rect 70000 865237 73866 865242
rect 70000 865181 70047 865237
rect 70103 865181 70171 865237
rect 70227 865181 70295 865237
rect 70351 865181 70419 865237
rect 70475 865186 73866 865237
rect 73922 865186 74008 865242
rect 74064 865186 74150 865242
rect 74206 865186 74292 865242
rect 74348 865186 74434 865242
rect 74490 865186 74576 865242
rect 74632 865186 74718 865242
rect 74774 865186 74860 865242
rect 74916 865186 75002 865242
rect 75058 865186 75144 865242
rect 75200 865186 75286 865242
rect 75342 865186 75428 865242
rect 75484 865186 75570 865242
rect 75626 865186 75712 865242
rect 75768 865186 75816 865242
rect 70475 865181 75816 865186
rect 70000 865113 75816 865181
rect 70000 865057 70047 865113
rect 70103 865057 70171 865113
rect 70227 865057 70295 865113
rect 70351 865057 70419 865113
rect 70475 865100 75816 865113
rect 70475 865057 73866 865100
rect 70000 865044 73866 865057
rect 73922 865044 74008 865100
rect 74064 865044 74150 865100
rect 74206 865044 74292 865100
rect 74348 865044 74434 865100
rect 74490 865044 74576 865100
rect 74632 865044 74718 865100
rect 74774 865044 74860 865100
rect 74916 865044 75002 865100
rect 75058 865044 75144 865100
rect 75200 865044 75286 865100
rect 75342 865044 75428 865100
rect 75484 865044 75570 865100
rect 75626 865044 75712 865100
rect 75768 865044 75816 865100
rect 70000 864989 75816 865044
rect 70000 864933 70047 864989
rect 70103 864933 70171 864989
rect 70227 864933 70295 864989
rect 70351 864933 70419 864989
rect 70475 864958 75816 864989
rect 70475 864933 73866 864958
rect 70000 864902 73866 864933
rect 73922 864902 74008 864958
rect 74064 864902 74150 864958
rect 74206 864902 74292 864958
rect 74348 864902 74434 864958
rect 74490 864902 74576 864958
rect 74632 864902 74718 864958
rect 74774 864902 74860 864958
rect 74916 864902 75002 864958
rect 75058 864902 75144 864958
rect 75200 864902 75286 864958
rect 75342 864902 75428 864958
rect 75484 864902 75570 864958
rect 75626 864902 75712 864958
rect 75768 864902 75816 864958
rect 70000 864865 75816 864902
rect 70000 864809 70047 864865
rect 70103 864809 70171 864865
rect 70227 864809 70295 864865
rect 70351 864809 70419 864865
rect 70475 864816 75816 864865
rect 70475 864809 73866 864816
rect 70000 864760 73866 864809
rect 73922 864760 74008 864816
rect 74064 864760 74150 864816
rect 74206 864760 74292 864816
rect 74348 864760 74434 864816
rect 74490 864760 74576 864816
rect 74632 864760 74718 864816
rect 74774 864760 74860 864816
rect 74916 864760 75002 864816
rect 75058 864760 75144 864816
rect 75200 864760 75286 864816
rect 75342 864760 75428 864816
rect 75484 864760 75570 864816
rect 75626 864760 75712 864816
rect 75768 864760 75816 864816
rect 70000 864741 75816 864760
rect 70000 864685 70047 864741
rect 70103 864685 70171 864741
rect 70227 864685 70295 864741
rect 70351 864685 70419 864741
rect 70475 864685 75816 864741
rect 70000 864674 75816 864685
rect 70000 864618 73866 864674
rect 73922 864618 74008 864674
rect 74064 864618 74150 864674
rect 74206 864618 74292 864674
rect 74348 864618 74434 864674
rect 74490 864618 74576 864674
rect 74632 864618 74718 864674
rect 74774 864618 74860 864674
rect 74916 864618 75002 864674
rect 75058 864618 75144 864674
rect 75200 864618 75286 864674
rect 75342 864618 75428 864674
rect 75484 864618 75570 864674
rect 75626 864618 75712 864674
rect 75768 864618 75816 864674
rect 70000 864617 75816 864618
rect 70000 864561 70047 864617
rect 70103 864561 70171 864617
rect 70227 864561 70295 864617
rect 70351 864561 70419 864617
rect 70475 864561 75816 864617
rect 70000 864532 75816 864561
rect 70000 864493 73866 864532
rect 70000 864437 70047 864493
rect 70103 864437 70171 864493
rect 70227 864437 70295 864493
rect 70351 864437 70419 864493
rect 70475 864476 73866 864493
rect 73922 864476 74008 864532
rect 74064 864476 74150 864532
rect 74206 864476 74292 864532
rect 74348 864476 74434 864532
rect 74490 864476 74576 864532
rect 74632 864476 74718 864532
rect 74774 864476 74860 864532
rect 74916 864476 75002 864532
rect 75058 864476 75144 864532
rect 75200 864476 75286 864532
rect 75342 864476 75428 864532
rect 75484 864476 75570 864532
rect 75626 864476 75712 864532
rect 75768 864476 75816 864532
rect 70475 864437 75816 864476
rect 70000 864390 75816 864437
rect 70000 864369 73866 864390
rect 70000 864313 70047 864369
rect 70103 864313 70171 864369
rect 70227 864313 70295 864369
rect 70351 864313 70419 864369
rect 70475 864334 73866 864369
rect 73922 864334 74008 864390
rect 74064 864334 74150 864390
rect 74206 864334 74292 864390
rect 74348 864334 74434 864390
rect 74490 864334 74576 864390
rect 74632 864334 74718 864390
rect 74774 864334 74860 864390
rect 74916 864334 75002 864390
rect 75058 864334 75144 864390
rect 75200 864334 75286 864390
rect 75342 864334 75428 864390
rect 75484 864334 75570 864390
rect 75626 864334 75712 864390
rect 75768 864334 75816 864390
rect 70475 864313 75816 864334
rect 70000 864272 75816 864313
rect 699992 865131 706000 865172
rect 699992 865110 705525 865131
rect 699992 865054 700040 865110
rect 700096 865054 700182 865110
rect 700238 865054 700324 865110
rect 700380 865054 700466 865110
rect 700522 865054 700608 865110
rect 700664 865054 700750 865110
rect 700806 865054 700892 865110
rect 700948 865054 701034 865110
rect 701090 865054 701176 865110
rect 701232 865054 701318 865110
rect 701374 865054 701460 865110
rect 701516 865054 701602 865110
rect 701658 865054 701744 865110
rect 701800 865054 701886 865110
rect 701942 865075 705525 865110
rect 705581 865075 705649 865131
rect 705705 865075 705773 865131
rect 705829 865075 705897 865131
rect 705953 865075 706000 865131
rect 701942 865054 706000 865075
rect 699992 865007 706000 865054
rect 699992 864968 705525 865007
rect 699992 864912 700040 864968
rect 700096 864912 700182 864968
rect 700238 864912 700324 864968
rect 700380 864912 700466 864968
rect 700522 864912 700608 864968
rect 700664 864912 700750 864968
rect 700806 864912 700892 864968
rect 700948 864912 701034 864968
rect 701090 864912 701176 864968
rect 701232 864912 701318 864968
rect 701374 864912 701460 864968
rect 701516 864912 701602 864968
rect 701658 864912 701744 864968
rect 701800 864912 701886 864968
rect 701942 864951 705525 864968
rect 705581 864951 705649 865007
rect 705705 864951 705773 865007
rect 705829 864951 705897 865007
rect 705953 864951 706000 865007
rect 701942 864912 706000 864951
rect 699992 864883 706000 864912
rect 699992 864827 705525 864883
rect 705581 864827 705649 864883
rect 705705 864827 705773 864883
rect 705829 864827 705897 864883
rect 705953 864827 706000 864883
rect 699992 864826 706000 864827
rect 699992 864770 700040 864826
rect 700096 864770 700182 864826
rect 700238 864770 700324 864826
rect 700380 864770 700466 864826
rect 700522 864770 700608 864826
rect 700664 864770 700750 864826
rect 700806 864770 700892 864826
rect 700948 864770 701034 864826
rect 701090 864770 701176 864826
rect 701232 864770 701318 864826
rect 701374 864770 701460 864826
rect 701516 864770 701602 864826
rect 701658 864770 701744 864826
rect 701800 864770 701886 864826
rect 701942 864770 706000 864826
rect 699992 864759 706000 864770
rect 699992 864703 705525 864759
rect 705581 864703 705649 864759
rect 705705 864703 705773 864759
rect 705829 864703 705897 864759
rect 705953 864703 706000 864759
rect 699992 864684 706000 864703
rect 699992 864628 700040 864684
rect 700096 864628 700182 864684
rect 700238 864628 700324 864684
rect 700380 864628 700466 864684
rect 700522 864628 700608 864684
rect 700664 864628 700750 864684
rect 700806 864628 700892 864684
rect 700948 864628 701034 864684
rect 701090 864628 701176 864684
rect 701232 864628 701318 864684
rect 701374 864628 701460 864684
rect 701516 864628 701602 864684
rect 701658 864628 701744 864684
rect 701800 864628 701886 864684
rect 701942 864635 706000 864684
rect 701942 864628 705525 864635
rect 699992 864579 705525 864628
rect 705581 864579 705649 864635
rect 705705 864579 705773 864635
rect 705829 864579 705897 864635
rect 705953 864579 706000 864635
rect 699992 864542 706000 864579
rect 699992 864486 700040 864542
rect 700096 864486 700182 864542
rect 700238 864486 700324 864542
rect 700380 864486 700466 864542
rect 700522 864486 700608 864542
rect 700664 864486 700750 864542
rect 700806 864486 700892 864542
rect 700948 864486 701034 864542
rect 701090 864486 701176 864542
rect 701232 864486 701318 864542
rect 701374 864486 701460 864542
rect 701516 864486 701602 864542
rect 701658 864486 701744 864542
rect 701800 864486 701886 864542
rect 701942 864511 706000 864542
rect 701942 864486 705525 864511
rect 699992 864455 705525 864486
rect 705581 864455 705649 864511
rect 705705 864455 705773 864511
rect 705829 864455 705897 864511
rect 705953 864455 706000 864511
rect 699992 864400 706000 864455
rect 699992 864344 700040 864400
rect 700096 864344 700182 864400
rect 700238 864344 700324 864400
rect 700380 864344 700466 864400
rect 700522 864344 700608 864400
rect 700664 864344 700750 864400
rect 700806 864344 700892 864400
rect 700948 864344 701034 864400
rect 701090 864344 701176 864400
rect 701232 864344 701318 864400
rect 701374 864344 701460 864400
rect 701516 864344 701602 864400
rect 701658 864344 701744 864400
rect 701800 864344 701886 864400
rect 701942 864387 706000 864400
rect 701942 864344 705525 864387
rect 699992 864331 705525 864344
rect 705581 864331 705649 864387
rect 705705 864331 705773 864387
rect 705829 864331 705897 864387
rect 705953 864331 706000 864387
rect 699992 864263 706000 864331
rect 699992 864258 705525 864263
rect 699992 864202 700040 864258
rect 700096 864202 700182 864258
rect 700238 864202 700324 864258
rect 700380 864202 700466 864258
rect 700522 864202 700608 864258
rect 700664 864202 700750 864258
rect 700806 864202 700892 864258
rect 700948 864202 701034 864258
rect 701090 864202 701176 864258
rect 701232 864202 701318 864258
rect 701374 864202 701460 864258
rect 701516 864202 701602 864258
rect 701658 864202 701744 864258
rect 701800 864202 701886 864258
rect 701942 864207 705525 864258
rect 705581 864207 705649 864263
rect 705705 864207 705773 864263
rect 705829 864207 705897 864263
rect 705953 864207 706000 864263
rect 701942 864202 706000 864207
rect 699992 864139 706000 864202
rect 699992 864116 705525 864139
rect 699992 864060 700040 864116
rect 700096 864060 700182 864116
rect 700238 864060 700324 864116
rect 700380 864060 700466 864116
rect 700522 864060 700608 864116
rect 700664 864060 700750 864116
rect 700806 864060 700892 864116
rect 700948 864060 701034 864116
rect 701090 864060 701176 864116
rect 701232 864060 701318 864116
rect 701374 864060 701460 864116
rect 701516 864060 701602 864116
rect 701658 864060 701744 864116
rect 701800 864060 701886 864116
rect 701942 864083 705525 864116
rect 705581 864083 705649 864139
rect 705705 864083 705773 864139
rect 705829 864083 705897 864139
rect 705953 864083 706000 864139
rect 701942 864060 706000 864083
rect 699992 864015 706000 864060
rect 699992 863974 705525 864015
rect 699992 863918 700040 863974
rect 700096 863918 700182 863974
rect 700238 863918 700324 863974
rect 700380 863918 700466 863974
rect 700522 863918 700608 863974
rect 700664 863918 700750 863974
rect 700806 863918 700892 863974
rect 700948 863918 701034 863974
rect 701090 863918 701176 863974
rect 701232 863918 701318 863974
rect 701374 863918 701460 863974
rect 701516 863918 701602 863974
rect 701658 863918 701744 863974
rect 701800 863918 701886 863974
rect 701942 863959 705525 863974
rect 705581 863959 705649 864015
rect 705705 863959 705773 864015
rect 705829 863959 705897 864015
rect 705953 863959 706000 864015
rect 701942 863918 706000 863959
rect 699992 863891 706000 863918
rect 699992 863835 705525 863891
rect 705581 863835 705649 863891
rect 705705 863835 705773 863891
rect 705829 863835 705897 863891
rect 705953 863835 706000 863891
rect 699992 863832 706000 863835
rect 699992 863776 700040 863832
rect 700096 863776 700182 863832
rect 700238 863776 700324 863832
rect 700380 863776 700466 863832
rect 700522 863776 700608 863832
rect 700664 863776 700750 863832
rect 700806 863776 700892 863832
rect 700948 863776 701034 863832
rect 701090 863776 701176 863832
rect 701232 863776 701318 863832
rect 701374 863776 701460 863832
rect 701516 863776 701602 863832
rect 701658 863776 701744 863832
rect 701800 863776 701886 863832
rect 701942 863776 706000 863832
rect 699992 863767 706000 863776
rect 699992 863711 705525 863767
rect 705581 863711 705649 863767
rect 705705 863711 705773 863767
rect 705829 863711 705897 863767
rect 705953 863711 706000 863767
rect 699992 863690 706000 863711
rect 699992 863634 700040 863690
rect 700096 863634 700182 863690
rect 700238 863634 700324 863690
rect 700380 863634 700466 863690
rect 700522 863634 700608 863690
rect 700664 863634 700750 863690
rect 700806 863634 700892 863690
rect 700948 863634 701034 863690
rect 701090 863634 701176 863690
rect 701232 863634 701318 863690
rect 701374 863634 701460 863690
rect 701516 863634 701602 863690
rect 701658 863634 701744 863690
rect 701800 863634 701886 863690
rect 701942 863643 706000 863690
rect 701942 863634 705525 863643
rect 699992 863587 705525 863634
rect 705581 863587 705649 863643
rect 705705 863587 705773 863643
rect 705829 863587 705897 863643
rect 705953 863587 706000 863643
rect 699992 863548 706000 863587
rect 699992 863492 700040 863548
rect 700096 863492 700182 863548
rect 700238 863492 700324 863548
rect 700380 863492 700466 863548
rect 700522 863492 700608 863548
rect 700664 863492 700750 863548
rect 700806 863492 700892 863548
rect 700948 863492 701034 863548
rect 701090 863492 701176 863548
rect 701232 863492 701318 863548
rect 701374 863492 701460 863548
rect 701516 863492 701602 863548
rect 701658 863492 701744 863548
rect 701800 863492 701886 863548
rect 701942 863519 706000 863548
rect 701942 863492 705525 863519
rect 699992 863463 705525 863492
rect 705581 863463 705649 863519
rect 705705 863463 705773 863519
rect 705829 863463 705897 863519
rect 705953 863463 706000 863519
rect 699992 863406 706000 863463
rect 699992 863350 700040 863406
rect 700096 863350 700182 863406
rect 700238 863350 700324 863406
rect 700380 863350 700466 863406
rect 700522 863350 700608 863406
rect 700664 863350 700750 863406
rect 700806 863350 700892 863406
rect 700948 863350 701034 863406
rect 701090 863350 701176 863406
rect 701232 863350 701318 863406
rect 701374 863350 701460 863406
rect 701516 863350 701602 863406
rect 701658 863350 701744 863406
rect 701800 863350 701886 863406
rect 701942 863395 706000 863406
rect 701942 863350 705525 863395
rect 699992 863339 705525 863350
rect 705581 863339 705649 863395
rect 705705 863339 705773 863395
rect 705829 863339 705897 863395
rect 705953 863339 706000 863395
rect 699992 863272 706000 863339
rect 70000 837661 75416 837728
rect 70000 837605 70047 837661
rect 70103 837605 70171 837661
rect 70227 837605 70295 837661
rect 70351 837605 70419 837661
rect 70475 837650 75416 837661
rect 70475 837605 73866 837650
rect 70000 837594 73866 837605
rect 73922 837594 74008 837650
rect 74064 837594 74150 837650
rect 74206 837594 74292 837650
rect 74348 837594 74434 837650
rect 74490 837594 74576 837650
rect 74632 837594 74718 837650
rect 74774 837594 74860 837650
rect 74916 837594 75002 837650
rect 75058 837594 75144 837650
rect 75200 837594 75286 837650
rect 75342 837594 75416 837650
rect 70000 837537 75416 837594
rect 70000 837481 70047 837537
rect 70103 837481 70171 837537
rect 70227 837481 70295 837537
rect 70351 837481 70419 837537
rect 70475 837508 75416 837537
rect 70475 837481 73866 837508
rect 70000 837452 73866 837481
rect 73922 837452 74008 837508
rect 74064 837452 74150 837508
rect 74206 837452 74292 837508
rect 74348 837452 74434 837508
rect 74490 837452 74576 837508
rect 74632 837452 74718 837508
rect 74774 837452 74860 837508
rect 74916 837452 75002 837508
rect 75058 837452 75144 837508
rect 75200 837452 75286 837508
rect 75342 837452 75416 837508
rect 70000 837413 75416 837452
rect 70000 837357 70047 837413
rect 70103 837357 70171 837413
rect 70227 837357 70295 837413
rect 70351 837357 70419 837413
rect 70475 837366 75416 837413
rect 70475 837357 73866 837366
rect 70000 837310 73866 837357
rect 73922 837310 74008 837366
rect 74064 837310 74150 837366
rect 74206 837310 74292 837366
rect 74348 837310 74434 837366
rect 74490 837310 74576 837366
rect 74632 837310 74718 837366
rect 74774 837310 74860 837366
rect 74916 837310 75002 837366
rect 75058 837310 75144 837366
rect 75200 837310 75286 837366
rect 75342 837310 75416 837366
rect 70000 837289 75416 837310
rect 70000 837233 70047 837289
rect 70103 837233 70171 837289
rect 70227 837233 70295 837289
rect 70351 837233 70419 837289
rect 70475 837233 75416 837289
rect 70000 837224 75416 837233
rect 70000 837168 73866 837224
rect 73922 837168 74008 837224
rect 74064 837168 74150 837224
rect 74206 837168 74292 837224
rect 74348 837168 74434 837224
rect 74490 837168 74576 837224
rect 74632 837168 74718 837224
rect 74774 837168 74860 837224
rect 74916 837168 75002 837224
rect 75058 837168 75144 837224
rect 75200 837168 75286 837224
rect 75342 837168 75416 837224
rect 70000 837165 75416 837168
rect 70000 837109 70047 837165
rect 70103 837109 70171 837165
rect 70227 837109 70295 837165
rect 70351 837109 70419 837165
rect 70475 837109 75416 837165
rect 70000 837082 75416 837109
rect 70000 837041 73866 837082
rect 70000 836985 70047 837041
rect 70103 836985 70171 837041
rect 70227 836985 70295 837041
rect 70351 836985 70419 837041
rect 70475 837026 73866 837041
rect 73922 837026 74008 837082
rect 74064 837026 74150 837082
rect 74206 837026 74292 837082
rect 74348 837026 74434 837082
rect 74490 837026 74576 837082
rect 74632 837026 74718 837082
rect 74774 837026 74860 837082
rect 74916 837026 75002 837082
rect 75058 837026 75144 837082
rect 75200 837026 75286 837082
rect 75342 837026 75416 837082
rect 70475 836985 75416 837026
rect 70000 836940 75416 836985
rect 70000 836917 73866 836940
rect 70000 836861 70047 836917
rect 70103 836861 70171 836917
rect 70227 836861 70295 836917
rect 70351 836861 70419 836917
rect 70475 836884 73866 836917
rect 73922 836884 74008 836940
rect 74064 836884 74150 836940
rect 74206 836884 74292 836940
rect 74348 836884 74434 836940
rect 74490 836884 74576 836940
rect 74632 836884 74718 836940
rect 74774 836884 74860 836940
rect 74916 836884 75002 836940
rect 75058 836884 75144 836940
rect 75200 836884 75286 836940
rect 75342 836884 75416 836940
rect 70475 836861 75416 836884
rect 70000 836798 75416 836861
rect 70000 836793 73866 836798
rect 70000 836737 70047 836793
rect 70103 836737 70171 836793
rect 70227 836737 70295 836793
rect 70351 836737 70419 836793
rect 70475 836742 73866 836793
rect 73922 836742 74008 836798
rect 74064 836742 74150 836798
rect 74206 836742 74292 836798
rect 74348 836742 74434 836798
rect 74490 836742 74576 836798
rect 74632 836742 74718 836798
rect 74774 836742 74860 836798
rect 74916 836742 75002 836798
rect 75058 836742 75144 836798
rect 75200 836742 75286 836798
rect 75342 836742 75416 836798
rect 70475 836737 75416 836742
rect 70000 836669 75416 836737
rect 70000 836613 70047 836669
rect 70103 836613 70171 836669
rect 70227 836613 70295 836669
rect 70351 836613 70419 836669
rect 70475 836656 75416 836669
rect 70475 836613 73866 836656
rect 70000 836600 73866 836613
rect 73922 836600 74008 836656
rect 74064 836600 74150 836656
rect 74206 836600 74292 836656
rect 74348 836600 74434 836656
rect 74490 836600 74576 836656
rect 74632 836600 74718 836656
rect 74774 836600 74860 836656
rect 74916 836600 75002 836656
rect 75058 836600 75144 836656
rect 75200 836600 75286 836656
rect 75342 836600 75416 836656
rect 70000 836545 75416 836600
rect 70000 836489 70047 836545
rect 70103 836489 70171 836545
rect 70227 836489 70295 836545
rect 70351 836489 70419 836545
rect 70475 836514 75416 836545
rect 70475 836489 73866 836514
rect 70000 836458 73866 836489
rect 73922 836458 74008 836514
rect 74064 836458 74150 836514
rect 74206 836458 74292 836514
rect 74348 836458 74434 836514
rect 74490 836458 74576 836514
rect 74632 836458 74718 836514
rect 74774 836458 74860 836514
rect 74916 836458 75002 836514
rect 75058 836458 75144 836514
rect 75200 836458 75286 836514
rect 75342 836458 75416 836514
rect 70000 836421 75416 836458
rect 70000 836365 70047 836421
rect 70103 836365 70171 836421
rect 70227 836365 70295 836421
rect 70351 836365 70419 836421
rect 70475 836372 75416 836421
rect 70475 836365 73866 836372
rect 70000 836316 73866 836365
rect 73922 836316 74008 836372
rect 74064 836316 74150 836372
rect 74206 836316 74292 836372
rect 74348 836316 74434 836372
rect 74490 836316 74576 836372
rect 74632 836316 74718 836372
rect 74774 836316 74860 836372
rect 74916 836316 75002 836372
rect 75058 836316 75144 836372
rect 75200 836316 75286 836372
rect 75342 836316 75416 836372
rect 70000 836297 75416 836316
rect 70000 836241 70047 836297
rect 70103 836241 70171 836297
rect 70227 836241 70295 836297
rect 70351 836241 70419 836297
rect 70475 836241 75416 836297
rect 70000 836230 75416 836241
rect 70000 836174 73866 836230
rect 73922 836174 74008 836230
rect 74064 836174 74150 836230
rect 74206 836174 74292 836230
rect 74348 836174 74434 836230
rect 74490 836174 74576 836230
rect 74632 836174 74718 836230
rect 74774 836174 74860 836230
rect 74916 836174 75002 836230
rect 75058 836174 75144 836230
rect 75200 836174 75286 836230
rect 75342 836174 75416 836230
rect 70000 836173 75416 836174
rect 70000 836117 70047 836173
rect 70103 836117 70171 836173
rect 70227 836117 70295 836173
rect 70351 836117 70419 836173
rect 70475 836117 75416 836173
rect 70000 836088 75416 836117
rect 70000 836049 73866 836088
rect 70000 835993 70047 836049
rect 70103 835993 70171 836049
rect 70227 835993 70295 836049
rect 70351 835993 70419 836049
rect 70475 836032 73866 836049
rect 73922 836032 74008 836088
rect 74064 836032 74150 836088
rect 74206 836032 74292 836088
rect 74348 836032 74434 836088
rect 74490 836032 74576 836088
rect 74632 836032 74718 836088
rect 74774 836032 74860 836088
rect 74916 836032 75002 836088
rect 75058 836032 75144 836088
rect 75200 836032 75286 836088
rect 75342 836032 75416 836088
rect 70475 835993 75416 836032
rect 70000 835946 75416 835993
rect 70000 835925 73866 835946
rect 70000 835869 70047 835925
rect 70103 835869 70171 835925
rect 70227 835869 70295 835925
rect 70351 835869 70419 835925
rect 70475 835890 73866 835925
rect 73922 835890 74008 835946
rect 74064 835890 74150 835946
rect 74206 835890 74292 835946
rect 74348 835890 74434 835946
rect 74490 835890 74576 835946
rect 74632 835890 74718 835946
rect 74774 835890 74860 835946
rect 74916 835890 75002 835946
rect 75058 835890 75144 835946
rect 75200 835890 75286 835946
rect 75342 835890 75416 835946
rect 70475 835869 75416 835890
rect 70000 835828 75416 835869
rect 70000 835181 75416 835248
rect 70000 835125 70047 835181
rect 70103 835125 70171 835181
rect 70227 835125 70295 835181
rect 70351 835125 70419 835181
rect 70475 835169 75416 835181
rect 70475 835125 73855 835169
rect 70000 835113 73855 835125
rect 73911 835113 73997 835169
rect 74053 835113 74139 835169
rect 74195 835113 74281 835169
rect 74337 835113 74423 835169
rect 74479 835113 74565 835169
rect 74621 835113 74707 835169
rect 74763 835113 74849 835169
rect 74905 835113 74991 835169
rect 75047 835113 75133 835169
rect 75189 835113 75275 835169
rect 75331 835113 75416 835169
rect 70000 835057 75416 835113
rect 70000 835001 70047 835057
rect 70103 835001 70171 835057
rect 70227 835001 70295 835057
rect 70351 835001 70419 835057
rect 70475 835027 75416 835057
rect 70475 835001 73855 835027
rect 70000 834971 73855 835001
rect 73911 834971 73997 835027
rect 74053 834971 74139 835027
rect 74195 834971 74281 835027
rect 74337 834971 74423 835027
rect 74479 834971 74565 835027
rect 74621 834971 74707 835027
rect 74763 834971 74849 835027
rect 74905 834971 74991 835027
rect 75047 834971 75133 835027
rect 75189 834971 75275 835027
rect 75331 834971 75416 835027
rect 70000 834933 75416 834971
rect 70000 834877 70047 834933
rect 70103 834877 70171 834933
rect 70227 834877 70295 834933
rect 70351 834877 70419 834933
rect 70475 834885 75416 834933
rect 70475 834877 73855 834885
rect 70000 834829 73855 834877
rect 73911 834829 73997 834885
rect 74053 834829 74139 834885
rect 74195 834829 74281 834885
rect 74337 834829 74423 834885
rect 74479 834829 74565 834885
rect 74621 834829 74707 834885
rect 74763 834829 74849 834885
rect 74905 834829 74991 834885
rect 75047 834829 75133 834885
rect 75189 834829 75275 834885
rect 75331 834829 75416 834885
rect 70000 834809 75416 834829
rect 70000 834753 70047 834809
rect 70103 834753 70171 834809
rect 70227 834753 70295 834809
rect 70351 834753 70419 834809
rect 70475 834753 75416 834809
rect 70000 834743 75416 834753
rect 70000 834687 73855 834743
rect 73911 834687 73997 834743
rect 74053 834687 74139 834743
rect 74195 834687 74281 834743
rect 74337 834687 74423 834743
rect 74479 834687 74565 834743
rect 74621 834687 74707 834743
rect 74763 834687 74849 834743
rect 74905 834687 74991 834743
rect 75047 834687 75133 834743
rect 75189 834687 75275 834743
rect 75331 834687 75416 834743
rect 70000 834685 75416 834687
rect 70000 834629 70047 834685
rect 70103 834629 70171 834685
rect 70227 834629 70295 834685
rect 70351 834629 70419 834685
rect 70475 834629 75416 834685
rect 70000 834601 75416 834629
rect 70000 834561 73855 834601
rect 70000 834505 70047 834561
rect 70103 834505 70171 834561
rect 70227 834505 70295 834561
rect 70351 834505 70419 834561
rect 70475 834545 73855 834561
rect 73911 834545 73997 834601
rect 74053 834545 74139 834601
rect 74195 834545 74281 834601
rect 74337 834545 74423 834601
rect 74479 834545 74565 834601
rect 74621 834545 74707 834601
rect 74763 834545 74849 834601
rect 74905 834545 74991 834601
rect 75047 834545 75133 834601
rect 75189 834545 75275 834601
rect 75331 834545 75416 834601
rect 70475 834505 75416 834545
rect 70000 834459 75416 834505
rect 70000 834437 73855 834459
rect 70000 834381 70047 834437
rect 70103 834381 70171 834437
rect 70227 834381 70295 834437
rect 70351 834381 70419 834437
rect 70475 834403 73855 834437
rect 73911 834403 73997 834459
rect 74053 834403 74139 834459
rect 74195 834403 74281 834459
rect 74337 834403 74423 834459
rect 74479 834403 74565 834459
rect 74621 834403 74707 834459
rect 74763 834403 74849 834459
rect 74905 834403 74991 834459
rect 75047 834403 75133 834459
rect 75189 834403 75275 834459
rect 75331 834403 75416 834459
rect 70475 834381 75416 834403
rect 70000 834317 75416 834381
rect 70000 834313 73855 834317
rect 70000 834257 70047 834313
rect 70103 834257 70171 834313
rect 70227 834257 70295 834313
rect 70351 834257 70419 834313
rect 70475 834261 73855 834313
rect 73911 834261 73997 834317
rect 74053 834261 74139 834317
rect 74195 834261 74281 834317
rect 74337 834261 74423 834317
rect 74479 834261 74565 834317
rect 74621 834261 74707 834317
rect 74763 834261 74849 834317
rect 74905 834261 74991 834317
rect 75047 834261 75133 834317
rect 75189 834261 75275 834317
rect 75331 834261 75416 834317
rect 70475 834257 75416 834261
rect 70000 834189 75416 834257
rect 70000 834133 70047 834189
rect 70103 834133 70171 834189
rect 70227 834133 70295 834189
rect 70351 834133 70419 834189
rect 70475 834175 75416 834189
rect 70475 834133 73855 834175
rect 70000 834119 73855 834133
rect 73911 834119 73997 834175
rect 74053 834119 74139 834175
rect 74195 834119 74281 834175
rect 74337 834119 74423 834175
rect 74479 834119 74565 834175
rect 74621 834119 74707 834175
rect 74763 834119 74849 834175
rect 74905 834119 74991 834175
rect 75047 834119 75133 834175
rect 75189 834119 75275 834175
rect 75331 834119 75416 834175
rect 70000 834065 75416 834119
rect 70000 834009 70047 834065
rect 70103 834009 70171 834065
rect 70227 834009 70295 834065
rect 70351 834009 70419 834065
rect 70475 834033 75416 834065
rect 70475 834009 73855 834033
rect 70000 833977 73855 834009
rect 73911 833977 73997 834033
rect 74053 833977 74139 834033
rect 74195 833977 74281 834033
rect 74337 833977 74423 834033
rect 74479 833977 74565 834033
rect 74621 833977 74707 834033
rect 74763 833977 74849 834033
rect 74905 833977 74991 834033
rect 75047 833977 75133 834033
rect 75189 833977 75275 834033
rect 75331 833977 75416 834033
rect 70000 833941 75416 833977
rect 70000 833885 70047 833941
rect 70103 833885 70171 833941
rect 70227 833885 70295 833941
rect 70351 833885 70419 833941
rect 70475 833891 75416 833941
rect 70475 833885 73855 833891
rect 70000 833835 73855 833885
rect 73911 833835 73997 833891
rect 74053 833835 74139 833891
rect 74195 833835 74281 833891
rect 74337 833835 74423 833891
rect 74479 833835 74565 833891
rect 74621 833835 74707 833891
rect 74763 833835 74849 833891
rect 74905 833835 74991 833891
rect 75047 833835 75133 833891
rect 75189 833835 75275 833891
rect 75331 833835 75416 833891
rect 70000 833817 75416 833835
rect 70000 833761 70047 833817
rect 70103 833761 70171 833817
rect 70227 833761 70295 833817
rect 70351 833761 70419 833817
rect 70475 833761 75416 833817
rect 70000 833749 75416 833761
rect 70000 833693 73855 833749
rect 73911 833693 73997 833749
rect 74053 833693 74139 833749
rect 74195 833693 74281 833749
rect 74337 833693 74423 833749
rect 74479 833693 74565 833749
rect 74621 833693 74707 833749
rect 74763 833693 74849 833749
rect 74905 833693 74991 833749
rect 75047 833693 75133 833749
rect 75189 833693 75275 833749
rect 75331 833693 75416 833749
rect 70000 833637 70047 833693
rect 70103 833637 70171 833693
rect 70227 833637 70295 833693
rect 70351 833637 70419 833693
rect 70475 833637 75416 833693
rect 70000 833607 75416 833637
rect 70000 833569 73855 833607
rect 70000 833513 70047 833569
rect 70103 833513 70171 833569
rect 70227 833513 70295 833569
rect 70351 833513 70419 833569
rect 70475 833551 73855 833569
rect 73911 833551 73997 833607
rect 74053 833551 74139 833607
rect 74195 833551 74281 833607
rect 74337 833551 74423 833607
rect 74479 833551 74565 833607
rect 74621 833551 74707 833607
rect 74763 833551 74849 833607
rect 74905 833551 74991 833607
rect 75047 833551 75133 833607
rect 75189 833551 75275 833607
rect 75331 833551 75416 833607
rect 70475 833513 75416 833551
rect 70000 833465 75416 833513
rect 70000 833445 73855 833465
rect 70000 833389 70047 833445
rect 70103 833389 70171 833445
rect 70227 833389 70295 833445
rect 70351 833389 70419 833445
rect 70475 833409 73855 833445
rect 73911 833409 73997 833465
rect 74053 833409 74139 833465
rect 74195 833409 74281 833465
rect 74337 833409 74423 833465
rect 74479 833409 74565 833465
rect 74621 833409 74707 833465
rect 74763 833409 74849 833465
rect 74905 833409 74991 833465
rect 75047 833409 75133 833465
rect 75189 833409 75275 833465
rect 75331 833409 75416 833465
rect 70475 833389 75416 833409
rect 70000 833323 75416 833389
rect 70000 833321 73855 833323
rect 70000 833265 70047 833321
rect 70103 833265 70171 833321
rect 70227 833265 70295 833321
rect 70351 833265 70419 833321
rect 70475 833267 73855 833321
rect 73911 833267 73997 833323
rect 74053 833267 74139 833323
rect 74195 833267 74281 833323
rect 74337 833267 74423 833323
rect 74479 833267 74565 833323
rect 74621 833267 74707 833323
rect 74763 833267 74849 833323
rect 74905 833267 74991 833323
rect 75047 833267 75133 833323
rect 75189 833267 75275 833323
rect 75331 833267 75416 833323
rect 70475 833265 75416 833267
rect 70000 833198 75416 833265
rect 70000 832811 75416 832878
rect 70000 832755 70047 832811
rect 70103 832755 70171 832811
rect 70227 832755 70295 832811
rect 70351 832755 70419 832811
rect 70475 832799 75416 832811
rect 70475 832755 73855 832799
rect 70000 832743 73855 832755
rect 73911 832743 73997 832799
rect 74053 832743 74139 832799
rect 74195 832743 74281 832799
rect 74337 832743 74423 832799
rect 74479 832743 74565 832799
rect 74621 832743 74707 832799
rect 74763 832743 74849 832799
rect 74905 832743 74991 832799
rect 75047 832743 75133 832799
rect 75189 832743 75275 832799
rect 75331 832743 75416 832799
rect 70000 832687 75416 832743
rect 70000 832631 70047 832687
rect 70103 832631 70171 832687
rect 70227 832631 70295 832687
rect 70351 832631 70419 832687
rect 70475 832657 75416 832687
rect 70475 832631 73855 832657
rect 70000 832601 73855 832631
rect 73911 832601 73997 832657
rect 74053 832601 74139 832657
rect 74195 832601 74281 832657
rect 74337 832601 74423 832657
rect 74479 832601 74565 832657
rect 74621 832601 74707 832657
rect 74763 832601 74849 832657
rect 74905 832601 74991 832657
rect 75047 832601 75133 832657
rect 75189 832601 75275 832657
rect 75331 832601 75416 832657
rect 70000 832563 75416 832601
rect 70000 832507 70047 832563
rect 70103 832507 70171 832563
rect 70227 832507 70295 832563
rect 70351 832507 70419 832563
rect 70475 832515 75416 832563
rect 70475 832507 73855 832515
rect 70000 832459 73855 832507
rect 73911 832459 73997 832515
rect 74053 832459 74139 832515
rect 74195 832459 74281 832515
rect 74337 832459 74423 832515
rect 74479 832459 74565 832515
rect 74621 832459 74707 832515
rect 74763 832459 74849 832515
rect 74905 832459 74991 832515
rect 75047 832459 75133 832515
rect 75189 832459 75275 832515
rect 75331 832459 75416 832515
rect 70000 832439 75416 832459
rect 70000 832383 70047 832439
rect 70103 832383 70171 832439
rect 70227 832383 70295 832439
rect 70351 832383 70419 832439
rect 70475 832383 75416 832439
rect 70000 832373 75416 832383
rect 70000 832317 73855 832373
rect 73911 832317 73997 832373
rect 74053 832317 74139 832373
rect 74195 832317 74281 832373
rect 74337 832317 74423 832373
rect 74479 832317 74565 832373
rect 74621 832317 74707 832373
rect 74763 832317 74849 832373
rect 74905 832317 74991 832373
rect 75047 832317 75133 832373
rect 75189 832317 75275 832373
rect 75331 832317 75416 832373
rect 70000 832315 75416 832317
rect 70000 832259 70047 832315
rect 70103 832259 70171 832315
rect 70227 832259 70295 832315
rect 70351 832259 70419 832315
rect 70475 832259 75416 832315
rect 70000 832231 75416 832259
rect 70000 832191 73855 832231
rect 70000 832135 70047 832191
rect 70103 832135 70171 832191
rect 70227 832135 70295 832191
rect 70351 832135 70419 832191
rect 70475 832175 73855 832191
rect 73911 832175 73997 832231
rect 74053 832175 74139 832231
rect 74195 832175 74281 832231
rect 74337 832175 74423 832231
rect 74479 832175 74565 832231
rect 74621 832175 74707 832231
rect 74763 832175 74849 832231
rect 74905 832175 74991 832231
rect 75047 832175 75133 832231
rect 75189 832175 75275 832231
rect 75331 832175 75416 832231
rect 70475 832135 75416 832175
rect 70000 832089 75416 832135
rect 70000 832067 73855 832089
rect 70000 832011 70047 832067
rect 70103 832011 70171 832067
rect 70227 832011 70295 832067
rect 70351 832011 70419 832067
rect 70475 832033 73855 832067
rect 73911 832033 73997 832089
rect 74053 832033 74139 832089
rect 74195 832033 74281 832089
rect 74337 832033 74423 832089
rect 74479 832033 74565 832089
rect 74621 832033 74707 832089
rect 74763 832033 74849 832089
rect 74905 832033 74991 832089
rect 75047 832033 75133 832089
rect 75189 832033 75275 832089
rect 75331 832033 75416 832089
rect 70475 832011 75416 832033
rect 70000 831947 75416 832011
rect 70000 831943 73855 831947
rect 70000 831887 70047 831943
rect 70103 831887 70171 831943
rect 70227 831887 70295 831943
rect 70351 831887 70419 831943
rect 70475 831891 73855 831943
rect 73911 831891 73997 831947
rect 74053 831891 74139 831947
rect 74195 831891 74281 831947
rect 74337 831891 74423 831947
rect 74479 831891 74565 831947
rect 74621 831891 74707 831947
rect 74763 831891 74849 831947
rect 74905 831891 74991 831947
rect 75047 831891 75133 831947
rect 75189 831891 75275 831947
rect 75331 831891 75416 831947
rect 70475 831887 75416 831891
rect 70000 831819 75416 831887
rect 70000 831763 70047 831819
rect 70103 831763 70171 831819
rect 70227 831763 70295 831819
rect 70351 831763 70419 831819
rect 70475 831805 75416 831819
rect 70475 831763 73855 831805
rect 70000 831749 73855 831763
rect 73911 831749 73997 831805
rect 74053 831749 74139 831805
rect 74195 831749 74281 831805
rect 74337 831749 74423 831805
rect 74479 831749 74565 831805
rect 74621 831749 74707 831805
rect 74763 831749 74849 831805
rect 74905 831749 74991 831805
rect 75047 831749 75133 831805
rect 75189 831749 75275 831805
rect 75331 831749 75416 831805
rect 70000 831695 75416 831749
rect 70000 831639 70047 831695
rect 70103 831639 70171 831695
rect 70227 831639 70295 831695
rect 70351 831639 70419 831695
rect 70475 831663 75416 831695
rect 70475 831639 73855 831663
rect 70000 831607 73855 831639
rect 73911 831607 73997 831663
rect 74053 831607 74139 831663
rect 74195 831607 74281 831663
rect 74337 831607 74423 831663
rect 74479 831607 74565 831663
rect 74621 831607 74707 831663
rect 74763 831607 74849 831663
rect 74905 831607 74991 831663
rect 75047 831607 75133 831663
rect 75189 831607 75275 831663
rect 75331 831607 75416 831663
rect 70000 831571 75416 831607
rect 70000 831515 70047 831571
rect 70103 831515 70171 831571
rect 70227 831515 70295 831571
rect 70351 831515 70419 831571
rect 70475 831521 75416 831571
rect 70475 831515 73855 831521
rect 70000 831465 73855 831515
rect 73911 831465 73997 831521
rect 74053 831465 74139 831521
rect 74195 831465 74281 831521
rect 74337 831465 74423 831521
rect 74479 831465 74565 831521
rect 74621 831465 74707 831521
rect 74763 831465 74849 831521
rect 74905 831465 74991 831521
rect 75047 831465 75133 831521
rect 75189 831465 75275 831521
rect 75331 831465 75416 831521
rect 70000 831447 75416 831465
rect 70000 831391 70047 831447
rect 70103 831391 70171 831447
rect 70227 831391 70295 831447
rect 70351 831391 70419 831447
rect 70475 831391 75416 831447
rect 70000 831379 75416 831391
rect 70000 831323 73855 831379
rect 73911 831323 73997 831379
rect 74053 831323 74139 831379
rect 74195 831323 74281 831379
rect 74337 831323 74423 831379
rect 74479 831323 74565 831379
rect 74621 831323 74707 831379
rect 74763 831323 74849 831379
rect 74905 831323 74991 831379
rect 75047 831323 75133 831379
rect 75189 831323 75275 831379
rect 75331 831323 75416 831379
rect 70000 831267 70047 831323
rect 70103 831267 70171 831323
rect 70227 831267 70295 831323
rect 70351 831267 70419 831323
rect 70475 831267 75416 831323
rect 70000 831237 75416 831267
rect 70000 831199 73855 831237
rect 70000 831143 70047 831199
rect 70103 831143 70171 831199
rect 70227 831143 70295 831199
rect 70351 831143 70419 831199
rect 70475 831181 73855 831199
rect 73911 831181 73997 831237
rect 74053 831181 74139 831237
rect 74195 831181 74281 831237
rect 74337 831181 74423 831237
rect 74479 831181 74565 831237
rect 74621 831181 74707 831237
rect 74763 831181 74849 831237
rect 74905 831181 74991 831237
rect 75047 831181 75133 831237
rect 75189 831181 75275 831237
rect 75331 831181 75416 831237
rect 70475 831143 75416 831181
rect 70000 831095 75416 831143
rect 70000 831075 73855 831095
rect 70000 831019 70047 831075
rect 70103 831019 70171 831075
rect 70227 831019 70295 831075
rect 70351 831019 70419 831075
rect 70475 831039 73855 831075
rect 73911 831039 73997 831095
rect 74053 831039 74139 831095
rect 74195 831039 74281 831095
rect 74337 831039 74423 831095
rect 74479 831039 74565 831095
rect 74621 831039 74707 831095
rect 74763 831039 74849 831095
rect 74905 831039 74991 831095
rect 75047 831039 75133 831095
rect 75189 831039 75275 831095
rect 75331 831039 75416 831095
rect 70475 831019 75416 831039
rect 70000 830953 75416 831019
rect 70000 830951 73855 830953
rect 70000 830895 70047 830951
rect 70103 830895 70171 830951
rect 70227 830895 70295 830951
rect 70351 830895 70419 830951
rect 70475 830897 73855 830951
rect 73911 830897 73997 830953
rect 74053 830897 74139 830953
rect 74195 830897 74281 830953
rect 74337 830897 74423 830953
rect 74479 830897 74565 830953
rect 74621 830897 74707 830953
rect 74763 830897 74849 830953
rect 74905 830897 74991 830953
rect 75047 830897 75133 830953
rect 75189 830897 75275 830953
rect 75331 830897 75416 830953
rect 70475 830895 75416 830897
rect 70000 830828 75416 830895
rect 70000 830105 75416 830172
rect 70000 830049 70047 830105
rect 70103 830049 70171 830105
rect 70227 830049 70295 830105
rect 70351 830049 70419 830105
rect 70475 830093 75416 830105
rect 70475 830049 73855 830093
rect 70000 830037 73855 830049
rect 73911 830037 73997 830093
rect 74053 830037 74139 830093
rect 74195 830037 74281 830093
rect 74337 830037 74423 830093
rect 74479 830037 74565 830093
rect 74621 830037 74707 830093
rect 74763 830037 74849 830093
rect 74905 830037 74991 830093
rect 75047 830037 75133 830093
rect 75189 830037 75275 830093
rect 75331 830037 75416 830093
rect 70000 829981 75416 830037
rect 70000 829925 70047 829981
rect 70103 829925 70171 829981
rect 70227 829925 70295 829981
rect 70351 829925 70419 829981
rect 70475 829951 75416 829981
rect 70475 829925 73855 829951
rect 70000 829895 73855 829925
rect 73911 829895 73997 829951
rect 74053 829895 74139 829951
rect 74195 829895 74281 829951
rect 74337 829895 74423 829951
rect 74479 829895 74565 829951
rect 74621 829895 74707 829951
rect 74763 829895 74849 829951
rect 74905 829895 74991 829951
rect 75047 829895 75133 829951
rect 75189 829895 75275 829951
rect 75331 829895 75416 829951
rect 70000 829857 75416 829895
rect 70000 829801 70047 829857
rect 70103 829801 70171 829857
rect 70227 829801 70295 829857
rect 70351 829801 70419 829857
rect 70475 829809 75416 829857
rect 70475 829801 73855 829809
rect 70000 829753 73855 829801
rect 73911 829753 73997 829809
rect 74053 829753 74139 829809
rect 74195 829753 74281 829809
rect 74337 829753 74423 829809
rect 74479 829753 74565 829809
rect 74621 829753 74707 829809
rect 74763 829753 74849 829809
rect 74905 829753 74991 829809
rect 75047 829753 75133 829809
rect 75189 829753 75275 829809
rect 75331 829753 75416 829809
rect 70000 829733 75416 829753
rect 70000 829677 70047 829733
rect 70103 829677 70171 829733
rect 70227 829677 70295 829733
rect 70351 829677 70419 829733
rect 70475 829677 75416 829733
rect 70000 829667 75416 829677
rect 70000 829611 73855 829667
rect 73911 829611 73997 829667
rect 74053 829611 74139 829667
rect 74195 829611 74281 829667
rect 74337 829611 74423 829667
rect 74479 829611 74565 829667
rect 74621 829611 74707 829667
rect 74763 829611 74849 829667
rect 74905 829611 74991 829667
rect 75047 829611 75133 829667
rect 75189 829611 75275 829667
rect 75331 829611 75416 829667
rect 70000 829609 75416 829611
rect 70000 829553 70047 829609
rect 70103 829553 70171 829609
rect 70227 829553 70295 829609
rect 70351 829553 70419 829609
rect 70475 829553 75416 829609
rect 70000 829525 75416 829553
rect 70000 829485 73855 829525
rect 70000 829429 70047 829485
rect 70103 829429 70171 829485
rect 70227 829429 70295 829485
rect 70351 829429 70419 829485
rect 70475 829469 73855 829485
rect 73911 829469 73997 829525
rect 74053 829469 74139 829525
rect 74195 829469 74281 829525
rect 74337 829469 74423 829525
rect 74479 829469 74565 829525
rect 74621 829469 74707 829525
rect 74763 829469 74849 829525
rect 74905 829469 74991 829525
rect 75047 829469 75133 829525
rect 75189 829469 75275 829525
rect 75331 829469 75416 829525
rect 70475 829429 75416 829469
rect 70000 829383 75416 829429
rect 70000 829361 73855 829383
rect 70000 829305 70047 829361
rect 70103 829305 70171 829361
rect 70227 829305 70295 829361
rect 70351 829305 70419 829361
rect 70475 829327 73855 829361
rect 73911 829327 73997 829383
rect 74053 829327 74139 829383
rect 74195 829327 74281 829383
rect 74337 829327 74423 829383
rect 74479 829327 74565 829383
rect 74621 829327 74707 829383
rect 74763 829327 74849 829383
rect 74905 829327 74991 829383
rect 75047 829327 75133 829383
rect 75189 829327 75275 829383
rect 75331 829327 75416 829383
rect 70475 829305 75416 829327
rect 70000 829241 75416 829305
rect 70000 829237 73855 829241
rect 70000 829181 70047 829237
rect 70103 829181 70171 829237
rect 70227 829181 70295 829237
rect 70351 829181 70419 829237
rect 70475 829185 73855 829237
rect 73911 829185 73997 829241
rect 74053 829185 74139 829241
rect 74195 829185 74281 829241
rect 74337 829185 74423 829241
rect 74479 829185 74565 829241
rect 74621 829185 74707 829241
rect 74763 829185 74849 829241
rect 74905 829185 74991 829241
rect 75047 829185 75133 829241
rect 75189 829185 75275 829241
rect 75331 829185 75416 829241
rect 70475 829181 75416 829185
rect 70000 829113 75416 829181
rect 70000 829057 70047 829113
rect 70103 829057 70171 829113
rect 70227 829057 70295 829113
rect 70351 829057 70419 829113
rect 70475 829099 75416 829113
rect 70475 829057 73855 829099
rect 70000 829043 73855 829057
rect 73911 829043 73997 829099
rect 74053 829043 74139 829099
rect 74195 829043 74281 829099
rect 74337 829043 74423 829099
rect 74479 829043 74565 829099
rect 74621 829043 74707 829099
rect 74763 829043 74849 829099
rect 74905 829043 74991 829099
rect 75047 829043 75133 829099
rect 75189 829043 75275 829099
rect 75331 829043 75416 829099
rect 70000 828989 75416 829043
rect 70000 828933 70047 828989
rect 70103 828933 70171 828989
rect 70227 828933 70295 828989
rect 70351 828933 70419 828989
rect 70475 828957 75416 828989
rect 70475 828933 73855 828957
rect 70000 828901 73855 828933
rect 73911 828901 73997 828957
rect 74053 828901 74139 828957
rect 74195 828901 74281 828957
rect 74337 828901 74423 828957
rect 74479 828901 74565 828957
rect 74621 828901 74707 828957
rect 74763 828901 74849 828957
rect 74905 828901 74991 828957
rect 75047 828901 75133 828957
rect 75189 828901 75275 828957
rect 75331 828901 75416 828957
rect 70000 828865 75416 828901
rect 70000 828809 70047 828865
rect 70103 828809 70171 828865
rect 70227 828809 70295 828865
rect 70351 828809 70419 828865
rect 70475 828815 75416 828865
rect 70475 828809 73855 828815
rect 70000 828759 73855 828809
rect 73911 828759 73997 828815
rect 74053 828759 74139 828815
rect 74195 828759 74281 828815
rect 74337 828759 74423 828815
rect 74479 828759 74565 828815
rect 74621 828759 74707 828815
rect 74763 828759 74849 828815
rect 74905 828759 74991 828815
rect 75047 828759 75133 828815
rect 75189 828759 75275 828815
rect 75331 828759 75416 828815
rect 70000 828741 75416 828759
rect 70000 828685 70047 828741
rect 70103 828685 70171 828741
rect 70227 828685 70295 828741
rect 70351 828685 70419 828741
rect 70475 828685 75416 828741
rect 70000 828673 75416 828685
rect 70000 828617 73855 828673
rect 73911 828617 73997 828673
rect 74053 828617 74139 828673
rect 74195 828617 74281 828673
rect 74337 828617 74423 828673
rect 74479 828617 74565 828673
rect 74621 828617 74707 828673
rect 74763 828617 74849 828673
rect 74905 828617 74991 828673
rect 75047 828617 75133 828673
rect 75189 828617 75275 828673
rect 75331 828617 75416 828673
rect 70000 828561 70047 828617
rect 70103 828561 70171 828617
rect 70227 828561 70295 828617
rect 70351 828561 70419 828617
rect 70475 828561 75416 828617
rect 70000 828531 75416 828561
rect 70000 828493 73855 828531
rect 70000 828437 70047 828493
rect 70103 828437 70171 828493
rect 70227 828437 70295 828493
rect 70351 828437 70419 828493
rect 70475 828475 73855 828493
rect 73911 828475 73997 828531
rect 74053 828475 74139 828531
rect 74195 828475 74281 828531
rect 74337 828475 74423 828531
rect 74479 828475 74565 828531
rect 74621 828475 74707 828531
rect 74763 828475 74849 828531
rect 74905 828475 74991 828531
rect 75047 828475 75133 828531
rect 75189 828475 75275 828531
rect 75331 828475 75416 828531
rect 70475 828437 75416 828475
rect 70000 828389 75416 828437
rect 70000 828369 73855 828389
rect 70000 828313 70047 828369
rect 70103 828313 70171 828369
rect 70227 828313 70295 828369
rect 70351 828313 70419 828369
rect 70475 828333 73855 828369
rect 73911 828333 73997 828389
rect 74053 828333 74139 828389
rect 74195 828333 74281 828389
rect 74337 828333 74423 828389
rect 74479 828333 74565 828389
rect 74621 828333 74707 828389
rect 74763 828333 74849 828389
rect 74905 828333 74991 828389
rect 75047 828333 75133 828389
rect 75189 828333 75275 828389
rect 75331 828333 75416 828389
rect 70475 828313 75416 828333
rect 70000 828247 75416 828313
rect 70000 828245 73855 828247
rect 70000 828189 70047 828245
rect 70103 828189 70171 828245
rect 70227 828189 70295 828245
rect 70351 828189 70419 828245
rect 70475 828191 73855 828245
rect 73911 828191 73997 828247
rect 74053 828191 74139 828247
rect 74195 828191 74281 828247
rect 74337 828191 74423 828247
rect 74479 828191 74565 828247
rect 74621 828191 74707 828247
rect 74763 828191 74849 828247
rect 74905 828191 74991 828247
rect 75047 828191 75133 828247
rect 75189 828191 75275 828247
rect 75331 828191 75416 828247
rect 70475 828189 75416 828191
rect 70000 828122 75416 828189
rect 70000 827735 75416 827802
rect 70000 827679 70047 827735
rect 70103 827679 70171 827735
rect 70227 827679 70295 827735
rect 70351 827679 70419 827735
rect 70475 827723 75416 827735
rect 70475 827679 73855 827723
rect 70000 827667 73855 827679
rect 73911 827667 73997 827723
rect 74053 827667 74139 827723
rect 74195 827667 74281 827723
rect 74337 827667 74423 827723
rect 74479 827667 74565 827723
rect 74621 827667 74707 827723
rect 74763 827667 74849 827723
rect 74905 827667 74991 827723
rect 75047 827667 75133 827723
rect 75189 827667 75275 827723
rect 75331 827667 75416 827723
rect 70000 827611 75416 827667
rect 70000 827555 70047 827611
rect 70103 827555 70171 827611
rect 70227 827555 70295 827611
rect 70351 827555 70419 827611
rect 70475 827581 75416 827611
rect 70475 827555 73855 827581
rect 70000 827525 73855 827555
rect 73911 827525 73997 827581
rect 74053 827525 74139 827581
rect 74195 827525 74281 827581
rect 74337 827525 74423 827581
rect 74479 827525 74565 827581
rect 74621 827525 74707 827581
rect 74763 827525 74849 827581
rect 74905 827525 74991 827581
rect 75047 827525 75133 827581
rect 75189 827525 75275 827581
rect 75331 827525 75416 827581
rect 70000 827487 75416 827525
rect 70000 827431 70047 827487
rect 70103 827431 70171 827487
rect 70227 827431 70295 827487
rect 70351 827431 70419 827487
rect 70475 827439 75416 827487
rect 70475 827431 73855 827439
rect 70000 827383 73855 827431
rect 73911 827383 73997 827439
rect 74053 827383 74139 827439
rect 74195 827383 74281 827439
rect 74337 827383 74423 827439
rect 74479 827383 74565 827439
rect 74621 827383 74707 827439
rect 74763 827383 74849 827439
rect 74905 827383 74991 827439
rect 75047 827383 75133 827439
rect 75189 827383 75275 827439
rect 75331 827383 75416 827439
rect 70000 827363 75416 827383
rect 70000 827307 70047 827363
rect 70103 827307 70171 827363
rect 70227 827307 70295 827363
rect 70351 827307 70419 827363
rect 70475 827307 75416 827363
rect 70000 827297 75416 827307
rect 70000 827241 73855 827297
rect 73911 827241 73997 827297
rect 74053 827241 74139 827297
rect 74195 827241 74281 827297
rect 74337 827241 74423 827297
rect 74479 827241 74565 827297
rect 74621 827241 74707 827297
rect 74763 827241 74849 827297
rect 74905 827241 74991 827297
rect 75047 827241 75133 827297
rect 75189 827241 75275 827297
rect 75331 827241 75416 827297
rect 70000 827239 75416 827241
rect 70000 827183 70047 827239
rect 70103 827183 70171 827239
rect 70227 827183 70295 827239
rect 70351 827183 70419 827239
rect 70475 827183 75416 827239
rect 70000 827155 75416 827183
rect 70000 827115 73855 827155
rect 70000 827059 70047 827115
rect 70103 827059 70171 827115
rect 70227 827059 70295 827115
rect 70351 827059 70419 827115
rect 70475 827099 73855 827115
rect 73911 827099 73997 827155
rect 74053 827099 74139 827155
rect 74195 827099 74281 827155
rect 74337 827099 74423 827155
rect 74479 827099 74565 827155
rect 74621 827099 74707 827155
rect 74763 827099 74849 827155
rect 74905 827099 74991 827155
rect 75047 827099 75133 827155
rect 75189 827099 75275 827155
rect 75331 827099 75416 827155
rect 70475 827059 75416 827099
rect 70000 827013 75416 827059
rect 70000 826991 73855 827013
rect 70000 826935 70047 826991
rect 70103 826935 70171 826991
rect 70227 826935 70295 826991
rect 70351 826935 70419 826991
rect 70475 826957 73855 826991
rect 73911 826957 73997 827013
rect 74053 826957 74139 827013
rect 74195 826957 74281 827013
rect 74337 826957 74423 827013
rect 74479 826957 74565 827013
rect 74621 826957 74707 827013
rect 74763 826957 74849 827013
rect 74905 826957 74991 827013
rect 75047 826957 75133 827013
rect 75189 826957 75275 827013
rect 75331 826957 75416 827013
rect 70475 826935 75416 826957
rect 70000 826871 75416 826935
rect 70000 826867 73855 826871
rect 70000 826811 70047 826867
rect 70103 826811 70171 826867
rect 70227 826811 70295 826867
rect 70351 826811 70419 826867
rect 70475 826815 73855 826867
rect 73911 826815 73997 826871
rect 74053 826815 74139 826871
rect 74195 826815 74281 826871
rect 74337 826815 74423 826871
rect 74479 826815 74565 826871
rect 74621 826815 74707 826871
rect 74763 826815 74849 826871
rect 74905 826815 74991 826871
rect 75047 826815 75133 826871
rect 75189 826815 75275 826871
rect 75331 826815 75416 826871
rect 70475 826811 75416 826815
rect 70000 826743 75416 826811
rect 70000 826687 70047 826743
rect 70103 826687 70171 826743
rect 70227 826687 70295 826743
rect 70351 826687 70419 826743
rect 70475 826729 75416 826743
rect 70475 826687 73855 826729
rect 70000 826673 73855 826687
rect 73911 826673 73997 826729
rect 74053 826673 74139 826729
rect 74195 826673 74281 826729
rect 74337 826673 74423 826729
rect 74479 826673 74565 826729
rect 74621 826673 74707 826729
rect 74763 826673 74849 826729
rect 74905 826673 74991 826729
rect 75047 826673 75133 826729
rect 75189 826673 75275 826729
rect 75331 826673 75416 826729
rect 70000 826619 75416 826673
rect 70000 826563 70047 826619
rect 70103 826563 70171 826619
rect 70227 826563 70295 826619
rect 70351 826563 70419 826619
rect 70475 826587 75416 826619
rect 70475 826563 73855 826587
rect 70000 826531 73855 826563
rect 73911 826531 73997 826587
rect 74053 826531 74139 826587
rect 74195 826531 74281 826587
rect 74337 826531 74423 826587
rect 74479 826531 74565 826587
rect 74621 826531 74707 826587
rect 74763 826531 74849 826587
rect 74905 826531 74991 826587
rect 75047 826531 75133 826587
rect 75189 826531 75275 826587
rect 75331 826531 75416 826587
rect 70000 826495 75416 826531
rect 70000 826439 70047 826495
rect 70103 826439 70171 826495
rect 70227 826439 70295 826495
rect 70351 826439 70419 826495
rect 70475 826445 75416 826495
rect 70475 826439 73855 826445
rect 70000 826389 73855 826439
rect 73911 826389 73997 826445
rect 74053 826389 74139 826445
rect 74195 826389 74281 826445
rect 74337 826389 74423 826445
rect 74479 826389 74565 826445
rect 74621 826389 74707 826445
rect 74763 826389 74849 826445
rect 74905 826389 74991 826445
rect 75047 826389 75133 826445
rect 75189 826389 75275 826445
rect 75331 826389 75416 826445
rect 70000 826371 75416 826389
rect 70000 826315 70047 826371
rect 70103 826315 70171 826371
rect 70227 826315 70295 826371
rect 70351 826315 70419 826371
rect 70475 826315 75416 826371
rect 70000 826303 75416 826315
rect 70000 826247 73855 826303
rect 73911 826247 73997 826303
rect 74053 826247 74139 826303
rect 74195 826247 74281 826303
rect 74337 826247 74423 826303
rect 74479 826247 74565 826303
rect 74621 826247 74707 826303
rect 74763 826247 74849 826303
rect 74905 826247 74991 826303
rect 75047 826247 75133 826303
rect 75189 826247 75275 826303
rect 75331 826247 75416 826303
rect 70000 826191 70047 826247
rect 70103 826191 70171 826247
rect 70227 826191 70295 826247
rect 70351 826191 70419 826247
rect 70475 826191 75416 826247
rect 70000 826161 75416 826191
rect 70000 826123 73855 826161
rect 70000 826067 70047 826123
rect 70103 826067 70171 826123
rect 70227 826067 70295 826123
rect 70351 826067 70419 826123
rect 70475 826105 73855 826123
rect 73911 826105 73997 826161
rect 74053 826105 74139 826161
rect 74195 826105 74281 826161
rect 74337 826105 74423 826161
rect 74479 826105 74565 826161
rect 74621 826105 74707 826161
rect 74763 826105 74849 826161
rect 74905 826105 74991 826161
rect 75047 826105 75133 826161
rect 75189 826105 75275 826161
rect 75331 826105 75416 826161
rect 70475 826067 75416 826105
rect 70000 826019 75416 826067
rect 70000 825999 73855 826019
rect 70000 825943 70047 825999
rect 70103 825943 70171 825999
rect 70227 825943 70295 825999
rect 70351 825943 70419 825999
rect 70475 825963 73855 825999
rect 73911 825963 73997 826019
rect 74053 825963 74139 826019
rect 74195 825963 74281 826019
rect 74337 825963 74423 826019
rect 74479 825963 74565 826019
rect 74621 825963 74707 826019
rect 74763 825963 74849 826019
rect 74905 825963 74991 826019
rect 75047 825963 75133 826019
rect 75189 825963 75275 826019
rect 75331 825963 75416 826019
rect 70475 825943 75416 825963
rect 70000 825877 75416 825943
rect 70000 825875 73855 825877
rect 70000 825819 70047 825875
rect 70103 825819 70171 825875
rect 70227 825819 70295 825875
rect 70351 825819 70419 825875
rect 70475 825821 73855 825875
rect 73911 825821 73997 825877
rect 74053 825821 74139 825877
rect 74195 825821 74281 825877
rect 74337 825821 74423 825877
rect 74479 825821 74565 825877
rect 74621 825821 74707 825877
rect 74763 825821 74849 825877
rect 74905 825821 74991 825877
rect 75047 825821 75133 825877
rect 75189 825821 75275 825877
rect 75331 825821 75416 825877
rect 70475 825819 75416 825821
rect 70000 825752 75416 825819
rect 70000 825105 75416 825172
rect 70000 825049 70047 825105
rect 70103 825049 70171 825105
rect 70227 825049 70295 825105
rect 70351 825049 70419 825105
rect 70475 825094 75416 825105
rect 70475 825049 73866 825094
rect 70000 825038 73866 825049
rect 73922 825038 74008 825094
rect 74064 825038 74150 825094
rect 74206 825038 74292 825094
rect 74348 825038 74434 825094
rect 74490 825038 74576 825094
rect 74632 825038 74718 825094
rect 74774 825038 74860 825094
rect 74916 825038 75002 825094
rect 75058 825038 75144 825094
rect 75200 825038 75286 825094
rect 75342 825038 75416 825094
rect 70000 824981 75416 825038
rect 70000 824925 70047 824981
rect 70103 824925 70171 824981
rect 70227 824925 70295 824981
rect 70351 824925 70419 824981
rect 70475 824952 75416 824981
rect 70475 824925 73866 824952
rect 70000 824896 73866 824925
rect 73922 824896 74008 824952
rect 74064 824896 74150 824952
rect 74206 824896 74292 824952
rect 74348 824896 74434 824952
rect 74490 824896 74576 824952
rect 74632 824896 74718 824952
rect 74774 824896 74860 824952
rect 74916 824896 75002 824952
rect 75058 824896 75144 824952
rect 75200 824896 75286 824952
rect 75342 824896 75416 824952
rect 70000 824857 75416 824896
rect 70000 824801 70047 824857
rect 70103 824801 70171 824857
rect 70227 824801 70295 824857
rect 70351 824801 70419 824857
rect 70475 824810 75416 824857
rect 70475 824801 73866 824810
rect 70000 824754 73866 824801
rect 73922 824754 74008 824810
rect 74064 824754 74150 824810
rect 74206 824754 74292 824810
rect 74348 824754 74434 824810
rect 74490 824754 74576 824810
rect 74632 824754 74718 824810
rect 74774 824754 74860 824810
rect 74916 824754 75002 824810
rect 75058 824754 75144 824810
rect 75200 824754 75286 824810
rect 75342 824754 75416 824810
rect 70000 824733 75416 824754
rect 70000 824677 70047 824733
rect 70103 824677 70171 824733
rect 70227 824677 70295 824733
rect 70351 824677 70419 824733
rect 70475 824677 75416 824733
rect 70000 824668 75416 824677
rect 70000 824612 73866 824668
rect 73922 824612 74008 824668
rect 74064 824612 74150 824668
rect 74206 824612 74292 824668
rect 74348 824612 74434 824668
rect 74490 824612 74576 824668
rect 74632 824612 74718 824668
rect 74774 824612 74860 824668
rect 74916 824612 75002 824668
rect 75058 824612 75144 824668
rect 75200 824612 75286 824668
rect 75342 824612 75416 824668
rect 70000 824609 75416 824612
rect 70000 824553 70047 824609
rect 70103 824553 70171 824609
rect 70227 824553 70295 824609
rect 70351 824553 70419 824609
rect 70475 824553 75416 824609
rect 70000 824526 75416 824553
rect 70000 824485 73866 824526
rect 70000 824429 70047 824485
rect 70103 824429 70171 824485
rect 70227 824429 70295 824485
rect 70351 824429 70419 824485
rect 70475 824470 73866 824485
rect 73922 824470 74008 824526
rect 74064 824470 74150 824526
rect 74206 824470 74292 824526
rect 74348 824470 74434 824526
rect 74490 824470 74576 824526
rect 74632 824470 74718 824526
rect 74774 824470 74860 824526
rect 74916 824470 75002 824526
rect 75058 824470 75144 824526
rect 75200 824470 75286 824526
rect 75342 824470 75416 824526
rect 70475 824429 75416 824470
rect 70000 824384 75416 824429
rect 70000 824361 73866 824384
rect 70000 824305 70047 824361
rect 70103 824305 70171 824361
rect 70227 824305 70295 824361
rect 70351 824305 70419 824361
rect 70475 824328 73866 824361
rect 73922 824328 74008 824384
rect 74064 824328 74150 824384
rect 74206 824328 74292 824384
rect 74348 824328 74434 824384
rect 74490 824328 74576 824384
rect 74632 824328 74718 824384
rect 74774 824328 74860 824384
rect 74916 824328 75002 824384
rect 75058 824328 75144 824384
rect 75200 824328 75286 824384
rect 75342 824328 75416 824384
rect 70475 824305 75416 824328
rect 70000 824242 75416 824305
rect 70000 824237 73866 824242
rect 70000 824181 70047 824237
rect 70103 824181 70171 824237
rect 70227 824181 70295 824237
rect 70351 824181 70419 824237
rect 70475 824186 73866 824237
rect 73922 824186 74008 824242
rect 74064 824186 74150 824242
rect 74206 824186 74292 824242
rect 74348 824186 74434 824242
rect 74490 824186 74576 824242
rect 74632 824186 74718 824242
rect 74774 824186 74860 824242
rect 74916 824186 75002 824242
rect 75058 824186 75144 824242
rect 75200 824186 75286 824242
rect 75342 824186 75416 824242
rect 70475 824181 75416 824186
rect 70000 824113 75416 824181
rect 70000 824057 70047 824113
rect 70103 824057 70171 824113
rect 70227 824057 70295 824113
rect 70351 824057 70419 824113
rect 70475 824100 75416 824113
rect 70475 824057 73866 824100
rect 70000 824044 73866 824057
rect 73922 824044 74008 824100
rect 74064 824044 74150 824100
rect 74206 824044 74292 824100
rect 74348 824044 74434 824100
rect 74490 824044 74576 824100
rect 74632 824044 74718 824100
rect 74774 824044 74860 824100
rect 74916 824044 75002 824100
rect 75058 824044 75144 824100
rect 75200 824044 75286 824100
rect 75342 824044 75416 824100
rect 70000 823989 75416 824044
rect 70000 823933 70047 823989
rect 70103 823933 70171 823989
rect 70227 823933 70295 823989
rect 70351 823933 70419 823989
rect 70475 823958 75416 823989
rect 70475 823933 73866 823958
rect 70000 823902 73866 823933
rect 73922 823902 74008 823958
rect 74064 823902 74150 823958
rect 74206 823902 74292 823958
rect 74348 823902 74434 823958
rect 74490 823902 74576 823958
rect 74632 823902 74718 823958
rect 74774 823902 74860 823958
rect 74916 823902 75002 823958
rect 75058 823902 75144 823958
rect 75200 823902 75286 823958
rect 75342 823902 75416 823958
rect 70000 823865 75416 823902
rect 70000 823809 70047 823865
rect 70103 823809 70171 823865
rect 70227 823809 70295 823865
rect 70351 823809 70419 823865
rect 70475 823816 75416 823865
rect 70475 823809 73866 823816
rect 70000 823760 73866 823809
rect 73922 823760 74008 823816
rect 74064 823760 74150 823816
rect 74206 823760 74292 823816
rect 74348 823760 74434 823816
rect 74490 823760 74576 823816
rect 74632 823760 74718 823816
rect 74774 823760 74860 823816
rect 74916 823760 75002 823816
rect 75058 823760 75144 823816
rect 75200 823760 75286 823816
rect 75342 823760 75416 823816
rect 70000 823741 75416 823760
rect 70000 823685 70047 823741
rect 70103 823685 70171 823741
rect 70227 823685 70295 823741
rect 70351 823685 70419 823741
rect 70475 823685 75416 823741
rect 70000 823674 75416 823685
rect 70000 823618 73866 823674
rect 73922 823618 74008 823674
rect 74064 823618 74150 823674
rect 74206 823618 74292 823674
rect 74348 823618 74434 823674
rect 74490 823618 74576 823674
rect 74632 823618 74718 823674
rect 74774 823618 74860 823674
rect 74916 823618 75002 823674
rect 75058 823618 75144 823674
rect 75200 823618 75286 823674
rect 75342 823618 75416 823674
rect 70000 823617 75416 823618
rect 70000 823561 70047 823617
rect 70103 823561 70171 823617
rect 70227 823561 70295 823617
rect 70351 823561 70419 823617
rect 70475 823561 75416 823617
rect 70000 823532 75416 823561
rect 70000 823493 73866 823532
rect 70000 823437 70047 823493
rect 70103 823437 70171 823493
rect 70227 823437 70295 823493
rect 70351 823437 70419 823493
rect 70475 823476 73866 823493
rect 73922 823476 74008 823532
rect 74064 823476 74150 823532
rect 74206 823476 74292 823532
rect 74348 823476 74434 823532
rect 74490 823476 74576 823532
rect 74632 823476 74718 823532
rect 74774 823476 74860 823532
rect 74916 823476 75002 823532
rect 75058 823476 75144 823532
rect 75200 823476 75286 823532
rect 75342 823476 75416 823532
rect 70475 823437 75416 823476
rect 70000 823390 75416 823437
rect 70000 823369 73866 823390
rect 70000 823313 70047 823369
rect 70103 823313 70171 823369
rect 70227 823313 70295 823369
rect 70351 823313 70419 823369
rect 70475 823334 73866 823369
rect 73922 823334 74008 823390
rect 74064 823334 74150 823390
rect 74206 823334 74292 823390
rect 74348 823334 74434 823390
rect 74490 823334 74576 823390
rect 74632 823334 74718 823390
rect 74774 823334 74860 823390
rect 74916 823334 75002 823390
rect 75058 823334 75144 823390
rect 75200 823334 75286 823390
rect 75342 823334 75416 823390
rect 70475 823313 75416 823334
rect 70000 823272 75416 823313
rect 70000 796661 73416 796728
rect 70000 796605 70047 796661
rect 70103 796605 70171 796661
rect 70227 796605 70295 796661
rect 70351 796605 70419 796661
rect 70475 796650 73416 796661
rect 70475 796605 71466 796650
rect 70000 796594 71466 796605
rect 71522 796594 71608 796650
rect 71664 796594 71750 796650
rect 71806 796594 71892 796650
rect 71948 796594 72034 796650
rect 72090 796594 72176 796650
rect 72232 796594 72318 796650
rect 72374 796594 72460 796650
rect 72516 796594 72602 796650
rect 72658 796594 72744 796650
rect 72800 796594 72886 796650
rect 72942 796594 73028 796650
rect 73084 796594 73170 796650
rect 73226 796594 73312 796650
rect 73368 796594 73416 796650
rect 70000 796537 73416 796594
rect 70000 796481 70047 796537
rect 70103 796481 70171 796537
rect 70227 796481 70295 796537
rect 70351 796481 70419 796537
rect 70475 796508 73416 796537
rect 70475 796481 71466 796508
rect 70000 796452 71466 796481
rect 71522 796452 71608 796508
rect 71664 796452 71750 796508
rect 71806 796452 71892 796508
rect 71948 796452 72034 796508
rect 72090 796452 72176 796508
rect 72232 796452 72318 796508
rect 72374 796452 72460 796508
rect 72516 796452 72602 796508
rect 72658 796452 72744 796508
rect 72800 796452 72886 796508
rect 72942 796452 73028 796508
rect 73084 796452 73170 796508
rect 73226 796452 73312 796508
rect 73368 796452 73416 796508
rect 70000 796413 73416 796452
rect 70000 796357 70047 796413
rect 70103 796357 70171 796413
rect 70227 796357 70295 796413
rect 70351 796357 70419 796413
rect 70475 796366 73416 796413
rect 70475 796357 71466 796366
rect 70000 796310 71466 796357
rect 71522 796310 71608 796366
rect 71664 796310 71750 796366
rect 71806 796310 71892 796366
rect 71948 796310 72034 796366
rect 72090 796310 72176 796366
rect 72232 796310 72318 796366
rect 72374 796310 72460 796366
rect 72516 796310 72602 796366
rect 72658 796310 72744 796366
rect 72800 796310 72886 796366
rect 72942 796310 73028 796366
rect 73084 796310 73170 796366
rect 73226 796310 73312 796366
rect 73368 796310 73416 796366
rect 70000 796289 73416 796310
rect 70000 796233 70047 796289
rect 70103 796233 70171 796289
rect 70227 796233 70295 796289
rect 70351 796233 70419 796289
rect 70475 796233 73416 796289
rect 70000 796224 73416 796233
rect 70000 796168 71466 796224
rect 71522 796168 71608 796224
rect 71664 796168 71750 796224
rect 71806 796168 71892 796224
rect 71948 796168 72034 796224
rect 72090 796168 72176 796224
rect 72232 796168 72318 796224
rect 72374 796168 72460 796224
rect 72516 796168 72602 796224
rect 72658 796168 72744 796224
rect 72800 796168 72886 796224
rect 72942 796168 73028 796224
rect 73084 796168 73170 796224
rect 73226 796168 73312 796224
rect 73368 796168 73416 796224
rect 70000 796165 73416 796168
rect 70000 796109 70047 796165
rect 70103 796109 70171 796165
rect 70227 796109 70295 796165
rect 70351 796109 70419 796165
rect 70475 796109 73416 796165
rect 70000 796082 73416 796109
rect 70000 796041 71466 796082
rect 70000 795985 70047 796041
rect 70103 795985 70171 796041
rect 70227 795985 70295 796041
rect 70351 795985 70419 796041
rect 70475 796026 71466 796041
rect 71522 796026 71608 796082
rect 71664 796026 71750 796082
rect 71806 796026 71892 796082
rect 71948 796026 72034 796082
rect 72090 796026 72176 796082
rect 72232 796026 72318 796082
rect 72374 796026 72460 796082
rect 72516 796026 72602 796082
rect 72658 796026 72744 796082
rect 72800 796026 72886 796082
rect 72942 796026 73028 796082
rect 73084 796026 73170 796082
rect 73226 796026 73312 796082
rect 73368 796026 73416 796082
rect 70475 795985 73416 796026
rect 70000 795940 73416 795985
rect 70000 795917 71466 795940
rect 70000 795861 70047 795917
rect 70103 795861 70171 795917
rect 70227 795861 70295 795917
rect 70351 795861 70419 795917
rect 70475 795884 71466 795917
rect 71522 795884 71608 795940
rect 71664 795884 71750 795940
rect 71806 795884 71892 795940
rect 71948 795884 72034 795940
rect 72090 795884 72176 795940
rect 72232 795884 72318 795940
rect 72374 795884 72460 795940
rect 72516 795884 72602 795940
rect 72658 795884 72744 795940
rect 72800 795884 72886 795940
rect 72942 795884 73028 795940
rect 73084 795884 73170 795940
rect 73226 795884 73312 795940
rect 73368 795884 73416 795940
rect 70475 795861 73416 795884
rect 70000 795798 73416 795861
rect 70000 795793 71466 795798
rect 70000 795737 70047 795793
rect 70103 795737 70171 795793
rect 70227 795737 70295 795793
rect 70351 795737 70419 795793
rect 70475 795742 71466 795793
rect 71522 795742 71608 795798
rect 71664 795742 71750 795798
rect 71806 795742 71892 795798
rect 71948 795742 72034 795798
rect 72090 795742 72176 795798
rect 72232 795742 72318 795798
rect 72374 795742 72460 795798
rect 72516 795742 72602 795798
rect 72658 795742 72744 795798
rect 72800 795742 72886 795798
rect 72942 795742 73028 795798
rect 73084 795742 73170 795798
rect 73226 795742 73312 795798
rect 73368 795742 73416 795798
rect 70475 795737 73416 795742
rect 70000 795669 73416 795737
rect 70000 795613 70047 795669
rect 70103 795613 70171 795669
rect 70227 795613 70295 795669
rect 70351 795613 70419 795669
rect 70475 795656 73416 795669
rect 70475 795613 71466 795656
rect 70000 795600 71466 795613
rect 71522 795600 71608 795656
rect 71664 795600 71750 795656
rect 71806 795600 71892 795656
rect 71948 795600 72034 795656
rect 72090 795600 72176 795656
rect 72232 795600 72318 795656
rect 72374 795600 72460 795656
rect 72516 795600 72602 795656
rect 72658 795600 72744 795656
rect 72800 795600 72886 795656
rect 72942 795600 73028 795656
rect 73084 795600 73170 795656
rect 73226 795600 73312 795656
rect 73368 795600 73416 795656
rect 70000 795545 73416 795600
rect 70000 795489 70047 795545
rect 70103 795489 70171 795545
rect 70227 795489 70295 795545
rect 70351 795489 70419 795545
rect 70475 795514 73416 795545
rect 70475 795489 71466 795514
rect 70000 795458 71466 795489
rect 71522 795458 71608 795514
rect 71664 795458 71750 795514
rect 71806 795458 71892 795514
rect 71948 795458 72034 795514
rect 72090 795458 72176 795514
rect 72232 795458 72318 795514
rect 72374 795458 72460 795514
rect 72516 795458 72602 795514
rect 72658 795458 72744 795514
rect 72800 795458 72886 795514
rect 72942 795458 73028 795514
rect 73084 795458 73170 795514
rect 73226 795458 73312 795514
rect 73368 795458 73416 795514
rect 70000 795421 73416 795458
rect 70000 795365 70047 795421
rect 70103 795365 70171 795421
rect 70227 795365 70295 795421
rect 70351 795365 70419 795421
rect 70475 795372 73416 795421
rect 70475 795365 71466 795372
rect 70000 795316 71466 795365
rect 71522 795316 71608 795372
rect 71664 795316 71750 795372
rect 71806 795316 71892 795372
rect 71948 795316 72034 795372
rect 72090 795316 72176 795372
rect 72232 795316 72318 795372
rect 72374 795316 72460 795372
rect 72516 795316 72602 795372
rect 72658 795316 72744 795372
rect 72800 795316 72886 795372
rect 72942 795316 73028 795372
rect 73084 795316 73170 795372
rect 73226 795316 73312 795372
rect 73368 795316 73416 795372
rect 70000 795297 73416 795316
rect 70000 795241 70047 795297
rect 70103 795241 70171 795297
rect 70227 795241 70295 795297
rect 70351 795241 70419 795297
rect 70475 795241 73416 795297
rect 70000 795230 73416 795241
rect 70000 795174 71466 795230
rect 71522 795174 71608 795230
rect 71664 795174 71750 795230
rect 71806 795174 71892 795230
rect 71948 795174 72034 795230
rect 72090 795174 72176 795230
rect 72232 795174 72318 795230
rect 72374 795174 72460 795230
rect 72516 795174 72602 795230
rect 72658 795174 72744 795230
rect 72800 795174 72886 795230
rect 72942 795174 73028 795230
rect 73084 795174 73170 795230
rect 73226 795174 73312 795230
rect 73368 795174 73416 795230
rect 70000 795173 73416 795174
rect 70000 795117 70047 795173
rect 70103 795117 70171 795173
rect 70227 795117 70295 795173
rect 70351 795117 70419 795173
rect 70475 795117 73416 795173
rect 70000 795088 73416 795117
rect 70000 795049 71466 795088
rect 70000 794993 70047 795049
rect 70103 794993 70171 795049
rect 70227 794993 70295 795049
rect 70351 794993 70419 795049
rect 70475 795032 71466 795049
rect 71522 795032 71608 795088
rect 71664 795032 71750 795088
rect 71806 795032 71892 795088
rect 71948 795032 72034 795088
rect 72090 795032 72176 795088
rect 72232 795032 72318 795088
rect 72374 795032 72460 795088
rect 72516 795032 72602 795088
rect 72658 795032 72744 795088
rect 72800 795032 72886 795088
rect 72942 795032 73028 795088
rect 73084 795032 73170 795088
rect 73226 795032 73312 795088
rect 73368 795032 73416 795088
rect 70475 794993 73416 795032
rect 70000 794946 73416 794993
rect 70000 794925 71466 794946
rect 70000 794869 70047 794925
rect 70103 794869 70171 794925
rect 70227 794869 70295 794925
rect 70351 794869 70419 794925
rect 70475 794890 71466 794925
rect 71522 794890 71608 794946
rect 71664 794890 71750 794946
rect 71806 794890 71892 794946
rect 71948 794890 72034 794946
rect 72090 794890 72176 794946
rect 72232 794890 72318 794946
rect 72374 794890 72460 794946
rect 72516 794890 72602 794946
rect 72658 794890 72744 794946
rect 72800 794890 72886 794946
rect 72942 794890 73028 794946
rect 73084 794890 73170 794946
rect 73226 794890 73312 794946
rect 73368 794890 73416 794946
rect 70475 794869 73416 794890
rect 70000 794828 73416 794869
rect 70000 794181 73416 794248
rect 70000 794125 70047 794181
rect 70103 794125 70171 794181
rect 70227 794125 70295 794181
rect 70351 794125 70419 794181
rect 70475 794169 73416 794181
rect 70475 794125 71455 794169
rect 70000 794113 71455 794125
rect 71511 794113 71597 794169
rect 71653 794113 71739 794169
rect 71795 794113 71881 794169
rect 71937 794113 72023 794169
rect 72079 794113 72165 794169
rect 72221 794113 72307 794169
rect 72363 794113 72449 794169
rect 72505 794113 72591 794169
rect 72647 794113 72733 794169
rect 72789 794113 72875 794169
rect 72931 794113 73017 794169
rect 73073 794113 73159 794169
rect 73215 794113 73301 794169
rect 73357 794113 73416 794169
rect 70000 794057 73416 794113
rect 70000 794001 70047 794057
rect 70103 794001 70171 794057
rect 70227 794001 70295 794057
rect 70351 794001 70419 794057
rect 70475 794027 73416 794057
rect 70475 794001 71455 794027
rect 70000 793971 71455 794001
rect 71511 793971 71597 794027
rect 71653 793971 71739 794027
rect 71795 793971 71881 794027
rect 71937 793971 72023 794027
rect 72079 793971 72165 794027
rect 72221 793971 72307 794027
rect 72363 793971 72449 794027
rect 72505 793971 72591 794027
rect 72647 793971 72733 794027
rect 72789 793971 72875 794027
rect 72931 793971 73017 794027
rect 73073 793971 73159 794027
rect 73215 793971 73301 794027
rect 73357 793971 73416 794027
rect 70000 793933 73416 793971
rect 70000 793877 70047 793933
rect 70103 793877 70171 793933
rect 70227 793877 70295 793933
rect 70351 793877 70419 793933
rect 70475 793885 73416 793933
rect 70475 793877 71455 793885
rect 70000 793829 71455 793877
rect 71511 793829 71597 793885
rect 71653 793829 71739 793885
rect 71795 793829 71881 793885
rect 71937 793829 72023 793885
rect 72079 793829 72165 793885
rect 72221 793829 72307 793885
rect 72363 793829 72449 793885
rect 72505 793829 72591 793885
rect 72647 793829 72733 793885
rect 72789 793829 72875 793885
rect 72931 793829 73017 793885
rect 73073 793829 73159 793885
rect 73215 793829 73301 793885
rect 73357 793829 73416 793885
rect 70000 793809 73416 793829
rect 70000 793753 70047 793809
rect 70103 793753 70171 793809
rect 70227 793753 70295 793809
rect 70351 793753 70419 793809
rect 70475 793753 73416 793809
rect 70000 793743 73416 793753
rect 70000 793687 71455 793743
rect 71511 793687 71597 793743
rect 71653 793687 71739 793743
rect 71795 793687 71881 793743
rect 71937 793687 72023 793743
rect 72079 793687 72165 793743
rect 72221 793687 72307 793743
rect 72363 793687 72449 793743
rect 72505 793687 72591 793743
rect 72647 793687 72733 793743
rect 72789 793687 72875 793743
rect 72931 793687 73017 793743
rect 73073 793687 73159 793743
rect 73215 793687 73301 793743
rect 73357 793687 73416 793743
rect 70000 793685 73416 793687
rect 70000 793629 70047 793685
rect 70103 793629 70171 793685
rect 70227 793629 70295 793685
rect 70351 793629 70419 793685
rect 70475 793629 73416 793685
rect 70000 793601 73416 793629
rect 70000 793561 71455 793601
rect 70000 793505 70047 793561
rect 70103 793505 70171 793561
rect 70227 793505 70295 793561
rect 70351 793505 70419 793561
rect 70475 793545 71455 793561
rect 71511 793545 71597 793601
rect 71653 793545 71739 793601
rect 71795 793545 71881 793601
rect 71937 793545 72023 793601
rect 72079 793545 72165 793601
rect 72221 793545 72307 793601
rect 72363 793545 72449 793601
rect 72505 793545 72591 793601
rect 72647 793545 72733 793601
rect 72789 793545 72875 793601
rect 72931 793545 73017 793601
rect 73073 793545 73159 793601
rect 73215 793545 73301 793601
rect 73357 793545 73416 793601
rect 70475 793505 73416 793545
rect 70000 793459 73416 793505
rect 70000 793437 71455 793459
rect 70000 793381 70047 793437
rect 70103 793381 70171 793437
rect 70227 793381 70295 793437
rect 70351 793381 70419 793437
rect 70475 793403 71455 793437
rect 71511 793403 71597 793459
rect 71653 793403 71739 793459
rect 71795 793403 71881 793459
rect 71937 793403 72023 793459
rect 72079 793403 72165 793459
rect 72221 793403 72307 793459
rect 72363 793403 72449 793459
rect 72505 793403 72591 793459
rect 72647 793403 72733 793459
rect 72789 793403 72875 793459
rect 72931 793403 73017 793459
rect 73073 793403 73159 793459
rect 73215 793403 73301 793459
rect 73357 793403 73416 793459
rect 70475 793381 73416 793403
rect 70000 793317 73416 793381
rect 70000 793313 71455 793317
rect 70000 793257 70047 793313
rect 70103 793257 70171 793313
rect 70227 793257 70295 793313
rect 70351 793257 70419 793313
rect 70475 793261 71455 793313
rect 71511 793261 71597 793317
rect 71653 793261 71739 793317
rect 71795 793261 71881 793317
rect 71937 793261 72023 793317
rect 72079 793261 72165 793317
rect 72221 793261 72307 793317
rect 72363 793261 72449 793317
rect 72505 793261 72591 793317
rect 72647 793261 72733 793317
rect 72789 793261 72875 793317
rect 72931 793261 73017 793317
rect 73073 793261 73159 793317
rect 73215 793261 73301 793317
rect 73357 793261 73416 793317
rect 70475 793257 73416 793261
rect 70000 793189 73416 793257
rect 70000 793133 70047 793189
rect 70103 793133 70171 793189
rect 70227 793133 70295 793189
rect 70351 793133 70419 793189
rect 70475 793175 73416 793189
rect 70475 793133 71455 793175
rect 70000 793119 71455 793133
rect 71511 793119 71597 793175
rect 71653 793119 71739 793175
rect 71795 793119 71881 793175
rect 71937 793119 72023 793175
rect 72079 793119 72165 793175
rect 72221 793119 72307 793175
rect 72363 793119 72449 793175
rect 72505 793119 72591 793175
rect 72647 793119 72733 793175
rect 72789 793119 72875 793175
rect 72931 793119 73017 793175
rect 73073 793119 73159 793175
rect 73215 793119 73301 793175
rect 73357 793119 73416 793175
rect 70000 793065 73416 793119
rect 70000 793009 70047 793065
rect 70103 793009 70171 793065
rect 70227 793009 70295 793065
rect 70351 793009 70419 793065
rect 70475 793033 73416 793065
rect 70475 793009 71455 793033
rect 70000 792977 71455 793009
rect 71511 792977 71597 793033
rect 71653 792977 71739 793033
rect 71795 792977 71881 793033
rect 71937 792977 72023 793033
rect 72079 792977 72165 793033
rect 72221 792977 72307 793033
rect 72363 792977 72449 793033
rect 72505 792977 72591 793033
rect 72647 792977 72733 793033
rect 72789 792977 72875 793033
rect 72931 792977 73017 793033
rect 73073 792977 73159 793033
rect 73215 792977 73301 793033
rect 73357 792977 73416 793033
rect 70000 792941 73416 792977
rect 70000 792885 70047 792941
rect 70103 792885 70171 792941
rect 70227 792885 70295 792941
rect 70351 792885 70419 792941
rect 70475 792891 73416 792941
rect 70475 792885 71455 792891
rect 70000 792835 71455 792885
rect 71511 792835 71597 792891
rect 71653 792835 71739 792891
rect 71795 792835 71881 792891
rect 71937 792835 72023 792891
rect 72079 792835 72165 792891
rect 72221 792835 72307 792891
rect 72363 792835 72449 792891
rect 72505 792835 72591 792891
rect 72647 792835 72733 792891
rect 72789 792835 72875 792891
rect 72931 792835 73017 792891
rect 73073 792835 73159 792891
rect 73215 792835 73301 792891
rect 73357 792835 73416 792891
rect 70000 792817 73416 792835
rect 70000 792761 70047 792817
rect 70103 792761 70171 792817
rect 70227 792761 70295 792817
rect 70351 792761 70419 792817
rect 70475 792761 73416 792817
rect 70000 792749 73416 792761
rect 70000 792693 71455 792749
rect 71511 792693 71597 792749
rect 71653 792693 71739 792749
rect 71795 792693 71881 792749
rect 71937 792693 72023 792749
rect 72079 792693 72165 792749
rect 72221 792693 72307 792749
rect 72363 792693 72449 792749
rect 72505 792693 72591 792749
rect 72647 792693 72733 792749
rect 72789 792693 72875 792749
rect 72931 792693 73017 792749
rect 73073 792693 73159 792749
rect 73215 792693 73301 792749
rect 73357 792693 73416 792749
rect 70000 792637 70047 792693
rect 70103 792637 70171 792693
rect 70227 792637 70295 792693
rect 70351 792637 70419 792693
rect 70475 792637 73416 792693
rect 70000 792607 73416 792637
rect 70000 792569 71455 792607
rect 70000 792513 70047 792569
rect 70103 792513 70171 792569
rect 70227 792513 70295 792569
rect 70351 792513 70419 792569
rect 70475 792551 71455 792569
rect 71511 792551 71597 792607
rect 71653 792551 71739 792607
rect 71795 792551 71881 792607
rect 71937 792551 72023 792607
rect 72079 792551 72165 792607
rect 72221 792551 72307 792607
rect 72363 792551 72449 792607
rect 72505 792551 72591 792607
rect 72647 792551 72733 792607
rect 72789 792551 72875 792607
rect 72931 792551 73017 792607
rect 73073 792551 73159 792607
rect 73215 792551 73301 792607
rect 73357 792551 73416 792607
rect 70475 792513 73416 792551
rect 70000 792465 73416 792513
rect 70000 792445 71455 792465
rect 70000 792389 70047 792445
rect 70103 792389 70171 792445
rect 70227 792389 70295 792445
rect 70351 792389 70419 792445
rect 70475 792409 71455 792445
rect 71511 792409 71597 792465
rect 71653 792409 71739 792465
rect 71795 792409 71881 792465
rect 71937 792409 72023 792465
rect 72079 792409 72165 792465
rect 72221 792409 72307 792465
rect 72363 792409 72449 792465
rect 72505 792409 72591 792465
rect 72647 792409 72733 792465
rect 72789 792409 72875 792465
rect 72931 792409 73017 792465
rect 73073 792409 73159 792465
rect 73215 792409 73301 792465
rect 73357 792409 73416 792465
rect 70475 792389 73416 792409
rect 70000 792323 73416 792389
rect 70000 792321 71455 792323
rect 70000 792265 70047 792321
rect 70103 792265 70171 792321
rect 70227 792265 70295 792321
rect 70351 792265 70419 792321
rect 70475 792267 71455 792321
rect 71511 792267 71597 792323
rect 71653 792267 71739 792323
rect 71795 792267 71881 792323
rect 71937 792267 72023 792323
rect 72079 792267 72165 792323
rect 72221 792267 72307 792323
rect 72363 792267 72449 792323
rect 72505 792267 72591 792323
rect 72647 792267 72733 792323
rect 72789 792267 72875 792323
rect 72931 792267 73017 792323
rect 73073 792267 73159 792323
rect 73215 792267 73301 792323
rect 73357 792267 73416 792323
rect 70475 792265 73416 792267
rect 70000 792198 73416 792265
rect 70000 791811 73416 791878
rect 70000 791755 70047 791811
rect 70103 791755 70171 791811
rect 70227 791755 70295 791811
rect 70351 791755 70419 791811
rect 70475 791799 73416 791811
rect 70475 791755 71455 791799
rect 70000 791743 71455 791755
rect 71511 791743 71597 791799
rect 71653 791743 71739 791799
rect 71795 791743 71881 791799
rect 71937 791743 72023 791799
rect 72079 791743 72165 791799
rect 72221 791743 72307 791799
rect 72363 791743 72449 791799
rect 72505 791743 72591 791799
rect 72647 791743 72733 791799
rect 72789 791743 72875 791799
rect 72931 791743 73017 791799
rect 73073 791743 73159 791799
rect 73215 791743 73301 791799
rect 73357 791743 73416 791799
rect 70000 791687 73416 791743
rect 70000 791631 70047 791687
rect 70103 791631 70171 791687
rect 70227 791631 70295 791687
rect 70351 791631 70419 791687
rect 70475 791657 73416 791687
rect 70475 791631 71455 791657
rect 70000 791601 71455 791631
rect 71511 791601 71597 791657
rect 71653 791601 71739 791657
rect 71795 791601 71881 791657
rect 71937 791601 72023 791657
rect 72079 791601 72165 791657
rect 72221 791601 72307 791657
rect 72363 791601 72449 791657
rect 72505 791601 72591 791657
rect 72647 791601 72733 791657
rect 72789 791601 72875 791657
rect 72931 791601 73017 791657
rect 73073 791601 73159 791657
rect 73215 791601 73301 791657
rect 73357 791601 73416 791657
rect 70000 791563 73416 791601
rect 70000 791507 70047 791563
rect 70103 791507 70171 791563
rect 70227 791507 70295 791563
rect 70351 791507 70419 791563
rect 70475 791515 73416 791563
rect 70475 791507 71455 791515
rect 70000 791459 71455 791507
rect 71511 791459 71597 791515
rect 71653 791459 71739 791515
rect 71795 791459 71881 791515
rect 71937 791459 72023 791515
rect 72079 791459 72165 791515
rect 72221 791459 72307 791515
rect 72363 791459 72449 791515
rect 72505 791459 72591 791515
rect 72647 791459 72733 791515
rect 72789 791459 72875 791515
rect 72931 791459 73017 791515
rect 73073 791459 73159 791515
rect 73215 791459 73301 791515
rect 73357 791459 73416 791515
rect 70000 791439 73416 791459
rect 70000 791383 70047 791439
rect 70103 791383 70171 791439
rect 70227 791383 70295 791439
rect 70351 791383 70419 791439
rect 70475 791383 73416 791439
rect 70000 791373 73416 791383
rect 70000 791317 71455 791373
rect 71511 791317 71597 791373
rect 71653 791317 71739 791373
rect 71795 791317 71881 791373
rect 71937 791317 72023 791373
rect 72079 791317 72165 791373
rect 72221 791317 72307 791373
rect 72363 791317 72449 791373
rect 72505 791317 72591 791373
rect 72647 791317 72733 791373
rect 72789 791317 72875 791373
rect 72931 791317 73017 791373
rect 73073 791317 73159 791373
rect 73215 791317 73301 791373
rect 73357 791317 73416 791373
rect 70000 791315 73416 791317
rect 70000 791259 70047 791315
rect 70103 791259 70171 791315
rect 70227 791259 70295 791315
rect 70351 791259 70419 791315
rect 70475 791259 73416 791315
rect 70000 791231 73416 791259
rect 70000 791191 71455 791231
rect 70000 791135 70047 791191
rect 70103 791135 70171 791191
rect 70227 791135 70295 791191
rect 70351 791135 70419 791191
rect 70475 791175 71455 791191
rect 71511 791175 71597 791231
rect 71653 791175 71739 791231
rect 71795 791175 71881 791231
rect 71937 791175 72023 791231
rect 72079 791175 72165 791231
rect 72221 791175 72307 791231
rect 72363 791175 72449 791231
rect 72505 791175 72591 791231
rect 72647 791175 72733 791231
rect 72789 791175 72875 791231
rect 72931 791175 73017 791231
rect 73073 791175 73159 791231
rect 73215 791175 73301 791231
rect 73357 791175 73416 791231
rect 70475 791135 73416 791175
rect 70000 791089 73416 791135
rect 70000 791067 71455 791089
rect 70000 791011 70047 791067
rect 70103 791011 70171 791067
rect 70227 791011 70295 791067
rect 70351 791011 70419 791067
rect 70475 791033 71455 791067
rect 71511 791033 71597 791089
rect 71653 791033 71739 791089
rect 71795 791033 71881 791089
rect 71937 791033 72023 791089
rect 72079 791033 72165 791089
rect 72221 791033 72307 791089
rect 72363 791033 72449 791089
rect 72505 791033 72591 791089
rect 72647 791033 72733 791089
rect 72789 791033 72875 791089
rect 72931 791033 73017 791089
rect 73073 791033 73159 791089
rect 73215 791033 73301 791089
rect 73357 791033 73416 791089
rect 70475 791011 73416 791033
rect 70000 790947 73416 791011
rect 70000 790943 71455 790947
rect 70000 790887 70047 790943
rect 70103 790887 70171 790943
rect 70227 790887 70295 790943
rect 70351 790887 70419 790943
rect 70475 790891 71455 790943
rect 71511 790891 71597 790947
rect 71653 790891 71739 790947
rect 71795 790891 71881 790947
rect 71937 790891 72023 790947
rect 72079 790891 72165 790947
rect 72221 790891 72307 790947
rect 72363 790891 72449 790947
rect 72505 790891 72591 790947
rect 72647 790891 72733 790947
rect 72789 790891 72875 790947
rect 72931 790891 73017 790947
rect 73073 790891 73159 790947
rect 73215 790891 73301 790947
rect 73357 790891 73416 790947
rect 70475 790887 73416 790891
rect 70000 790819 73416 790887
rect 70000 790763 70047 790819
rect 70103 790763 70171 790819
rect 70227 790763 70295 790819
rect 70351 790763 70419 790819
rect 70475 790805 73416 790819
rect 70475 790763 71455 790805
rect 70000 790749 71455 790763
rect 71511 790749 71597 790805
rect 71653 790749 71739 790805
rect 71795 790749 71881 790805
rect 71937 790749 72023 790805
rect 72079 790749 72165 790805
rect 72221 790749 72307 790805
rect 72363 790749 72449 790805
rect 72505 790749 72591 790805
rect 72647 790749 72733 790805
rect 72789 790749 72875 790805
rect 72931 790749 73017 790805
rect 73073 790749 73159 790805
rect 73215 790749 73301 790805
rect 73357 790749 73416 790805
rect 70000 790695 73416 790749
rect 70000 790639 70047 790695
rect 70103 790639 70171 790695
rect 70227 790639 70295 790695
rect 70351 790639 70419 790695
rect 70475 790663 73416 790695
rect 70475 790639 71455 790663
rect 70000 790607 71455 790639
rect 71511 790607 71597 790663
rect 71653 790607 71739 790663
rect 71795 790607 71881 790663
rect 71937 790607 72023 790663
rect 72079 790607 72165 790663
rect 72221 790607 72307 790663
rect 72363 790607 72449 790663
rect 72505 790607 72591 790663
rect 72647 790607 72733 790663
rect 72789 790607 72875 790663
rect 72931 790607 73017 790663
rect 73073 790607 73159 790663
rect 73215 790607 73301 790663
rect 73357 790607 73416 790663
rect 70000 790571 73416 790607
rect 70000 790515 70047 790571
rect 70103 790515 70171 790571
rect 70227 790515 70295 790571
rect 70351 790515 70419 790571
rect 70475 790521 73416 790571
rect 70475 790515 71455 790521
rect 70000 790465 71455 790515
rect 71511 790465 71597 790521
rect 71653 790465 71739 790521
rect 71795 790465 71881 790521
rect 71937 790465 72023 790521
rect 72079 790465 72165 790521
rect 72221 790465 72307 790521
rect 72363 790465 72449 790521
rect 72505 790465 72591 790521
rect 72647 790465 72733 790521
rect 72789 790465 72875 790521
rect 72931 790465 73017 790521
rect 73073 790465 73159 790521
rect 73215 790465 73301 790521
rect 73357 790465 73416 790521
rect 70000 790447 73416 790465
rect 70000 790391 70047 790447
rect 70103 790391 70171 790447
rect 70227 790391 70295 790447
rect 70351 790391 70419 790447
rect 70475 790391 73416 790447
rect 70000 790379 73416 790391
rect 70000 790323 71455 790379
rect 71511 790323 71597 790379
rect 71653 790323 71739 790379
rect 71795 790323 71881 790379
rect 71937 790323 72023 790379
rect 72079 790323 72165 790379
rect 72221 790323 72307 790379
rect 72363 790323 72449 790379
rect 72505 790323 72591 790379
rect 72647 790323 72733 790379
rect 72789 790323 72875 790379
rect 72931 790323 73017 790379
rect 73073 790323 73159 790379
rect 73215 790323 73301 790379
rect 73357 790323 73416 790379
rect 70000 790267 70047 790323
rect 70103 790267 70171 790323
rect 70227 790267 70295 790323
rect 70351 790267 70419 790323
rect 70475 790267 73416 790323
rect 70000 790237 73416 790267
rect 70000 790199 71455 790237
rect 70000 790143 70047 790199
rect 70103 790143 70171 790199
rect 70227 790143 70295 790199
rect 70351 790143 70419 790199
rect 70475 790181 71455 790199
rect 71511 790181 71597 790237
rect 71653 790181 71739 790237
rect 71795 790181 71881 790237
rect 71937 790181 72023 790237
rect 72079 790181 72165 790237
rect 72221 790181 72307 790237
rect 72363 790181 72449 790237
rect 72505 790181 72591 790237
rect 72647 790181 72733 790237
rect 72789 790181 72875 790237
rect 72931 790181 73017 790237
rect 73073 790181 73159 790237
rect 73215 790181 73301 790237
rect 73357 790181 73416 790237
rect 70475 790143 73416 790181
rect 70000 790095 73416 790143
rect 70000 790075 71455 790095
rect 70000 790019 70047 790075
rect 70103 790019 70171 790075
rect 70227 790019 70295 790075
rect 70351 790019 70419 790075
rect 70475 790039 71455 790075
rect 71511 790039 71597 790095
rect 71653 790039 71739 790095
rect 71795 790039 71881 790095
rect 71937 790039 72023 790095
rect 72079 790039 72165 790095
rect 72221 790039 72307 790095
rect 72363 790039 72449 790095
rect 72505 790039 72591 790095
rect 72647 790039 72733 790095
rect 72789 790039 72875 790095
rect 72931 790039 73017 790095
rect 73073 790039 73159 790095
rect 73215 790039 73301 790095
rect 73357 790039 73416 790095
rect 70475 790019 73416 790039
rect 70000 789953 73416 790019
rect 70000 789951 71455 789953
rect 70000 789895 70047 789951
rect 70103 789895 70171 789951
rect 70227 789895 70295 789951
rect 70351 789895 70419 789951
rect 70475 789897 71455 789951
rect 71511 789897 71597 789953
rect 71653 789897 71739 789953
rect 71795 789897 71881 789953
rect 71937 789897 72023 789953
rect 72079 789897 72165 789953
rect 72221 789897 72307 789953
rect 72363 789897 72449 789953
rect 72505 789897 72591 789953
rect 72647 789897 72733 789953
rect 72789 789897 72875 789953
rect 72931 789897 73017 789953
rect 73073 789897 73159 789953
rect 73215 789897 73301 789953
rect 73357 789897 73416 789953
rect 70475 789895 73416 789897
rect 70000 789828 73416 789895
rect 699992 791687 706000 791728
rect 699992 791666 705525 791687
rect 699992 791610 700040 791666
rect 700096 791610 700182 791666
rect 700238 791610 700324 791666
rect 700380 791610 700466 791666
rect 700522 791610 700608 791666
rect 700664 791610 700750 791666
rect 700806 791610 700892 791666
rect 700948 791610 701034 791666
rect 701090 791610 701176 791666
rect 701232 791610 701318 791666
rect 701374 791610 701460 791666
rect 701516 791610 701602 791666
rect 701658 791610 701744 791666
rect 701800 791610 701886 791666
rect 701942 791631 705525 791666
rect 705581 791631 705649 791687
rect 705705 791631 705773 791687
rect 705829 791631 705897 791687
rect 705953 791631 706000 791687
rect 701942 791610 706000 791631
rect 699992 791563 706000 791610
rect 699992 791524 705525 791563
rect 699992 791468 700040 791524
rect 700096 791468 700182 791524
rect 700238 791468 700324 791524
rect 700380 791468 700466 791524
rect 700522 791468 700608 791524
rect 700664 791468 700750 791524
rect 700806 791468 700892 791524
rect 700948 791468 701034 791524
rect 701090 791468 701176 791524
rect 701232 791468 701318 791524
rect 701374 791468 701460 791524
rect 701516 791468 701602 791524
rect 701658 791468 701744 791524
rect 701800 791468 701886 791524
rect 701942 791507 705525 791524
rect 705581 791507 705649 791563
rect 705705 791507 705773 791563
rect 705829 791507 705897 791563
rect 705953 791507 706000 791563
rect 701942 791468 706000 791507
rect 699992 791439 706000 791468
rect 699992 791383 705525 791439
rect 705581 791383 705649 791439
rect 705705 791383 705773 791439
rect 705829 791383 705897 791439
rect 705953 791383 706000 791439
rect 699992 791382 706000 791383
rect 699992 791326 700040 791382
rect 700096 791326 700182 791382
rect 700238 791326 700324 791382
rect 700380 791326 700466 791382
rect 700522 791326 700608 791382
rect 700664 791326 700750 791382
rect 700806 791326 700892 791382
rect 700948 791326 701034 791382
rect 701090 791326 701176 791382
rect 701232 791326 701318 791382
rect 701374 791326 701460 791382
rect 701516 791326 701602 791382
rect 701658 791326 701744 791382
rect 701800 791326 701886 791382
rect 701942 791326 706000 791382
rect 699992 791315 706000 791326
rect 699992 791259 705525 791315
rect 705581 791259 705649 791315
rect 705705 791259 705773 791315
rect 705829 791259 705897 791315
rect 705953 791259 706000 791315
rect 699992 791240 706000 791259
rect 699992 791184 700040 791240
rect 700096 791184 700182 791240
rect 700238 791184 700324 791240
rect 700380 791184 700466 791240
rect 700522 791184 700608 791240
rect 700664 791184 700750 791240
rect 700806 791184 700892 791240
rect 700948 791184 701034 791240
rect 701090 791184 701176 791240
rect 701232 791184 701318 791240
rect 701374 791184 701460 791240
rect 701516 791184 701602 791240
rect 701658 791184 701744 791240
rect 701800 791184 701886 791240
rect 701942 791191 706000 791240
rect 701942 791184 705525 791191
rect 699992 791135 705525 791184
rect 705581 791135 705649 791191
rect 705705 791135 705773 791191
rect 705829 791135 705897 791191
rect 705953 791135 706000 791191
rect 699992 791098 706000 791135
rect 699992 791042 700040 791098
rect 700096 791042 700182 791098
rect 700238 791042 700324 791098
rect 700380 791042 700466 791098
rect 700522 791042 700608 791098
rect 700664 791042 700750 791098
rect 700806 791042 700892 791098
rect 700948 791042 701034 791098
rect 701090 791042 701176 791098
rect 701232 791042 701318 791098
rect 701374 791042 701460 791098
rect 701516 791042 701602 791098
rect 701658 791042 701744 791098
rect 701800 791042 701886 791098
rect 701942 791067 706000 791098
rect 701942 791042 705525 791067
rect 699992 791011 705525 791042
rect 705581 791011 705649 791067
rect 705705 791011 705773 791067
rect 705829 791011 705897 791067
rect 705953 791011 706000 791067
rect 699992 790956 706000 791011
rect 699992 790900 700040 790956
rect 700096 790900 700182 790956
rect 700238 790900 700324 790956
rect 700380 790900 700466 790956
rect 700522 790900 700608 790956
rect 700664 790900 700750 790956
rect 700806 790900 700892 790956
rect 700948 790900 701034 790956
rect 701090 790900 701176 790956
rect 701232 790900 701318 790956
rect 701374 790900 701460 790956
rect 701516 790900 701602 790956
rect 701658 790900 701744 790956
rect 701800 790900 701886 790956
rect 701942 790943 706000 790956
rect 701942 790900 705525 790943
rect 699992 790887 705525 790900
rect 705581 790887 705649 790943
rect 705705 790887 705773 790943
rect 705829 790887 705897 790943
rect 705953 790887 706000 790943
rect 699992 790819 706000 790887
rect 699992 790814 705525 790819
rect 699992 790758 700040 790814
rect 700096 790758 700182 790814
rect 700238 790758 700324 790814
rect 700380 790758 700466 790814
rect 700522 790758 700608 790814
rect 700664 790758 700750 790814
rect 700806 790758 700892 790814
rect 700948 790758 701034 790814
rect 701090 790758 701176 790814
rect 701232 790758 701318 790814
rect 701374 790758 701460 790814
rect 701516 790758 701602 790814
rect 701658 790758 701744 790814
rect 701800 790758 701886 790814
rect 701942 790763 705525 790814
rect 705581 790763 705649 790819
rect 705705 790763 705773 790819
rect 705829 790763 705897 790819
rect 705953 790763 706000 790819
rect 701942 790758 706000 790763
rect 699992 790695 706000 790758
rect 699992 790672 705525 790695
rect 699992 790616 700040 790672
rect 700096 790616 700182 790672
rect 700238 790616 700324 790672
rect 700380 790616 700466 790672
rect 700522 790616 700608 790672
rect 700664 790616 700750 790672
rect 700806 790616 700892 790672
rect 700948 790616 701034 790672
rect 701090 790616 701176 790672
rect 701232 790616 701318 790672
rect 701374 790616 701460 790672
rect 701516 790616 701602 790672
rect 701658 790616 701744 790672
rect 701800 790616 701886 790672
rect 701942 790639 705525 790672
rect 705581 790639 705649 790695
rect 705705 790639 705773 790695
rect 705829 790639 705897 790695
rect 705953 790639 706000 790695
rect 701942 790616 706000 790639
rect 699992 790571 706000 790616
rect 699992 790530 705525 790571
rect 699992 790474 700040 790530
rect 700096 790474 700182 790530
rect 700238 790474 700324 790530
rect 700380 790474 700466 790530
rect 700522 790474 700608 790530
rect 700664 790474 700750 790530
rect 700806 790474 700892 790530
rect 700948 790474 701034 790530
rect 701090 790474 701176 790530
rect 701232 790474 701318 790530
rect 701374 790474 701460 790530
rect 701516 790474 701602 790530
rect 701658 790474 701744 790530
rect 701800 790474 701886 790530
rect 701942 790515 705525 790530
rect 705581 790515 705649 790571
rect 705705 790515 705773 790571
rect 705829 790515 705897 790571
rect 705953 790515 706000 790571
rect 701942 790474 706000 790515
rect 699992 790447 706000 790474
rect 699992 790391 705525 790447
rect 705581 790391 705649 790447
rect 705705 790391 705773 790447
rect 705829 790391 705897 790447
rect 705953 790391 706000 790447
rect 699992 790388 706000 790391
rect 699992 790332 700040 790388
rect 700096 790332 700182 790388
rect 700238 790332 700324 790388
rect 700380 790332 700466 790388
rect 700522 790332 700608 790388
rect 700664 790332 700750 790388
rect 700806 790332 700892 790388
rect 700948 790332 701034 790388
rect 701090 790332 701176 790388
rect 701232 790332 701318 790388
rect 701374 790332 701460 790388
rect 701516 790332 701602 790388
rect 701658 790332 701744 790388
rect 701800 790332 701886 790388
rect 701942 790332 706000 790388
rect 699992 790323 706000 790332
rect 699992 790267 705525 790323
rect 705581 790267 705649 790323
rect 705705 790267 705773 790323
rect 705829 790267 705897 790323
rect 705953 790267 706000 790323
rect 699992 790246 706000 790267
rect 699992 790190 700040 790246
rect 700096 790190 700182 790246
rect 700238 790190 700324 790246
rect 700380 790190 700466 790246
rect 700522 790190 700608 790246
rect 700664 790190 700750 790246
rect 700806 790190 700892 790246
rect 700948 790190 701034 790246
rect 701090 790190 701176 790246
rect 701232 790190 701318 790246
rect 701374 790190 701460 790246
rect 701516 790190 701602 790246
rect 701658 790190 701744 790246
rect 701800 790190 701886 790246
rect 701942 790199 706000 790246
rect 701942 790190 705525 790199
rect 699992 790143 705525 790190
rect 705581 790143 705649 790199
rect 705705 790143 705773 790199
rect 705829 790143 705897 790199
rect 705953 790143 706000 790199
rect 699992 790104 706000 790143
rect 699992 790048 700040 790104
rect 700096 790048 700182 790104
rect 700238 790048 700324 790104
rect 700380 790048 700466 790104
rect 700522 790048 700608 790104
rect 700664 790048 700750 790104
rect 700806 790048 700892 790104
rect 700948 790048 701034 790104
rect 701090 790048 701176 790104
rect 701232 790048 701318 790104
rect 701374 790048 701460 790104
rect 701516 790048 701602 790104
rect 701658 790048 701744 790104
rect 701800 790048 701886 790104
rect 701942 790075 706000 790104
rect 701942 790048 705525 790075
rect 699992 790019 705525 790048
rect 705581 790019 705649 790075
rect 705705 790019 705773 790075
rect 705829 790019 705897 790075
rect 705953 790019 706000 790075
rect 699992 789962 706000 790019
rect 699992 789906 700040 789962
rect 700096 789906 700182 789962
rect 700238 789906 700324 789962
rect 700380 789906 700466 789962
rect 700522 789906 700608 789962
rect 700664 789906 700750 789962
rect 700806 789906 700892 789962
rect 700948 789906 701034 789962
rect 701090 789906 701176 789962
rect 701232 789906 701318 789962
rect 701374 789906 701460 789962
rect 701516 789906 701602 789962
rect 701658 789906 701744 789962
rect 701800 789906 701886 789962
rect 701942 789951 706000 789962
rect 701942 789906 705525 789951
rect 699992 789895 705525 789906
rect 705581 789895 705649 789951
rect 705705 789895 705773 789951
rect 705829 789895 705897 789951
rect 705953 789895 706000 789951
rect 699992 789828 706000 789895
rect 699992 789181 706000 789248
rect 699992 789179 705525 789181
rect 70000 789105 73416 789172
rect 70000 789049 70047 789105
rect 70103 789049 70171 789105
rect 70227 789049 70295 789105
rect 70351 789049 70419 789105
rect 70475 789093 73416 789105
rect 70475 789049 71455 789093
rect 70000 789037 71455 789049
rect 71511 789037 71597 789093
rect 71653 789037 71739 789093
rect 71795 789037 71881 789093
rect 71937 789037 72023 789093
rect 72079 789037 72165 789093
rect 72221 789037 72307 789093
rect 72363 789037 72449 789093
rect 72505 789037 72591 789093
rect 72647 789037 72733 789093
rect 72789 789037 72875 789093
rect 72931 789037 73017 789093
rect 73073 789037 73159 789093
rect 73215 789037 73301 789093
rect 73357 789037 73416 789093
rect 70000 788981 73416 789037
rect 70000 788925 70047 788981
rect 70103 788925 70171 788981
rect 70227 788925 70295 788981
rect 70351 788925 70419 788981
rect 70475 788951 73416 788981
rect 70475 788925 71455 788951
rect 70000 788895 71455 788925
rect 71511 788895 71597 788951
rect 71653 788895 71739 788951
rect 71795 788895 71881 788951
rect 71937 788895 72023 788951
rect 72079 788895 72165 788951
rect 72221 788895 72307 788951
rect 72363 788895 72449 788951
rect 72505 788895 72591 788951
rect 72647 788895 72733 788951
rect 72789 788895 72875 788951
rect 72931 788895 73017 788951
rect 73073 788895 73159 788951
rect 73215 788895 73301 788951
rect 73357 788895 73416 788951
rect 70000 788857 73416 788895
rect 70000 788801 70047 788857
rect 70103 788801 70171 788857
rect 70227 788801 70295 788857
rect 70351 788801 70419 788857
rect 70475 788809 73416 788857
rect 70475 788801 71455 788809
rect 70000 788753 71455 788801
rect 71511 788753 71597 788809
rect 71653 788753 71739 788809
rect 71795 788753 71881 788809
rect 71937 788753 72023 788809
rect 72079 788753 72165 788809
rect 72221 788753 72307 788809
rect 72363 788753 72449 788809
rect 72505 788753 72591 788809
rect 72647 788753 72733 788809
rect 72789 788753 72875 788809
rect 72931 788753 73017 788809
rect 73073 788753 73159 788809
rect 73215 788753 73301 788809
rect 73357 788753 73416 788809
rect 70000 788733 73416 788753
rect 70000 788677 70047 788733
rect 70103 788677 70171 788733
rect 70227 788677 70295 788733
rect 70351 788677 70419 788733
rect 70475 788677 73416 788733
rect 70000 788667 73416 788677
rect 70000 788611 71455 788667
rect 71511 788611 71597 788667
rect 71653 788611 71739 788667
rect 71795 788611 71881 788667
rect 71937 788611 72023 788667
rect 72079 788611 72165 788667
rect 72221 788611 72307 788667
rect 72363 788611 72449 788667
rect 72505 788611 72591 788667
rect 72647 788611 72733 788667
rect 72789 788611 72875 788667
rect 72931 788611 73017 788667
rect 73073 788611 73159 788667
rect 73215 788611 73301 788667
rect 73357 788611 73416 788667
rect 70000 788609 73416 788611
rect 70000 788553 70047 788609
rect 70103 788553 70171 788609
rect 70227 788553 70295 788609
rect 70351 788553 70419 788609
rect 70475 788553 73416 788609
rect 70000 788525 73416 788553
rect 70000 788485 71455 788525
rect 70000 788429 70047 788485
rect 70103 788429 70171 788485
rect 70227 788429 70295 788485
rect 70351 788429 70419 788485
rect 70475 788469 71455 788485
rect 71511 788469 71597 788525
rect 71653 788469 71739 788525
rect 71795 788469 71881 788525
rect 71937 788469 72023 788525
rect 72079 788469 72165 788525
rect 72221 788469 72307 788525
rect 72363 788469 72449 788525
rect 72505 788469 72591 788525
rect 72647 788469 72733 788525
rect 72789 788469 72875 788525
rect 72931 788469 73017 788525
rect 73073 788469 73159 788525
rect 73215 788469 73301 788525
rect 73357 788469 73416 788525
rect 70475 788429 73416 788469
rect 70000 788383 73416 788429
rect 70000 788361 71455 788383
rect 70000 788305 70047 788361
rect 70103 788305 70171 788361
rect 70227 788305 70295 788361
rect 70351 788305 70419 788361
rect 70475 788327 71455 788361
rect 71511 788327 71597 788383
rect 71653 788327 71739 788383
rect 71795 788327 71881 788383
rect 71937 788327 72023 788383
rect 72079 788327 72165 788383
rect 72221 788327 72307 788383
rect 72363 788327 72449 788383
rect 72505 788327 72591 788383
rect 72647 788327 72733 788383
rect 72789 788327 72875 788383
rect 72931 788327 73017 788383
rect 73073 788327 73159 788383
rect 73215 788327 73301 788383
rect 73357 788327 73416 788383
rect 70475 788305 73416 788327
rect 70000 788241 73416 788305
rect 70000 788237 71455 788241
rect 70000 788181 70047 788237
rect 70103 788181 70171 788237
rect 70227 788181 70295 788237
rect 70351 788181 70419 788237
rect 70475 788185 71455 788237
rect 71511 788185 71597 788241
rect 71653 788185 71739 788241
rect 71795 788185 71881 788241
rect 71937 788185 72023 788241
rect 72079 788185 72165 788241
rect 72221 788185 72307 788241
rect 72363 788185 72449 788241
rect 72505 788185 72591 788241
rect 72647 788185 72733 788241
rect 72789 788185 72875 788241
rect 72931 788185 73017 788241
rect 73073 788185 73159 788241
rect 73215 788185 73301 788241
rect 73357 788185 73416 788241
rect 70475 788181 73416 788185
rect 70000 788113 73416 788181
rect 70000 788057 70047 788113
rect 70103 788057 70171 788113
rect 70227 788057 70295 788113
rect 70351 788057 70419 788113
rect 70475 788099 73416 788113
rect 70475 788057 71455 788099
rect 70000 788043 71455 788057
rect 71511 788043 71597 788099
rect 71653 788043 71739 788099
rect 71795 788043 71881 788099
rect 71937 788043 72023 788099
rect 72079 788043 72165 788099
rect 72221 788043 72307 788099
rect 72363 788043 72449 788099
rect 72505 788043 72591 788099
rect 72647 788043 72733 788099
rect 72789 788043 72875 788099
rect 72931 788043 73017 788099
rect 73073 788043 73159 788099
rect 73215 788043 73301 788099
rect 73357 788043 73416 788099
rect 70000 787989 73416 788043
rect 70000 787933 70047 787989
rect 70103 787933 70171 787989
rect 70227 787933 70295 787989
rect 70351 787933 70419 787989
rect 70475 787957 73416 787989
rect 70475 787933 71455 787957
rect 70000 787901 71455 787933
rect 71511 787901 71597 787957
rect 71653 787901 71739 787957
rect 71795 787901 71881 787957
rect 71937 787901 72023 787957
rect 72079 787901 72165 787957
rect 72221 787901 72307 787957
rect 72363 787901 72449 787957
rect 72505 787901 72591 787957
rect 72647 787901 72733 787957
rect 72789 787901 72875 787957
rect 72931 787901 73017 787957
rect 73073 787901 73159 787957
rect 73215 787901 73301 787957
rect 73357 787901 73416 787957
rect 70000 787865 73416 787901
rect 70000 787809 70047 787865
rect 70103 787809 70171 787865
rect 70227 787809 70295 787865
rect 70351 787809 70419 787865
rect 70475 787815 73416 787865
rect 70475 787809 71455 787815
rect 70000 787759 71455 787809
rect 71511 787759 71597 787815
rect 71653 787759 71739 787815
rect 71795 787759 71881 787815
rect 71937 787759 72023 787815
rect 72079 787759 72165 787815
rect 72221 787759 72307 787815
rect 72363 787759 72449 787815
rect 72505 787759 72591 787815
rect 72647 787759 72733 787815
rect 72789 787759 72875 787815
rect 72931 787759 73017 787815
rect 73073 787759 73159 787815
rect 73215 787759 73301 787815
rect 73357 787759 73416 787815
rect 70000 787741 73416 787759
rect 70000 787685 70047 787741
rect 70103 787685 70171 787741
rect 70227 787685 70295 787741
rect 70351 787685 70419 787741
rect 70475 787685 73416 787741
rect 70000 787673 73416 787685
rect 70000 787617 71455 787673
rect 71511 787617 71597 787673
rect 71653 787617 71739 787673
rect 71795 787617 71881 787673
rect 71937 787617 72023 787673
rect 72079 787617 72165 787673
rect 72221 787617 72307 787673
rect 72363 787617 72449 787673
rect 72505 787617 72591 787673
rect 72647 787617 72733 787673
rect 72789 787617 72875 787673
rect 72931 787617 73017 787673
rect 73073 787617 73159 787673
rect 73215 787617 73301 787673
rect 73357 787617 73416 787673
rect 70000 787561 70047 787617
rect 70103 787561 70171 787617
rect 70227 787561 70295 787617
rect 70351 787561 70419 787617
rect 70475 787561 73416 787617
rect 70000 787531 73416 787561
rect 70000 787493 71455 787531
rect 70000 787437 70047 787493
rect 70103 787437 70171 787493
rect 70227 787437 70295 787493
rect 70351 787437 70419 787493
rect 70475 787475 71455 787493
rect 71511 787475 71597 787531
rect 71653 787475 71739 787531
rect 71795 787475 71881 787531
rect 71937 787475 72023 787531
rect 72079 787475 72165 787531
rect 72221 787475 72307 787531
rect 72363 787475 72449 787531
rect 72505 787475 72591 787531
rect 72647 787475 72733 787531
rect 72789 787475 72875 787531
rect 72931 787475 73017 787531
rect 73073 787475 73159 787531
rect 73215 787475 73301 787531
rect 73357 787475 73416 787531
rect 70475 787437 73416 787475
rect 70000 787389 73416 787437
rect 70000 787369 71455 787389
rect 70000 787313 70047 787369
rect 70103 787313 70171 787369
rect 70227 787313 70295 787369
rect 70351 787313 70419 787369
rect 70475 787333 71455 787369
rect 71511 787333 71597 787389
rect 71653 787333 71739 787389
rect 71795 787333 71881 787389
rect 71937 787333 72023 787389
rect 72079 787333 72165 787389
rect 72221 787333 72307 787389
rect 72363 787333 72449 787389
rect 72505 787333 72591 787389
rect 72647 787333 72733 787389
rect 72789 787333 72875 787389
rect 72931 787333 73017 787389
rect 73073 787333 73159 787389
rect 73215 787333 73301 787389
rect 73357 787333 73416 787389
rect 70475 787313 73416 787333
rect 70000 787247 73416 787313
rect 70000 787245 71455 787247
rect 70000 787189 70047 787245
rect 70103 787189 70171 787245
rect 70227 787189 70295 787245
rect 70351 787189 70419 787245
rect 70475 787191 71455 787245
rect 71511 787191 71597 787247
rect 71653 787191 71739 787247
rect 71795 787191 71881 787247
rect 71937 787191 72023 787247
rect 72079 787191 72165 787247
rect 72221 787191 72307 787247
rect 72363 787191 72449 787247
rect 72505 787191 72591 787247
rect 72647 787191 72733 787247
rect 72789 787191 72875 787247
rect 72931 787191 73017 787247
rect 73073 787191 73159 787247
rect 73215 787191 73301 787247
rect 73357 787191 73416 787247
rect 699992 789123 700051 789179
rect 700107 789123 700193 789179
rect 700249 789123 700335 789179
rect 700391 789123 700477 789179
rect 700533 789123 700619 789179
rect 700675 789123 700761 789179
rect 700817 789123 700903 789179
rect 700959 789123 701045 789179
rect 701101 789123 701187 789179
rect 701243 789123 701329 789179
rect 701385 789123 701471 789179
rect 701527 789123 701613 789179
rect 701669 789123 701755 789179
rect 701811 789123 701897 789179
rect 701953 789125 705525 789179
rect 705581 789125 705649 789181
rect 705705 789125 705773 789181
rect 705829 789125 705897 789181
rect 705953 789125 706000 789181
rect 701953 789123 706000 789125
rect 699992 789057 706000 789123
rect 699992 789037 705525 789057
rect 699992 788981 700051 789037
rect 700107 788981 700193 789037
rect 700249 788981 700335 789037
rect 700391 788981 700477 789037
rect 700533 788981 700619 789037
rect 700675 788981 700761 789037
rect 700817 788981 700903 789037
rect 700959 788981 701045 789037
rect 701101 788981 701187 789037
rect 701243 788981 701329 789037
rect 701385 788981 701471 789037
rect 701527 788981 701613 789037
rect 701669 788981 701755 789037
rect 701811 788981 701897 789037
rect 701953 789001 705525 789037
rect 705581 789001 705649 789057
rect 705705 789001 705773 789057
rect 705829 789001 705897 789057
rect 705953 789001 706000 789057
rect 701953 788981 706000 789001
rect 699992 788933 706000 788981
rect 699992 788895 705525 788933
rect 699992 788839 700051 788895
rect 700107 788839 700193 788895
rect 700249 788839 700335 788895
rect 700391 788839 700477 788895
rect 700533 788839 700619 788895
rect 700675 788839 700761 788895
rect 700817 788839 700903 788895
rect 700959 788839 701045 788895
rect 701101 788839 701187 788895
rect 701243 788839 701329 788895
rect 701385 788839 701471 788895
rect 701527 788839 701613 788895
rect 701669 788839 701755 788895
rect 701811 788839 701897 788895
rect 701953 788877 705525 788895
rect 705581 788877 705649 788933
rect 705705 788877 705773 788933
rect 705829 788877 705897 788933
rect 705953 788877 706000 788933
rect 701953 788839 706000 788877
rect 699992 788809 706000 788839
rect 699992 788753 705525 788809
rect 705581 788753 705649 788809
rect 705705 788753 705773 788809
rect 705829 788753 705897 788809
rect 705953 788753 706000 788809
rect 699992 788697 700051 788753
rect 700107 788697 700193 788753
rect 700249 788697 700335 788753
rect 700391 788697 700477 788753
rect 700533 788697 700619 788753
rect 700675 788697 700761 788753
rect 700817 788697 700903 788753
rect 700959 788697 701045 788753
rect 701101 788697 701187 788753
rect 701243 788697 701329 788753
rect 701385 788697 701471 788753
rect 701527 788697 701613 788753
rect 701669 788697 701755 788753
rect 701811 788697 701897 788753
rect 701953 788697 706000 788753
rect 699992 788685 706000 788697
rect 699992 788629 705525 788685
rect 705581 788629 705649 788685
rect 705705 788629 705773 788685
rect 705829 788629 705897 788685
rect 705953 788629 706000 788685
rect 699992 788611 706000 788629
rect 699992 788555 700051 788611
rect 700107 788555 700193 788611
rect 700249 788555 700335 788611
rect 700391 788555 700477 788611
rect 700533 788555 700619 788611
rect 700675 788555 700761 788611
rect 700817 788555 700903 788611
rect 700959 788555 701045 788611
rect 701101 788555 701187 788611
rect 701243 788555 701329 788611
rect 701385 788555 701471 788611
rect 701527 788555 701613 788611
rect 701669 788555 701755 788611
rect 701811 788555 701897 788611
rect 701953 788561 706000 788611
rect 701953 788555 705525 788561
rect 699992 788505 705525 788555
rect 705581 788505 705649 788561
rect 705705 788505 705773 788561
rect 705829 788505 705897 788561
rect 705953 788505 706000 788561
rect 699992 788469 706000 788505
rect 699992 788413 700051 788469
rect 700107 788413 700193 788469
rect 700249 788413 700335 788469
rect 700391 788413 700477 788469
rect 700533 788413 700619 788469
rect 700675 788413 700761 788469
rect 700817 788413 700903 788469
rect 700959 788413 701045 788469
rect 701101 788413 701187 788469
rect 701243 788413 701329 788469
rect 701385 788413 701471 788469
rect 701527 788413 701613 788469
rect 701669 788413 701755 788469
rect 701811 788413 701897 788469
rect 701953 788437 706000 788469
rect 701953 788413 705525 788437
rect 699992 788381 705525 788413
rect 705581 788381 705649 788437
rect 705705 788381 705773 788437
rect 705829 788381 705897 788437
rect 705953 788381 706000 788437
rect 699992 788327 706000 788381
rect 699992 788271 700051 788327
rect 700107 788271 700193 788327
rect 700249 788271 700335 788327
rect 700391 788271 700477 788327
rect 700533 788271 700619 788327
rect 700675 788271 700761 788327
rect 700817 788271 700903 788327
rect 700959 788271 701045 788327
rect 701101 788271 701187 788327
rect 701243 788271 701329 788327
rect 701385 788271 701471 788327
rect 701527 788271 701613 788327
rect 701669 788271 701755 788327
rect 701811 788271 701897 788327
rect 701953 788313 706000 788327
rect 701953 788271 705525 788313
rect 699992 788257 705525 788271
rect 705581 788257 705649 788313
rect 705705 788257 705773 788313
rect 705829 788257 705897 788313
rect 705953 788257 706000 788313
rect 699992 788189 706000 788257
rect 699992 788185 705525 788189
rect 699992 788129 700051 788185
rect 700107 788129 700193 788185
rect 700249 788129 700335 788185
rect 700391 788129 700477 788185
rect 700533 788129 700619 788185
rect 700675 788129 700761 788185
rect 700817 788129 700903 788185
rect 700959 788129 701045 788185
rect 701101 788129 701187 788185
rect 701243 788129 701329 788185
rect 701385 788129 701471 788185
rect 701527 788129 701613 788185
rect 701669 788129 701755 788185
rect 701811 788129 701897 788185
rect 701953 788133 705525 788185
rect 705581 788133 705649 788189
rect 705705 788133 705773 788189
rect 705829 788133 705897 788189
rect 705953 788133 706000 788189
rect 701953 788129 706000 788133
rect 699992 788065 706000 788129
rect 699992 788043 705525 788065
rect 699992 787987 700051 788043
rect 700107 787987 700193 788043
rect 700249 787987 700335 788043
rect 700391 787987 700477 788043
rect 700533 787987 700619 788043
rect 700675 787987 700761 788043
rect 700817 787987 700903 788043
rect 700959 787987 701045 788043
rect 701101 787987 701187 788043
rect 701243 787987 701329 788043
rect 701385 787987 701471 788043
rect 701527 787987 701613 788043
rect 701669 787987 701755 788043
rect 701811 787987 701897 788043
rect 701953 788009 705525 788043
rect 705581 788009 705649 788065
rect 705705 788009 705773 788065
rect 705829 788009 705897 788065
rect 705953 788009 706000 788065
rect 701953 787987 706000 788009
rect 699992 787941 706000 787987
rect 699992 787901 705525 787941
rect 699992 787845 700051 787901
rect 700107 787845 700193 787901
rect 700249 787845 700335 787901
rect 700391 787845 700477 787901
rect 700533 787845 700619 787901
rect 700675 787845 700761 787901
rect 700817 787845 700903 787901
rect 700959 787845 701045 787901
rect 701101 787845 701187 787901
rect 701243 787845 701329 787901
rect 701385 787845 701471 787901
rect 701527 787845 701613 787901
rect 701669 787845 701755 787901
rect 701811 787845 701897 787901
rect 701953 787885 705525 787901
rect 705581 787885 705649 787941
rect 705705 787885 705773 787941
rect 705829 787885 705897 787941
rect 705953 787885 706000 787941
rect 701953 787845 706000 787885
rect 699992 787817 706000 787845
rect 699992 787761 705525 787817
rect 705581 787761 705649 787817
rect 705705 787761 705773 787817
rect 705829 787761 705897 787817
rect 705953 787761 706000 787817
rect 699992 787759 706000 787761
rect 699992 787703 700051 787759
rect 700107 787703 700193 787759
rect 700249 787703 700335 787759
rect 700391 787703 700477 787759
rect 700533 787703 700619 787759
rect 700675 787703 700761 787759
rect 700817 787703 700903 787759
rect 700959 787703 701045 787759
rect 701101 787703 701187 787759
rect 701243 787703 701329 787759
rect 701385 787703 701471 787759
rect 701527 787703 701613 787759
rect 701669 787703 701755 787759
rect 701811 787703 701897 787759
rect 701953 787703 706000 787759
rect 699992 787693 706000 787703
rect 699992 787637 705525 787693
rect 705581 787637 705649 787693
rect 705705 787637 705773 787693
rect 705829 787637 705897 787693
rect 705953 787637 706000 787693
rect 699992 787617 706000 787637
rect 699992 787561 700051 787617
rect 700107 787561 700193 787617
rect 700249 787561 700335 787617
rect 700391 787561 700477 787617
rect 700533 787561 700619 787617
rect 700675 787561 700761 787617
rect 700817 787561 700903 787617
rect 700959 787561 701045 787617
rect 701101 787561 701187 787617
rect 701243 787561 701329 787617
rect 701385 787561 701471 787617
rect 701527 787561 701613 787617
rect 701669 787561 701755 787617
rect 701811 787561 701897 787617
rect 701953 787569 706000 787617
rect 701953 787561 705525 787569
rect 699992 787513 705525 787561
rect 705581 787513 705649 787569
rect 705705 787513 705773 787569
rect 705829 787513 705897 787569
rect 705953 787513 706000 787569
rect 699992 787475 706000 787513
rect 699992 787419 700051 787475
rect 700107 787419 700193 787475
rect 700249 787419 700335 787475
rect 700391 787419 700477 787475
rect 700533 787419 700619 787475
rect 700675 787419 700761 787475
rect 700817 787419 700903 787475
rect 700959 787419 701045 787475
rect 701101 787419 701187 787475
rect 701243 787419 701329 787475
rect 701385 787419 701471 787475
rect 701527 787419 701613 787475
rect 701669 787419 701755 787475
rect 701811 787419 701897 787475
rect 701953 787445 706000 787475
rect 701953 787419 705525 787445
rect 699992 787389 705525 787419
rect 705581 787389 705649 787445
rect 705705 787389 705773 787445
rect 705829 787389 705897 787445
rect 705953 787389 706000 787445
rect 699992 787333 706000 787389
rect 699992 787277 700051 787333
rect 700107 787277 700193 787333
rect 700249 787277 700335 787333
rect 700391 787277 700477 787333
rect 700533 787277 700619 787333
rect 700675 787277 700761 787333
rect 700817 787277 700903 787333
rect 700959 787277 701045 787333
rect 701101 787277 701187 787333
rect 701243 787277 701329 787333
rect 701385 787277 701471 787333
rect 701527 787277 701613 787333
rect 701669 787277 701755 787333
rect 701811 787277 701897 787333
rect 701953 787321 706000 787333
rect 701953 787277 705525 787321
rect 699992 787265 705525 787277
rect 705581 787265 705649 787321
rect 705705 787265 705773 787321
rect 705829 787265 705897 787321
rect 705953 787265 706000 787321
rect 699992 787198 706000 787265
rect 70475 787189 73416 787191
rect 70000 787122 73416 787189
rect 699992 786811 706000 786878
rect 699992 786809 705525 786811
rect 70000 786735 73416 786802
rect 70000 786679 70047 786735
rect 70103 786679 70171 786735
rect 70227 786679 70295 786735
rect 70351 786679 70419 786735
rect 70475 786723 73416 786735
rect 70475 786679 71455 786723
rect 70000 786667 71455 786679
rect 71511 786667 71597 786723
rect 71653 786667 71739 786723
rect 71795 786667 71881 786723
rect 71937 786667 72023 786723
rect 72079 786667 72165 786723
rect 72221 786667 72307 786723
rect 72363 786667 72449 786723
rect 72505 786667 72591 786723
rect 72647 786667 72733 786723
rect 72789 786667 72875 786723
rect 72931 786667 73017 786723
rect 73073 786667 73159 786723
rect 73215 786667 73301 786723
rect 73357 786667 73416 786723
rect 70000 786611 73416 786667
rect 70000 786555 70047 786611
rect 70103 786555 70171 786611
rect 70227 786555 70295 786611
rect 70351 786555 70419 786611
rect 70475 786581 73416 786611
rect 70475 786555 71455 786581
rect 70000 786525 71455 786555
rect 71511 786525 71597 786581
rect 71653 786525 71739 786581
rect 71795 786525 71881 786581
rect 71937 786525 72023 786581
rect 72079 786525 72165 786581
rect 72221 786525 72307 786581
rect 72363 786525 72449 786581
rect 72505 786525 72591 786581
rect 72647 786525 72733 786581
rect 72789 786525 72875 786581
rect 72931 786525 73017 786581
rect 73073 786525 73159 786581
rect 73215 786525 73301 786581
rect 73357 786525 73416 786581
rect 70000 786487 73416 786525
rect 70000 786431 70047 786487
rect 70103 786431 70171 786487
rect 70227 786431 70295 786487
rect 70351 786431 70419 786487
rect 70475 786439 73416 786487
rect 70475 786431 71455 786439
rect 70000 786383 71455 786431
rect 71511 786383 71597 786439
rect 71653 786383 71739 786439
rect 71795 786383 71881 786439
rect 71937 786383 72023 786439
rect 72079 786383 72165 786439
rect 72221 786383 72307 786439
rect 72363 786383 72449 786439
rect 72505 786383 72591 786439
rect 72647 786383 72733 786439
rect 72789 786383 72875 786439
rect 72931 786383 73017 786439
rect 73073 786383 73159 786439
rect 73215 786383 73301 786439
rect 73357 786383 73416 786439
rect 70000 786363 73416 786383
rect 70000 786307 70047 786363
rect 70103 786307 70171 786363
rect 70227 786307 70295 786363
rect 70351 786307 70419 786363
rect 70475 786307 73416 786363
rect 70000 786297 73416 786307
rect 70000 786241 71455 786297
rect 71511 786241 71597 786297
rect 71653 786241 71739 786297
rect 71795 786241 71881 786297
rect 71937 786241 72023 786297
rect 72079 786241 72165 786297
rect 72221 786241 72307 786297
rect 72363 786241 72449 786297
rect 72505 786241 72591 786297
rect 72647 786241 72733 786297
rect 72789 786241 72875 786297
rect 72931 786241 73017 786297
rect 73073 786241 73159 786297
rect 73215 786241 73301 786297
rect 73357 786241 73416 786297
rect 70000 786239 73416 786241
rect 70000 786183 70047 786239
rect 70103 786183 70171 786239
rect 70227 786183 70295 786239
rect 70351 786183 70419 786239
rect 70475 786183 73416 786239
rect 70000 786155 73416 786183
rect 70000 786115 71455 786155
rect 70000 786059 70047 786115
rect 70103 786059 70171 786115
rect 70227 786059 70295 786115
rect 70351 786059 70419 786115
rect 70475 786099 71455 786115
rect 71511 786099 71597 786155
rect 71653 786099 71739 786155
rect 71795 786099 71881 786155
rect 71937 786099 72023 786155
rect 72079 786099 72165 786155
rect 72221 786099 72307 786155
rect 72363 786099 72449 786155
rect 72505 786099 72591 786155
rect 72647 786099 72733 786155
rect 72789 786099 72875 786155
rect 72931 786099 73017 786155
rect 73073 786099 73159 786155
rect 73215 786099 73301 786155
rect 73357 786099 73416 786155
rect 70475 786059 73416 786099
rect 70000 786013 73416 786059
rect 70000 785991 71455 786013
rect 70000 785935 70047 785991
rect 70103 785935 70171 785991
rect 70227 785935 70295 785991
rect 70351 785935 70419 785991
rect 70475 785957 71455 785991
rect 71511 785957 71597 786013
rect 71653 785957 71739 786013
rect 71795 785957 71881 786013
rect 71937 785957 72023 786013
rect 72079 785957 72165 786013
rect 72221 785957 72307 786013
rect 72363 785957 72449 786013
rect 72505 785957 72591 786013
rect 72647 785957 72733 786013
rect 72789 785957 72875 786013
rect 72931 785957 73017 786013
rect 73073 785957 73159 786013
rect 73215 785957 73301 786013
rect 73357 785957 73416 786013
rect 70475 785935 73416 785957
rect 70000 785871 73416 785935
rect 70000 785867 71455 785871
rect 70000 785811 70047 785867
rect 70103 785811 70171 785867
rect 70227 785811 70295 785867
rect 70351 785811 70419 785867
rect 70475 785815 71455 785867
rect 71511 785815 71597 785871
rect 71653 785815 71739 785871
rect 71795 785815 71881 785871
rect 71937 785815 72023 785871
rect 72079 785815 72165 785871
rect 72221 785815 72307 785871
rect 72363 785815 72449 785871
rect 72505 785815 72591 785871
rect 72647 785815 72733 785871
rect 72789 785815 72875 785871
rect 72931 785815 73017 785871
rect 73073 785815 73159 785871
rect 73215 785815 73301 785871
rect 73357 785815 73416 785871
rect 70475 785811 73416 785815
rect 70000 785743 73416 785811
rect 70000 785687 70047 785743
rect 70103 785687 70171 785743
rect 70227 785687 70295 785743
rect 70351 785687 70419 785743
rect 70475 785729 73416 785743
rect 70475 785687 71455 785729
rect 70000 785673 71455 785687
rect 71511 785673 71597 785729
rect 71653 785673 71739 785729
rect 71795 785673 71881 785729
rect 71937 785673 72023 785729
rect 72079 785673 72165 785729
rect 72221 785673 72307 785729
rect 72363 785673 72449 785729
rect 72505 785673 72591 785729
rect 72647 785673 72733 785729
rect 72789 785673 72875 785729
rect 72931 785673 73017 785729
rect 73073 785673 73159 785729
rect 73215 785673 73301 785729
rect 73357 785673 73416 785729
rect 70000 785619 73416 785673
rect 70000 785563 70047 785619
rect 70103 785563 70171 785619
rect 70227 785563 70295 785619
rect 70351 785563 70419 785619
rect 70475 785587 73416 785619
rect 70475 785563 71455 785587
rect 70000 785531 71455 785563
rect 71511 785531 71597 785587
rect 71653 785531 71739 785587
rect 71795 785531 71881 785587
rect 71937 785531 72023 785587
rect 72079 785531 72165 785587
rect 72221 785531 72307 785587
rect 72363 785531 72449 785587
rect 72505 785531 72591 785587
rect 72647 785531 72733 785587
rect 72789 785531 72875 785587
rect 72931 785531 73017 785587
rect 73073 785531 73159 785587
rect 73215 785531 73301 785587
rect 73357 785531 73416 785587
rect 70000 785495 73416 785531
rect 70000 785439 70047 785495
rect 70103 785439 70171 785495
rect 70227 785439 70295 785495
rect 70351 785439 70419 785495
rect 70475 785445 73416 785495
rect 70475 785439 71455 785445
rect 70000 785389 71455 785439
rect 71511 785389 71597 785445
rect 71653 785389 71739 785445
rect 71795 785389 71881 785445
rect 71937 785389 72023 785445
rect 72079 785389 72165 785445
rect 72221 785389 72307 785445
rect 72363 785389 72449 785445
rect 72505 785389 72591 785445
rect 72647 785389 72733 785445
rect 72789 785389 72875 785445
rect 72931 785389 73017 785445
rect 73073 785389 73159 785445
rect 73215 785389 73301 785445
rect 73357 785389 73416 785445
rect 70000 785371 73416 785389
rect 70000 785315 70047 785371
rect 70103 785315 70171 785371
rect 70227 785315 70295 785371
rect 70351 785315 70419 785371
rect 70475 785315 73416 785371
rect 70000 785303 73416 785315
rect 70000 785247 71455 785303
rect 71511 785247 71597 785303
rect 71653 785247 71739 785303
rect 71795 785247 71881 785303
rect 71937 785247 72023 785303
rect 72079 785247 72165 785303
rect 72221 785247 72307 785303
rect 72363 785247 72449 785303
rect 72505 785247 72591 785303
rect 72647 785247 72733 785303
rect 72789 785247 72875 785303
rect 72931 785247 73017 785303
rect 73073 785247 73159 785303
rect 73215 785247 73301 785303
rect 73357 785247 73416 785303
rect 70000 785191 70047 785247
rect 70103 785191 70171 785247
rect 70227 785191 70295 785247
rect 70351 785191 70419 785247
rect 70475 785191 73416 785247
rect 70000 785161 73416 785191
rect 70000 785123 71455 785161
rect 70000 785067 70047 785123
rect 70103 785067 70171 785123
rect 70227 785067 70295 785123
rect 70351 785067 70419 785123
rect 70475 785105 71455 785123
rect 71511 785105 71597 785161
rect 71653 785105 71739 785161
rect 71795 785105 71881 785161
rect 71937 785105 72023 785161
rect 72079 785105 72165 785161
rect 72221 785105 72307 785161
rect 72363 785105 72449 785161
rect 72505 785105 72591 785161
rect 72647 785105 72733 785161
rect 72789 785105 72875 785161
rect 72931 785105 73017 785161
rect 73073 785105 73159 785161
rect 73215 785105 73301 785161
rect 73357 785105 73416 785161
rect 70475 785067 73416 785105
rect 70000 785019 73416 785067
rect 70000 784999 71455 785019
rect 70000 784943 70047 784999
rect 70103 784943 70171 784999
rect 70227 784943 70295 784999
rect 70351 784943 70419 784999
rect 70475 784963 71455 784999
rect 71511 784963 71597 785019
rect 71653 784963 71739 785019
rect 71795 784963 71881 785019
rect 71937 784963 72023 785019
rect 72079 784963 72165 785019
rect 72221 784963 72307 785019
rect 72363 784963 72449 785019
rect 72505 784963 72591 785019
rect 72647 784963 72733 785019
rect 72789 784963 72875 785019
rect 72931 784963 73017 785019
rect 73073 784963 73159 785019
rect 73215 784963 73301 785019
rect 73357 784963 73416 785019
rect 70475 784943 73416 784963
rect 70000 784877 73416 784943
rect 70000 784875 71455 784877
rect 70000 784819 70047 784875
rect 70103 784819 70171 784875
rect 70227 784819 70295 784875
rect 70351 784819 70419 784875
rect 70475 784821 71455 784875
rect 71511 784821 71597 784877
rect 71653 784821 71739 784877
rect 71795 784821 71881 784877
rect 71937 784821 72023 784877
rect 72079 784821 72165 784877
rect 72221 784821 72307 784877
rect 72363 784821 72449 784877
rect 72505 784821 72591 784877
rect 72647 784821 72733 784877
rect 72789 784821 72875 784877
rect 72931 784821 73017 784877
rect 73073 784821 73159 784877
rect 73215 784821 73301 784877
rect 73357 784821 73416 784877
rect 699992 786753 700051 786809
rect 700107 786753 700193 786809
rect 700249 786753 700335 786809
rect 700391 786753 700477 786809
rect 700533 786753 700619 786809
rect 700675 786753 700761 786809
rect 700817 786753 700903 786809
rect 700959 786753 701045 786809
rect 701101 786753 701187 786809
rect 701243 786753 701329 786809
rect 701385 786753 701471 786809
rect 701527 786753 701613 786809
rect 701669 786753 701755 786809
rect 701811 786753 701897 786809
rect 701953 786755 705525 786809
rect 705581 786755 705649 786811
rect 705705 786755 705773 786811
rect 705829 786755 705897 786811
rect 705953 786755 706000 786811
rect 701953 786753 706000 786755
rect 699992 786687 706000 786753
rect 699992 786667 705525 786687
rect 699992 786611 700051 786667
rect 700107 786611 700193 786667
rect 700249 786611 700335 786667
rect 700391 786611 700477 786667
rect 700533 786611 700619 786667
rect 700675 786611 700761 786667
rect 700817 786611 700903 786667
rect 700959 786611 701045 786667
rect 701101 786611 701187 786667
rect 701243 786611 701329 786667
rect 701385 786611 701471 786667
rect 701527 786611 701613 786667
rect 701669 786611 701755 786667
rect 701811 786611 701897 786667
rect 701953 786631 705525 786667
rect 705581 786631 705649 786687
rect 705705 786631 705773 786687
rect 705829 786631 705897 786687
rect 705953 786631 706000 786687
rect 701953 786611 706000 786631
rect 699992 786563 706000 786611
rect 699992 786525 705525 786563
rect 699992 786469 700051 786525
rect 700107 786469 700193 786525
rect 700249 786469 700335 786525
rect 700391 786469 700477 786525
rect 700533 786469 700619 786525
rect 700675 786469 700761 786525
rect 700817 786469 700903 786525
rect 700959 786469 701045 786525
rect 701101 786469 701187 786525
rect 701243 786469 701329 786525
rect 701385 786469 701471 786525
rect 701527 786469 701613 786525
rect 701669 786469 701755 786525
rect 701811 786469 701897 786525
rect 701953 786507 705525 786525
rect 705581 786507 705649 786563
rect 705705 786507 705773 786563
rect 705829 786507 705897 786563
rect 705953 786507 706000 786563
rect 701953 786469 706000 786507
rect 699992 786439 706000 786469
rect 699992 786383 705525 786439
rect 705581 786383 705649 786439
rect 705705 786383 705773 786439
rect 705829 786383 705897 786439
rect 705953 786383 706000 786439
rect 699992 786327 700051 786383
rect 700107 786327 700193 786383
rect 700249 786327 700335 786383
rect 700391 786327 700477 786383
rect 700533 786327 700619 786383
rect 700675 786327 700761 786383
rect 700817 786327 700903 786383
rect 700959 786327 701045 786383
rect 701101 786327 701187 786383
rect 701243 786327 701329 786383
rect 701385 786327 701471 786383
rect 701527 786327 701613 786383
rect 701669 786327 701755 786383
rect 701811 786327 701897 786383
rect 701953 786327 706000 786383
rect 699992 786315 706000 786327
rect 699992 786259 705525 786315
rect 705581 786259 705649 786315
rect 705705 786259 705773 786315
rect 705829 786259 705897 786315
rect 705953 786259 706000 786315
rect 699992 786241 706000 786259
rect 699992 786185 700051 786241
rect 700107 786185 700193 786241
rect 700249 786185 700335 786241
rect 700391 786185 700477 786241
rect 700533 786185 700619 786241
rect 700675 786185 700761 786241
rect 700817 786185 700903 786241
rect 700959 786185 701045 786241
rect 701101 786185 701187 786241
rect 701243 786185 701329 786241
rect 701385 786185 701471 786241
rect 701527 786185 701613 786241
rect 701669 786185 701755 786241
rect 701811 786185 701897 786241
rect 701953 786191 706000 786241
rect 701953 786185 705525 786191
rect 699992 786135 705525 786185
rect 705581 786135 705649 786191
rect 705705 786135 705773 786191
rect 705829 786135 705897 786191
rect 705953 786135 706000 786191
rect 699992 786099 706000 786135
rect 699992 786043 700051 786099
rect 700107 786043 700193 786099
rect 700249 786043 700335 786099
rect 700391 786043 700477 786099
rect 700533 786043 700619 786099
rect 700675 786043 700761 786099
rect 700817 786043 700903 786099
rect 700959 786043 701045 786099
rect 701101 786043 701187 786099
rect 701243 786043 701329 786099
rect 701385 786043 701471 786099
rect 701527 786043 701613 786099
rect 701669 786043 701755 786099
rect 701811 786043 701897 786099
rect 701953 786067 706000 786099
rect 701953 786043 705525 786067
rect 699992 786011 705525 786043
rect 705581 786011 705649 786067
rect 705705 786011 705773 786067
rect 705829 786011 705897 786067
rect 705953 786011 706000 786067
rect 699992 785957 706000 786011
rect 699992 785901 700051 785957
rect 700107 785901 700193 785957
rect 700249 785901 700335 785957
rect 700391 785901 700477 785957
rect 700533 785901 700619 785957
rect 700675 785901 700761 785957
rect 700817 785901 700903 785957
rect 700959 785901 701045 785957
rect 701101 785901 701187 785957
rect 701243 785901 701329 785957
rect 701385 785901 701471 785957
rect 701527 785901 701613 785957
rect 701669 785901 701755 785957
rect 701811 785901 701897 785957
rect 701953 785943 706000 785957
rect 701953 785901 705525 785943
rect 699992 785887 705525 785901
rect 705581 785887 705649 785943
rect 705705 785887 705773 785943
rect 705829 785887 705897 785943
rect 705953 785887 706000 785943
rect 699992 785819 706000 785887
rect 699992 785815 705525 785819
rect 699992 785759 700051 785815
rect 700107 785759 700193 785815
rect 700249 785759 700335 785815
rect 700391 785759 700477 785815
rect 700533 785759 700619 785815
rect 700675 785759 700761 785815
rect 700817 785759 700903 785815
rect 700959 785759 701045 785815
rect 701101 785759 701187 785815
rect 701243 785759 701329 785815
rect 701385 785759 701471 785815
rect 701527 785759 701613 785815
rect 701669 785759 701755 785815
rect 701811 785759 701897 785815
rect 701953 785763 705525 785815
rect 705581 785763 705649 785819
rect 705705 785763 705773 785819
rect 705829 785763 705897 785819
rect 705953 785763 706000 785819
rect 701953 785759 706000 785763
rect 699992 785695 706000 785759
rect 699992 785673 705525 785695
rect 699992 785617 700051 785673
rect 700107 785617 700193 785673
rect 700249 785617 700335 785673
rect 700391 785617 700477 785673
rect 700533 785617 700619 785673
rect 700675 785617 700761 785673
rect 700817 785617 700903 785673
rect 700959 785617 701045 785673
rect 701101 785617 701187 785673
rect 701243 785617 701329 785673
rect 701385 785617 701471 785673
rect 701527 785617 701613 785673
rect 701669 785617 701755 785673
rect 701811 785617 701897 785673
rect 701953 785639 705525 785673
rect 705581 785639 705649 785695
rect 705705 785639 705773 785695
rect 705829 785639 705897 785695
rect 705953 785639 706000 785695
rect 701953 785617 706000 785639
rect 699992 785571 706000 785617
rect 699992 785531 705525 785571
rect 699992 785475 700051 785531
rect 700107 785475 700193 785531
rect 700249 785475 700335 785531
rect 700391 785475 700477 785531
rect 700533 785475 700619 785531
rect 700675 785475 700761 785531
rect 700817 785475 700903 785531
rect 700959 785475 701045 785531
rect 701101 785475 701187 785531
rect 701243 785475 701329 785531
rect 701385 785475 701471 785531
rect 701527 785475 701613 785531
rect 701669 785475 701755 785531
rect 701811 785475 701897 785531
rect 701953 785515 705525 785531
rect 705581 785515 705649 785571
rect 705705 785515 705773 785571
rect 705829 785515 705897 785571
rect 705953 785515 706000 785571
rect 701953 785475 706000 785515
rect 699992 785447 706000 785475
rect 699992 785391 705525 785447
rect 705581 785391 705649 785447
rect 705705 785391 705773 785447
rect 705829 785391 705897 785447
rect 705953 785391 706000 785447
rect 699992 785389 706000 785391
rect 699992 785333 700051 785389
rect 700107 785333 700193 785389
rect 700249 785333 700335 785389
rect 700391 785333 700477 785389
rect 700533 785333 700619 785389
rect 700675 785333 700761 785389
rect 700817 785333 700903 785389
rect 700959 785333 701045 785389
rect 701101 785333 701187 785389
rect 701243 785333 701329 785389
rect 701385 785333 701471 785389
rect 701527 785333 701613 785389
rect 701669 785333 701755 785389
rect 701811 785333 701897 785389
rect 701953 785333 706000 785389
rect 699992 785323 706000 785333
rect 699992 785267 705525 785323
rect 705581 785267 705649 785323
rect 705705 785267 705773 785323
rect 705829 785267 705897 785323
rect 705953 785267 706000 785323
rect 699992 785247 706000 785267
rect 699992 785191 700051 785247
rect 700107 785191 700193 785247
rect 700249 785191 700335 785247
rect 700391 785191 700477 785247
rect 700533 785191 700619 785247
rect 700675 785191 700761 785247
rect 700817 785191 700903 785247
rect 700959 785191 701045 785247
rect 701101 785191 701187 785247
rect 701243 785191 701329 785247
rect 701385 785191 701471 785247
rect 701527 785191 701613 785247
rect 701669 785191 701755 785247
rect 701811 785191 701897 785247
rect 701953 785199 706000 785247
rect 701953 785191 705525 785199
rect 699992 785143 705525 785191
rect 705581 785143 705649 785199
rect 705705 785143 705773 785199
rect 705829 785143 705897 785199
rect 705953 785143 706000 785199
rect 699992 785105 706000 785143
rect 699992 785049 700051 785105
rect 700107 785049 700193 785105
rect 700249 785049 700335 785105
rect 700391 785049 700477 785105
rect 700533 785049 700619 785105
rect 700675 785049 700761 785105
rect 700817 785049 700903 785105
rect 700959 785049 701045 785105
rect 701101 785049 701187 785105
rect 701243 785049 701329 785105
rect 701385 785049 701471 785105
rect 701527 785049 701613 785105
rect 701669 785049 701755 785105
rect 701811 785049 701897 785105
rect 701953 785075 706000 785105
rect 701953 785049 705525 785075
rect 699992 785019 705525 785049
rect 705581 785019 705649 785075
rect 705705 785019 705773 785075
rect 705829 785019 705897 785075
rect 705953 785019 706000 785075
rect 699992 784963 706000 785019
rect 699992 784907 700051 784963
rect 700107 784907 700193 784963
rect 700249 784907 700335 784963
rect 700391 784907 700477 784963
rect 700533 784907 700619 784963
rect 700675 784907 700761 784963
rect 700817 784907 700903 784963
rect 700959 784907 701045 784963
rect 701101 784907 701187 784963
rect 701243 784907 701329 784963
rect 701385 784907 701471 784963
rect 701527 784907 701613 784963
rect 701669 784907 701755 784963
rect 701811 784907 701897 784963
rect 701953 784951 706000 784963
rect 701953 784907 705525 784951
rect 699992 784895 705525 784907
rect 705581 784895 705649 784951
rect 705705 784895 705773 784951
rect 705829 784895 705897 784951
rect 705953 784895 706000 784951
rect 699992 784828 706000 784895
rect 70475 784819 73416 784821
rect 70000 784752 73416 784819
rect 70000 784105 73416 784172
rect 70000 784049 70047 784105
rect 70103 784049 70171 784105
rect 70227 784049 70295 784105
rect 70351 784049 70419 784105
rect 70475 784094 73416 784105
rect 70475 784049 71466 784094
rect 70000 784038 71466 784049
rect 71522 784038 71608 784094
rect 71664 784038 71750 784094
rect 71806 784038 71892 784094
rect 71948 784038 72034 784094
rect 72090 784038 72176 784094
rect 72232 784038 72318 784094
rect 72374 784038 72460 784094
rect 72516 784038 72602 784094
rect 72658 784038 72744 784094
rect 72800 784038 72886 784094
rect 72942 784038 73028 784094
rect 73084 784038 73170 784094
rect 73226 784038 73312 784094
rect 73368 784038 73416 784094
rect 70000 783981 73416 784038
rect 70000 783925 70047 783981
rect 70103 783925 70171 783981
rect 70227 783925 70295 783981
rect 70351 783925 70419 783981
rect 70475 783952 73416 783981
rect 70475 783925 71466 783952
rect 70000 783896 71466 783925
rect 71522 783896 71608 783952
rect 71664 783896 71750 783952
rect 71806 783896 71892 783952
rect 71948 783896 72034 783952
rect 72090 783896 72176 783952
rect 72232 783896 72318 783952
rect 72374 783896 72460 783952
rect 72516 783896 72602 783952
rect 72658 783896 72744 783952
rect 72800 783896 72886 783952
rect 72942 783896 73028 783952
rect 73084 783896 73170 783952
rect 73226 783896 73312 783952
rect 73368 783896 73416 783952
rect 70000 783857 73416 783896
rect 70000 783801 70047 783857
rect 70103 783801 70171 783857
rect 70227 783801 70295 783857
rect 70351 783801 70419 783857
rect 70475 783810 73416 783857
rect 70475 783801 71466 783810
rect 70000 783754 71466 783801
rect 71522 783754 71608 783810
rect 71664 783754 71750 783810
rect 71806 783754 71892 783810
rect 71948 783754 72034 783810
rect 72090 783754 72176 783810
rect 72232 783754 72318 783810
rect 72374 783754 72460 783810
rect 72516 783754 72602 783810
rect 72658 783754 72744 783810
rect 72800 783754 72886 783810
rect 72942 783754 73028 783810
rect 73084 783754 73170 783810
rect 73226 783754 73312 783810
rect 73368 783754 73416 783810
rect 70000 783733 73416 783754
rect 70000 783677 70047 783733
rect 70103 783677 70171 783733
rect 70227 783677 70295 783733
rect 70351 783677 70419 783733
rect 70475 783677 73416 783733
rect 70000 783668 73416 783677
rect 70000 783612 71466 783668
rect 71522 783612 71608 783668
rect 71664 783612 71750 783668
rect 71806 783612 71892 783668
rect 71948 783612 72034 783668
rect 72090 783612 72176 783668
rect 72232 783612 72318 783668
rect 72374 783612 72460 783668
rect 72516 783612 72602 783668
rect 72658 783612 72744 783668
rect 72800 783612 72886 783668
rect 72942 783612 73028 783668
rect 73084 783612 73170 783668
rect 73226 783612 73312 783668
rect 73368 783612 73416 783668
rect 70000 783609 73416 783612
rect 70000 783553 70047 783609
rect 70103 783553 70171 783609
rect 70227 783553 70295 783609
rect 70351 783553 70419 783609
rect 70475 783553 73416 783609
rect 70000 783526 73416 783553
rect 70000 783485 71466 783526
rect 70000 783429 70047 783485
rect 70103 783429 70171 783485
rect 70227 783429 70295 783485
rect 70351 783429 70419 783485
rect 70475 783470 71466 783485
rect 71522 783470 71608 783526
rect 71664 783470 71750 783526
rect 71806 783470 71892 783526
rect 71948 783470 72034 783526
rect 72090 783470 72176 783526
rect 72232 783470 72318 783526
rect 72374 783470 72460 783526
rect 72516 783470 72602 783526
rect 72658 783470 72744 783526
rect 72800 783470 72886 783526
rect 72942 783470 73028 783526
rect 73084 783470 73170 783526
rect 73226 783470 73312 783526
rect 73368 783470 73416 783526
rect 70475 783429 73416 783470
rect 70000 783384 73416 783429
rect 70000 783361 71466 783384
rect 70000 783305 70047 783361
rect 70103 783305 70171 783361
rect 70227 783305 70295 783361
rect 70351 783305 70419 783361
rect 70475 783328 71466 783361
rect 71522 783328 71608 783384
rect 71664 783328 71750 783384
rect 71806 783328 71892 783384
rect 71948 783328 72034 783384
rect 72090 783328 72176 783384
rect 72232 783328 72318 783384
rect 72374 783328 72460 783384
rect 72516 783328 72602 783384
rect 72658 783328 72744 783384
rect 72800 783328 72886 783384
rect 72942 783328 73028 783384
rect 73084 783328 73170 783384
rect 73226 783328 73312 783384
rect 73368 783328 73416 783384
rect 70475 783305 73416 783328
rect 70000 783242 73416 783305
rect 70000 783237 71466 783242
rect 70000 783181 70047 783237
rect 70103 783181 70171 783237
rect 70227 783181 70295 783237
rect 70351 783181 70419 783237
rect 70475 783186 71466 783237
rect 71522 783186 71608 783242
rect 71664 783186 71750 783242
rect 71806 783186 71892 783242
rect 71948 783186 72034 783242
rect 72090 783186 72176 783242
rect 72232 783186 72318 783242
rect 72374 783186 72460 783242
rect 72516 783186 72602 783242
rect 72658 783186 72744 783242
rect 72800 783186 72886 783242
rect 72942 783186 73028 783242
rect 73084 783186 73170 783242
rect 73226 783186 73312 783242
rect 73368 783186 73416 783242
rect 70475 783181 73416 783186
rect 70000 783113 73416 783181
rect 70000 783057 70047 783113
rect 70103 783057 70171 783113
rect 70227 783057 70295 783113
rect 70351 783057 70419 783113
rect 70475 783100 73416 783113
rect 70475 783057 71466 783100
rect 70000 783044 71466 783057
rect 71522 783044 71608 783100
rect 71664 783044 71750 783100
rect 71806 783044 71892 783100
rect 71948 783044 72034 783100
rect 72090 783044 72176 783100
rect 72232 783044 72318 783100
rect 72374 783044 72460 783100
rect 72516 783044 72602 783100
rect 72658 783044 72744 783100
rect 72800 783044 72886 783100
rect 72942 783044 73028 783100
rect 73084 783044 73170 783100
rect 73226 783044 73312 783100
rect 73368 783044 73416 783100
rect 70000 782989 73416 783044
rect 70000 782933 70047 782989
rect 70103 782933 70171 782989
rect 70227 782933 70295 782989
rect 70351 782933 70419 782989
rect 70475 782958 73416 782989
rect 70475 782933 71466 782958
rect 70000 782902 71466 782933
rect 71522 782902 71608 782958
rect 71664 782902 71750 782958
rect 71806 782902 71892 782958
rect 71948 782902 72034 782958
rect 72090 782902 72176 782958
rect 72232 782902 72318 782958
rect 72374 782902 72460 782958
rect 72516 782902 72602 782958
rect 72658 782902 72744 782958
rect 72800 782902 72886 782958
rect 72942 782902 73028 782958
rect 73084 782902 73170 782958
rect 73226 782902 73312 782958
rect 73368 782902 73416 782958
rect 70000 782865 73416 782902
rect 70000 782809 70047 782865
rect 70103 782809 70171 782865
rect 70227 782809 70295 782865
rect 70351 782809 70419 782865
rect 70475 782816 73416 782865
rect 70475 782809 71466 782816
rect 70000 782760 71466 782809
rect 71522 782760 71608 782816
rect 71664 782760 71750 782816
rect 71806 782760 71892 782816
rect 71948 782760 72034 782816
rect 72090 782760 72176 782816
rect 72232 782760 72318 782816
rect 72374 782760 72460 782816
rect 72516 782760 72602 782816
rect 72658 782760 72744 782816
rect 72800 782760 72886 782816
rect 72942 782760 73028 782816
rect 73084 782760 73170 782816
rect 73226 782760 73312 782816
rect 73368 782760 73416 782816
rect 70000 782741 73416 782760
rect 70000 782685 70047 782741
rect 70103 782685 70171 782741
rect 70227 782685 70295 782741
rect 70351 782685 70419 782741
rect 70475 782685 73416 782741
rect 70000 782674 73416 782685
rect 70000 782618 71466 782674
rect 71522 782618 71608 782674
rect 71664 782618 71750 782674
rect 71806 782618 71892 782674
rect 71948 782618 72034 782674
rect 72090 782618 72176 782674
rect 72232 782618 72318 782674
rect 72374 782618 72460 782674
rect 72516 782618 72602 782674
rect 72658 782618 72744 782674
rect 72800 782618 72886 782674
rect 72942 782618 73028 782674
rect 73084 782618 73170 782674
rect 73226 782618 73312 782674
rect 73368 782618 73416 782674
rect 70000 782617 73416 782618
rect 70000 782561 70047 782617
rect 70103 782561 70171 782617
rect 70227 782561 70295 782617
rect 70351 782561 70419 782617
rect 70475 782561 73416 782617
rect 70000 782532 73416 782561
rect 70000 782493 71466 782532
rect 70000 782437 70047 782493
rect 70103 782437 70171 782493
rect 70227 782437 70295 782493
rect 70351 782437 70419 782493
rect 70475 782476 71466 782493
rect 71522 782476 71608 782532
rect 71664 782476 71750 782532
rect 71806 782476 71892 782532
rect 71948 782476 72034 782532
rect 72090 782476 72176 782532
rect 72232 782476 72318 782532
rect 72374 782476 72460 782532
rect 72516 782476 72602 782532
rect 72658 782476 72744 782532
rect 72800 782476 72886 782532
rect 72942 782476 73028 782532
rect 73084 782476 73170 782532
rect 73226 782476 73312 782532
rect 73368 782476 73416 782532
rect 70475 782437 73416 782476
rect 70000 782390 73416 782437
rect 70000 782369 71466 782390
rect 70000 782313 70047 782369
rect 70103 782313 70171 782369
rect 70227 782313 70295 782369
rect 70351 782313 70419 782369
rect 70475 782334 71466 782369
rect 71522 782334 71608 782390
rect 71664 782334 71750 782390
rect 71806 782334 71892 782390
rect 71948 782334 72034 782390
rect 72090 782334 72176 782390
rect 72232 782334 72318 782390
rect 72374 782334 72460 782390
rect 72516 782334 72602 782390
rect 72658 782334 72744 782390
rect 72800 782334 72886 782390
rect 72942 782334 73028 782390
rect 73084 782334 73170 782390
rect 73226 782334 73312 782390
rect 73368 782334 73416 782390
rect 70475 782313 73416 782334
rect 70000 782272 73416 782313
rect 699992 784105 706000 784172
rect 699992 784103 705525 784105
rect 699992 784047 700051 784103
rect 700107 784047 700193 784103
rect 700249 784047 700335 784103
rect 700391 784047 700477 784103
rect 700533 784047 700619 784103
rect 700675 784047 700761 784103
rect 700817 784047 700903 784103
rect 700959 784047 701045 784103
rect 701101 784047 701187 784103
rect 701243 784047 701329 784103
rect 701385 784047 701471 784103
rect 701527 784047 701613 784103
rect 701669 784047 701755 784103
rect 701811 784047 701897 784103
rect 701953 784049 705525 784103
rect 705581 784049 705649 784105
rect 705705 784049 705773 784105
rect 705829 784049 705897 784105
rect 705953 784049 706000 784105
rect 701953 784047 706000 784049
rect 699992 783981 706000 784047
rect 699992 783961 705525 783981
rect 699992 783905 700051 783961
rect 700107 783905 700193 783961
rect 700249 783905 700335 783961
rect 700391 783905 700477 783961
rect 700533 783905 700619 783961
rect 700675 783905 700761 783961
rect 700817 783905 700903 783961
rect 700959 783905 701045 783961
rect 701101 783905 701187 783961
rect 701243 783905 701329 783961
rect 701385 783905 701471 783961
rect 701527 783905 701613 783961
rect 701669 783905 701755 783961
rect 701811 783905 701897 783961
rect 701953 783925 705525 783961
rect 705581 783925 705649 783981
rect 705705 783925 705773 783981
rect 705829 783925 705897 783981
rect 705953 783925 706000 783981
rect 701953 783905 706000 783925
rect 699992 783857 706000 783905
rect 699992 783819 705525 783857
rect 699992 783763 700051 783819
rect 700107 783763 700193 783819
rect 700249 783763 700335 783819
rect 700391 783763 700477 783819
rect 700533 783763 700619 783819
rect 700675 783763 700761 783819
rect 700817 783763 700903 783819
rect 700959 783763 701045 783819
rect 701101 783763 701187 783819
rect 701243 783763 701329 783819
rect 701385 783763 701471 783819
rect 701527 783763 701613 783819
rect 701669 783763 701755 783819
rect 701811 783763 701897 783819
rect 701953 783801 705525 783819
rect 705581 783801 705649 783857
rect 705705 783801 705773 783857
rect 705829 783801 705897 783857
rect 705953 783801 706000 783857
rect 701953 783763 706000 783801
rect 699992 783733 706000 783763
rect 699992 783677 705525 783733
rect 705581 783677 705649 783733
rect 705705 783677 705773 783733
rect 705829 783677 705897 783733
rect 705953 783677 706000 783733
rect 699992 783621 700051 783677
rect 700107 783621 700193 783677
rect 700249 783621 700335 783677
rect 700391 783621 700477 783677
rect 700533 783621 700619 783677
rect 700675 783621 700761 783677
rect 700817 783621 700903 783677
rect 700959 783621 701045 783677
rect 701101 783621 701187 783677
rect 701243 783621 701329 783677
rect 701385 783621 701471 783677
rect 701527 783621 701613 783677
rect 701669 783621 701755 783677
rect 701811 783621 701897 783677
rect 701953 783621 706000 783677
rect 699992 783609 706000 783621
rect 699992 783553 705525 783609
rect 705581 783553 705649 783609
rect 705705 783553 705773 783609
rect 705829 783553 705897 783609
rect 705953 783553 706000 783609
rect 699992 783535 706000 783553
rect 699992 783479 700051 783535
rect 700107 783479 700193 783535
rect 700249 783479 700335 783535
rect 700391 783479 700477 783535
rect 700533 783479 700619 783535
rect 700675 783479 700761 783535
rect 700817 783479 700903 783535
rect 700959 783479 701045 783535
rect 701101 783479 701187 783535
rect 701243 783479 701329 783535
rect 701385 783479 701471 783535
rect 701527 783479 701613 783535
rect 701669 783479 701755 783535
rect 701811 783479 701897 783535
rect 701953 783485 706000 783535
rect 701953 783479 705525 783485
rect 699992 783429 705525 783479
rect 705581 783429 705649 783485
rect 705705 783429 705773 783485
rect 705829 783429 705897 783485
rect 705953 783429 706000 783485
rect 699992 783393 706000 783429
rect 699992 783337 700051 783393
rect 700107 783337 700193 783393
rect 700249 783337 700335 783393
rect 700391 783337 700477 783393
rect 700533 783337 700619 783393
rect 700675 783337 700761 783393
rect 700817 783337 700903 783393
rect 700959 783337 701045 783393
rect 701101 783337 701187 783393
rect 701243 783337 701329 783393
rect 701385 783337 701471 783393
rect 701527 783337 701613 783393
rect 701669 783337 701755 783393
rect 701811 783337 701897 783393
rect 701953 783361 706000 783393
rect 701953 783337 705525 783361
rect 699992 783305 705525 783337
rect 705581 783305 705649 783361
rect 705705 783305 705773 783361
rect 705829 783305 705897 783361
rect 705953 783305 706000 783361
rect 699992 783251 706000 783305
rect 699992 783195 700051 783251
rect 700107 783195 700193 783251
rect 700249 783195 700335 783251
rect 700391 783195 700477 783251
rect 700533 783195 700619 783251
rect 700675 783195 700761 783251
rect 700817 783195 700903 783251
rect 700959 783195 701045 783251
rect 701101 783195 701187 783251
rect 701243 783195 701329 783251
rect 701385 783195 701471 783251
rect 701527 783195 701613 783251
rect 701669 783195 701755 783251
rect 701811 783195 701897 783251
rect 701953 783237 706000 783251
rect 701953 783195 705525 783237
rect 699992 783181 705525 783195
rect 705581 783181 705649 783237
rect 705705 783181 705773 783237
rect 705829 783181 705897 783237
rect 705953 783181 706000 783237
rect 699992 783113 706000 783181
rect 699992 783109 705525 783113
rect 699992 783053 700051 783109
rect 700107 783053 700193 783109
rect 700249 783053 700335 783109
rect 700391 783053 700477 783109
rect 700533 783053 700619 783109
rect 700675 783053 700761 783109
rect 700817 783053 700903 783109
rect 700959 783053 701045 783109
rect 701101 783053 701187 783109
rect 701243 783053 701329 783109
rect 701385 783053 701471 783109
rect 701527 783053 701613 783109
rect 701669 783053 701755 783109
rect 701811 783053 701897 783109
rect 701953 783057 705525 783109
rect 705581 783057 705649 783113
rect 705705 783057 705773 783113
rect 705829 783057 705897 783113
rect 705953 783057 706000 783113
rect 701953 783053 706000 783057
rect 699992 782989 706000 783053
rect 699992 782967 705525 782989
rect 699992 782911 700051 782967
rect 700107 782911 700193 782967
rect 700249 782911 700335 782967
rect 700391 782911 700477 782967
rect 700533 782911 700619 782967
rect 700675 782911 700761 782967
rect 700817 782911 700903 782967
rect 700959 782911 701045 782967
rect 701101 782911 701187 782967
rect 701243 782911 701329 782967
rect 701385 782911 701471 782967
rect 701527 782911 701613 782967
rect 701669 782911 701755 782967
rect 701811 782911 701897 782967
rect 701953 782933 705525 782967
rect 705581 782933 705649 782989
rect 705705 782933 705773 782989
rect 705829 782933 705897 782989
rect 705953 782933 706000 782989
rect 701953 782911 706000 782933
rect 699992 782865 706000 782911
rect 699992 782825 705525 782865
rect 699992 782769 700051 782825
rect 700107 782769 700193 782825
rect 700249 782769 700335 782825
rect 700391 782769 700477 782825
rect 700533 782769 700619 782825
rect 700675 782769 700761 782825
rect 700817 782769 700903 782825
rect 700959 782769 701045 782825
rect 701101 782769 701187 782825
rect 701243 782769 701329 782825
rect 701385 782769 701471 782825
rect 701527 782769 701613 782825
rect 701669 782769 701755 782825
rect 701811 782769 701897 782825
rect 701953 782809 705525 782825
rect 705581 782809 705649 782865
rect 705705 782809 705773 782865
rect 705829 782809 705897 782865
rect 705953 782809 706000 782865
rect 701953 782769 706000 782809
rect 699992 782741 706000 782769
rect 699992 782685 705525 782741
rect 705581 782685 705649 782741
rect 705705 782685 705773 782741
rect 705829 782685 705897 782741
rect 705953 782685 706000 782741
rect 699992 782683 706000 782685
rect 699992 782627 700051 782683
rect 700107 782627 700193 782683
rect 700249 782627 700335 782683
rect 700391 782627 700477 782683
rect 700533 782627 700619 782683
rect 700675 782627 700761 782683
rect 700817 782627 700903 782683
rect 700959 782627 701045 782683
rect 701101 782627 701187 782683
rect 701243 782627 701329 782683
rect 701385 782627 701471 782683
rect 701527 782627 701613 782683
rect 701669 782627 701755 782683
rect 701811 782627 701897 782683
rect 701953 782627 706000 782683
rect 699992 782617 706000 782627
rect 699992 782561 705525 782617
rect 705581 782561 705649 782617
rect 705705 782561 705773 782617
rect 705829 782561 705897 782617
rect 705953 782561 706000 782617
rect 699992 782541 706000 782561
rect 699992 782485 700051 782541
rect 700107 782485 700193 782541
rect 700249 782485 700335 782541
rect 700391 782485 700477 782541
rect 700533 782485 700619 782541
rect 700675 782485 700761 782541
rect 700817 782485 700903 782541
rect 700959 782485 701045 782541
rect 701101 782485 701187 782541
rect 701243 782485 701329 782541
rect 701385 782485 701471 782541
rect 701527 782485 701613 782541
rect 701669 782485 701755 782541
rect 701811 782485 701897 782541
rect 701953 782493 706000 782541
rect 701953 782485 705525 782493
rect 699992 782437 705525 782485
rect 705581 782437 705649 782493
rect 705705 782437 705773 782493
rect 705829 782437 705897 782493
rect 705953 782437 706000 782493
rect 699992 782399 706000 782437
rect 699992 782343 700051 782399
rect 700107 782343 700193 782399
rect 700249 782343 700335 782399
rect 700391 782343 700477 782399
rect 700533 782343 700619 782399
rect 700675 782343 700761 782399
rect 700817 782343 700903 782399
rect 700959 782343 701045 782399
rect 701101 782343 701187 782399
rect 701243 782343 701329 782399
rect 701385 782343 701471 782399
rect 701527 782343 701613 782399
rect 701669 782343 701755 782399
rect 701811 782343 701897 782399
rect 701953 782369 706000 782399
rect 701953 782343 705525 782369
rect 699992 782313 705525 782343
rect 705581 782313 705649 782369
rect 705705 782313 705773 782369
rect 705829 782313 705897 782369
rect 705953 782313 706000 782369
rect 699992 782257 706000 782313
rect 699992 782201 700051 782257
rect 700107 782201 700193 782257
rect 700249 782201 700335 782257
rect 700391 782201 700477 782257
rect 700533 782201 700619 782257
rect 700675 782201 700761 782257
rect 700817 782201 700903 782257
rect 700959 782201 701045 782257
rect 701101 782201 701187 782257
rect 701243 782201 701329 782257
rect 701385 782201 701471 782257
rect 701527 782201 701613 782257
rect 701669 782201 701755 782257
rect 701811 782201 701897 782257
rect 701953 782245 706000 782257
rect 701953 782201 705525 782245
rect 699992 782189 705525 782201
rect 705581 782189 705649 782245
rect 705705 782189 705773 782245
rect 705829 782189 705897 782245
rect 705953 782189 706000 782245
rect 699992 782122 706000 782189
rect 699992 781735 706000 781802
rect 699992 781733 705525 781735
rect 699992 781677 700051 781733
rect 700107 781677 700193 781733
rect 700249 781677 700335 781733
rect 700391 781677 700477 781733
rect 700533 781677 700619 781733
rect 700675 781677 700761 781733
rect 700817 781677 700903 781733
rect 700959 781677 701045 781733
rect 701101 781677 701187 781733
rect 701243 781677 701329 781733
rect 701385 781677 701471 781733
rect 701527 781677 701613 781733
rect 701669 781677 701755 781733
rect 701811 781677 701897 781733
rect 701953 781679 705525 781733
rect 705581 781679 705649 781735
rect 705705 781679 705773 781735
rect 705829 781679 705897 781735
rect 705953 781679 706000 781735
rect 701953 781677 706000 781679
rect 699992 781611 706000 781677
rect 699992 781591 705525 781611
rect 699992 781535 700051 781591
rect 700107 781535 700193 781591
rect 700249 781535 700335 781591
rect 700391 781535 700477 781591
rect 700533 781535 700619 781591
rect 700675 781535 700761 781591
rect 700817 781535 700903 781591
rect 700959 781535 701045 781591
rect 701101 781535 701187 781591
rect 701243 781535 701329 781591
rect 701385 781535 701471 781591
rect 701527 781535 701613 781591
rect 701669 781535 701755 781591
rect 701811 781535 701897 781591
rect 701953 781555 705525 781591
rect 705581 781555 705649 781611
rect 705705 781555 705773 781611
rect 705829 781555 705897 781611
rect 705953 781555 706000 781611
rect 701953 781535 706000 781555
rect 699992 781487 706000 781535
rect 699992 781449 705525 781487
rect 699992 781393 700051 781449
rect 700107 781393 700193 781449
rect 700249 781393 700335 781449
rect 700391 781393 700477 781449
rect 700533 781393 700619 781449
rect 700675 781393 700761 781449
rect 700817 781393 700903 781449
rect 700959 781393 701045 781449
rect 701101 781393 701187 781449
rect 701243 781393 701329 781449
rect 701385 781393 701471 781449
rect 701527 781393 701613 781449
rect 701669 781393 701755 781449
rect 701811 781393 701897 781449
rect 701953 781431 705525 781449
rect 705581 781431 705649 781487
rect 705705 781431 705773 781487
rect 705829 781431 705897 781487
rect 705953 781431 706000 781487
rect 701953 781393 706000 781431
rect 699992 781363 706000 781393
rect 699992 781307 705525 781363
rect 705581 781307 705649 781363
rect 705705 781307 705773 781363
rect 705829 781307 705897 781363
rect 705953 781307 706000 781363
rect 699992 781251 700051 781307
rect 700107 781251 700193 781307
rect 700249 781251 700335 781307
rect 700391 781251 700477 781307
rect 700533 781251 700619 781307
rect 700675 781251 700761 781307
rect 700817 781251 700903 781307
rect 700959 781251 701045 781307
rect 701101 781251 701187 781307
rect 701243 781251 701329 781307
rect 701385 781251 701471 781307
rect 701527 781251 701613 781307
rect 701669 781251 701755 781307
rect 701811 781251 701897 781307
rect 701953 781251 706000 781307
rect 699992 781239 706000 781251
rect 699992 781183 705525 781239
rect 705581 781183 705649 781239
rect 705705 781183 705773 781239
rect 705829 781183 705897 781239
rect 705953 781183 706000 781239
rect 699992 781165 706000 781183
rect 699992 781109 700051 781165
rect 700107 781109 700193 781165
rect 700249 781109 700335 781165
rect 700391 781109 700477 781165
rect 700533 781109 700619 781165
rect 700675 781109 700761 781165
rect 700817 781109 700903 781165
rect 700959 781109 701045 781165
rect 701101 781109 701187 781165
rect 701243 781109 701329 781165
rect 701385 781109 701471 781165
rect 701527 781109 701613 781165
rect 701669 781109 701755 781165
rect 701811 781109 701897 781165
rect 701953 781115 706000 781165
rect 701953 781109 705525 781115
rect 699992 781059 705525 781109
rect 705581 781059 705649 781115
rect 705705 781059 705773 781115
rect 705829 781059 705897 781115
rect 705953 781059 706000 781115
rect 699992 781023 706000 781059
rect 699992 780967 700051 781023
rect 700107 780967 700193 781023
rect 700249 780967 700335 781023
rect 700391 780967 700477 781023
rect 700533 780967 700619 781023
rect 700675 780967 700761 781023
rect 700817 780967 700903 781023
rect 700959 780967 701045 781023
rect 701101 780967 701187 781023
rect 701243 780967 701329 781023
rect 701385 780967 701471 781023
rect 701527 780967 701613 781023
rect 701669 780967 701755 781023
rect 701811 780967 701897 781023
rect 701953 780991 706000 781023
rect 701953 780967 705525 780991
rect 699992 780935 705525 780967
rect 705581 780935 705649 780991
rect 705705 780935 705773 780991
rect 705829 780935 705897 780991
rect 705953 780935 706000 780991
rect 699992 780881 706000 780935
rect 699992 780825 700051 780881
rect 700107 780825 700193 780881
rect 700249 780825 700335 780881
rect 700391 780825 700477 780881
rect 700533 780825 700619 780881
rect 700675 780825 700761 780881
rect 700817 780825 700903 780881
rect 700959 780825 701045 780881
rect 701101 780825 701187 780881
rect 701243 780825 701329 780881
rect 701385 780825 701471 780881
rect 701527 780825 701613 780881
rect 701669 780825 701755 780881
rect 701811 780825 701897 780881
rect 701953 780867 706000 780881
rect 701953 780825 705525 780867
rect 699992 780811 705525 780825
rect 705581 780811 705649 780867
rect 705705 780811 705773 780867
rect 705829 780811 705897 780867
rect 705953 780811 706000 780867
rect 699992 780743 706000 780811
rect 699992 780739 705525 780743
rect 699992 780683 700051 780739
rect 700107 780683 700193 780739
rect 700249 780683 700335 780739
rect 700391 780683 700477 780739
rect 700533 780683 700619 780739
rect 700675 780683 700761 780739
rect 700817 780683 700903 780739
rect 700959 780683 701045 780739
rect 701101 780683 701187 780739
rect 701243 780683 701329 780739
rect 701385 780683 701471 780739
rect 701527 780683 701613 780739
rect 701669 780683 701755 780739
rect 701811 780683 701897 780739
rect 701953 780687 705525 780739
rect 705581 780687 705649 780743
rect 705705 780687 705773 780743
rect 705829 780687 705897 780743
rect 705953 780687 706000 780743
rect 701953 780683 706000 780687
rect 699992 780619 706000 780683
rect 699992 780597 705525 780619
rect 699992 780541 700051 780597
rect 700107 780541 700193 780597
rect 700249 780541 700335 780597
rect 700391 780541 700477 780597
rect 700533 780541 700619 780597
rect 700675 780541 700761 780597
rect 700817 780541 700903 780597
rect 700959 780541 701045 780597
rect 701101 780541 701187 780597
rect 701243 780541 701329 780597
rect 701385 780541 701471 780597
rect 701527 780541 701613 780597
rect 701669 780541 701755 780597
rect 701811 780541 701897 780597
rect 701953 780563 705525 780597
rect 705581 780563 705649 780619
rect 705705 780563 705773 780619
rect 705829 780563 705897 780619
rect 705953 780563 706000 780619
rect 701953 780541 706000 780563
rect 699992 780495 706000 780541
rect 699992 780455 705525 780495
rect 699992 780399 700051 780455
rect 700107 780399 700193 780455
rect 700249 780399 700335 780455
rect 700391 780399 700477 780455
rect 700533 780399 700619 780455
rect 700675 780399 700761 780455
rect 700817 780399 700903 780455
rect 700959 780399 701045 780455
rect 701101 780399 701187 780455
rect 701243 780399 701329 780455
rect 701385 780399 701471 780455
rect 701527 780399 701613 780455
rect 701669 780399 701755 780455
rect 701811 780399 701897 780455
rect 701953 780439 705525 780455
rect 705581 780439 705649 780495
rect 705705 780439 705773 780495
rect 705829 780439 705897 780495
rect 705953 780439 706000 780495
rect 701953 780399 706000 780439
rect 699992 780371 706000 780399
rect 699992 780315 705525 780371
rect 705581 780315 705649 780371
rect 705705 780315 705773 780371
rect 705829 780315 705897 780371
rect 705953 780315 706000 780371
rect 699992 780313 706000 780315
rect 699992 780257 700051 780313
rect 700107 780257 700193 780313
rect 700249 780257 700335 780313
rect 700391 780257 700477 780313
rect 700533 780257 700619 780313
rect 700675 780257 700761 780313
rect 700817 780257 700903 780313
rect 700959 780257 701045 780313
rect 701101 780257 701187 780313
rect 701243 780257 701329 780313
rect 701385 780257 701471 780313
rect 701527 780257 701613 780313
rect 701669 780257 701755 780313
rect 701811 780257 701897 780313
rect 701953 780257 706000 780313
rect 699992 780247 706000 780257
rect 699992 780191 705525 780247
rect 705581 780191 705649 780247
rect 705705 780191 705773 780247
rect 705829 780191 705897 780247
rect 705953 780191 706000 780247
rect 699992 780171 706000 780191
rect 699992 780115 700051 780171
rect 700107 780115 700193 780171
rect 700249 780115 700335 780171
rect 700391 780115 700477 780171
rect 700533 780115 700619 780171
rect 700675 780115 700761 780171
rect 700817 780115 700903 780171
rect 700959 780115 701045 780171
rect 701101 780115 701187 780171
rect 701243 780115 701329 780171
rect 701385 780115 701471 780171
rect 701527 780115 701613 780171
rect 701669 780115 701755 780171
rect 701811 780115 701897 780171
rect 701953 780123 706000 780171
rect 701953 780115 705525 780123
rect 699992 780067 705525 780115
rect 705581 780067 705649 780123
rect 705705 780067 705773 780123
rect 705829 780067 705897 780123
rect 705953 780067 706000 780123
rect 699992 780029 706000 780067
rect 699992 779973 700051 780029
rect 700107 779973 700193 780029
rect 700249 779973 700335 780029
rect 700391 779973 700477 780029
rect 700533 779973 700619 780029
rect 700675 779973 700761 780029
rect 700817 779973 700903 780029
rect 700959 779973 701045 780029
rect 701101 779973 701187 780029
rect 701243 779973 701329 780029
rect 701385 779973 701471 780029
rect 701527 779973 701613 780029
rect 701669 779973 701755 780029
rect 701811 779973 701897 780029
rect 701953 779999 706000 780029
rect 701953 779973 705525 779999
rect 699992 779943 705525 779973
rect 705581 779943 705649 779999
rect 705705 779943 705773 779999
rect 705829 779943 705897 779999
rect 705953 779943 706000 779999
rect 699992 779887 706000 779943
rect 699992 779831 700051 779887
rect 700107 779831 700193 779887
rect 700249 779831 700335 779887
rect 700391 779831 700477 779887
rect 700533 779831 700619 779887
rect 700675 779831 700761 779887
rect 700817 779831 700903 779887
rect 700959 779831 701045 779887
rect 701101 779831 701187 779887
rect 701243 779831 701329 779887
rect 701385 779831 701471 779887
rect 701527 779831 701613 779887
rect 701669 779831 701755 779887
rect 701811 779831 701897 779887
rect 701953 779875 706000 779887
rect 701953 779831 705525 779875
rect 699992 779819 705525 779831
rect 705581 779819 705649 779875
rect 705705 779819 705773 779875
rect 705829 779819 705897 779875
rect 705953 779819 706000 779875
rect 699992 779752 706000 779819
rect 699992 779131 706000 779172
rect 699992 779110 705525 779131
rect 699992 779054 700040 779110
rect 700096 779054 700182 779110
rect 700238 779054 700324 779110
rect 700380 779054 700466 779110
rect 700522 779054 700608 779110
rect 700664 779054 700750 779110
rect 700806 779054 700892 779110
rect 700948 779054 701034 779110
rect 701090 779054 701176 779110
rect 701232 779054 701318 779110
rect 701374 779054 701460 779110
rect 701516 779054 701602 779110
rect 701658 779054 701744 779110
rect 701800 779054 701886 779110
rect 701942 779075 705525 779110
rect 705581 779075 705649 779131
rect 705705 779075 705773 779131
rect 705829 779075 705897 779131
rect 705953 779075 706000 779131
rect 701942 779054 706000 779075
rect 699992 779007 706000 779054
rect 699992 778968 705525 779007
rect 699992 778912 700040 778968
rect 700096 778912 700182 778968
rect 700238 778912 700324 778968
rect 700380 778912 700466 778968
rect 700522 778912 700608 778968
rect 700664 778912 700750 778968
rect 700806 778912 700892 778968
rect 700948 778912 701034 778968
rect 701090 778912 701176 778968
rect 701232 778912 701318 778968
rect 701374 778912 701460 778968
rect 701516 778912 701602 778968
rect 701658 778912 701744 778968
rect 701800 778912 701886 778968
rect 701942 778951 705525 778968
rect 705581 778951 705649 779007
rect 705705 778951 705773 779007
rect 705829 778951 705897 779007
rect 705953 778951 706000 779007
rect 701942 778912 706000 778951
rect 699992 778883 706000 778912
rect 699992 778827 705525 778883
rect 705581 778827 705649 778883
rect 705705 778827 705773 778883
rect 705829 778827 705897 778883
rect 705953 778827 706000 778883
rect 699992 778826 706000 778827
rect 699992 778770 700040 778826
rect 700096 778770 700182 778826
rect 700238 778770 700324 778826
rect 700380 778770 700466 778826
rect 700522 778770 700608 778826
rect 700664 778770 700750 778826
rect 700806 778770 700892 778826
rect 700948 778770 701034 778826
rect 701090 778770 701176 778826
rect 701232 778770 701318 778826
rect 701374 778770 701460 778826
rect 701516 778770 701602 778826
rect 701658 778770 701744 778826
rect 701800 778770 701886 778826
rect 701942 778770 706000 778826
rect 699992 778759 706000 778770
rect 699992 778703 705525 778759
rect 705581 778703 705649 778759
rect 705705 778703 705773 778759
rect 705829 778703 705897 778759
rect 705953 778703 706000 778759
rect 699992 778684 706000 778703
rect 699992 778628 700040 778684
rect 700096 778628 700182 778684
rect 700238 778628 700324 778684
rect 700380 778628 700466 778684
rect 700522 778628 700608 778684
rect 700664 778628 700750 778684
rect 700806 778628 700892 778684
rect 700948 778628 701034 778684
rect 701090 778628 701176 778684
rect 701232 778628 701318 778684
rect 701374 778628 701460 778684
rect 701516 778628 701602 778684
rect 701658 778628 701744 778684
rect 701800 778628 701886 778684
rect 701942 778635 706000 778684
rect 701942 778628 705525 778635
rect 699992 778579 705525 778628
rect 705581 778579 705649 778635
rect 705705 778579 705773 778635
rect 705829 778579 705897 778635
rect 705953 778579 706000 778635
rect 699992 778542 706000 778579
rect 699992 778486 700040 778542
rect 700096 778486 700182 778542
rect 700238 778486 700324 778542
rect 700380 778486 700466 778542
rect 700522 778486 700608 778542
rect 700664 778486 700750 778542
rect 700806 778486 700892 778542
rect 700948 778486 701034 778542
rect 701090 778486 701176 778542
rect 701232 778486 701318 778542
rect 701374 778486 701460 778542
rect 701516 778486 701602 778542
rect 701658 778486 701744 778542
rect 701800 778486 701886 778542
rect 701942 778511 706000 778542
rect 701942 778486 705525 778511
rect 699992 778455 705525 778486
rect 705581 778455 705649 778511
rect 705705 778455 705773 778511
rect 705829 778455 705897 778511
rect 705953 778455 706000 778511
rect 699992 778400 706000 778455
rect 699992 778344 700040 778400
rect 700096 778344 700182 778400
rect 700238 778344 700324 778400
rect 700380 778344 700466 778400
rect 700522 778344 700608 778400
rect 700664 778344 700750 778400
rect 700806 778344 700892 778400
rect 700948 778344 701034 778400
rect 701090 778344 701176 778400
rect 701232 778344 701318 778400
rect 701374 778344 701460 778400
rect 701516 778344 701602 778400
rect 701658 778344 701744 778400
rect 701800 778344 701886 778400
rect 701942 778387 706000 778400
rect 701942 778344 705525 778387
rect 699992 778331 705525 778344
rect 705581 778331 705649 778387
rect 705705 778331 705773 778387
rect 705829 778331 705897 778387
rect 705953 778331 706000 778387
rect 699992 778263 706000 778331
rect 699992 778258 705525 778263
rect 699992 778202 700040 778258
rect 700096 778202 700182 778258
rect 700238 778202 700324 778258
rect 700380 778202 700466 778258
rect 700522 778202 700608 778258
rect 700664 778202 700750 778258
rect 700806 778202 700892 778258
rect 700948 778202 701034 778258
rect 701090 778202 701176 778258
rect 701232 778202 701318 778258
rect 701374 778202 701460 778258
rect 701516 778202 701602 778258
rect 701658 778202 701744 778258
rect 701800 778202 701886 778258
rect 701942 778207 705525 778258
rect 705581 778207 705649 778263
rect 705705 778207 705773 778263
rect 705829 778207 705897 778263
rect 705953 778207 706000 778263
rect 701942 778202 706000 778207
rect 699992 778139 706000 778202
rect 699992 778116 705525 778139
rect 699992 778060 700040 778116
rect 700096 778060 700182 778116
rect 700238 778060 700324 778116
rect 700380 778060 700466 778116
rect 700522 778060 700608 778116
rect 700664 778060 700750 778116
rect 700806 778060 700892 778116
rect 700948 778060 701034 778116
rect 701090 778060 701176 778116
rect 701232 778060 701318 778116
rect 701374 778060 701460 778116
rect 701516 778060 701602 778116
rect 701658 778060 701744 778116
rect 701800 778060 701886 778116
rect 701942 778083 705525 778116
rect 705581 778083 705649 778139
rect 705705 778083 705773 778139
rect 705829 778083 705897 778139
rect 705953 778083 706000 778139
rect 701942 778060 706000 778083
rect 699992 778015 706000 778060
rect 699992 777974 705525 778015
rect 699992 777918 700040 777974
rect 700096 777918 700182 777974
rect 700238 777918 700324 777974
rect 700380 777918 700466 777974
rect 700522 777918 700608 777974
rect 700664 777918 700750 777974
rect 700806 777918 700892 777974
rect 700948 777918 701034 777974
rect 701090 777918 701176 777974
rect 701232 777918 701318 777974
rect 701374 777918 701460 777974
rect 701516 777918 701602 777974
rect 701658 777918 701744 777974
rect 701800 777918 701886 777974
rect 701942 777959 705525 777974
rect 705581 777959 705649 778015
rect 705705 777959 705773 778015
rect 705829 777959 705897 778015
rect 705953 777959 706000 778015
rect 701942 777918 706000 777959
rect 699992 777891 706000 777918
rect 699992 777835 705525 777891
rect 705581 777835 705649 777891
rect 705705 777835 705773 777891
rect 705829 777835 705897 777891
rect 705953 777835 706000 777891
rect 699992 777832 706000 777835
rect 699992 777776 700040 777832
rect 700096 777776 700182 777832
rect 700238 777776 700324 777832
rect 700380 777776 700466 777832
rect 700522 777776 700608 777832
rect 700664 777776 700750 777832
rect 700806 777776 700892 777832
rect 700948 777776 701034 777832
rect 701090 777776 701176 777832
rect 701232 777776 701318 777832
rect 701374 777776 701460 777832
rect 701516 777776 701602 777832
rect 701658 777776 701744 777832
rect 701800 777776 701886 777832
rect 701942 777776 706000 777832
rect 699992 777767 706000 777776
rect 699992 777711 705525 777767
rect 705581 777711 705649 777767
rect 705705 777711 705773 777767
rect 705829 777711 705897 777767
rect 705953 777711 706000 777767
rect 699992 777690 706000 777711
rect 699992 777634 700040 777690
rect 700096 777634 700182 777690
rect 700238 777634 700324 777690
rect 700380 777634 700466 777690
rect 700522 777634 700608 777690
rect 700664 777634 700750 777690
rect 700806 777634 700892 777690
rect 700948 777634 701034 777690
rect 701090 777634 701176 777690
rect 701232 777634 701318 777690
rect 701374 777634 701460 777690
rect 701516 777634 701602 777690
rect 701658 777634 701744 777690
rect 701800 777634 701886 777690
rect 701942 777643 706000 777690
rect 701942 777634 705525 777643
rect 699992 777587 705525 777634
rect 705581 777587 705649 777643
rect 705705 777587 705773 777643
rect 705829 777587 705897 777643
rect 705953 777587 706000 777643
rect 699992 777548 706000 777587
rect 699992 777492 700040 777548
rect 700096 777492 700182 777548
rect 700238 777492 700324 777548
rect 700380 777492 700466 777548
rect 700522 777492 700608 777548
rect 700664 777492 700750 777548
rect 700806 777492 700892 777548
rect 700948 777492 701034 777548
rect 701090 777492 701176 777548
rect 701232 777492 701318 777548
rect 701374 777492 701460 777548
rect 701516 777492 701602 777548
rect 701658 777492 701744 777548
rect 701800 777492 701886 777548
rect 701942 777519 706000 777548
rect 701942 777492 705525 777519
rect 699992 777463 705525 777492
rect 705581 777463 705649 777519
rect 705705 777463 705773 777519
rect 705829 777463 705897 777519
rect 705953 777463 706000 777519
rect 699992 777406 706000 777463
rect 699992 777350 700040 777406
rect 700096 777350 700182 777406
rect 700238 777350 700324 777406
rect 700380 777350 700466 777406
rect 700522 777350 700608 777406
rect 700664 777350 700750 777406
rect 700806 777350 700892 777406
rect 700948 777350 701034 777406
rect 701090 777350 701176 777406
rect 701232 777350 701318 777406
rect 701374 777350 701460 777406
rect 701516 777350 701602 777406
rect 701658 777350 701744 777406
rect 701800 777350 701886 777406
rect 701942 777395 706000 777406
rect 701942 777350 705525 777395
rect 699992 777339 705525 777350
rect 705581 777339 705649 777395
rect 705705 777339 705773 777395
rect 705829 777339 705897 777395
rect 705953 777339 706000 777395
rect 699992 777272 706000 777339
rect 699992 490687 706000 490728
rect 699992 490666 705525 490687
rect 699992 490610 700040 490666
rect 700096 490610 700182 490666
rect 700238 490610 700324 490666
rect 700380 490610 700466 490666
rect 700522 490610 700608 490666
rect 700664 490610 700750 490666
rect 700806 490610 700892 490666
rect 700948 490610 701034 490666
rect 701090 490610 701176 490666
rect 701232 490610 701318 490666
rect 701374 490610 701460 490666
rect 701516 490610 701602 490666
rect 701658 490610 701744 490666
rect 701800 490610 701886 490666
rect 701942 490631 705525 490666
rect 705581 490631 705649 490687
rect 705705 490631 705773 490687
rect 705829 490631 705897 490687
rect 705953 490631 706000 490687
rect 701942 490610 706000 490631
rect 699992 490563 706000 490610
rect 699992 490524 705525 490563
rect 699992 490468 700040 490524
rect 700096 490468 700182 490524
rect 700238 490468 700324 490524
rect 700380 490468 700466 490524
rect 700522 490468 700608 490524
rect 700664 490468 700750 490524
rect 700806 490468 700892 490524
rect 700948 490468 701034 490524
rect 701090 490468 701176 490524
rect 701232 490468 701318 490524
rect 701374 490468 701460 490524
rect 701516 490468 701602 490524
rect 701658 490468 701744 490524
rect 701800 490468 701886 490524
rect 701942 490507 705525 490524
rect 705581 490507 705649 490563
rect 705705 490507 705773 490563
rect 705829 490507 705897 490563
rect 705953 490507 706000 490563
rect 701942 490468 706000 490507
rect 699992 490439 706000 490468
rect 699992 490383 705525 490439
rect 705581 490383 705649 490439
rect 705705 490383 705773 490439
rect 705829 490383 705897 490439
rect 705953 490383 706000 490439
rect 699992 490382 706000 490383
rect 699992 490326 700040 490382
rect 700096 490326 700182 490382
rect 700238 490326 700324 490382
rect 700380 490326 700466 490382
rect 700522 490326 700608 490382
rect 700664 490326 700750 490382
rect 700806 490326 700892 490382
rect 700948 490326 701034 490382
rect 701090 490326 701176 490382
rect 701232 490326 701318 490382
rect 701374 490326 701460 490382
rect 701516 490326 701602 490382
rect 701658 490326 701744 490382
rect 701800 490326 701886 490382
rect 701942 490326 706000 490382
rect 699992 490315 706000 490326
rect 699992 490259 705525 490315
rect 705581 490259 705649 490315
rect 705705 490259 705773 490315
rect 705829 490259 705897 490315
rect 705953 490259 706000 490315
rect 699992 490240 706000 490259
rect 699992 490184 700040 490240
rect 700096 490184 700182 490240
rect 700238 490184 700324 490240
rect 700380 490184 700466 490240
rect 700522 490184 700608 490240
rect 700664 490184 700750 490240
rect 700806 490184 700892 490240
rect 700948 490184 701034 490240
rect 701090 490184 701176 490240
rect 701232 490184 701318 490240
rect 701374 490184 701460 490240
rect 701516 490184 701602 490240
rect 701658 490184 701744 490240
rect 701800 490184 701886 490240
rect 701942 490191 706000 490240
rect 701942 490184 705525 490191
rect 699992 490135 705525 490184
rect 705581 490135 705649 490191
rect 705705 490135 705773 490191
rect 705829 490135 705897 490191
rect 705953 490135 706000 490191
rect 699992 490098 706000 490135
rect 699992 490042 700040 490098
rect 700096 490042 700182 490098
rect 700238 490042 700324 490098
rect 700380 490042 700466 490098
rect 700522 490042 700608 490098
rect 700664 490042 700750 490098
rect 700806 490042 700892 490098
rect 700948 490042 701034 490098
rect 701090 490042 701176 490098
rect 701232 490042 701318 490098
rect 701374 490042 701460 490098
rect 701516 490042 701602 490098
rect 701658 490042 701744 490098
rect 701800 490042 701886 490098
rect 701942 490067 706000 490098
rect 701942 490042 705525 490067
rect 699992 490011 705525 490042
rect 705581 490011 705649 490067
rect 705705 490011 705773 490067
rect 705829 490011 705897 490067
rect 705953 490011 706000 490067
rect 699992 489956 706000 490011
rect 699992 489900 700040 489956
rect 700096 489900 700182 489956
rect 700238 489900 700324 489956
rect 700380 489900 700466 489956
rect 700522 489900 700608 489956
rect 700664 489900 700750 489956
rect 700806 489900 700892 489956
rect 700948 489900 701034 489956
rect 701090 489900 701176 489956
rect 701232 489900 701318 489956
rect 701374 489900 701460 489956
rect 701516 489900 701602 489956
rect 701658 489900 701744 489956
rect 701800 489900 701886 489956
rect 701942 489943 706000 489956
rect 701942 489900 705525 489943
rect 699992 489887 705525 489900
rect 705581 489887 705649 489943
rect 705705 489887 705773 489943
rect 705829 489887 705897 489943
rect 705953 489887 706000 489943
rect 699992 489819 706000 489887
rect 699992 489814 705525 489819
rect 699992 489758 700040 489814
rect 700096 489758 700182 489814
rect 700238 489758 700324 489814
rect 700380 489758 700466 489814
rect 700522 489758 700608 489814
rect 700664 489758 700750 489814
rect 700806 489758 700892 489814
rect 700948 489758 701034 489814
rect 701090 489758 701176 489814
rect 701232 489758 701318 489814
rect 701374 489758 701460 489814
rect 701516 489758 701602 489814
rect 701658 489758 701744 489814
rect 701800 489758 701886 489814
rect 701942 489763 705525 489814
rect 705581 489763 705649 489819
rect 705705 489763 705773 489819
rect 705829 489763 705897 489819
rect 705953 489763 706000 489819
rect 701942 489758 706000 489763
rect 699992 489695 706000 489758
rect 699992 489672 705525 489695
rect 699992 489616 700040 489672
rect 700096 489616 700182 489672
rect 700238 489616 700324 489672
rect 700380 489616 700466 489672
rect 700522 489616 700608 489672
rect 700664 489616 700750 489672
rect 700806 489616 700892 489672
rect 700948 489616 701034 489672
rect 701090 489616 701176 489672
rect 701232 489616 701318 489672
rect 701374 489616 701460 489672
rect 701516 489616 701602 489672
rect 701658 489616 701744 489672
rect 701800 489616 701886 489672
rect 701942 489639 705525 489672
rect 705581 489639 705649 489695
rect 705705 489639 705773 489695
rect 705829 489639 705897 489695
rect 705953 489639 706000 489695
rect 701942 489616 706000 489639
rect 699992 489571 706000 489616
rect 699992 489530 705525 489571
rect 699992 489474 700040 489530
rect 700096 489474 700182 489530
rect 700238 489474 700324 489530
rect 700380 489474 700466 489530
rect 700522 489474 700608 489530
rect 700664 489474 700750 489530
rect 700806 489474 700892 489530
rect 700948 489474 701034 489530
rect 701090 489474 701176 489530
rect 701232 489474 701318 489530
rect 701374 489474 701460 489530
rect 701516 489474 701602 489530
rect 701658 489474 701744 489530
rect 701800 489474 701886 489530
rect 701942 489515 705525 489530
rect 705581 489515 705649 489571
rect 705705 489515 705773 489571
rect 705829 489515 705897 489571
rect 705953 489515 706000 489571
rect 701942 489474 706000 489515
rect 699992 489447 706000 489474
rect 699992 489391 705525 489447
rect 705581 489391 705649 489447
rect 705705 489391 705773 489447
rect 705829 489391 705897 489447
rect 705953 489391 706000 489447
rect 699992 489388 706000 489391
rect 699992 489332 700040 489388
rect 700096 489332 700182 489388
rect 700238 489332 700324 489388
rect 700380 489332 700466 489388
rect 700522 489332 700608 489388
rect 700664 489332 700750 489388
rect 700806 489332 700892 489388
rect 700948 489332 701034 489388
rect 701090 489332 701176 489388
rect 701232 489332 701318 489388
rect 701374 489332 701460 489388
rect 701516 489332 701602 489388
rect 701658 489332 701744 489388
rect 701800 489332 701886 489388
rect 701942 489332 706000 489388
rect 699992 489323 706000 489332
rect 699992 489267 705525 489323
rect 705581 489267 705649 489323
rect 705705 489267 705773 489323
rect 705829 489267 705897 489323
rect 705953 489267 706000 489323
rect 699992 489246 706000 489267
rect 699992 489190 700040 489246
rect 700096 489190 700182 489246
rect 700238 489190 700324 489246
rect 700380 489190 700466 489246
rect 700522 489190 700608 489246
rect 700664 489190 700750 489246
rect 700806 489190 700892 489246
rect 700948 489190 701034 489246
rect 701090 489190 701176 489246
rect 701232 489190 701318 489246
rect 701374 489190 701460 489246
rect 701516 489190 701602 489246
rect 701658 489190 701744 489246
rect 701800 489190 701886 489246
rect 701942 489199 706000 489246
rect 701942 489190 705525 489199
rect 699992 489143 705525 489190
rect 705581 489143 705649 489199
rect 705705 489143 705773 489199
rect 705829 489143 705897 489199
rect 705953 489143 706000 489199
rect 699992 489104 706000 489143
rect 699992 489048 700040 489104
rect 700096 489048 700182 489104
rect 700238 489048 700324 489104
rect 700380 489048 700466 489104
rect 700522 489048 700608 489104
rect 700664 489048 700750 489104
rect 700806 489048 700892 489104
rect 700948 489048 701034 489104
rect 701090 489048 701176 489104
rect 701232 489048 701318 489104
rect 701374 489048 701460 489104
rect 701516 489048 701602 489104
rect 701658 489048 701744 489104
rect 701800 489048 701886 489104
rect 701942 489075 706000 489104
rect 701942 489048 705525 489075
rect 699992 489019 705525 489048
rect 705581 489019 705649 489075
rect 705705 489019 705773 489075
rect 705829 489019 705897 489075
rect 705953 489019 706000 489075
rect 699992 488962 706000 489019
rect 699992 488906 700040 488962
rect 700096 488906 700182 488962
rect 700238 488906 700324 488962
rect 700380 488906 700466 488962
rect 700522 488906 700608 488962
rect 700664 488906 700750 488962
rect 700806 488906 700892 488962
rect 700948 488906 701034 488962
rect 701090 488906 701176 488962
rect 701232 488906 701318 488962
rect 701374 488906 701460 488962
rect 701516 488906 701602 488962
rect 701658 488906 701744 488962
rect 701800 488906 701886 488962
rect 701942 488951 706000 488962
rect 701942 488906 705525 488951
rect 699992 488895 705525 488906
rect 705581 488895 705649 488951
rect 705705 488895 705773 488951
rect 705829 488895 705897 488951
rect 705953 488895 706000 488951
rect 699992 488828 706000 488895
rect 699992 488181 706000 488248
rect 699992 488179 705525 488181
rect 699992 488123 700051 488179
rect 700107 488123 700193 488179
rect 700249 488123 700335 488179
rect 700391 488123 700477 488179
rect 700533 488123 700619 488179
rect 700675 488123 700761 488179
rect 700817 488123 700903 488179
rect 700959 488123 701045 488179
rect 701101 488123 701187 488179
rect 701243 488123 701329 488179
rect 701385 488123 701471 488179
rect 701527 488123 701613 488179
rect 701669 488123 701755 488179
rect 701811 488123 701897 488179
rect 701953 488125 705525 488179
rect 705581 488125 705649 488181
rect 705705 488125 705773 488181
rect 705829 488125 705897 488181
rect 705953 488125 706000 488181
rect 701953 488123 706000 488125
rect 699992 488057 706000 488123
rect 699992 488037 705525 488057
rect 699992 487981 700051 488037
rect 700107 487981 700193 488037
rect 700249 487981 700335 488037
rect 700391 487981 700477 488037
rect 700533 487981 700619 488037
rect 700675 487981 700761 488037
rect 700817 487981 700903 488037
rect 700959 487981 701045 488037
rect 701101 487981 701187 488037
rect 701243 487981 701329 488037
rect 701385 487981 701471 488037
rect 701527 487981 701613 488037
rect 701669 487981 701755 488037
rect 701811 487981 701897 488037
rect 701953 488001 705525 488037
rect 705581 488001 705649 488057
rect 705705 488001 705773 488057
rect 705829 488001 705897 488057
rect 705953 488001 706000 488057
rect 701953 487981 706000 488001
rect 699992 487933 706000 487981
rect 699992 487895 705525 487933
rect 699992 487839 700051 487895
rect 700107 487839 700193 487895
rect 700249 487839 700335 487895
rect 700391 487839 700477 487895
rect 700533 487839 700619 487895
rect 700675 487839 700761 487895
rect 700817 487839 700903 487895
rect 700959 487839 701045 487895
rect 701101 487839 701187 487895
rect 701243 487839 701329 487895
rect 701385 487839 701471 487895
rect 701527 487839 701613 487895
rect 701669 487839 701755 487895
rect 701811 487839 701897 487895
rect 701953 487877 705525 487895
rect 705581 487877 705649 487933
rect 705705 487877 705773 487933
rect 705829 487877 705897 487933
rect 705953 487877 706000 487933
rect 701953 487839 706000 487877
rect 699992 487809 706000 487839
rect 699992 487753 705525 487809
rect 705581 487753 705649 487809
rect 705705 487753 705773 487809
rect 705829 487753 705897 487809
rect 705953 487753 706000 487809
rect 699992 487697 700051 487753
rect 700107 487697 700193 487753
rect 700249 487697 700335 487753
rect 700391 487697 700477 487753
rect 700533 487697 700619 487753
rect 700675 487697 700761 487753
rect 700817 487697 700903 487753
rect 700959 487697 701045 487753
rect 701101 487697 701187 487753
rect 701243 487697 701329 487753
rect 701385 487697 701471 487753
rect 701527 487697 701613 487753
rect 701669 487697 701755 487753
rect 701811 487697 701897 487753
rect 701953 487697 706000 487753
rect 699992 487685 706000 487697
rect 699992 487629 705525 487685
rect 705581 487629 705649 487685
rect 705705 487629 705773 487685
rect 705829 487629 705897 487685
rect 705953 487629 706000 487685
rect 699992 487611 706000 487629
rect 699992 487555 700051 487611
rect 700107 487555 700193 487611
rect 700249 487555 700335 487611
rect 700391 487555 700477 487611
rect 700533 487555 700619 487611
rect 700675 487555 700761 487611
rect 700817 487555 700903 487611
rect 700959 487555 701045 487611
rect 701101 487555 701187 487611
rect 701243 487555 701329 487611
rect 701385 487555 701471 487611
rect 701527 487555 701613 487611
rect 701669 487555 701755 487611
rect 701811 487555 701897 487611
rect 701953 487561 706000 487611
rect 701953 487555 705525 487561
rect 699992 487505 705525 487555
rect 705581 487505 705649 487561
rect 705705 487505 705773 487561
rect 705829 487505 705897 487561
rect 705953 487505 706000 487561
rect 699992 487469 706000 487505
rect 699992 487413 700051 487469
rect 700107 487413 700193 487469
rect 700249 487413 700335 487469
rect 700391 487413 700477 487469
rect 700533 487413 700619 487469
rect 700675 487413 700761 487469
rect 700817 487413 700903 487469
rect 700959 487413 701045 487469
rect 701101 487413 701187 487469
rect 701243 487413 701329 487469
rect 701385 487413 701471 487469
rect 701527 487413 701613 487469
rect 701669 487413 701755 487469
rect 701811 487413 701897 487469
rect 701953 487437 706000 487469
rect 701953 487413 705525 487437
rect 699992 487381 705525 487413
rect 705581 487381 705649 487437
rect 705705 487381 705773 487437
rect 705829 487381 705897 487437
rect 705953 487381 706000 487437
rect 699992 487327 706000 487381
rect 699992 487271 700051 487327
rect 700107 487271 700193 487327
rect 700249 487271 700335 487327
rect 700391 487271 700477 487327
rect 700533 487271 700619 487327
rect 700675 487271 700761 487327
rect 700817 487271 700903 487327
rect 700959 487271 701045 487327
rect 701101 487271 701187 487327
rect 701243 487271 701329 487327
rect 701385 487271 701471 487327
rect 701527 487271 701613 487327
rect 701669 487271 701755 487327
rect 701811 487271 701897 487327
rect 701953 487313 706000 487327
rect 701953 487271 705525 487313
rect 699992 487257 705525 487271
rect 705581 487257 705649 487313
rect 705705 487257 705773 487313
rect 705829 487257 705897 487313
rect 705953 487257 706000 487313
rect 699992 487189 706000 487257
rect 699992 487185 705525 487189
rect 699992 487129 700051 487185
rect 700107 487129 700193 487185
rect 700249 487129 700335 487185
rect 700391 487129 700477 487185
rect 700533 487129 700619 487185
rect 700675 487129 700761 487185
rect 700817 487129 700903 487185
rect 700959 487129 701045 487185
rect 701101 487129 701187 487185
rect 701243 487129 701329 487185
rect 701385 487129 701471 487185
rect 701527 487129 701613 487185
rect 701669 487129 701755 487185
rect 701811 487129 701897 487185
rect 701953 487133 705525 487185
rect 705581 487133 705649 487189
rect 705705 487133 705773 487189
rect 705829 487133 705897 487189
rect 705953 487133 706000 487189
rect 701953 487129 706000 487133
rect 699992 487065 706000 487129
rect 699992 487043 705525 487065
rect 699992 486987 700051 487043
rect 700107 486987 700193 487043
rect 700249 486987 700335 487043
rect 700391 486987 700477 487043
rect 700533 486987 700619 487043
rect 700675 486987 700761 487043
rect 700817 486987 700903 487043
rect 700959 486987 701045 487043
rect 701101 486987 701187 487043
rect 701243 486987 701329 487043
rect 701385 486987 701471 487043
rect 701527 486987 701613 487043
rect 701669 486987 701755 487043
rect 701811 486987 701897 487043
rect 701953 487009 705525 487043
rect 705581 487009 705649 487065
rect 705705 487009 705773 487065
rect 705829 487009 705897 487065
rect 705953 487009 706000 487065
rect 701953 486987 706000 487009
rect 699992 486941 706000 486987
rect 699992 486901 705525 486941
rect 699992 486845 700051 486901
rect 700107 486845 700193 486901
rect 700249 486845 700335 486901
rect 700391 486845 700477 486901
rect 700533 486845 700619 486901
rect 700675 486845 700761 486901
rect 700817 486845 700903 486901
rect 700959 486845 701045 486901
rect 701101 486845 701187 486901
rect 701243 486845 701329 486901
rect 701385 486845 701471 486901
rect 701527 486845 701613 486901
rect 701669 486845 701755 486901
rect 701811 486845 701897 486901
rect 701953 486885 705525 486901
rect 705581 486885 705649 486941
rect 705705 486885 705773 486941
rect 705829 486885 705897 486941
rect 705953 486885 706000 486941
rect 701953 486845 706000 486885
rect 699992 486817 706000 486845
rect 699992 486761 705525 486817
rect 705581 486761 705649 486817
rect 705705 486761 705773 486817
rect 705829 486761 705897 486817
rect 705953 486761 706000 486817
rect 699992 486759 706000 486761
rect 699992 486703 700051 486759
rect 700107 486703 700193 486759
rect 700249 486703 700335 486759
rect 700391 486703 700477 486759
rect 700533 486703 700619 486759
rect 700675 486703 700761 486759
rect 700817 486703 700903 486759
rect 700959 486703 701045 486759
rect 701101 486703 701187 486759
rect 701243 486703 701329 486759
rect 701385 486703 701471 486759
rect 701527 486703 701613 486759
rect 701669 486703 701755 486759
rect 701811 486703 701897 486759
rect 701953 486703 706000 486759
rect 699992 486693 706000 486703
rect 699992 486637 705525 486693
rect 705581 486637 705649 486693
rect 705705 486637 705773 486693
rect 705829 486637 705897 486693
rect 705953 486637 706000 486693
rect 699992 486617 706000 486637
rect 699992 486561 700051 486617
rect 700107 486561 700193 486617
rect 700249 486561 700335 486617
rect 700391 486561 700477 486617
rect 700533 486561 700619 486617
rect 700675 486561 700761 486617
rect 700817 486561 700903 486617
rect 700959 486561 701045 486617
rect 701101 486561 701187 486617
rect 701243 486561 701329 486617
rect 701385 486561 701471 486617
rect 701527 486561 701613 486617
rect 701669 486561 701755 486617
rect 701811 486561 701897 486617
rect 701953 486569 706000 486617
rect 701953 486561 705525 486569
rect 699992 486513 705525 486561
rect 705581 486513 705649 486569
rect 705705 486513 705773 486569
rect 705829 486513 705897 486569
rect 705953 486513 706000 486569
rect 699992 486475 706000 486513
rect 699992 486419 700051 486475
rect 700107 486419 700193 486475
rect 700249 486419 700335 486475
rect 700391 486419 700477 486475
rect 700533 486419 700619 486475
rect 700675 486419 700761 486475
rect 700817 486419 700903 486475
rect 700959 486419 701045 486475
rect 701101 486419 701187 486475
rect 701243 486419 701329 486475
rect 701385 486419 701471 486475
rect 701527 486419 701613 486475
rect 701669 486419 701755 486475
rect 701811 486419 701897 486475
rect 701953 486445 706000 486475
rect 701953 486419 705525 486445
rect 699992 486389 705525 486419
rect 705581 486389 705649 486445
rect 705705 486389 705773 486445
rect 705829 486389 705897 486445
rect 705953 486389 706000 486445
rect 699992 486333 706000 486389
rect 699992 486277 700051 486333
rect 700107 486277 700193 486333
rect 700249 486277 700335 486333
rect 700391 486277 700477 486333
rect 700533 486277 700619 486333
rect 700675 486277 700761 486333
rect 700817 486277 700903 486333
rect 700959 486277 701045 486333
rect 701101 486277 701187 486333
rect 701243 486277 701329 486333
rect 701385 486277 701471 486333
rect 701527 486277 701613 486333
rect 701669 486277 701755 486333
rect 701811 486277 701897 486333
rect 701953 486321 706000 486333
rect 701953 486277 705525 486321
rect 699992 486265 705525 486277
rect 705581 486265 705649 486321
rect 705705 486265 705773 486321
rect 705829 486265 705897 486321
rect 705953 486265 706000 486321
rect 699992 486198 706000 486265
rect 699992 485811 706000 485878
rect 699992 485809 705525 485811
rect 699992 485753 700051 485809
rect 700107 485753 700193 485809
rect 700249 485753 700335 485809
rect 700391 485753 700477 485809
rect 700533 485753 700619 485809
rect 700675 485753 700761 485809
rect 700817 485753 700903 485809
rect 700959 485753 701045 485809
rect 701101 485753 701187 485809
rect 701243 485753 701329 485809
rect 701385 485753 701471 485809
rect 701527 485753 701613 485809
rect 701669 485753 701755 485809
rect 701811 485753 701897 485809
rect 701953 485755 705525 485809
rect 705581 485755 705649 485811
rect 705705 485755 705773 485811
rect 705829 485755 705897 485811
rect 705953 485755 706000 485811
rect 701953 485753 706000 485755
rect 699992 485687 706000 485753
rect 699992 485667 705525 485687
rect 699992 485611 700051 485667
rect 700107 485611 700193 485667
rect 700249 485611 700335 485667
rect 700391 485611 700477 485667
rect 700533 485611 700619 485667
rect 700675 485611 700761 485667
rect 700817 485611 700903 485667
rect 700959 485611 701045 485667
rect 701101 485611 701187 485667
rect 701243 485611 701329 485667
rect 701385 485611 701471 485667
rect 701527 485611 701613 485667
rect 701669 485611 701755 485667
rect 701811 485611 701897 485667
rect 701953 485631 705525 485667
rect 705581 485631 705649 485687
rect 705705 485631 705773 485687
rect 705829 485631 705897 485687
rect 705953 485631 706000 485687
rect 701953 485611 706000 485631
rect 699992 485563 706000 485611
rect 699992 485525 705525 485563
rect 699992 485469 700051 485525
rect 700107 485469 700193 485525
rect 700249 485469 700335 485525
rect 700391 485469 700477 485525
rect 700533 485469 700619 485525
rect 700675 485469 700761 485525
rect 700817 485469 700903 485525
rect 700959 485469 701045 485525
rect 701101 485469 701187 485525
rect 701243 485469 701329 485525
rect 701385 485469 701471 485525
rect 701527 485469 701613 485525
rect 701669 485469 701755 485525
rect 701811 485469 701897 485525
rect 701953 485507 705525 485525
rect 705581 485507 705649 485563
rect 705705 485507 705773 485563
rect 705829 485507 705897 485563
rect 705953 485507 706000 485563
rect 701953 485469 706000 485507
rect 699992 485439 706000 485469
rect 699992 485383 705525 485439
rect 705581 485383 705649 485439
rect 705705 485383 705773 485439
rect 705829 485383 705897 485439
rect 705953 485383 706000 485439
rect 699992 485327 700051 485383
rect 700107 485327 700193 485383
rect 700249 485327 700335 485383
rect 700391 485327 700477 485383
rect 700533 485327 700619 485383
rect 700675 485327 700761 485383
rect 700817 485327 700903 485383
rect 700959 485327 701045 485383
rect 701101 485327 701187 485383
rect 701243 485327 701329 485383
rect 701385 485327 701471 485383
rect 701527 485327 701613 485383
rect 701669 485327 701755 485383
rect 701811 485327 701897 485383
rect 701953 485327 706000 485383
rect 699992 485315 706000 485327
rect 699992 485259 705525 485315
rect 705581 485259 705649 485315
rect 705705 485259 705773 485315
rect 705829 485259 705897 485315
rect 705953 485259 706000 485315
rect 699992 485241 706000 485259
rect 699992 485185 700051 485241
rect 700107 485185 700193 485241
rect 700249 485185 700335 485241
rect 700391 485185 700477 485241
rect 700533 485185 700619 485241
rect 700675 485185 700761 485241
rect 700817 485185 700903 485241
rect 700959 485185 701045 485241
rect 701101 485185 701187 485241
rect 701243 485185 701329 485241
rect 701385 485185 701471 485241
rect 701527 485185 701613 485241
rect 701669 485185 701755 485241
rect 701811 485185 701897 485241
rect 701953 485191 706000 485241
rect 701953 485185 705525 485191
rect 699992 485135 705525 485185
rect 705581 485135 705649 485191
rect 705705 485135 705773 485191
rect 705829 485135 705897 485191
rect 705953 485135 706000 485191
rect 699992 485099 706000 485135
rect 699992 485043 700051 485099
rect 700107 485043 700193 485099
rect 700249 485043 700335 485099
rect 700391 485043 700477 485099
rect 700533 485043 700619 485099
rect 700675 485043 700761 485099
rect 700817 485043 700903 485099
rect 700959 485043 701045 485099
rect 701101 485043 701187 485099
rect 701243 485043 701329 485099
rect 701385 485043 701471 485099
rect 701527 485043 701613 485099
rect 701669 485043 701755 485099
rect 701811 485043 701897 485099
rect 701953 485067 706000 485099
rect 701953 485043 705525 485067
rect 699992 485011 705525 485043
rect 705581 485011 705649 485067
rect 705705 485011 705773 485067
rect 705829 485011 705897 485067
rect 705953 485011 706000 485067
rect 699992 484957 706000 485011
rect 699992 484901 700051 484957
rect 700107 484901 700193 484957
rect 700249 484901 700335 484957
rect 700391 484901 700477 484957
rect 700533 484901 700619 484957
rect 700675 484901 700761 484957
rect 700817 484901 700903 484957
rect 700959 484901 701045 484957
rect 701101 484901 701187 484957
rect 701243 484901 701329 484957
rect 701385 484901 701471 484957
rect 701527 484901 701613 484957
rect 701669 484901 701755 484957
rect 701811 484901 701897 484957
rect 701953 484943 706000 484957
rect 701953 484901 705525 484943
rect 699992 484887 705525 484901
rect 705581 484887 705649 484943
rect 705705 484887 705773 484943
rect 705829 484887 705897 484943
rect 705953 484887 706000 484943
rect 699992 484819 706000 484887
rect 699992 484815 705525 484819
rect 699992 484759 700051 484815
rect 700107 484759 700193 484815
rect 700249 484759 700335 484815
rect 700391 484759 700477 484815
rect 700533 484759 700619 484815
rect 700675 484759 700761 484815
rect 700817 484759 700903 484815
rect 700959 484759 701045 484815
rect 701101 484759 701187 484815
rect 701243 484759 701329 484815
rect 701385 484759 701471 484815
rect 701527 484759 701613 484815
rect 701669 484759 701755 484815
rect 701811 484759 701897 484815
rect 701953 484763 705525 484815
rect 705581 484763 705649 484819
rect 705705 484763 705773 484819
rect 705829 484763 705897 484819
rect 705953 484763 706000 484819
rect 701953 484759 706000 484763
rect 699992 484695 706000 484759
rect 699992 484673 705525 484695
rect 699992 484617 700051 484673
rect 700107 484617 700193 484673
rect 700249 484617 700335 484673
rect 700391 484617 700477 484673
rect 700533 484617 700619 484673
rect 700675 484617 700761 484673
rect 700817 484617 700903 484673
rect 700959 484617 701045 484673
rect 701101 484617 701187 484673
rect 701243 484617 701329 484673
rect 701385 484617 701471 484673
rect 701527 484617 701613 484673
rect 701669 484617 701755 484673
rect 701811 484617 701897 484673
rect 701953 484639 705525 484673
rect 705581 484639 705649 484695
rect 705705 484639 705773 484695
rect 705829 484639 705897 484695
rect 705953 484639 706000 484695
rect 701953 484617 706000 484639
rect 699992 484571 706000 484617
rect 699992 484531 705525 484571
rect 699992 484475 700051 484531
rect 700107 484475 700193 484531
rect 700249 484475 700335 484531
rect 700391 484475 700477 484531
rect 700533 484475 700619 484531
rect 700675 484475 700761 484531
rect 700817 484475 700903 484531
rect 700959 484475 701045 484531
rect 701101 484475 701187 484531
rect 701243 484475 701329 484531
rect 701385 484475 701471 484531
rect 701527 484475 701613 484531
rect 701669 484475 701755 484531
rect 701811 484475 701897 484531
rect 701953 484515 705525 484531
rect 705581 484515 705649 484571
rect 705705 484515 705773 484571
rect 705829 484515 705897 484571
rect 705953 484515 706000 484571
rect 701953 484475 706000 484515
rect 699992 484447 706000 484475
rect 699992 484391 705525 484447
rect 705581 484391 705649 484447
rect 705705 484391 705773 484447
rect 705829 484391 705897 484447
rect 705953 484391 706000 484447
rect 699992 484389 706000 484391
rect 699992 484333 700051 484389
rect 700107 484333 700193 484389
rect 700249 484333 700335 484389
rect 700391 484333 700477 484389
rect 700533 484333 700619 484389
rect 700675 484333 700761 484389
rect 700817 484333 700903 484389
rect 700959 484333 701045 484389
rect 701101 484333 701187 484389
rect 701243 484333 701329 484389
rect 701385 484333 701471 484389
rect 701527 484333 701613 484389
rect 701669 484333 701755 484389
rect 701811 484333 701897 484389
rect 701953 484333 706000 484389
rect 699992 484323 706000 484333
rect 699992 484267 705525 484323
rect 705581 484267 705649 484323
rect 705705 484267 705773 484323
rect 705829 484267 705897 484323
rect 705953 484267 706000 484323
rect 699992 484247 706000 484267
rect 699992 484191 700051 484247
rect 700107 484191 700193 484247
rect 700249 484191 700335 484247
rect 700391 484191 700477 484247
rect 700533 484191 700619 484247
rect 700675 484191 700761 484247
rect 700817 484191 700903 484247
rect 700959 484191 701045 484247
rect 701101 484191 701187 484247
rect 701243 484191 701329 484247
rect 701385 484191 701471 484247
rect 701527 484191 701613 484247
rect 701669 484191 701755 484247
rect 701811 484191 701897 484247
rect 701953 484199 706000 484247
rect 701953 484191 705525 484199
rect 699992 484143 705525 484191
rect 705581 484143 705649 484199
rect 705705 484143 705773 484199
rect 705829 484143 705897 484199
rect 705953 484143 706000 484199
rect 699992 484105 706000 484143
rect 699992 484049 700051 484105
rect 700107 484049 700193 484105
rect 700249 484049 700335 484105
rect 700391 484049 700477 484105
rect 700533 484049 700619 484105
rect 700675 484049 700761 484105
rect 700817 484049 700903 484105
rect 700959 484049 701045 484105
rect 701101 484049 701187 484105
rect 701243 484049 701329 484105
rect 701385 484049 701471 484105
rect 701527 484049 701613 484105
rect 701669 484049 701755 484105
rect 701811 484049 701897 484105
rect 701953 484075 706000 484105
rect 701953 484049 705525 484075
rect 699992 484019 705525 484049
rect 705581 484019 705649 484075
rect 705705 484019 705773 484075
rect 705829 484019 705897 484075
rect 705953 484019 706000 484075
rect 699992 483963 706000 484019
rect 699992 483907 700051 483963
rect 700107 483907 700193 483963
rect 700249 483907 700335 483963
rect 700391 483907 700477 483963
rect 700533 483907 700619 483963
rect 700675 483907 700761 483963
rect 700817 483907 700903 483963
rect 700959 483907 701045 483963
rect 701101 483907 701187 483963
rect 701243 483907 701329 483963
rect 701385 483907 701471 483963
rect 701527 483907 701613 483963
rect 701669 483907 701755 483963
rect 701811 483907 701897 483963
rect 701953 483951 706000 483963
rect 701953 483907 705525 483951
rect 699992 483895 705525 483907
rect 705581 483895 705649 483951
rect 705705 483895 705773 483951
rect 705829 483895 705897 483951
rect 705953 483895 706000 483951
rect 699992 483828 706000 483895
rect 699992 483105 706000 483172
rect 699992 483103 705525 483105
rect 699992 483047 700051 483103
rect 700107 483047 700193 483103
rect 700249 483047 700335 483103
rect 700391 483047 700477 483103
rect 700533 483047 700619 483103
rect 700675 483047 700761 483103
rect 700817 483047 700903 483103
rect 700959 483047 701045 483103
rect 701101 483047 701187 483103
rect 701243 483047 701329 483103
rect 701385 483047 701471 483103
rect 701527 483047 701613 483103
rect 701669 483047 701755 483103
rect 701811 483047 701897 483103
rect 701953 483049 705525 483103
rect 705581 483049 705649 483105
rect 705705 483049 705773 483105
rect 705829 483049 705897 483105
rect 705953 483049 706000 483105
rect 701953 483047 706000 483049
rect 699992 482981 706000 483047
rect 699992 482961 705525 482981
rect 699992 482905 700051 482961
rect 700107 482905 700193 482961
rect 700249 482905 700335 482961
rect 700391 482905 700477 482961
rect 700533 482905 700619 482961
rect 700675 482905 700761 482961
rect 700817 482905 700903 482961
rect 700959 482905 701045 482961
rect 701101 482905 701187 482961
rect 701243 482905 701329 482961
rect 701385 482905 701471 482961
rect 701527 482905 701613 482961
rect 701669 482905 701755 482961
rect 701811 482905 701897 482961
rect 701953 482925 705525 482961
rect 705581 482925 705649 482981
rect 705705 482925 705773 482981
rect 705829 482925 705897 482981
rect 705953 482925 706000 482981
rect 701953 482905 706000 482925
rect 699992 482857 706000 482905
rect 699992 482819 705525 482857
rect 699992 482763 700051 482819
rect 700107 482763 700193 482819
rect 700249 482763 700335 482819
rect 700391 482763 700477 482819
rect 700533 482763 700619 482819
rect 700675 482763 700761 482819
rect 700817 482763 700903 482819
rect 700959 482763 701045 482819
rect 701101 482763 701187 482819
rect 701243 482763 701329 482819
rect 701385 482763 701471 482819
rect 701527 482763 701613 482819
rect 701669 482763 701755 482819
rect 701811 482763 701897 482819
rect 701953 482801 705525 482819
rect 705581 482801 705649 482857
rect 705705 482801 705773 482857
rect 705829 482801 705897 482857
rect 705953 482801 706000 482857
rect 701953 482763 706000 482801
rect 699992 482733 706000 482763
rect 699992 482677 705525 482733
rect 705581 482677 705649 482733
rect 705705 482677 705773 482733
rect 705829 482677 705897 482733
rect 705953 482677 706000 482733
rect 699992 482621 700051 482677
rect 700107 482621 700193 482677
rect 700249 482621 700335 482677
rect 700391 482621 700477 482677
rect 700533 482621 700619 482677
rect 700675 482621 700761 482677
rect 700817 482621 700903 482677
rect 700959 482621 701045 482677
rect 701101 482621 701187 482677
rect 701243 482621 701329 482677
rect 701385 482621 701471 482677
rect 701527 482621 701613 482677
rect 701669 482621 701755 482677
rect 701811 482621 701897 482677
rect 701953 482621 706000 482677
rect 699992 482609 706000 482621
rect 699992 482553 705525 482609
rect 705581 482553 705649 482609
rect 705705 482553 705773 482609
rect 705829 482553 705897 482609
rect 705953 482553 706000 482609
rect 699992 482535 706000 482553
rect 699992 482479 700051 482535
rect 700107 482479 700193 482535
rect 700249 482479 700335 482535
rect 700391 482479 700477 482535
rect 700533 482479 700619 482535
rect 700675 482479 700761 482535
rect 700817 482479 700903 482535
rect 700959 482479 701045 482535
rect 701101 482479 701187 482535
rect 701243 482479 701329 482535
rect 701385 482479 701471 482535
rect 701527 482479 701613 482535
rect 701669 482479 701755 482535
rect 701811 482479 701897 482535
rect 701953 482485 706000 482535
rect 701953 482479 705525 482485
rect 699992 482429 705525 482479
rect 705581 482429 705649 482485
rect 705705 482429 705773 482485
rect 705829 482429 705897 482485
rect 705953 482429 706000 482485
rect 699992 482393 706000 482429
rect 699992 482337 700051 482393
rect 700107 482337 700193 482393
rect 700249 482337 700335 482393
rect 700391 482337 700477 482393
rect 700533 482337 700619 482393
rect 700675 482337 700761 482393
rect 700817 482337 700903 482393
rect 700959 482337 701045 482393
rect 701101 482337 701187 482393
rect 701243 482337 701329 482393
rect 701385 482337 701471 482393
rect 701527 482337 701613 482393
rect 701669 482337 701755 482393
rect 701811 482337 701897 482393
rect 701953 482361 706000 482393
rect 701953 482337 705525 482361
rect 699992 482305 705525 482337
rect 705581 482305 705649 482361
rect 705705 482305 705773 482361
rect 705829 482305 705897 482361
rect 705953 482305 706000 482361
rect 699992 482251 706000 482305
rect 699992 482195 700051 482251
rect 700107 482195 700193 482251
rect 700249 482195 700335 482251
rect 700391 482195 700477 482251
rect 700533 482195 700619 482251
rect 700675 482195 700761 482251
rect 700817 482195 700903 482251
rect 700959 482195 701045 482251
rect 701101 482195 701187 482251
rect 701243 482195 701329 482251
rect 701385 482195 701471 482251
rect 701527 482195 701613 482251
rect 701669 482195 701755 482251
rect 701811 482195 701897 482251
rect 701953 482237 706000 482251
rect 701953 482195 705525 482237
rect 699992 482181 705525 482195
rect 705581 482181 705649 482237
rect 705705 482181 705773 482237
rect 705829 482181 705897 482237
rect 705953 482181 706000 482237
rect 699992 482113 706000 482181
rect 699992 482109 705525 482113
rect 699992 482053 700051 482109
rect 700107 482053 700193 482109
rect 700249 482053 700335 482109
rect 700391 482053 700477 482109
rect 700533 482053 700619 482109
rect 700675 482053 700761 482109
rect 700817 482053 700903 482109
rect 700959 482053 701045 482109
rect 701101 482053 701187 482109
rect 701243 482053 701329 482109
rect 701385 482053 701471 482109
rect 701527 482053 701613 482109
rect 701669 482053 701755 482109
rect 701811 482053 701897 482109
rect 701953 482057 705525 482109
rect 705581 482057 705649 482113
rect 705705 482057 705773 482113
rect 705829 482057 705897 482113
rect 705953 482057 706000 482113
rect 701953 482053 706000 482057
rect 699992 481989 706000 482053
rect 699992 481967 705525 481989
rect 699992 481911 700051 481967
rect 700107 481911 700193 481967
rect 700249 481911 700335 481967
rect 700391 481911 700477 481967
rect 700533 481911 700619 481967
rect 700675 481911 700761 481967
rect 700817 481911 700903 481967
rect 700959 481911 701045 481967
rect 701101 481911 701187 481967
rect 701243 481911 701329 481967
rect 701385 481911 701471 481967
rect 701527 481911 701613 481967
rect 701669 481911 701755 481967
rect 701811 481911 701897 481967
rect 701953 481933 705525 481967
rect 705581 481933 705649 481989
rect 705705 481933 705773 481989
rect 705829 481933 705897 481989
rect 705953 481933 706000 481989
rect 701953 481911 706000 481933
rect 699992 481865 706000 481911
rect 699992 481825 705525 481865
rect 699992 481769 700051 481825
rect 700107 481769 700193 481825
rect 700249 481769 700335 481825
rect 700391 481769 700477 481825
rect 700533 481769 700619 481825
rect 700675 481769 700761 481825
rect 700817 481769 700903 481825
rect 700959 481769 701045 481825
rect 701101 481769 701187 481825
rect 701243 481769 701329 481825
rect 701385 481769 701471 481825
rect 701527 481769 701613 481825
rect 701669 481769 701755 481825
rect 701811 481769 701897 481825
rect 701953 481809 705525 481825
rect 705581 481809 705649 481865
rect 705705 481809 705773 481865
rect 705829 481809 705897 481865
rect 705953 481809 706000 481865
rect 701953 481769 706000 481809
rect 699992 481741 706000 481769
rect 699992 481685 705525 481741
rect 705581 481685 705649 481741
rect 705705 481685 705773 481741
rect 705829 481685 705897 481741
rect 705953 481685 706000 481741
rect 699992 481683 706000 481685
rect 699992 481627 700051 481683
rect 700107 481627 700193 481683
rect 700249 481627 700335 481683
rect 700391 481627 700477 481683
rect 700533 481627 700619 481683
rect 700675 481627 700761 481683
rect 700817 481627 700903 481683
rect 700959 481627 701045 481683
rect 701101 481627 701187 481683
rect 701243 481627 701329 481683
rect 701385 481627 701471 481683
rect 701527 481627 701613 481683
rect 701669 481627 701755 481683
rect 701811 481627 701897 481683
rect 701953 481627 706000 481683
rect 699992 481617 706000 481627
rect 699992 481561 705525 481617
rect 705581 481561 705649 481617
rect 705705 481561 705773 481617
rect 705829 481561 705897 481617
rect 705953 481561 706000 481617
rect 699992 481541 706000 481561
rect 699992 481485 700051 481541
rect 700107 481485 700193 481541
rect 700249 481485 700335 481541
rect 700391 481485 700477 481541
rect 700533 481485 700619 481541
rect 700675 481485 700761 481541
rect 700817 481485 700903 481541
rect 700959 481485 701045 481541
rect 701101 481485 701187 481541
rect 701243 481485 701329 481541
rect 701385 481485 701471 481541
rect 701527 481485 701613 481541
rect 701669 481485 701755 481541
rect 701811 481485 701897 481541
rect 701953 481493 706000 481541
rect 701953 481485 705525 481493
rect 699992 481437 705525 481485
rect 705581 481437 705649 481493
rect 705705 481437 705773 481493
rect 705829 481437 705897 481493
rect 705953 481437 706000 481493
rect 699992 481399 706000 481437
rect 699992 481343 700051 481399
rect 700107 481343 700193 481399
rect 700249 481343 700335 481399
rect 700391 481343 700477 481399
rect 700533 481343 700619 481399
rect 700675 481343 700761 481399
rect 700817 481343 700903 481399
rect 700959 481343 701045 481399
rect 701101 481343 701187 481399
rect 701243 481343 701329 481399
rect 701385 481343 701471 481399
rect 701527 481343 701613 481399
rect 701669 481343 701755 481399
rect 701811 481343 701897 481399
rect 701953 481369 706000 481399
rect 701953 481343 705525 481369
rect 699992 481313 705525 481343
rect 705581 481313 705649 481369
rect 705705 481313 705773 481369
rect 705829 481313 705897 481369
rect 705953 481313 706000 481369
rect 699992 481257 706000 481313
rect 699992 481201 700051 481257
rect 700107 481201 700193 481257
rect 700249 481201 700335 481257
rect 700391 481201 700477 481257
rect 700533 481201 700619 481257
rect 700675 481201 700761 481257
rect 700817 481201 700903 481257
rect 700959 481201 701045 481257
rect 701101 481201 701187 481257
rect 701243 481201 701329 481257
rect 701385 481201 701471 481257
rect 701527 481201 701613 481257
rect 701669 481201 701755 481257
rect 701811 481201 701897 481257
rect 701953 481245 706000 481257
rect 701953 481201 705525 481245
rect 699992 481189 705525 481201
rect 705581 481189 705649 481245
rect 705705 481189 705773 481245
rect 705829 481189 705897 481245
rect 705953 481189 706000 481245
rect 699992 481122 706000 481189
rect 699992 480735 706000 480802
rect 699992 480733 705525 480735
rect 699992 480677 700051 480733
rect 700107 480677 700193 480733
rect 700249 480677 700335 480733
rect 700391 480677 700477 480733
rect 700533 480677 700619 480733
rect 700675 480677 700761 480733
rect 700817 480677 700903 480733
rect 700959 480677 701045 480733
rect 701101 480677 701187 480733
rect 701243 480677 701329 480733
rect 701385 480677 701471 480733
rect 701527 480677 701613 480733
rect 701669 480677 701755 480733
rect 701811 480677 701897 480733
rect 701953 480679 705525 480733
rect 705581 480679 705649 480735
rect 705705 480679 705773 480735
rect 705829 480679 705897 480735
rect 705953 480679 706000 480735
rect 701953 480677 706000 480679
rect 699992 480611 706000 480677
rect 699992 480591 705525 480611
rect 699992 480535 700051 480591
rect 700107 480535 700193 480591
rect 700249 480535 700335 480591
rect 700391 480535 700477 480591
rect 700533 480535 700619 480591
rect 700675 480535 700761 480591
rect 700817 480535 700903 480591
rect 700959 480535 701045 480591
rect 701101 480535 701187 480591
rect 701243 480535 701329 480591
rect 701385 480535 701471 480591
rect 701527 480535 701613 480591
rect 701669 480535 701755 480591
rect 701811 480535 701897 480591
rect 701953 480555 705525 480591
rect 705581 480555 705649 480611
rect 705705 480555 705773 480611
rect 705829 480555 705897 480611
rect 705953 480555 706000 480611
rect 701953 480535 706000 480555
rect 699992 480487 706000 480535
rect 699992 480449 705525 480487
rect 699992 480393 700051 480449
rect 700107 480393 700193 480449
rect 700249 480393 700335 480449
rect 700391 480393 700477 480449
rect 700533 480393 700619 480449
rect 700675 480393 700761 480449
rect 700817 480393 700903 480449
rect 700959 480393 701045 480449
rect 701101 480393 701187 480449
rect 701243 480393 701329 480449
rect 701385 480393 701471 480449
rect 701527 480393 701613 480449
rect 701669 480393 701755 480449
rect 701811 480393 701897 480449
rect 701953 480431 705525 480449
rect 705581 480431 705649 480487
rect 705705 480431 705773 480487
rect 705829 480431 705897 480487
rect 705953 480431 706000 480487
rect 701953 480393 706000 480431
rect 699992 480363 706000 480393
rect 699992 480307 705525 480363
rect 705581 480307 705649 480363
rect 705705 480307 705773 480363
rect 705829 480307 705897 480363
rect 705953 480307 706000 480363
rect 699992 480251 700051 480307
rect 700107 480251 700193 480307
rect 700249 480251 700335 480307
rect 700391 480251 700477 480307
rect 700533 480251 700619 480307
rect 700675 480251 700761 480307
rect 700817 480251 700903 480307
rect 700959 480251 701045 480307
rect 701101 480251 701187 480307
rect 701243 480251 701329 480307
rect 701385 480251 701471 480307
rect 701527 480251 701613 480307
rect 701669 480251 701755 480307
rect 701811 480251 701897 480307
rect 701953 480251 706000 480307
rect 699992 480239 706000 480251
rect 699992 480183 705525 480239
rect 705581 480183 705649 480239
rect 705705 480183 705773 480239
rect 705829 480183 705897 480239
rect 705953 480183 706000 480239
rect 699992 480165 706000 480183
rect 699992 480109 700051 480165
rect 700107 480109 700193 480165
rect 700249 480109 700335 480165
rect 700391 480109 700477 480165
rect 700533 480109 700619 480165
rect 700675 480109 700761 480165
rect 700817 480109 700903 480165
rect 700959 480109 701045 480165
rect 701101 480109 701187 480165
rect 701243 480109 701329 480165
rect 701385 480109 701471 480165
rect 701527 480109 701613 480165
rect 701669 480109 701755 480165
rect 701811 480109 701897 480165
rect 701953 480115 706000 480165
rect 701953 480109 705525 480115
rect 699992 480059 705525 480109
rect 705581 480059 705649 480115
rect 705705 480059 705773 480115
rect 705829 480059 705897 480115
rect 705953 480059 706000 480115
rect 699992 480023 706000 480059
rect 699992 479967 700051 480023
rect 700107 479967 700193 480023
rect 700249 479967 700335 480023
rect 700391 479967 700477 480023
rect 700533 479967 700619 480023
rect 700675 479967 700761 480023
rect 700817 479967 700903 480023
rect 700959 479967 701045 480023
rect 701101 479967 701187 480023
rect 701243 479967 701329 480023
rect 701385 479967 701471 480023
rect 701527 479967 701613 480023
rect 701669 479967 701755 480023
rect 701811 479967 701897 480023
rect 701953 479991 706000 480023
rect 701953 479967 705525 479991
rect 699992 479935 705525 479967
rect 705581 479935 705649 479991
rect 705705 479935 705773 479991
rect 705829 479935 705897 479991
rect 705953 479935 706000 479991
rect 699992 479881 706000 479935
rect 699992 479825 700051 479881
rect 700107 479825 700193 479881
rect 700249 479825 700335 479881
rect 700391 479825 700477 479881
rect 700533 479825 700619 479881
rect 700675 479825 700761 479881
rect 700817 479825 700903 479881
rect 700959 479825 701045 479881
rect 701101 479825 701187 479881
rect 701243 479825 701329 479881
rect 701385 479825 701471 479881
rect 701527 479825 701613 479881
rect 701669 479825 701755 479881
rect 701811 479825 701897 479881
rect 701953 479867 706000 479881
rect 701953 479825 705525 479867
rect 699992 479811 705525 479825
rect 705581 479811 705649 479867
rect 705705 479811 705773 479867
rect 705829 479811 705897 479867
rect 705953 479811 706000 479867
rect 699992 479743 706000 479811
rect 699992 479739 705525 479743
rect 699992 479683 700051 479739
rect 700107 479683 700193 479739
rect 700249 479683 700335 479739
rect 700391 479683 700477 479739
rect 700533 479683 700619 479739
rect 700675 479683 700761 479739
rect 700817 479683 700903 479739
rect 700959 479683 701045 479739
rect 701101 479683 701187 479739
rect 701243 479683 701329 479739
rect 701385 479683 701471 479739
rect 701527 479683 701613 479739
rect 701669 479683 701755 479739
rect 701811 479683 701897 479739
rect 701953 479687 705525 479739
rect 705581 479687 705649 479743
rect 705705 479687 705773 479743
rect 705829 479687 705897 479743
rect 705953 479687 706000 479743
rect 701953 479683 706000 479687
rect 699992 479619 706000 479683
rect 699992 479597 705525 479619
rect 699992 479541 700051 479597
rect 700107 479541 700193 479597
rect 700249 479541 700335 479597
rect 700391 479541 700477 479597
rect 700533 479541 700619 479597
rect 700675 479541 700761 479597
rect 700817 479541 700903 479597
rect 700959 479541 701045 479597
rect 701101 479541 701187 479597
rect 701243 479541 701329 479597
rect 701385 479541 701471 479597
rect 701527 479541 701613 479597
rect 701669 479541 701755 479597
rect 701811 479541 701897 479597
rect 701953 479563 705525 479597
rect 705581 479563 705649 479619
rect 705705 479563 705773 479619
rect 705829 479563 705897 479619
rect 705953 479563 706000 479619
rect 701953 479541 706000 479563
rect 699992 479495 706000 479541
rect 699992 479455 705525 479495
rect 699992 479399 700051 479455
rect 700107 479399 700193 479455
rect 700249 479399 700335 479455
rect 700391 479399 700477 479455
rect 700533 479399 700619 479455
rect 700675 479399 700761 479455
rect 700817 479399 700903 479455
rect 700959 479399 701045 479455
rect 701101 479399 701187 479455
rect 701243 479399 701329 479455
rect 701385 479399 701471 479455
rect 701527 479399 701613 479455
rect 701669 479399 701755 479455
rect 701811 479399 701897 479455
rect 701953 479439 705525 479455
rect 705581 479439 705649 479495
rect 705705 479439 705773 479495
rect 705829 479439 705897 479495
rect 705953 479439 706000 479495
rect 701953 479399 706000 479439
rect 699992 479371 706000 479399
rect 699992 479315 705525 479371
rect 705581 479315 705649 479371
rect 705705 479315 705773 479371
rect 705829 479315 705897 479371
rect 705953 479315 706000 479371
rect 699992 479313 706000 479315
rect 699992 479257 700051 479313
rect 700107 479257 700193 479313
rect 700249 479257 700335 479313
rect 700391 479257 700477 479313
rect 700533 479257 700619 479313
rect 700675 479257 700761 479313
rect 700817 479257 700903 479313
rect 700959 479257 701045 479313
rect 701101 479257 701187 479313
rect 701243 479257 701329 479313
rect 701385 479257 701471 479313
rect 701527 479257 701613 479313
rect 701669 479257 701755 479313
rect 701811 479257 701897 479313
rect 701953 479257 706000 479313
rect 699992 479247 706000 479257
rect 699992 479191 705525 479247
rect 705581 479191 705649 479247
rect 705705 479191 705773 479247
rect 705829 479191 705897 479247
rect 705953 479191 706000 479247
rect 699992 479171 706000 479191
rect 699992 479115 700051 479171
rect 700107 479115 700193 479171
rect 700249 479115 700335 479171
rect 700391 479115 700477 479171
rect 700533 479115 700619 479171
rect 700675 479115 700761 479171
rect 700817 479115 700903 479171
rect 700959 479115 701045 479171
rect 701101 479115 701187 479171
rect 701243 479115 701329 479171
rect 701385 479115 701471 479171
rect 701527 479115 701613 479171
rect 701669 479115 701755 479171
rect 701811 479115 701897 479171
rect 701953 479123 706000 479171
rect 701953 479115 705525 479123
rect 699992 479067 705525 479115
rect 705581 479067 705649 479123
rect 705705 479067 705773 479123
rect 705829 479067 705897 479123
rect 705953 479067 706000 479123
rect 699992 479029 706000 479067
rect 699992 478973 700051 479029
rect 700107 478973 700193 479029
rect 700249 478973 700335 479029
rect 700391 478973 700477 479029
rect 700533 478973 700619 479029
rect 700675 478973 700761 479029
rect 700817 478973 700903 479029
rect 700959 478973 701045 479029
rect 701101 478973 701187 479029
rect 701243 478973 701329 479029
rect 701385 478973 701471 479029
rect 701527 478973 701613 479029
rect 701669 478973 701755 479029
rect 701811 478973 701897 479029
rect 701953 478999 706000 479029
rect 701953 478973 705525 478999
rect 699992 478943 705525 478973
rect 705581 478943 705649 478999
rect 705705 478943 705773 478999
rect 705829 478943 705897 478999
rect 705953 478943 706000 478999
rect 699992 478887 706000 478943
rect 699992 478831 700051 478887
rect 700107 478831 700193 478887
rect 700249 478831 700335 478887
rect 700391 478831 700477 478887
rect 700533 478831 700619 478887
rect 700675 478831 700761 478887
rect 700817 478831 700903 478887
rect 700959 478831 701045 478887
rect 701101 478831 701187 478887
rect 701243 478831 701329 478887
rect 701385 478831 701471 478887
rect 701527 478831 701613 478887
rect 701669 478831 701755 478887
rect 701811 478831 701897 478887
rect 701953 478875 706000 478887
rect 701953 478831 705525 478875
rect 699992 478819 705525 478831
rect 705581 478819 705649 478875
rect 705705 478819 705773 478875
rect 705829 478819 705897 478875
rect 705953 478819 706000 478875
rect 699992 478752 706000 478819
rect 699992 478131 706000 478172
rect 699992 478110 705525 478131
rect 699992 478054 700040 478110
rect 700096 478054 700182 478110
rect 700238 478054 700324 478110
rect 700380 478054 700466 478110
rect 700522 478054 700608 478110
rect 700664 478054 700750 478110
rect 700806 478054 700892 478110
rect 700948 478054 701034 478110
rect 701090 478054 701176 478110
rect 701232 478054 701318 478110
rect 701374 478054 701460 478110
rect 701516 478054 701602 478110
rect 701658 478054 701744 478110
rect 701800 478054 701886 478110
rect 701942 478075 705525 478110
rect 705581 478075 705649 478131
rect 705705 478075 705773 478131
rect 705829 478075 705897 478131
rect 705953 478075 706000 478131
rect 701942 478054 706000 478075
rect 699992 478007 706000 478054
rect 699992 477968 705525 478007
rect 699992 477912 700040 477968
rect 700096 477912 700182 477968
rect 700238 477912 700324 477968
rect 700380 477912 700466 477968
rect 700522 477912 700608 477968
rect 700664 477912 700750 477968
rect 700806 477912 700892 477968
rect 700948 477912 701034 477968
rect 701090 477912 701176 477968
rect 701232 477912 701318 477968
rect 701374 477912 701460 477968
rect 701516 477912 701602 477968
rect 701658 477912 701744 477968
rect 701800 477912 701886 477968
rect 701942 477951 705525 477968
rect 705581 477951 705649 478007
rect 705705 477951 705773 478007
rect 705829 477951 705897 478007
rect 705953 477951 706000 478007
rect 701942 477912 706000 477951
rect 699992 477883 706000 477912
rect 699992 477827 705525 477883
rect 705581 477827 705649 477883
rect 705705 477827 705773 477883
rect 705829 477827 705897 477883
rect 705953 477827 706000 477883
rect 699992 477826 706000 477827
rect 699992 477770 700040 477826
rect 700096 477770 700182 477826
rect 700238 477770 700324 477826
rect 700380 477770 700466 477826
rect 700522 477770 700608 477826
rect 700664 477770 700750 477826
rect 700806 477770 700892 477826
rect 700948 477770 701034 477826
rect 701090 477770 701176 477826
rect 701232 477770 701318 477826
rect 701374 477770 701460 477826
rect 701516 477770 701602 477826
rect 701658 477770 701744 477826
rect 701800 477770 701886 477826
rect 701942 477770 706000 477826
rect 699992 477759 706000 477770
rect 699992 477703 705525 477759
rect 705581 477703 705649 477759
rect 705705 477703 705773 477759
rect 705829 477703 705897 477759
rect 705953 477703 706000 477759
rect 699992 477684 706000 477703
rect 699992 477628 700040 477684
rect 700096 477628 700182 477684
rect 700238 477628 700324 477684
rect 700380 477628 700466 477684
rect 700522 477628 700608 477684
rect 700664 477628 700750 477684
rect 700806 477628 700892 477684
rect 700948 477628 701034 477684
rect 701090 477628 701176 477684
rect 701232 477628 701318 477684
rect 701374 477628 701460 477684
rect 701516 477628 701602 477684
rect 701658 477628 701744 477684
rect 701800 477628 701886 477684
rect 701942 477635 706000 477684
rect 701942 477628 705525 477635
rect 699992 477579 705525 477628
rect 705581 477579 705649 477635
rect 705705 477579 705773 477635
rect 705829 477579 705897 477635
rect 705953 477579 706000 477635
rect 699992 477542 706000 477579
rect 699992 477486 700040 477542
rect 700096 477486 700182 477542
rect 700238 477486 700324 477542
rect 700380 477486 700466 477542
rect 700522 477486 700608 477542
rect 700664 477486 700750 477542
rect 700806 477486 700892 477542
rect 700948 477486 701034 477542
rect 701090 477486 701176 477542
rect 701232 477486 701318 477542
rect 701374 477486 701460 477542
rect 701516 477486 701602 477542
rect 701658 477486 701744 477542
rect 701800 477486 701886 477542
rect 701942 477511 706000 477542
rect 701942 477486 705525 477511
rect 699992 477455 705525 477486
rect 705581 477455 705649 477511
rect 705705 477455 705773 477511
rect 705829 477455 705897 477511
rect 705953 477455 706000 477511
rect 699992 477400 706000 477455
rect 699992 477344 700040 477400
rect 700096 477344 700182 477400
rect 700238 477344 700324 477400
rect 700380 477344 700466 477400
rect 700522 477344 700608 477400
rect 700664 477344 700750 477400
rect 700806 477344 700892 477400
rect 700948 477344 701034 477400
rect 701090 477344 701176 477400
rect 701232 477344 701318 477400
rect 701374 477344 701460 477400
rect 701516 477344 701602 477400
rect 701658 477344 701744 477400
rect 701800 477344 701886 477400
rect 701942 477387 706000 477400
rect 701942 477344 705525 477387
rect 699992 477331 705525 477344
rect 705581 477331 705649 477387
rect 705705 477331 705773 477387
rect 705829 477331 705897 477387
rect 705953 477331 706000 477387
rect 699992 477263 706000 477331
rect 699992 477258 705525 477263
rect 699992 477202 700040 477258
rect 700096 477202 700182 477258
rect 700238 477202 700324 477258
rect 700380 477202 700466 477258
rect 700522 477202 700608 477258
rect 700664 477202 700750 477258
rect 700806 477202 700892 477258
rect 700948 477202 701034 477258
rect 701090 477202 701176 477258
rect 701232 477202 701318 477258
rect 701374 477202 701460 477258
rect 701516 477202 701602 477258
rect 701658 477202 701744 477258
rect 701800 477202 701886 477258
rect 701942 477207 705525 477258
rect 705581 477207 705649 477263
rect 705705 477207 705773 477263
rect 705829 477207 705897 477263
rect 705953 477207 706000 477263
rect 701942 477202 706000 477207
rect 699992 477139 706000 477202
rect 699992 477116 705525 477139
rect 699992 477060 700040 477116
rect 700096 477060 700182 477116
rect 700238 477060 700324 477116
rect 700380 477060 700466 477116
rect 700522 477060 700608 477116
rect 700664 477060 700750 477116
rect 700806 477060 700892 477116
rect 700948 477060 701034 477116
rect 701090 477060 701176 477116
rect 701232 477060 701318 477116
rect 701374 477060 701460 477116
rect 701516 477060 701602 477116
rect 701658 477060 701744 477116
rect 701800 477060 701886 477116
rect 701942 477083 705525 477116
rect 705581 477083 705649 477139
rect 705705 477083 705773 477139
rect 705829 477083 705897 477139
rect 705953 477083 706000 477139
rect 701942 477060 706000 477083
rect 699992 477015 706000 477060
rect 699992 476974 705525 477015
rect 699992 476918 700040 476974
rect 700096 476918 700182 476974
rect 700238 476918 700324 476974
rect 700380 476918 700466 476974
rect 700522 476918 700608 476974
rect 700664 476918 700750 476974
rect 700806 476918 700892 476974
rect 700948 476918 701034 476974
rect 701090 476918 701176 476974
rect 701232 476918 701318 476974
rect 701374 476918 701460 476974
rect 701516 476918 701602 476974
rect 701658 476918 701744 476974
rect 701800 476918 701886 476974
rect 701942 476959 705525 476974
rect 705581 476959 705649 477015
rect 705705 476959 705773 477015
rect 705829 476959 705897 477015
rect 705953 476959 706000 477015
rect 701942 476918 706000 476959
rect 699992 476891 706000 476918
rect 699992 476835 705525 476891
rect 705581 476835 705649 476891
rect 705705 476835 705773 476891
rect 705829 476835 705897 476891
rect 705953 476835 706000 476891
rect 699992 476832 706000 476835
rect 699992 476776 700040 476832
rect 700096 476776 700182 476832
rect 700238 476776 700324 476832
rect 700380 476776 700466 476832
rect 700522 476776 700608 476832
rect 700664 476776 700750 476832
rect 700806 476776 700892 476832
rect 700948 476776 701034 476832
rect 701090 476776 701176 476832
rect 701232 476776 701318 476832
rect 701374 476776 701460 476832
rect 701516 476776 701602 476832
rect 701658 476776 701744 476832
rect 701800 476776 701886 476832
rect 701942 476776 706000 476832
rect 699992 476767 706000 476776
rect 699992 476711 705525 476767
rect 705581 476711 705649 476767
rect 705705 476711 705773 476767
rect 705829 476711 705897 476767
rect 705953 476711 706000 476767
rect 699992 476690 706000 476711
rect 699992 476634 700040 476690
rect 700096 476634 700182 476690
rect 700238 476634 700324 476690
rect 700380 476634 700466 476690
rect 700522 476634 700608 476690
rect 700664 476634 700750 476690
rect 700806 476634 700892 476690
rect 700948 476634 701034 476690
rect 701090 476634 701176 476690
rect 701232 476634 701318 476690
rect 701374 476634 701460 476690
rect 701516 476634 701602 476690
rect 701658 476634 701744 476690
rect 701800 476634 701886 476690
rect 701942 476643 706000 476690
rect 701942 476634 705525 476643
rect 699992 476587 705525 476634
rect 705581 476587 705649 476643
rect 705705 476587 705773 476643
rect 705829 476587 705897 476643
rect 705953 476587 706000 476643
rect 699992 476548 706000 476587
rect 699992 476492 700040 476548
rect 700096 476492 700182 476548
rect 700238 476492 700324 476548
rect 700380 476492 700466 476548
rect 700522 476492 700608 476548
rect 700664 476492 700750 476548
rect 700806 476492 700892 476548
rect 700948 476492 701034 476548
rect 701090 476492 701176 476548
rect 701232 476492 701318 476548
rect 701374 476492 701460 476548
rect 701516 476492 701602 476548
rect 701658 476492 701744 476548
rect 701800 476492 701886 476548
rect 701942 476519 706000 476548
rect 701942 476492 705525 476519
rect 699992 476463 705525 476492
rect 705581 476463 705649 476519
rect 705705 476463 705773 476519
rect 705829 476463 705897 476519
rect 705953 476463 706000 476519
rect 699992 476406 706000 476463
rect 699992 476350 700040 476406
rect 700096 476350 700182 476406
rect 700238 476350 700324 476406
rect 700380 476350 700466 476406
rect 700522 476350 700608 476406
rect 700664 476350 700750 476406
rect 700806 476350 700892 476406
rect 700948 476350 701034 476406
rect 701090 476350 701176 476406
rect 701232 476350 701318 476406
rect 701374 476350 701460 476406
rect 701516 476350 701602 476406
rect 701658 476350 701744 476406
rect 701800 476350 701886 476406
rect 701942 476395 706000 476406
rect 701942 476350 705525 476395
rect 699992 476339 705525 476350
rect 705581 476339 705649 476395
rect 705705 476339 705773 476395
rect 705829 476339 705897 476395
rect 705953 476339 706000 476395
rect 699992 476272 706000 476339
rect 70000 468661 75416 468728
rect 70000 468605 70047 468661
rect 70103 468605 70171 468661
rect 70227 468605 70295 468661
rect 70351 468605 70419 468661
rect 70475 468650 75416 468661
rect 70475 468605 73866 468650
rect 70000 468594 73866 468605
rect 73922 468594 74008 468650
rect 74064 468594 74150 468650
rect 74206 468594 74292 468650
rect 74348 468594 74434 468650
rect 74490 468594 74576 468650
rect 74632 468594 74718 468650
rect 74774 468594 74860 468650
rect 74916 468594 75002 468650
rect 75058 468594 75144 468650
rect 75200 468594 75286 468650
rect 75342 468594 75416 468650
rect 70000 468537 75416 468594
rect 70000 468481 70047 468537
rect 70103 468481 70171 468537
rect 70227 468481 70295 468537
rect 70351 468481 70419 468537
rect 70475 468508 75416 468537
rect 70475 468481 73866 468508
rect 70000 468452 73866 468481
rect 73922 468452 74008 468508
rect 74064 468452 74150 468508
rect 74206 468452 74292 468508
rect 74348 468452 74434 468508
rect 74490 468452 74576 468508
rect 74632 468452 74718 468508
rect 74774 468452 74860 468508
rect 74916 468452 75002 468508
rect 75058 468452 75144 468508
rect 75200 468452 75286 468508
rect 75342 468452 75416 468508
rect 70000 468413 75416 468452
rect 70000 468357 70047 468413
rect 70103 468357 70171 468413
rect 70227 468357 70295 468413
rect 70351 468357 70419 468413
rect 70475 468366 75416 468413
rect 70475 468357 73866 468366
rect 70000 468310 73866 468357
rect 73922 468310 74008 468366
rect 74064 468310 74150 468366
rect 74206 468310 74292 468366
rect 74348 468310 74434 468366
rect 74490 468310 74576 468366
rect 74632 468310 74718 468366
rect 74774 468310 74860 468366
rect 74916 468310 75002 468366
rect 75058 468310 75144 468366
rect 75200 468310 75286 468366
rect 75342 468310 75416 468366
rect 70000 468289 75416 468310
rect 70000 468233 70047 468289
rect 70103 468233 70171 468289
rect 70227 468233 70295 468289
rect 70351 468233 70419 468289
rect 70475 468233 75416 468289
rect 70000 468224 75416 468233
rect 70000 468168 73866 468224
rect 73922 468168 74008 468224
rect 74064 468168 74150 468224
rect 74206 468168 74292 468224
rect 74348 468168 74434 468224
rect 74490 468168 74576 468224
rect 74632 468168 74718 468224
rect 74774 468168 74860 468224
rect 74916 468168 75002 468224
rect 75058 468168 75144 468224
rect 75200 468168 75286 468224
rect 75342 468168 75416 468224
rect 70000 468165 75416 468168
rect 70000 468109 70047 468165
rect 70103 468109 70171 468165
rect 70227 468109 70295 468165
rect 70351 468109 70419 468165
rect 70475 468109 75416 468165
rect 70000 468082 75416 468109
rect 70000 468041 73866 468082
rect 70000 467985 70047 468041
rect 70103 467985 70171 468041
rect 70227 467985 70295 468041
rect 70351 467985 70419 468041
rect 70475 468026 73866 468041
rect 73922 468026 74008 468082
rect 74064 468026 74150 468082
rect 74206 468026 74292 468082
rect 74348 468026 74434 468082
rect 74490 468026 74576 468082
rect 74632 468026 74718 468082
rect 74774 468026 74860 468082
rect 74916 468026 75002 468082
rect 75058 468026 75144 468082
rect 75200 468026 75286 468082
rect 75342 468026 75416 468082
rect 70475 467985 75416 468026
rect 70000 467940 75416 467985
rect 70000 467917 73866 467940
rect 70000 467861 70047 467917
rect 70103 467861 70171 467917
rect 70227 467861 70295 467917
rect 70351 467861 70419 467917
rect 70475 467884 73866 467917
rect 73922 467884 74008 467940
rect 74064 467884 74150 467940
rect 74206 467884 74292 467940
rect 74348 467884 74434 467940
rect 74490 467884 74576 467940
rect 74632 467884 74718 467940
rect 74774 467884 74860 467940
rect 74916 467884 75002 467940
rect 75058 467884 75144 467940
rect 75200 467884 75286 467940
rect 75342 467884 75416 467940
rect 70475 467861 75416 467884
rect 70000 467798 75416 467861
rect 70000 467793 73866 467798
rect 70000 467737 70047 467793
rect 70103 467737 70171 467793
rect 70227 467737 70295 467793
rect 70351 467737 70419 467793
rect 70475 467742 73866 467793
rect 73922 467742 74008 467798
rect 74064 467742 74150 467798
rect 74206 467742 74292 467798
rect 74348 467742 74434 467798
rect 74490 467742 74576 467798
rect 74632 467742 74718 467798
rect 74774 467742 74860 467798
rect 74916 467742 75002 467798
rect 75058 467742 75144 467798
rect 75200 467742 75286 467798
rect 75342 467742 75416 467798
rect 70475 467737 75416 467742
rect 70000 467669 75416 467737
rect 70000 467613 70047 467669
rect 70103 467613 70171 467669
rect 70227 467613 70295 467669
rect 70351 467613 70419 467669
rect 70475 467656 75416 467669
rect 70475 467613 73866 467656
rect 70000 467600 73866 467613
rect 73922 467600 74008 467656
rect 74064 467600 74150 467656
rect 74206 467600 74292 467656
rect 74348 467600 74434 467656
rect 74490 467600 74576 467656
rect 74632 467600 74718 467656
rect 74774 467600 74860 467656
rect 74916 467600 75002 467656
rect 75058 467600 75144 467656
rect 75200 467600 75286 467656
rect 75342 467600 75416 467656
rect 70000 467545 75416 467600
rect 70000 467489 70047 467545
rect 70103 467489 70171 467545
rect 70227 467489 70295 467545
rect 70351 467489 70419 467545
rect 70475 467514 75416 467545
rect 70475 467489 73866 467514
rect 70000 467458 73866 467489
rect 73922 467458 74008 467514
rect 74064 467458 74150 467514
rect 74206 467458 74292 467514
rect 74348 467458 74434 467514
rect 74490 467458 74576 467514
rect 74632 467458 74718 467514
rect 74774 467458 74860 467514
rect 74916 467458 75002 467514
rect 75058 467458 75144 467514
rect 75200 467458 75286 467514
rect 75342 467458 75416 467514
rect 70000 467421 75416 467458
rect 70000 467365 70047 467421
rect 70103 467365 70171 467421
rect 70227 467365 70295 467421
rect 70351 467365 70419 467421
rect 70475 467372 75416 467421
rect 70475 467365 73866 467372
rect 70000 467316 73866 467365
rect 73922 467316 74008 467372
rect 74064 467316 74150 467372
rect 74206 467316 74292 467372
rect 74348 467316 74434 467372
rect 74490 467316 74576 467372
rect 74632 467316 74718 467372
rect 74774 467316 74860 467372
rect 74916 467316 75002 467372
rect 75058 467316 75144 467372
rect 75200 467316 75286 467372
rect 75342 467316 75416 467372
rect 70000 467297 75416 467316
rect 70000 467241 70047 467297
rect 70103 467241 70171 467297
rect 70227 467241 70295 467297
rect 70351 467241 70419 467297
rect 70475 467241 75416 467297
rect 70000 467230 75416 467241
rect 70000 467174 73866 467230
rect 73922 467174 74008 467230
rect 74064 467174 74150 467230
rect 74206 467174 74292 467230
rect 74348 467174 74434 467230
rect 74490 467174 74576 467230
rect 74632 467174 74718 467230
rect 74774 467174 74860 467230
rect 74916 467174 75002 467230
rect 75058 467174 75144 467230
rect 75200 467174 75286 467230
rect 75342 467174 75416 467230
rect 70000 467173 75416 467174
rect 70000 467117 70047 467173
rect 70103 467117 70171 467173
rect 70227 467117 70295 467173
rect 70351 467117 70419 467173
rect 70475 467117 75416 467173
rect 70000 467088 75416 467117
rect 70000 467049 73866 467088
rect 70000 466993 70047 467049
rect 70103 466993 70171 467049
rect 70227 466993 70295 467049
rect 70351 466993 70419 467049
rect 70475 467032 73866 467049
rect 73922 467032 74008 467088
rect 74064 467032 74150 467088
rect 74206 467032 74292 467088
rect 74348 467032 74434 467088
rect 74490 467032 74576 467088
rect 74632 467032 74718 467088
rect 74774 467032 74860 467088
rect 74916 467032 75002 467088
rect 75058 467032 75144 467088
rect 75200 467032 75286 467088
rect 75342 467032 75416 467088
rect 70475 466993 75416 467032
rect 70000 466946 75416 466993
rect 70000 466925 73866 466946
rect 70000 466869 70047 466925
rect 70103 466869 70171 466925
rect 70227 466869 70295 466925
rect 70351 466869 70419 466925
rect 70475 466890 73866 466925
rect 73922 466890 74008 466946
rect 74064 466890 74150 466946
rect 74206 466890 74292 466946
rect 74348 466890 74434 466946
rect 74490 466890 74576 466946
rect 74632 466890 74718 466946
rect 74774 466890 74860 466946
rect 74916 466890 75002 466946
rect 75058 466890 75144 466946
rect 75200 466890 75286 466946
rect 75342 466890 75416 466946
rect 70475 466869 75416 466890
rect 70000 466828 75416 466869
rect 70000 466181 75416 466248
rect 70000 466125 70047 466181
rect 70103 466125 70171 466181
rect 70227 466125 70295 466181
rect 70351 466125 70419 466181
rect 70475 466169 75416 466181
rect 70475 466125 73855 466169
rect 70000 466113 73855 466125
rect 73911 466113 73997 466169
rect 74053 466113 74139 466169
rect 74195 466113 74281 466169
rect 74337 466113 74423 466169
rect 74479 466113 74565 466169
rect 74621 466113 74707 466169
rect 74763 466113 74849 466169
rect 74905 466113 74991 466169
rect 75047 466113 75133 466169
rect 75189 466113 75275 466169
rect 75331 466113 75416 466169
rect 70000 466057 75416 466113
rect 70000 466001 70047 466057
rect 70103 466001 70171 466057
rect 70227 466001 70295 466057
rect 70351 466001 70419 466057
rect 70475 466027 75416 466057
rect 70475 466001 73855 466027
rect 70000 465971 73855 466001
rect 73911 465971 73997 466027
rect 74053 465971 74139 466027
rect 74195 465971 74281 466027
rect 74337 465971 74423 466027
rect 74479 465971 74565 466027
rect 74621 465971 74707 466027
rect 74763 465971 74849 466027
rect 74905 465971 74991 466027
rect 75047 465971 75133 466027
rect 75189 465971 75275 466027
rect 75331 465971 75416 466027
rect 70000 465933 75416 465971
rect 70000 465877 70047 465933
rect 70103 465877 70171 465933
rect 70227 465877 70295 465933
rect 70351 465877 70419 465933
rect 70475 465885 75416 465933
rect 70475 465877 73855 465885
rect 70000 465829 73855 465877
rect 73911 465829 73997 465885
rect 74053 465829 74139 465885
rect 74195 465829 74281 465885
rect 74337 465829 74423 465885
rect 74479 465829 74565 465885
rect 74621 465829 74707 465885
rect 74763 465829 74849 465885
rect 74905 465829 74991 465885
rect 75047 465829 75133 465885
rect 75189 465829 75275 465885
rect 75331 465829 75416 465885
rect 70000 465809 75416 465829
rect 70000 465753 70047 465809
rect 70103 465753 70171 465809
rect 70227 465753 70295 465809
rect 70351 465753 70419 465809
rect 70475 465753 75416 465809
rect 70000 465743 75416 465753
rect 70000 465687 73855 465743
rect 73911 465687 73997 465743
rect 74053 465687 74139 465743
rect 74195 465687 74281 465743
rect 74337 465687 74423 465743
rect 74479 465687 74565 465743
rect 74621 465687 74707 465743
rect 74763 465687 74849 465743
rect 74905 465687 74991 465743
rect 75047 465687 75133 465743
rect 75189 465687 75275 465743
rect 75331 465687 75416 465743
rect 70000 465685 75416 465687
rect 70000 465629 70047 465685
rect 70103 465629 70171 465685
rect 70227 465629 70295 465685
rect 70351 465629 70419 465685
rect 70475 465629 75416 465685
rect 70000 465601 75416 465629
rect 70000 465561 73855 465601
rect 70000 465505 70047 465561
rect 70103 465505 70171 465561
rect 70227 465505 70295 465561
rect 70351 465505 70419 465561
rect 70475 465545 73855 465561
rect 73911 465545 73997 465601
rect 74053 465545 74139 465601
rect 74195 465545 74281 465601
rect 74337 465545 74423 465601
rect 74479 465545 74565 465601
rect 74621 465545 74707 465601
rect 74763 465545 74849 465601
rect 74905 465545 74991 465601
rect 75047 465545 75133 465601
rect 75189 465545 75275 465601
rect 75331 465545 75416 465601
rect 70475 465505 75416 465545
rect 70000 465459 75416 465505
rect 70000 465437 73855 465459
rect 70000 465381 70047 465437
rect 70103 465381 70171 465437
rect 70227 465381 70295 465437
rect 70351 465381 70419 465437
rect 70475 465403 73855 465437
rect 73911 465403 73997 465459
rect 74053 465403 74139 465459
rect 74195 465403 74281 465459
rect 74337 465403 74423 465459
rect 74479 465403 74565 465459
rect 74621 465403 74707 465459
rect 74763 465403 74849 465459
rect 74905 465403 74991 465459
rect 75047 465403 75133 465459
rect 75189 465403 75275 465459
rect 75331 465403 75416 465459
rect 70475 465381 75416 465403
rect 70000 465317 75416 465381
rect 70000 465313 73855 465317
rect 70000 465257 70047 465313
rect 70103 465257 70171 465313
rect 70227 465257 70295 465313
rect 70351 465257 70419 465313
rect 70475 465261 73855 465313
rect 73911 465261 73997 465317
rect 74053 465261 74139 465317
rect 74195 465261 74281 465317
rect 74337 465261 74423 465317
rect 74479 465261 74565 465317
rect 74621 465261 74707 465317
rect 74763 465261 74849 465317
rect 74905 465261 74991 465317
rect 75047 465261 75133 465317
rect 75189 465261 75275 465317
rect 75331 465261 75416 465317
rect 70475 465257 75416 465261
rect 70000 465189 75416 465257
rect 70000 465133 70047 465189
rect 70103 465133 70171 465189
rect 70227 465133 70295 465189
rect 70351 465133 70419 465189
rect 70475 465175 75416 465189
rect 70475 465133 73855 465175
rect 70000 465119 73855 465133
rect 73911 465119 73997 465175
rect 74053 465119 74139 465175
rect 74195 465119 74281 465175
rect 74337 465119 74423 465175
rect 74479 465119 74565 465175
rect 74621 465119 74707 465175
rect 74763 465119 74849 465175
rect 74905 465119 74991 465175
rect 75047 465119 75133 465175
rect 75189 465119 75275 465175
rect 75331 465119 75416 465175
rect 70000 465065 75416 465119
rect 70000 465009 70047 465065
rect 70103 465009 70171 465065
rect 70227 465009 70295 465065
rect 70351 465009 70419 465065
rect 70475 465033 75416 465065
rect 70475 465009 73855 465033
rect 70000 464977 73855 465009
rect 73911 464977 73997 465033
rect 74053 464977 74139 465033
rect 74195 464977 74281 465033
rect 74337 464977 74423 465033
rect 74479 464977 74565 465033
rect 74621 464977 74707 465033
rect 74763 464977 74849 465033
rect 74905 464977 74991 465033
rect 75047 464977 75133 465033
rect 75189 464977 75275 465033
rect 75331 464977 75416 465033
rect 70000 464941 75416 464977
rect 70000 464885 70047 464941
rect 70103 464885 70171 464941
rect 70227 464885 70295 464941
rect 70351 464885 70419 464941
rect 70475 464891 75416 464941
rect 70475 464885 73855 464891
rect 70000 464835 73855 464885
rect 73911 464835 73997 464891
rect 74053 464835 74139 464891
rect 74195 464835 74281 464891
rect 74337 464835 74423 464891
rect 74479 464835 74565 464891
rect 74621 464835 74707 464891
rect 74763 464835 74849 464891
rect 74905 464835 74991 464891
rect 75047 464835 75133 464891
rect 75189 464835 75275 464891
rect 75331 464835 75416 464891
rect 70000 464817 75416 464835
rect 70000 464761 70047 464817
rect 70103 464761 70171 464817
rect 70227 464761 70295 464817
rect 70351 464761 70419 464817
rect 70475 464761 75416 464817
rect 70000 464749 75416 464761
rect 70000 464693 73855 464749
rect 73911 464693 73997 464749
rect 74053 464693 74139 464749
rect 74195 464693 74281 464749
rect 74337 464693 74423 464749
rect 74479 464693 74565 464749
rect 74621 464693 74707 464749
rect 74763 464693 74849 464749
rect 74905 464693 74991 464749
rect 75047 464693 75133 464749
rect 75189 464693 75275 464749
rect 75331 464693 75416 464749
rect 70000 464637 70047 464693
rect 70103 464637 70171 464693
rect 70227 464637 70295 464693
rect 70351 464637 70419 464693
rect 70475 464637 75416 464693
rect 70000 464607 75416 464637
rect 70000 464569 73855 464607
rect 70000 464513 70047 464569
rect 70103 464513 70171 464569
rect 70227 464513 70295 464569
rect 70351 464513 70419 464569
rect 70475 464551 73855 464569
rect 73911 464551 73997 464607
rect 74053 464551 74139 464607
rect 74195 464551 74281 464607
rect 74337 464551 74423 464607
rect 74479 464551 74565 464607
rect 74621 464551 74707 464607
rect 74763 464551 74849 464607
rect 74905 464551 74991 464607
rect 75047 464551 75133 464607
rect 75189 464551 75275 464607
rect 75331 464551 75416 464607
rect 70475 464513 75416 464551
rect 70000 464465 75416 464513
rect 70000 464445 73855 464465
rect 70000 464389 70047 464445
rect 70103 464389 70171 464445
rect 70227 464389 70295 464445
rect 70351 464389 70419 464445
rect 70475 464409 73855 464445
rect 73911 464409 73997 464465
rect 74053 464409 74139 464465
rect 74195 464409 74281 464465
rect 74337 464409 74423 464465
rect 74479 464409 74565 464465
rect 74621 464409 74707 464465
rect 74763 464409 74849 464465
rect 74905 464409 74991 464465
rect 75047 464409 75133 464465
rect 75189 464409 75275 464465
rect 75331 464409 75416 464465
rect 70475 464389 75416 464409
rect 70000 464323 75416 464389
rect 70000 464321 73855 464323
rect 70000 464265 70047 464321
rect 70103 464265 70171 464321
rect 70227 464265 70295 464321
rect 70351 464265 70419 464321
rect 70475 464267 73855 464321
rect 73911 464267 73997 464323
rect 74053 464267 74139 464323
rect 74195 464267 74281 464323
rect 74337 464267 74423 464323
rect 74479 464267 74565 464323
rect 74621 464267 74707 464323
rect 74763 464267 74849 464323
rect 74905 464267 74991 464323
rect 75047 464267 75133 464323
rect 75189 464267 75275 464323
rect 75331 464267 75416 464323
rect 70475 464265 75416 464267
rect 70000 464198 75416 464265
rect 70000 463811 75416 463878
rect 70000 463755 70047 463811
rect 70103 463755 70171 463811
rect 70227 463755 70295 463811
rect 70351 463755 70419 463811
rect 70475 463799 75416 463811
rect 70475 463755 73855 463799
rect 70000 463743 73855 463755
rect 73911 463743 73997 463799
rect 74053 463743 74139 463799
rect 74195 463743 74281 463799
rect 74337 463743 74423 463799
rect 74479 463743 74565 463799
rect 74621 463743 74707 463799
rect 74763 463743 74849 463799
rect 74905 463743 74991 463799
rect 75047 463743 75133 463799
rect 75189 463743 75275 463799
rect 75331 463743 75416 463799
rect 70000 463687 75416 463743
rect 70000 463631 70047 463687
rect 70103 463631 70171 463687
rect 70227 463631 70295 463687
rect 70351 463631 70419 463687
rect 70475 463657 75416 463687
rect 70475 463631 73855 463657
rect 70000 463601 73855 463631
rect 73911 463601 73997 463657
rect 74053 463601 74139 463657
rect 74195 463601 74281 463657
rect 74337 463601 74423 463657
rect 74479 463601 74565 463657
rect 74621 463601 74707 463657
rect 74763 463601 74849 463657
rect 74905 463601 74991 463657
rect 75047 463601 75133 463657
rect 75189 463601 75275 463657
rect 75331 463601 75416 463657
rect 70000 463563 75416 463601
rect 70000 463507 70047 463563
rect 70103 463507 70171 463563
rect 70227 463507 70295 463563
rect 70351 463507 70419 463563
rect 70475 463515 75416 463563
rect 70475 463507 73855 463515
rect 70000 463459 73855 463507
rect 73911 463459 73997 463515
rect 74053 463459 74139 463515
rect 74195 463459 74281 463515
rect 74337 463459 74423 463515
rect 74479 463459 74565 463515
rect 74621 463459 74707 463515
rect 74763 463459 74849 463515
rect 74905 463459 74991 463515
rect 75047 463459 75133 463515
rect 75189 463459 75275 463515
rect 75331 463459 75416 463515
rect 70000 463439 75416 463459
rect 70000 463383 70047 463439
rect 70103 463383 70171 463439
rect 70227 463383 70295 463439
rect 70351 463383 70419 463439
rect 70475 463383 75416 463439
rect 70000 463373 75416 463383
rect 70000 463317 73855 463373
rect 73911 463317 73997 463373
rect 74053 463317 74139 463373
rect 74195 463317 74281 463373
rect 74337 463317 74423 463373
rect 74479 463317 74565 463373
rect 74621 463317 74707 463373
rect 74763 463317 74849 463373
rect 74905 463317 74991 463373
rect 75047 463317 75133 463373
rect 75189 463317 75275 463373
rect 75331 463317 75416 463373
rect 70000 463315 75416 463317
rect 70000 463259 70047 463315
rect 70103 463259 70171 463315
rect 70227 463259 70295 463315
rect 70351 463259 70419 463315
rect 70475 463259 75416 463315
rect 70000 463231 75416 463259
rect 70000 463191 73855 463231
rect 70000 463135 70047 463191
rect 70103 463135 70171 463191
rect 70227 463135 70295 463191
rect 70351 463135 70419 463191
rect 70475 463175 73855 463191
rect 73911 463175 73997 463231
rect 74053 463175 74139 463231
rect 74195 463175 74281 463231
rect 74337 463175 74423 463231
rect 74479 463175 74565 463231
rect 74621 463175 74707 463231
rect 74763 463175 74849 463231
rect 74905 463175 74991 463231
rect 75047 463175 75133 463231
rect 75189 463175 75275 463231
rect 75331 463175 75416 463231
rect 70475 463135 75416 463175
rect 70000 463089 75416 463135
rect 70000 463067 73855 463089
rect 70000 463011 70047 463067
rect 70103 463011 70171 463067
rect 70227 463011 70295 463067
rect 70351 463011 70419 463067
rect 70475 463033 73855 463067
rect 73911 463033 73997 463089
rect 74053 463033 74139 463089
rect 74195 463033 74281 463089
rect 74337 463033 74423 463089
rect 74479 463033 74565 463089
rect 74621 463033 74707 463089
rect 74763 463033 74849 463089
rect 74905 463033 74991 463089
rect 75047 463033 75133 463089
rect 75189 463033 75275 463089
rect 75331 463033 75416 463089
rect 70475 463011 75416 463033
rect 70000 462947 75416 463011
rect 70000 462943 73855 462947
rect 70000 462887 70047 462943
rect 70103 462887 70171 462943
rect 70227 462887 70295 462943
rect 70351 462887 70419 462943
rect 70475 462891 73855 462943
rect 73911 462891 73997 462947
rect 74053 462891 74139 462947
rect 74195 462891 74281 462947
rect 74337 462891 74423 462947
rect 74479 462891 74565 462947
rect 74621 462891 74707 462947
rect 74763 462891 74849 462947
rect 74905 462891 74991 462947
rect 75047 462891 75133 462947
rect 75189 462891 75275 462947
rect 75331 462891 75416 462947
rect 70475 462887 75416 462891
rect 70000 462819 75416 462887
rect 70000 462763 70047 462819
rect 70103 462763 70171 462819
rect 70227 462763 70295 462819
rect 70351 462763 70419 462819
rect 70475 462805 75416 462819
rect 70475 462763 73855 462805
rect 70000 462749 73855 462763
rect 73911 462749 73997 462805
rect 74053 462749 74139 462805
rect 74195 462749 74281 462805
rect 74337 462749 74423 462805
rect 74479 462749 74565 462805
rect 74621 462749 74707 462805
rect 74763 462749 74849 462805
rect 74905 462749 74991 462805
rect 75047 462749 75133 462805
rect 75189 462749 75275 462805
rect 75331 462749 75416 462805
rect 70000 462695 75416 462749
rect 70000 462639 70047 462695
rect 70103 462639 70171 462695
rect 70227 462639 70295 462695
rect 70351 462639 70419 462695
rect 70475 462663 75416 462695
rect 70475 462639 73855 462663
rect 70000 462607 73855 462639
rect 73911 462607 73997 462663
rect 74053 462607 74139 462663
rect 74195 462607 74281 462663
rect 74337 462607 74423 462663
rect 74479 462607 74565 462663
rect 74621 462607 74707 462663
rect 74763 462607 74849 462663
rect 74905 462607 74991 462663
rect 75047 462607 75133 462663
rect 75189 462607 75275 462663
rect 75331 462607 75416 462663
rect 70000 462571 75416 462607
rect 70000 462515 70047 462571
rect 70103 462515 70171 462571
rect 70227 462515 70295 462571
rect 70351 462515 70419 462571
rect 70475 462521 75416 462571
rect 70475 462515 73855 462521
rect 70000 462465 73855 462515
rect 73911 462465 73997 462521
rect 74053 462465 74139 462521
rect 74195 462465 74281 462521
rect 74337 462465 74423 462521
rect 74479 462465 74565 462521
rect 74621 462465 74707 462521
rect 74763 462465 74849 462521
rect 74905 462465 74991 462521
rect 75047 462465 75133 462521
rect 75189 462465 75275 462521
rect 75331 462465 75416 462521
rect 70000 462447 75416 462465
rect 70000 462391 70047 462447
rect 70103 462391 70171 462447
rect 70227 462391 70295 462447
rect 70351 462391 70419 462447
rect 70475 462391 75416 462447
rect 70000 462379 75416 462391
rect 70000 462323 73855 462379
rect 73911 462323 73997 462379
rect 74053 462323 74139 462379
rect 74195 462323 74281 462379
rect 74337 462323 74423 462379
rect 74479 462323 74565 462379
rect 74621 462323 74707 462379
rect 74763 462323 74849 462379
rect 74905 462323 74991 462379
rect 75047 462323 75133 462379
rect 75189 462323 75275 462379
rect 75331 462323 75416 462379
rect 70000 462267 70047 462323
rect 70103 462267 70171 462323
rect 70227 462267 70295 462323
rect 70351 462267 70419 462323
rect 70475 462267 75416 462323
rect 70000 462237 75416 462267
rect 70000 462199 73855 462237
rect 70000 462143 70047 462199
rect 70103 462143 70171 462199
rect 70227 462143 70295 462199
rect 70351 462143 70419 462199
rect 70475 462181 73855 462199
rect 73911 462181 73997 462237
rect 74053 462181 74139 462237
rect 74195 462181 74281 462237
rect 74337 462181 74423 462237
rect 74479 462181 74565 462237
rect 74621 462181 74707 462237
rect 74763 462181 74849 462237
rect 74905 462181 74991 462237
rect 75047 462181 75133 462237
rect 75189 462181 75275 462237
rect 75331 462181 75416 462237
rect 70475 462143 75416 462181
rect 70000 462095 75416 462143
rect 70000 462075 73855 462095
rect 70000 462019 70047 462075
rect 70103 462019 70171 462075
rect 70227 462019 70295 462075
rect 70351 462019 70419 462075
rect 70475 462039 73855 462075
rect 73911 462039 73997 462095
rect 74053 462039 74139 462095
rect 74195 462039 74281 462095
rect 74337 462039 74423 462095
rect 74479 462039 74565 462095
rect 74621 462039 74707 462095
rect 74763 462039 74849 462095
rect 74905 462039 74991 462095
rect 75047 462039 75133 462095
rect 75189 462039 75275 462095
rect 75331 462039 75416 462095
rect 70475 462019 75416 462039
rect 70000 461953 75416 462019
rect 70000 461951 73855 461953
rect 70000 461895 70047 461951
rect 70103 461895 70171 461951
rect 70227 461895 70295 461951
rect 70351 461895 70419 461951
rect 70475 461897 73855 461951
rect 73911 461897 73997 461953
rect 74053 461897 74139 461953
rect 74195 461897 74281 461953
rect 74337 461897 74423 461953
rect 74479 461897 74565 461953
rect 74621 461897 74707 461953
rect 74763 461897 74849 461953
rect 74905 461897 74991 461953
rect 75047 461897 75133 461953
rect 75189 461897 75275 461953
rect 75331 461897 75416 461953
rect 70475 461895 75416 461897
rect 70000 461828 75416 461895
rect 70000 461105 75416 461172
rect 70000 461049 70047 461105
rect 70103 461049 70171 461105
rect 70227 461049 70295 461105
rect 70351 461049 70419 461105
rect 70475 461093 75416 461105
rect 70475 461049 73855 461093
rect 70000 461037 73855 461049
rect 73911 461037 73997 461093
rect 74053 461037 74139 461093
rect 74195 461037 74281 461093
rect 74337 461037 74423 461093
rect 74479 461037 74565 461093
rect 74621 461037 74707 461093
rect 74763 461037 74849 461093
rect 74905 461037 74991 461093
rect 75047 461037 75133 461093
rect 75189 461037 75275 461093
rect 75331 461037 75416 461093
rect 70000 460981 75416 461037
rect 70000 460925 70047 460981
rect 70103 460925 70171 460981
rect 70227 460925 70295 460981
rect 70351 460925 70419 460981
rect 70475 460951 75416 460981
rect 70475 460925 73855 460951
rect 70000 460895 73855 460925
rect 73911 460895 73997 460951
rect 74053 460895 74139 460951
rect 74195 460895 74281 460951
rect 74337 460895 74423 460951
rect 74479 460895 74565 460951
rect 74621 460895 74707 460951
rect 74763 460895 74849 460951
rect 74905 460895 74991 460951
rect 75047 460895 75133 460951
rect 75189 460895 75275 460951
rect 75331 460895 75416 460951
rect 70000 460857 75416 460895
rect 70000 460801 70047 460857
rect 70103 460801 70171 460857
rect 70227 460801 70295 460857
rect 70351 460801 70419 460857
rect 70475 460809 75416 460857
rect 70475 460801 73855 460809
rect 70000 460753 73855 460801
rect 73911 460753 73997 460809
rect 74053 460753 74139 460809
rect 74195 460753 74281 460809
rect 74337 460753 74423 460809
rect 74479 460753 74565 460809
rect 74621 460753 74707 460809
rect 74763 460753 74849 460809
rect 74905 460753 74991 460809
rect 75047 460753 75133 460809
rect 75189 460753 75275 460809
rect 75331 460753 75416 460809
rect 70000 460733 75416 460753
rect 70000 460677 70047 460733
rect 70103 460677 70171 460733
rect 70227 460677 70295 460733
rect 70351 460677 70419 460733
rect 70475 460677 75416 460733
rect 70000 460667 75416 460677
rect 70000 460611 73855 460667
rect 73911 460611 73997 460667
rect 74053 460611 74139 460667
rect 74195 460611 74281 460667
rect 74337 460611 74423 460667
rect 74479 460611 74565 460667
rect 74621 460611 74707 460667
rect 74763 460611 74849 460667
rect 74905 460611 74991 460667
rect 75047 460611 75133 460667
rect 75189 460611 75275 460667
rect 75331 460611 75416 460667
rect 70000 460609 75416 460611
rect 70000 460553 70047 460609
rect 70103 460553 70171 460609
rect 70227 460553 70295 460609
rect 70351 460553 70419 460609
rect 70475 460553 75416 460609
rect 70000 460525 75416 460553
rect 70000 460485 73855 460525
rect 70000 460429 70047 460485
rect 70103 460429 70171 460485
rect 70227 460429 70295 460485
rect 70351 460429 70419 460485
rect 70475 460469 73855 460485
rect 73911 460469 73997 460525
rect 74053 460469 74139 460525
rect 74195 460469 74281 460525
rect 74337 460469 74423 460525
rect 74479 460469 74565 460525
rect 74621 460469 74707 460525
rect 74763 460469 74849 460525
rect 74905 460469 74991 460525
rect 75047 460469 75133 460525
rect 75189 460469 75275 460525
rect 75331 460469 75416 460525
rect 70475 460429 75416 460469
rect 70000 460383 75416 460429
rect 70000 460361 73855 460383
rect 70000 460305 70047 460361
rect 70103 460305 70171 460361
rect 70227 460305 70295 460361
rect 70351 460305 70419 460361
rect 70475 460327 73855 460361
rect 73911 460327 73997 460383
rect 74053 460327 74139 460383
rect 74195 460327 74281 460383
rect 74337 460327 74423 460383
rect 74479 460327 74565 460383
rect 74621 460327 74707 460383
rect 74763 460327 74849 460383
rect 74905 460327 74991 460383
rect 75047 460327 75133 460383
rect 75189 460327 75275 460383
rect 75331 460327 75416 460383
rect 70475 460305 75416 460327
rect 70000 460241 75416 460305
rect 70000 460237 73855 460241
rect 70000 460181 70047 460237
rect 70103 460181 70171 460237
rect 70227 460181 70295 460237
rect 70351 460181 70419 460237
rect 70475 460185 73855 460237
rect 73911 460185 73997 460241
rect 74053 460185 74139 460241
rect 74195 460185 74281 460241
rect 74337 460185 74423 460241
rect 74479 460185 74565 460241
rect 74621 460185 74707 460241
rect 74763 460185 74849 460241
rect 74905 460185 74991 460241
rect 75047 460185 75133 460241
rect 75189 460185 75275 460241
rect 75331 460185 75416 460241
rect 70475 460181 75416 460185
rect 70000 460113 75416 460181
rect 70000 460057 70047 460113
rect 70103 460057 70171 460113
rect 70227 460057 70295 460113
rect 70351 460057 70419 460113
rect 70475 460099 75416 460113
rect 70475 460057 73855 460099
rect 70000 460043 73855 460057
rect 73911 460043 73997 460099
rect 74053 460043 74139 460099
rect 74195 460043 74281 460099
rect 74337 460043 74423 460099
rect 74479 460043 74565 460099
rect 74621 460043 74707 460099
rect 74763 460043 74849 460099
rect 74905 460043 74991 460099
rect 75047 460043 75133 460099
rect 75189 460043 75275 460099
rect 75331 460043 75416 460099
rect 70000 459989 75416 460043
rect 70000 459933 70047 459989
rect 70103 459933 70171 459989
rect 70227 459933 70295 459989
rect 70351 459933 70419 459989
rect 70475 459957 75416 459989
rect 70475 459933 73855 459957
rect 70000 459901 73855 459933
rect 73911 459901 73997 459957
rect 74053 459901 74139 459957
rect 74195 459901 74281 459957
rect 74337 459901 74423 459957
rect 74479 459901 74565 459957
rect 74621 459901 74707 459957
rect 74763 459901 74849 459957
rect 74905 459901 74991 459957
rect 75047 459901 75133 459957
rect 75189 459901 75275 459957
rect 75331 459901 75416 459957
rect 70000 459865 75416 459901
rect 70000 459809 70047 459865
rect 70103 459809 70171 459865
rect 70227 459809 70295 459865
rect 70351 459809 70419 459865
rect 70475 459815 75416 459865
rect 70475 459809 73855 459815
rect 70000 459759 73855 459809
rect 73911 459759 73997 459815
rect 74053 459759 74139 459815
rect 74195 459759 74281 459815
rect 74337 459759 74423 459815
rect 74479 459759 74565 459815
rect 74621 459759 74707 459815
rect 74763 459759 74849 459815
rect 74905 459759 74991 459815
rect 75047 459759 75133 459815
rect 75189 459759 75275 459815
rect 75331 459759 75416 459815
rect 70000 459741 75416 459759
rect 70000 459685 70047 459741
rect 70103 459685 70171 459741
rect 70227 459685 70295 459741
rect 70351 459685 70419 459741
rect 70475 459685 75416 459741
rect 70000 459673 75416 459685
rect 70000 459617 73855 459673
rect 73911 459617 73997 459673
rect 74053 459617 74139 459673
rect 74195 459617 74281 459673
rect 74337 459617 74423 459673
rect 74479 459617 74565 459673
rect 74621 459617 74707 459673
rect 74763 459617 74849 459673
rect 74905 459617 74991 459673
rect 75047 459617 75133 459673
rect 75189 459617 75275 459673
rect 75331 459617 75416 459673
rect 70000 459561 70047 459617
rect 70103 459561 70171 459617
rect 70227 459561 70295 459617
rect 70351 459561 70419 459617
rect 70475 459561 75416 459617
rect 70000 459531 75416 459561
rect 70000 459493 73855 459531
rect 70000 459437 70047 459493
rect 70103 459437 70171 459493
rect 70227 459437 70295 459493
rect 70351 459437 70419 459493
rect 70475 459475 73855 459493
rect 73911 459475 73997 459531
rect 74053 459475 74139 459531
rect 74195 459475 74281 459531
rect 74337 459475 74423 459531
rect 74479 459475 74565 459531
rect 74621 459475 74707 459531
rect 74763 459475 74849 459531
rect 74905 459475 74991 459531
rect 75047 459475 75133 459531
rect 75189 459475 75275 459531
rect 75331 459475 75416 459531
rect 70475 459437 75416 459475
rect 70000 459389 75416 459437
rect 70000 459369 73855 459389
rect 70000 459313 70047 459369
rect 70103 459313 70171 459369
rect 70227 459313 70295 459369
rect 70351 459313 70419 459369
rect 70475 459333 73855 459369
rect 73911 459333 73997 459389
rect 74053 459333 74139 459389
rect 74195 459333 74281 459389
rect 74337 459333 74423 459389
rect 74479 459333 74565 459389
rect 74621 459333 74707 459389
rect 74763 459333 74849 459389
rect 74905 459333 74991 459389
rect 75047 459333 75133 459389
rect 75189 459333 75275 459389
rect 75331 459333 75416 459389
rect 70475 459313 75416 459333
rect 70000 459247 75416 459313
rect 70000 459245 73855 459247
rect 70000 459189 70047 459245
rect 70103 459189 70171 459245
rect 70227 459189 70295 459245
rect 70351 459189 70419 459245
rect 70475 459191 73855 459245
rect 73911 459191 73997 459247
rect 74053 459191 74139 459247
rect 74195 459191 74281 459247
rect 74337 459191 74423 459247
rect 74479 459191 74565 459247
rect 74621 459191 74707 459247
rect 74763 459191 74849 459247
rect 74905 459191 74991 459247
rect 75047 459191 75133 459247
rect 75189 459191 75275 459247
rect 75331 459191 75416 459247
rect 70475 459189 75416 459191
rect 70000 459122 75416 459189
rect 70000 458735 75416 458802
rect 70000 458679 70047 458735
rect 70103 458679 70171 458735
rect 70227 458679 70295 458735
rect 70351 458679 70419 458735
rect 70475 458723 75416 458735
rect 70475 458679 73855 458723
rect 70000 458667 73855 458679
rect 73911 458667 73997 458723
rect 74053 458667 74139 458723
rect 74195 458667 74281 458723
rect 74337 458667 74423 458723
rect 74479 458667 74565 458723
rect 74621 458667 74707 458723
rect 74763 458667 74849 458723
rect 74905 458667 74991 458723
rect 75047 458667 75133 458723
rect 75189 458667 75275 458723
rect 75331 458667 75416 458723
rect 70000 458611 75416 458667
rect 70000 458555 70047 458611
rect 70103 458555 70171 458611
rect 70227 458555 70295 458611
rect 70351 458555 70419 458611
rect 70475 458581 75416 458611
rect 70475 458555 73855 458581
rect 70000 458525 73855 458555
rect 73911 458525 73997 458581
rect 74053 458525 74139 458581
rect 74195 458525 74281 458581
rect 74337 458525 74423 458581
rect 74479 458525 74565 458581
rect 74621 458525 74707 458581
rect 74763 458525 74849 458581
rect 74905 458525 74991 458581
rect 75047 458525 75133 458581
rect 75189 458525 75275 458581
rect 75331 458525 75416 458581
rect 70000 458487 75416 458525
rect 70000 458431 70047 458487
rect 70103 458431 70171 458487
rect 70227 458431 70295 458487
rect 70351 458431 70419 458487
rect 70475 458439 75416 458487
rect 70475 458431 73855 458439
rect 70000 458383 73855 458431
rect 73911 458383 73997 458439
rect 74053 458383 74139 458439
rect 74195 458383 74281 458439
rect 74337 458383 74423 458439
rect 74479 458383 74565 458439
rect 74621 458383 74707 458439
rect 74763 458383 74849 458439
rect 74905 458383 74991 458439
rect 75047 458383 75133 458439
rect 75189 458383 75275 458439
rect 75331 458383 75416 458439
rect 70000 458363 75416 458383
rect 70000 458307 70047 458363
rect 70103 458307 70171 458363
rect 70227 458307 70295 458363
rect 70351 458307 70419 458363
rect 70475 458307 75416 458363
rect 70000 458297 75416 458307
rect 70000 458241 73855 458297
rect 73911 458241 73997 458297
rect 74053 458241 74139 458297
rect 74195 458241 74281 458297
rect 74337 458241 74423 458297
rect 74479 458241 74565 458297
rect 74621 458241 74707 458297
rect 74763 458241 74849 458297
rect 74905 458241 74991 458297
rect 75047 458241 75133 458297
rect 75189 458241 75275 458297
rect 75331 458241 75416 458297
rect 70000 458239 75416 458241
rect 70000 458183 70047 458239
rect 70103 458183 70171 458239
rect 70227 458183 70295 458239
rect 70351 458183 70419 458239
rect 70475 458183 75416 458239
rect 70000 458155 75416 458183
rect 70000 458115 73855 458155
rect 70000 458059 70047 458115
rect 70103 458059 70171 458115
rect 70227 458059 70295 458115
rect 70351 458059 70419 458115
rect 70475 458099 73855 458115
rect 73911 458099 73997 458155
rect 74053 458099 74139 458155
rect 74195 458099 74281 458155
rect 74337 458099 74423 458155
rect 74479 458099 74565 458155
rect 74621 458099 74707 458155
rect 74763 458099 74849 458155
rect 74905 458099 74991 458155
rect 75047 458099 75133 458155
rect 75189 458099 75275 458155
rect 75331 458099 75416 458155
rect 70475 458059 75416 458099
rect 70000 458013 75416 458059
rect 70000 457991 73855 458013
rect 70000 457935 70047 457991
rect 70103 457935 70171 457991
rect 70227 457935 70295 457991
rect 70351 457935 70419 457991
rect 70475 457957 73855 457991
rect 73911 457957 73997 458013
rect 74053 457957 74139 458013
rect 74195 457957 74281 458013
rect 74337 457957 74423 458013
rect 74479 457957 74565 458013
rect 74621 457957 74707 458013
rect 74763 457957 74849 458013
rect 74905 457957 74991 458013
rect 75047 457957 75133 458013
rect 75189 457957 75275 458013
rect 75331 457957 75416 458013
rect 70475 457935 75416 457957
rect 70000 457871 75416 457935
rect 70000 457867 73855 457871
rect 70000 457811 70047 457867
rect 70103 457811 70171 457867
rect 70227 457811 70295 457867
rect 70351 457811 70419 457867
rect 70475 457815 73855 457867
rect 73911 457815 73997 457871
rect 74053 457815 74139 457871
rect 74195 457815 74281 457871
rect 74337 457815 74423 457871
rect 74479 457815 74565 457871
rect 74621 457815 74707 457871
rect 74763 457815 74849 457871
rect 74905 457815 74991 457871
rect 75047 457815 75133 457871
rect 75189 457815 75275 457871
rect 75331 457815 75416 457871
rect 70475 457811 75416 457815
rect 70000 457743 75416 457811
rect 70000 457687 70047 457743
rect 70103 457687 70171 457743
rect 70227 457687 70295 457743
rect 70351 457687 70419 457743
rect 70475 457729 75416 457743
rect 70475 457687 73855 457729
rect 70000 457673 73855 457687
rect 73911 457673 73997 457729
rect 74053 457673 74139 457729
rect 74195 457673 74281 457729
rect 74337 457673 74423 457729
rect 74479 457673 74565 457729
rect 74621 457673 74707 457729
rect 74763 457673 74849 457729
rect 74905 457673 74991 457729
rect 75047 457673 75133 457729
rect 75189 457673 75275 457729
rect 75331 457673 75416 457729
rect 70000 457619 75416 457673
rect 70000 457563 70047 457619
rect 70103 457563 70171 457619
rect 70227 457563 70295 457619
rect 70351 457563 70419 457619
rect 70475 457587 75416 457619
rect 70475 457563 73855 457587
rect 70000 457531 73855 457563
rect 73911 457531 73997 457587
rect 74053 457531 74139 457587
rect 74195 457531 74281 457587
rect 74337 457531 74423 457587
rect 74479 457531 74565 457587
rect 74621 457531 74707 457587
rect 74763 457531 74849 457587
rect 74905 457531 74991 457587
rect 75047 457531 75133 457587
rect 75189 457531 75275 457587
rect 75331 457531 75416 457587
rect 70000 457495 75416 457531
rect 70000 457439 70047 457495
rect 70103 457439 70171 457495
rect 70227 457439 70295 457495
rect 70351 457439 70419 457495
rect 70475 457445 75416 457495
rect 70475 457439 73855 457445
rect 70000 457389 73855 457439
rect 73911 457389 73997 457445
rect 74053 457389 74139 457445
rect 74195 457389 74281 457445
rect 74337 457389 74423 457445
rect 74479 457389 74565 457445
rect 74621 457389 74707 457445
rect 74763 457389 74849 457445
rect 74905 457389 74991 457445
rect 75047 457389 75133 457445
rect 75189 457389 75275 457445
rect 75331 457389 75416 457445
rect 70000 457371 75416 457389
rect 70000 457315 70047 457371
rect 70103 457315 70171 457371
rect 70227 457315 70295 457371
rect 70351 457315 70419 457371
rect 70475 457315 75416 457371
rect 70000 457303 75416 457315
rect 70000 457247 73855 457303
rect 73911 457247 73997 457303
rect 74053 457247 74139 457303
rect 74195 457247 74281 457303
rect 74337 457247 74423 457303
rect 74479 457247 74565 457303
rect 74621 457247 74707 457303
rect 74763 457247 74849 457303
rect 74905 457247 74991 457303
rect 75047 457247 75133 457303
rect 75189 457247 75275 457303
rect 75331 457247 75416 457303
rect 70000 457191 70047 457247
rect 70103 457191 70171 457247
rect 70227 457191 70295 457247
rect 70351 457191 70419 457247
rect 70475 457191 75416 457247
rect 70000 457161 75416 457191
rect 70000 457123 73855 457161
rect 70000 457067 70047 457123
rect 70103 457067 70171 457123
rect 70227 457067 70295 457123
rect 70351 457067 70419 457123
rect 70475 457105 73855 457123
rect 73911 457105 73997 457161
rect 74053 457105 74139 457161
rect 74195 457105 74281 457161
rect 74337 457105 74423 457161
rect 74479 457105 74565 457161
rect 74621 457105 74707 457161
rect 74763 457105 74849 457161
rect 74905 457105 74991 457161
rect 75047 457105 75133 457161
rect 75189 457105 75275 457161
rect 75331 457105 75416 457161
rect 70475 457067 75416 457105
rect 70000 457019 75416 457067
rect 70000 456999 73855 457019
rect 70000 456943 70047 456999
rect 70103 456943 70171 456999
rect 70227 456943 70295 456999
rect 70351 456943 70419 456999
rect 70475 456963 73855 456999
rect 73911 456963 73997 457019
rect 74053 456963 74139 457019
rect 74195 456963 74281 457019
rect 74337 456963 74423 457019
rect 74479 456963 74565 457019
rect 74621 456963 74707 457019
rect 74763 456963 74849 457019
rect 74905 456963 74991 457019
rect 75047 456963 75133 457019
rect 75189 456963 75275 457019
rect 75331 456963 75416 457019
rect 70475 456943 75416 456963
rect 70000 456877 75416 456943
rect 70000 456875 73855 456877
rect 70000 456819 70047 456875
rect 70103 456819 70171 456875
rect 70227 456819 70295 456875
rect 70351 456819 70419 456875
rect 70475 456821 73855 456875
rect 73911 456821 73997 456877
rect 74053 456821 74139 456877
rect 74195 456821 74281 456877
rect 74337 456821 74423 456877
rect 74479 456821 74565 456877
rect 74621 456821 74707 456877
rect 74763 456821 74849 456877
rect 74905 456821 74991 456877
rect 75047 456821 75133 456877
rect 75189 456821 75275 456877
rect 75331 456821 75416 456877
rect 70475 456819 75416 456821
rect 70000 456752 75416 456819
rect 70000 456105 75416 456172
rect 70000 456049 70047 456105
rect 70103 456049 70171 456105
rect 70227 456049 70295 456105
rect 70351 456049 70419 456105
rect 70475 456094 75416 456105
rect 70475 456049 73866 456094
rect 70000 456038 73866 456049
rect 73922 456038 74008 456094
rect 74064 456038 74150 456094
rect 74206 456038 74292 456094
rect 74348 456038 74434 456094
rect 74490 456038 74576 456094
rect 74632 456038 74718 456094
rect 74774 456038 74860 456094
rect 74916 456038 75002 456094
rect 75058 456038 75144 456094
rect 75200 456038 75286 456094
rect 75342 456038 75416 456094
rect 70000 455981 75416 456038
rect 70000 455925 70047 455981
rect 70103 455925 70171 455981
rect 70227 455925 70295 455981
rect 70351 455925 70419 455981
rect 70475 455952 75416 455981
rect 70475 455925 73866 455952
rect 70000 455896 73866 455925
rect 73922 455896 74008 455952
rect 74064 455896 74150 455952
rect 74206 455896 74292 455952
rect 74348 455896 74434 455952
rect 74490 455896 74576 455952
rect 74632 455896 74718 455952
rect 74774 455896 74860 455952
rect 74916 455896 75002 455952
rect 75058 455896 75144 455952
rect 75200 455896 75286 455952
rect 75342 455896 75416 455952
rect 70000 455857 75416 455896
rect 70000 455801 70047 455857
rect 70103 455801 70171 455857
rect 70227 455801 70295 455857
rect 70351 455801 70419 455857
rect 70475 455810 75416 455857
rect 70475 455801 73866 455810
rect 70000 455754 73866 455801
rect 73922 455754 74008 455810
rect 74064 455754 74150 455810
rect 74206 455754 74292 455810
rect 74348 455754 74434 455810
rect 74490 455754 74576 455810
rect 74632 455754 74718 455810
rect 74774 455754 74860 455810
rect 74916 455754 75002 455810
rect 75058 455754 75144 455810
rect 75200 455754 75286 455810
rect 75342 455754 75416 455810
rect 70000 455733 75416 455754
rect 70000 455677 70047 455733
rect 70103 455677 70171 455733
rect 70227 455677 70295 455733
rect 70351 455677 70419 455733
rect 70475 455677 75416 455733
rect 70000 455668 75416 455677
rect 70000 455612 73866 455668
rect 73922 455612 74008 455668
rect 74064 455612 74150 455668
rect 74206 455612 74292 455668
rect 74348 455612 74434 455668
rect 74490 455612 74576 455668
rect 74632 455612 74718 455668
rect 74774 455612 74860 455668
rect 74916 455612 75002 455668
rect 75058 455612 75144 455668
rect 75200 455612 75286 455668
rect 75342 455612 75416 455668
rect 70000 455609 75416 455612
rect 70000 455553 70047 455609
rect 70103 455553 70171 455609
rect 70227 455553 70295 455609
rect 70351 455553 70419 455609
rect 70475 455553 75416 455609
rect 70000 455526 75416 455553
rect 70000 455485 73866 455526
rect 70000 455429 70047 455485
rect 70103 455429 70171 455485
rect 70227 455429 70295 455485
rect 70351 455429 70419 455485
rect 70475 455470 73866 455485
rect 73922 455470 74008 455526
rect 74064 455470 74150 455526
rect 74206 455470 74292 455526
rect 74348 455470 74434 455526
rect 74490 455470 74576 455526
rect 74632 455470 74718 455526
rect 74774 455470 74860 455526
rect 74916 455470 75002 455526
rect 75058 455470 75144 455526
rect 75200 455470 75286 455526
rect 75342 455470 75416 455526
rect 70475 455429 75416 455470
rect 70000 455384 75416 455429
rect 70000 455361 73866 455384
rect 70000 455305 70047 455361
rect 70103 455305 70171 455361
rect 70227 455305 70295 455361
rect 70351 455305 70419 455361
rect 70475 455328 73866 455361
rect 73922 455328 74008 455384
rect 74064 455328 74150 455384
rect 74206 455328 74292 455384
rect 74348 455328 74434 455384
rect 74490 455328 74576 455384
rect 74632 455328 74718 455384
rect 74774 455328 74860 455384
rect 74916 455328 75002 455384
rect 75058 455328 75144 455384
rect 75200 455328 75286 455384
rect 75342 455328 75416 455384
rect 70475 455305 75416 455328
rect 70000 455242 75416 455305
rect 70000 455237 73866 455242
rect 70000 455181 70047 455237
rect 70103 455181 70171 455237
rect 70227 455181 70295 455237
rect 70351 455181 70419 455237
rect 70475 455186 73866 455237
rect 73922 455186 74008 455242
rect 74064 455186 74150 455242
rect 74206 455186 74292 455242
rect 74348 455186 74434 455242
rect 74490 455186 74576 455242
rect 74632 455186 74718 455242
rect 74774 455186 74860 455242
rect 74916 455186 75002 455242
rect 75058 455186 75144 455242
rect 75200 455186 75286 455242
rect 75342 455186 75416 455242
rect 70475 455181 75416 455186
rect 70000 455113 75416 455181
rect 70000 455057 70047 455113
rect 70103 455057 70171 455113
rect 70227 455057 70295 455113
rect 70351 455057 70419 455113
rect 70475 455100 75416 455113
rect 70475 455057 73866 455100
rect 70000 455044 73866 455057
rect 73922 455044 74008 455100
rect 74064 455044 74150 455100
rect 74206 455044 74292 455100
rect 74348 455044 74434 455100
rect 74490 455044 74576 455100
rect 74632 455044 74718 455100
rect 74774 455044 74860 455100
rect 74916 455044 75002 455100
rect 75058 455044 75144 455100
rect 75200 455044 75286 455100
rect 75342 455044 75416 455100
rect 70000 454989 75416 455044
rect 70000 454933 70047 454989
rect 70103 454933 70171 454989
rect 70227 454933 70295 454989
rect 70351 454933 70419 454989
rect 70475 454958 75416 454989
rect 70475 454933 73866 454958
rect 70000 454902 73866 454933
rect 73922 454902 74008 454958
rect 74064 454902 74150 454958
rect 74206 454902 74292 454958
rect 74348 454902 74434 454958
rect 74490 454902 74576 454958
rect 74632 454902 74718 454958
rect 74774 454902 74860 454958
rect 74916 454902 75002 454958
rect 75058 454902 75144 454958
rect 75200 454902 75286 454958
rect 75342 454902 75416 454958
rect 70000 454865 75416 454902
rect 70000 454809 70047 454865
rect 70103 454809 70171 454865
rect 70227 454809 70295 454865
rect 70351 454809 70419 454865
rect 70475 454816 75416 454865
rect 70475 454809 73866 454816
rect 70000 454760 73866 454809
rect 73922 454760 74008 454816
rect 74064 454760 74150 454816
rect 74206 454760 74292 454816
rect 74348 454760 74434 454816
rect 74490 454760 74576 454816
rect 74632 454760 74718 454816
rect 74774 454760 74860 454816
rect 74916 454760 75002 454816
rect 75058 454760 75144 454816
rect 75200 454760 75286 454816
rect 75342 454760 75416 454816
rect 70000 454741 75416 454760
rect 70000 454685 70047 454741
rect 70103 454685 70171 454741
rect 70227 454685 70295 454741
rect 70351 454685 70419 454741
rect 70475 454685 75416 454741
rect 70000 454674 75416 454685
rect 70000 454618 73866 454674
rect 73922 454618 74008 454674
rect 74064 454618 74150 454674
rect 74206 454618 74292 454674
rect 74348 454618 74434 454674
rect 74490 454618 74576 454674
rect 74632 454618 74718 454674
rect 74774 454618 74860 454674
rect 74916 454618 75002 454674
rect 75058 454618 75144 454674
rect 75200 454618 75286 454674
rect 75342 454618 75416 454674
rect 70000 454617 75416 454618
rect 70000 454561 70047 454617
rect 70103 454561 70171 454617
rect 70227 454561 70295 454617
rect 70351 454561 70419 454617
rect 70475 454561 75416 454617
rect 70000 454532 75416 454561
rect 70000 454493 73866 454532
rect 70000 454437 70047 454493
rect 70103 454437 70171 454493
rect 70227 454437 70295 454493
rect 70351 454437 70419 454493
rect 70475 454476 73866 454493
rect 73922 454476 74008 454532
rect 74064 454476 74150 454532
rect 74206 454476 74292 454532
rect 74348 454476 74434 454532
rect 74490 454476 74576 454532
rect 74632 454476 74718 454532
rect 74774 454476 74860 454532
rect 74916 454476 75002 454532
rect 75058 454476 75144 454532
rect 75200 454476 75286 454532
rect 75342 454476 75416 454532
rect 70475 454437 75416 454476
rect 70000 454390 75416 454437
rect 70000 454369 73866 454390
rect 70000 454313 70047 454369
rect 70103 454313 70171 454369
rect 70227 454313 70295 454369
rect 70351 454313 70419 454369
rect 70475 454334 73866 454369
rect 73922 454334 74008 454390
rect 74064 454334 74150 454390
rect 74206 454334 74292 454390
rect 74348 454334 74434 454390
rect 74490 454334 74576 454390
rect 74632 454334 74718 454390
rect 74774 454334 74860 454390
rect 74916 454334 75002 454390
rect 75058 454334 75144 454390
rect 75200 454334 75286 454390
rect 75342 454334 75416 454390
rect 70475 454313 75416 454334
rect 70000 454272 75416 454313
rect 702392 447687 706000 447728
rect 702392 447666 705525 447687
rect 702392 447610 702440 447666
rect 702496 447610 702582 447666
rect 702638 447610 702724 447666
rect 702780 447610 702866 447666
rect 702922 447610 703008 447666
rect 703064 447610 703150 447666
rect 703206 447610 703292 447666
rect 703348 447610 703434 447666
rect 703490 447610 703576 447666
rect 703632 447610 703718 447666
rect 703774 447610 703860 447666
rect 703916 447610 704002 447666
rect 704058 447610 704144 447666
rect 704200 447610 704286 447666
rect 704342 447631 705525 447666
rect 705581 447631 705649 447687
rect 705705 447631 705773 447687
rect 705829 447631 705897 447687
rect 705953 447631 706000 447687
rect 704342 447610 706000 447631
rect 702392 447563 706000 447610
rect 702392 447524 705525 447563
rect 702392 447468 702440 447524
rect 702496 447468 702582 447524
rect 702638 447468 702724 447524
rect 702780 447468 702866 447524
rect 702922 447468 703008 447524
rect 703064 447468 703150 447524
rect 703206 447468 703292 447524
rect 703348 447468 703434 447524
rect 703490 447468 703576 447524
rect 703632 447468 703718 447524
rect 703774 447468 703860 447524
rect 703916 447468 704002 447524
rect 704058 447468 704144 447524
rect 704200 447468 704286 447524
rect 704342 447507 705525 447524
rect 705581 447507 705649 447563
rect 705705 447507 705773 447563
rect 705829 447507 705897 447563
rect 705953 447507 706000 447563
rect 704342 447468 706000 447507
rect 702392 447439 706000 447468
rect 702392 447383 705525 447439
rect 705581 447383 705649 447439
rect 705705 447383 705773 447439
rect 705829 447383 705897 447439
rect 705953 447383 706000 447439
rect 702392 447382 706000 447383
rect 702392 447326 702440 447382
rect 702496 447326 702582 447382
rect 702638 447326 702724 447382
rect 702780 447326 702866 447382
rect 702922 447326 703008 447382
rect 703064 447326 703150 447382
rect 703206 447326 703292 447382
rect 703348 447326 703434 447382
rect 703490 447326 703576 447382
rect 703632 447326 703718 447382
rect 703774 447326 703860 447382
rect 703916 447326 704002 447382
rect 704058 447326 704144 447382
rect 704200 447326 704286 447382
rect 704342 447326 706000 447382
rect 702392 447315 706000 447326
rect 702392 447259 705525 447315
rect 705581 447259 705649 447315
rect 705705 447259 705773 447315
rect 705829 447259 705897 447315
rect 705953 447259 706000 447315
rect 702392 447240 706000 447259
rect 702392 447184 702440 447240
rect 702496 447184 702582 447240
rect 702638 447184 702724 447240
rect 702780 447184 702866 447240
rect 702922 447184 703008 447240
rect 703064 447184 703150 447240
rect 703206 447184 703292 447240
rect 703348 447184 703434 447240
rect 703490 447184 703576 447240
rect 703632 447184 703718 447240
rect 703774 447184 703860 447240
rect 703916 447184 704002 447240
rect 704058 447184 704144 447240
rect 704200 447184 704286 447240
rect 704342 447191 706000 447240
rect 704342 447184 705525 447191
rect 702392 447135 705525 447184
rect 705581 447135 705649 447191
rect 705705 447135 705773 447191
rect 705829 447135 705897 447191
rect 705953 447135 706000 447191
rect 702392 447098 706000 447135
rect 702392 447042 702440 447098
rect 702496 447042 702582 447098
rect 702638 447042 702724 447098
rect 702780 447042 702866 447098
rect 702922 447042 703008 447098
rect 703064 447042 703150 447098
rect 703206 447042 703292 447098
rect 703348 447042 703434 447098
rect 703490 447042 703576 447098
rect 703632 447042 703718 447098
rect 703774 447042 703860 447098
rect 703916 447042 704002 447098
rect 704058 447042 704144 447098
rect 704200 447042 704286 447098
rect 704342 447067 706000 447098
rect 704342 447042 705525 447067
rect 702392 447011 705525 447042
rect 705581 447011 705649 447067
rect 705705 447011 705773 447067
rect 705829 447011 705897 447067
rect 705953 447011 706000 447067
rect 702392 446956 706000 447011
rect 702392 446900 702440 446956
rect 702496 446900 702582 446956
rect 702638 446900 702724 446956
rect 702780 446900 702866 446956
rect 702922 446900 703008 446956
rect 703064 446900 703150 446956
rect 703206 446900 703292 446956
rect 703348 446900 703434 446956
rect 703490 446900 703576 446956
rect 703632 446900 703718 446956
rect 703774 446900 703860 446956
rect 703916 446900 704002 446956
rect 704058 446900 704144 446956
rect 704200 446900 704286 446956
rect 704342 446943 706000 446956
rect 704342 446900 705525 446943
rect 702392 446887 705525 446900
rect 705581 446887 705649 446943
rect 705705 446887 705773 446943
rect 705829 446887 705897 446943
rect 705953 446887 706000 446943
rect 702392 446819 706000 446887
rect 702392 446814 705525 446819
rect 702392 446758 702440 446814
rect 702496 446758 702582 446814
rect 702638 446758 702724 446814
rect 702780 446758 702866 446814
rect 702922 446758 703008 446814
rect 703064 446758 703150 446814
rect 703206 446758 703292 446814
rect 703348 446758 703434 446814
rect 703490 446758 703576 446814
rect 703632 446758 703718 446814
rect 703774 446758 703860 446814
rect 703916 446758 704002 446814
rect 704058 446758 704144 446814
rect 704200 446758 704286 446814
rect 704342 446763 705525 446814
rect 705581 446763 705649 446819
rect 705705 446763 705773 446819
rect 705829 446763 705897 446819
rect 705953 446763 706000 446819
rect 704342 446758 706000 446763
rect 702392 446695 706000 446758
rect 702392 446672 705525 446695
rect 702392 446616 702440 446672
rect 702496 446616 702582 446672
rect 702638 446616 702724 446672
rect 702780 446616 702866 446672
rect 702922 446616 703008 446672
rect 703064 446616 703150 446672
rect 703206 446616 703292 446672
rect 703348 446616 703434 446672
rect 703490 446616 703576 446672
rect 703632 446616 703718 446672
rect 703774 446616 703860 446672
rect 703916 446616 704002 446672
rect 704058 446616 704144 446672
rect 704200 446616 704286 446672
rect 704342 446639 705525 446672
rect 705581 446639 705649 446695
rect 705705 446639 705773 446695
rect 705829 446639 705897 446695
rect 705953 446639 706000 446695
rect 704342 446616 706000 446639
rect 702392 446571 706000 446616
rect 702392 446530 705525 446571
rect 702392 446474 702440 446530
rect 702496 446474 702582 446530
rect 702638 446474 702724 446530
rect 702780 446474 702866 446530
rect 702922 446474 703008 446530
rect 703064 446474 703150 446530
rect 703206 446474 703292 446530
rect 703348 446474 703434 446530
rect 703490 446474 703576 446530
rect 703632 446474 703718 446530
rect 703774 446474 703860 446530
rect 703916 446474 704002 446530
rect 704058 446474 704144 446530
rect 704200 446474 704286 446530
rect 704342 446515 705525 446530
rect 705581 446515 705649 446571
rect 705705 446515 705773 446571
rect 705829 446515 705897 446571
rect 705953 446515 706000 446571
rect 704342 446474 706000 446515
rect 702392 446447 706000 446474
rect 702392 446391 705525 446447
rect 705581 446391 705649 446447
rect 705705 446391 705773 446447
rect 705829 446391 705897 446447
rect 705953 446391 706000 446447
rect 702392 446388 706000 446391
rect 702392 446332 702440 446388
rect 702496 446332 702582 446388
rect 702638 446332 702724 446388
rect 702780 446332 702866 446388
rect 702922 446332 703008 446388
rect 703064 446332 703150 446388
rect 703206 446332 703292 446388
rect 703348 446332 703434 446388
rect 703490 446332 703576 446388
rect 703632 446332 703718 446388
rect 703774 446332 703860 446388
rect 703916 446332 704002 446388
rect 704058 446332 704144 446388
rect 704200 446332 704286 446388
rect 704342 446332 706000 446388
rect 702392 446323 706000 446332
rect 702392 446267 705525 446323
rect 705581 446267 705649 446323
rect 705705 446267 705773 446323
rect 705829 446267 705897 446323
rect 705953 446267 706000 446323
rect 702392 446246 706000 446267
rect 702392 446190 702440 446246
rect 702496 446190 702582 446246
rect 702638 446190 702724 446246
rect 702780 446190 702866 446246
rect 702922 446190 703008 446246
rect 703064 446190 703150 446246
rect 703206 446190 703292 446246
rect 703348 446190 703434 446246
rect 703490 446190 703576 446246
rect 703632 446190 703718 446246
rect 703774 446190 703860 446246
rect 703916 446190 704002 446246
rect 704058 446190 704144 446246
rect 704200 446190 704286 446246
rect 704342 446199 706000 446246
rect 704342 446190 705525 446199
rect 702392 446143 705525 446190
rect 705581 446143 705649 446199
rect 705705 446143 705773 446199
rect 705829 446143 705897 446199
rect 705953 446143 706000 446199
rect 702392 446104 706000 446143
rect 702392 446048 702440 446104
rect 702496 446048 702582 446104
rect 702638 446048 702724 446104
rect 702780 446048 702866 446104
rect 702922 446048 703008 446104
rect 703064 446048 703150 446104
rect 703206 446048 703292 446104
rect 703348 446048 703434 446104
rect 703490 446048 703576 446104
rect 703632 446048 703718 446104
rect 703774 446048 703860 446104
rect 703916 446048 704002 446104
rect 704058 446048 704144 446104
rect 704200 446048 704286 446104
rect 704342 446075 706000 446104
rect 704342 446048 705525 446075
rect 702392 446019 705525 446048
rect 705581 446019 705649 446075
rect 705705 446019 705773 446075
rect 705829 446019 705897 446075
rect 705953 446019 706000 446075
rect 702392 445962 706000 446019
rect 702392 445906 702440 445962
rect 702496 445906 702582 445962
rect 702638 445906 702724 445962
rect 702780 445906 702866 445962
rect 702922 445906 703008 445962
rect 703064 445906 703150 445962
rect 703206 445906 703292 445962
rect 703348 445906 703434 445962
rect 703490 445906 703576 445962
rect 703632 445906 703718 445962
rect 703774 445906 703860 445962
rect 703916 445906 704002 445962
rect 704058 445906 704144 445962
rect 704200 445906 704286 445962
rect 704342 445951 706000 445962
rect 704342 445906 705525 445951
rect 702392 445895 705525 445906
rect 705581 445895 705649 445951
rect 705705 445895 705773 445951
rect 705829 445895 705897 445951
rect 705953 445895 706000 445951
rect 702392 445828 706000 445895
rect 702392 445181 706000 445248
rect 702392 445179 705525 445181
rect 702392 445123 702451 445179
rect 702507 445123 702593 445179
rect 702649 445123 702735 445179
rect 702791 445123 702877 445179
rect 702933 445123 703019 445179
rect 703075 445123 703161 445179
rect 703217 445123 703303 445179
rect 703359 445123 703445 445179
rect 703501 445123 703587 445179
rect 703643 445123 703729 445179
rect 703785 445123 703871 445179
rect 703927 445123 704013 445179
rect 704069 445123 704155 445179
rect 704211 445123 704297 445179
rect 704353 445125 705525 445179
rect 705581 445125 705649 445181
rect 705705 445125 705773 445181
rect 705829 445125 705897 445181
rect 705953 445125 706000 445181
rect 704353 445123 706000 445125
rect 702392 445057 706000 445123
rect 702392 445037 705525 445057
rect 702392 444981 702451 445037
rect 702507 444981 702593 445037
rect 702649 444981 702735 445037
rect 702791 444981 702877 445037
rect 702933 444981 703019 445037
rect 703075 444981 703161 445037
rect 703217 444981 703303 445037
rect 703359 444981 703445 445037
rect 703501 444981 703587 445037
rect 703643 444981 703729 445037
rect 703785 444981 703871 445037
rect 703927 444981 704013 445037
rect 704069 444981 704155 445037
rect 704211 444981 704297 445037
rect 704353 445001 705525 445037
rect 705581 445001 705649 445057
rect 705705 445001 705773 445057
rect 705829 445001 705897 445057
rect 705953 445001 706000 445057
rect 704353 444981 706000 445001
rect 702392 444933 706000 444981
rect 702392 444895 705525 444933
rect 702392 444839 702451 444895
rect 702507 444839 702593 444895
rect 702649 444839 702735 444895
rect 702791 444839 702877 444895
rect 702933 444839 703019 444895
rect 703075 444839 703161 444895
rect 703217 444839 703303 444895
rect 703359 444839 703445 444895
rect 703501 444839 703587 444895
rect 703643 444839 703729 444895
rect 703785 444839 703871 444895
rect 703927 444839 704013 444895
rect 704069 444839 704155 444895
rect 704211 444839 704297 444895
rect 704353 444877 705525 444895
rect 705581 444877 705649 444933
rect 705705 444877 705773 444933
rect 705829 444877 705897 444933
rect 705953 444877 706000 444933
rect 704353 444839 706000 444877
rect 702392 444809 706000 444839
rect 702392 444753 705525 444809
rect 705581 444753 705649 444809
rect 705705 444753 705773 444809
rect 705829 444753 705897 444809
rect 705953 444753 706000 444809
rect 702392 444697 702451 444753
rect 702507 444697 702593 444753
rect 702649 444697 702735 444753
rect 702791 444697 702877 444753
rect 702933 444697 703019 444753
rect 703075 444697 703161 444753
rect 703217 444697 703303 444753
rect 703359 444697 703445 444753
rect 703501 444697 703587 444753
rect 703643 444697 703729 444753
rect 703785 444697 703871 444753
rect 703927 444697 704013 444753
rect 704069 444697 704155 444753
rect 704211 444697 704297 444753
rect 704353 444697 706000 444753
rect 702392 444685 706000 444697
rect 702392 444629 705525 444685
rect 705581 444629 705649 444685
rect 705705 444629 705773 444685
rect 705829 444629 705897 444685
rect 705953 444629 706000 444685
rect 702392 444611 706000 444629
rect 702392 444555 702451 444611
rect 702507 444555 702593 444611
rect 702649 444555 702735 444611
rect 702791 444555 702877 444611
rect 702933 444555 703019 444611
rect 703075 444555 703161 444611
rect 703217 444555 703303 444611
rect 703359 444555 703445 444611
rect 703501 444555 703587 444611
rect 703643 444555 703729 444611
rect 703785 444555 703871 444611
rect 703927 444555 704013 444611
rect 704069 444555 704155 444611
rect 704211 444555 704297 444611
rect 704353 444561 706000 444611
rect 704353 444555 705525 444561
rect 702392 444505 705525 444555
rect 705581 444505 705649 444561
rect 705705 444505 705773 444561
rect 705829 444505 705897 444561
rect 705953 444505 706000 444561
rect 702392 444469 706000 444505
rect 702392 444413 702451 444469
rect 702507 444413 702593 444469
rect 702649 444413 702735 444469
rect 702791 444413 702877 444469
rect 702933 444413 703019 444469
rect 703075 444413 703161 444469
rect 703217 444413 703303 444469
rect 703359 444413 703445 444469
rect 703501 444413 703587 444469
rect 703643 444413 703729 444469
rect 703785 444413 703871 444469
rect 703927 444413 704013 444469
rect 704069 444413 704155 444469
rect 704211 444413 704297 444469
rect 704353 444437 706000 444469
rect 704353 444413 705525 444437
rect 702392 444381 705525 444413
rect 705581 444381 705649 444437
rect 705705 444381 705773 444437
rect 705829 444381 705897 444437
rect 705953 444381 706000 444437
rect 702392 444327 706000 444381
rect 702392 444271 702451 444327
rect 702507 444271 702593 444327
rect 702649 444271 702735 444327
rect 702791 444271 702877 444327
rect 702933 444271 703019 444327
rect 703075 444271 703161 444327
rect 703217 444271 703303 444327
rect 703359 444271 703445 444327
rect 703501 444271 703587 444327
rect 703643 444271 703729 444327
rect 703785 444271 703871 444327
rect 703927 444271 704013 444327
rect 704069 444271 704155 444327
rect 704211 444271 704297 444327
rect 704353 444313 706000 444327
rect 704353 444271 705525 444313
rect 702392 444257 705525 444271
rect 705581 444257 705649 444313
rect 705705 444257 705773 444313
rect 705829 444257 705897 444313
rect 705953 444257 706000 444313
rect 702392 444189 706000 444257
rect 702392 444185 705525 444189
rect 702392 444129 702451 444185
rect 702507 444129 702593 444185
rect 702649 444129 702735 444185
rect 702791 444129 702877 444185
rect 702933 444129 703019 444185
rect 703075 444129 703161 444185
rect 703217 444129 703303 444185
rect 703359 444129 703445 444185
rect 703501 444129 703587 444185
rect 703643 444129 703729 444185
rect 703785 444129 703871 444185
rect 703927 444129 704013 444185
rect 704069 444129 704155 444185
rect 704211 444129 704297 444185
rect 704353 444133 705525 444185
rect 705581 444133 705649 444189
rect 705705 444133 705773 444189
rect 705829 444133 705897 444189
rect 705953 444133 706000 444189
rect 704353 444129 706000 444133
rect 702392 444065 706000 444129
rect 702392 444043 705525 444065
rect 702392 443987 702451 444043
rect 702507 443987 702593 444043
rect 702649 443987 702735 444043
rect 702791 443987 702877 444043
rect 702933 443987 703019 444043
rect 703075 443987 703161 444043
rect 703217 443987 703303 444043
rect 703359 443987 703445 444043
rect 703501 443987 703587 444043
rect 703643 443987 703729 444043
rect 703785 443987 703871 444043
rect 703927 443987 704013 444043
rect 704069 443987 704155 444043
rect 704211 443987 704297 444043
rect 704353 444009 705525 444043
rect 705581 444009 705649 444065
rect 705705 444009 705773 444065
rect 705829 444009 705897 444065
rect 705953 444009 706000 444065
rect 704353 443987 706000 444009
rect 702392 443941 706000 443987
rect 702392 443901 705525 443941
rect 702392 443845 702451 443901
rect 702507 443845 702593 443901
rect 702649 443845 702735 443901
rect 702791 443845 702877 443901
rect 702933 443845 703019 443901
rect 703075 443845 703161 443901
rect 703217 443845 703303 443901
rect 703359 443845 703445 443901
rect 703501 443845 703587 443901
rect 703643 443845 703729 443901
rect 703785 443845 703871 443901
rect 703927 443845 704013 443901
rect 704069 443845 704155 443901
rect 704211 443845 704297 443901
rect 704353 443885 705525 443901
rect 705581 443885 705649 443941
rect 705705 443885 705773 443941
rect 705829 443885 705897 443941
rect 705953 443885 706000 443941
rect 704353 443845 706000 443885
rect 702392 443817 706000 443845
rect 702392 443761 705525 443817
rect 705581 443761 705649 443817
rect 705705 443761 705773 443817
rect 705829 443761 705897 443817
rect 705953 443761 706000 443817
rect 702392 443759 706000 443761
rect 702392 443703 702451 443759
rect 702507 443703 702593 443759
rect 702649 443703 702735 443759
rect 702791 443703 702877 443759
rect 702933 443703 703019 443759
rect 703075 443703 703161 443759
rect 703217 443703 703303 443759
rect 703359 443703 703445 443759
rect 703501 443703 703587 443759
rect 703643 443703 703729 443759
rect 703785 443703 703871 443759
rect 703927 443703 704013 443759
rect 704069 443703 704155 443759
rect 704211 443703 704297 443759
rect 704353 443703 706000 443759
rect 702392 443693 706000 443703
rect 702392 443637 705525 443693
rect 705581 443637 705649 443693
rect 705705 443637 705773 443693
rect 705829 443637 705897 443693
rect 705953 443637 706000 443693
rect 702392 443617 706000 443637
rect 702392 443561 702451 443617
rect 702507 443561 702593 443617
rect 702649 443561 702735 443617
rect 702791 443561 702877 443617
rect 702933 443561 703019 443617
rect 703075 443561 703161 443617
rect 703217 443561 703303 443617
rect 703359 443561 703445 443617
rect 703501 443561 703587 443617
rect 703643 443561 703729 443617
rect 703785 443561 703871 443617
rect 703927 443561 704013 443617
rect 704069 443561 704155 443617
rect 704211 443561 704297 443617
rect 704353 443569 706000 443617
rect 704353 443561 705525 443569
rect 702392 443513 705525 443561
rect 705581 443513 705649 443569
rect 705705 443513 705773 443569
rect 705829 443513 705897 443569
rect 705953 443513 706000 443569
rect 702392 443475 706000 443513
rect 702392 443419 702451 443475
rect 702507 443419 702593 443475
rect 702649 443419 702735 443475
rect 702791 443419 702877 443475
rect 702933 443419 703019 443475
rect 703075 443419 703161 443475
rect 703217 443419 703303 443475
rect 703359 443419 703445 443475
rect 703501 443419 703587 443475
rect 703643 443419 703729 443475
rect 703785 443419 703871 443475
rect 703927 443419 704013 443475
rect 704069 443419 704155 443475
rect 704211 443419 704297 443475
rect 704353 443445 706000 443475
rect 704353 443419 705525 443445
rect 702392 443389 705525 443419
rect 705581 443389 705649 443445
rect 705705 443389 705773 443445
rect 705829 443389 705897 443445
rect 705953 443389 706000 443445
rect 702392 443333 706000 443389
rect 702392 443277 702451 443333
rect 702507 443277 702593 443333
rect 702649 443277 702735 443333
rect 702791 443277 702877 443333
rect 702933 443277 703019 443333
rect 703075 443277 703161 443333
rect 703217 443277 703303 443333
rect 703359 443277 703445 443333
rect 703501 443277 703587 443333
rect 703643 443277 703729 443333
rect 703785 443277 703871 443333
rect 703927 443277 704013 443333
rect 704069 443277 704155 443333
rect 704211 443277 704297 443333
rect 704353 443321 706000 443333
rect 704353 443277 705525 443321
rect 702392 443265 705525 443277
rect 705581 443265 705649 443321
rect 705705 443265 705773 443321
rect 705829 443265 705897 443321
rect 705953 443265 706000 443321
rect 702392 443198 706000 443265
rect 702392 442811 706000 442878
rect 702392 442809 705525 442811
rect 702392 442753 702451 442809
rect 702507 442753 702593 442809
rect 702649 442753 702735 442809
rect 702791 442753 702877 442809
rect 702933 442753 703019 442809
rect 703075 442753 703161 442809
rect 703217 442753 703303 442809
rect 703359 442753 703445 442809
rect 703501 442753 703587 442809
rect 703643 442753 703729 442809
rect 703785 442753 703871 442809
rect 703927 442753 704013 442809
rect 704069 442753 704155 442809
rect 704211 442753 704297 442809
rect 704353 442755 705525 442809
rect 705581 442755 705649 442811
rect 705705 442755 705773 442811
rect 705829 442755 705897 442811
rect 705953 442755 706000 442811
rect 704353 442753 706000 442755
rect 702392 442687 706000 442753
rect 702392 442667 705525 442687
rect 702392 442611 702451 442667
rect 702507 442611 702593 442667
rect 702649 442611 702735 442667
rect 702791 442611 702877 442667
rect 702933 442611 703019 442667
rect 703075 442611 703161 442667
rect 703217 442611 703303 442667
rect 703359 442611 703445 442667
rect 703501 442611 703587 442667
rect 703643 442611 703729 442667
rect 703785 442611 703871 442667
rect 703927 442611 704013 442667
rect 704069 442611 704155 442667
rect 704211 442611 704297 442667
rect 704353 442631 705525 442667
rect 705581 442631 705649 442687
rect 705705 442631 705773 442687
rect 705829 442631 705897 442687
rect 705953 442631 706000 442687
rect 704353 442611 706000 442631
rect 702392 442563 706000 442611
rect 702392 442525 705525 442563
rect 702392 442469 702451 442525
rect 702507 442469 702593 442525
rect 702649 442469 702735 442525
rect 702791 442469 702877 442525
rect 702933 442469 703019 442525
rect 703075 442469 703161 442525
rect 703217 442469 703303 442525
rect 703359 442469 703445 442525
rect 703501 442469 703587 442525
rect 703643 442469 703729 442525
rect 703785 442469 703871 442525
rect 703927 442469 704013 442525
rect 704069 442469 704155 442525
rect 704211 442469 704297 442525
rect 704353 442507 705525 442525
rect 705581 442507 705649 442563
rect 705705 442507 705773 442563
rect 705829 442507 705897 442563
rect 705953 442507 706000 442563
rect 704353 442469 706000 442507
rect 702392 442439 706000 442469
rect 702392 442383 705525 442439
rect 705581 442383 705649 442439
rect 705705 442383 705773 442439
rect 705829 442383 705897 442439
rect 705953 442383 706000 442439
rect 702392 442327 702451 442383
rect 702507 442327 702593 442383
rect 702649 442327 702735 442383
rect 702791 442327 702877 442383
rect 702933 442327 703019 442383
rect 703075 442327 703161 442383
rect 703217 442327 703303 442383
rect 703359 442327 703445 442383
rect 703501 442327 703587 442383
rect 703643 442327 703729 442383
rect 703785 442327 703871 442383
rect 703927 442327 704013 442383
rect 704069 442327 704155 442383
rect 704211 442327 704297 442383
rect 704353 442327 706000 442383
rect 702392 442315 706000 442327
rect 702392 442259 705525 442315
rect 705581 442259 705649 442315
rect 705705 442259 705773 442315
rect 705829 442259 705897 442315
rect 705953 442259 706000 442315
rect 702392 442241 706000 442259
rect 702392 442185 702451 442241
rect 702507 442185 702593 442241
rect 702649 442185 702735 442241
rect 702791 442185 702877 442241
rect 702933 442185 703019 442241
rect 703075 442185 703161 442241
rect 703217 442185 703303 442241
rect 703359 442185 703445 442241
rect 703501 442185 703587 442241
rect 703643 442185 703729 442241
rect 703785 442185 703871 442241
rect 703927 442185 704013 442241
rect 704069 442185 704155 442241
rect 704211 442185 704297 442241
rect 704353 442191 706000 442241
rect 704353 442185 705525 442191
rect 702392 442135 705525 442185
rect 705581 442135 705649 442191
rect 705705 442135 705773 442191
rect 705829 442135 705897 442191
rect 705953 442135 706000 442191
rect 702392 442099 706000 442135
rect 702392 442043 702451 442099
rect 702507 442043 702593 442099
rect 702649 442043 702735 442099
rect 702791 442043 702877 442099
rect 702933 442043 703019 442099
rect 703075 442043 703161 442099
rect 703217 442043 703303 442099
rect 703359 442043 703445 442099
rect 703501 442043 703587 442099
rect 703643 442043 703729 442099
rect 703785 442043 703871 442099
rect 703927 442043 704013 442099
rect 704069 442043 704155 442099
rect 704211 442043 704297 442099
rect 704353 442067 706000 442099
rect 704353 442043 705525 442067
rect 702392 442011 705525 442043
rect 705581 442011 705649 442067
rect 705705 442011 705773 442067
rect 705829 442011 705897 442067
rect 705953 442011 706000 442067
rect 702392 441957 706000 442011
rect 702392 441901 702451 441957
rect 702507 441901 702593 441957
rect 702649 441901 702735 441957
rect 702791 441901 702877 441957
rect 702933 441901 703019 441957
rect 703075 441901 703161 441957
rect 703217 441901 703303 441957
rect 703359 441901 703445 441957
rect 703501 441901 703587 441957
rect 703643 441901 703729 441957
rect 703785 441901 703871 441957
rect 703927 441901 704013 441957
rect 704069 441901 704155 441957
rect 704211 441901 704297 441957
rect 704353 441943 706000 441957
rect 704353 441901 705525 441943
rect 702392 441887 705525 441901
rect 705581 441887 705649 441943
rect 705705 441887 705773 441943
rect 705829 441887 705897 441943
rect 705953 441887 706000 441943
rect 702392 441819 706000 441887
rect 702392 441815 705525 441819
rect 702392 441759 702451 441815
rect 702507 441759 702593 441815
rect 702649 441759 702735 441815
rect 702791 441759 702877 441815
rect 702933 441759 703019 441815
rect 703075 441759 703161 441815
rect 703217 441759 703303 441815
rect 703359 441759 703445 441815
rect 703501 441759 703587 441815
rect 703643 441759 703729 441815
rect 703785 441759 703871 441815
rect 703927 441759 704013 441815
rect 704069 441759 704155 441815
rect 704211 441759 704297 441815
rect 704353 441763 705525 441815
rect 705581 441763 705649 441819
rect 705705 441763 705773 441819
rect 705829 441763 705897 441819
rect 705953 441763 706000 441819
rect 704353 441759 706000 441763
rect 702392 441695 706000 441759
rect 702392 441673 705525 441695
rect 702392 441617 702451 441673
rect 702507 441617 702593 441673
rect 702649 441617 702735 441673
rect 702791 441617 702877 441673
rect 702933 441617 703019 441673
rect 703075 441617 703161 441673
rect 703217 441617 703303 441673
rect 703359 441617 703445 441673
rect 703501 441617 703587 441673
rect 703643 441617 703729 441673
rect 703785 441617 703871 441673
rect 703927 441617 704013 441673
rect 704069 441617 704155 441673
rect 704211 441617 704297 441673
rect 704353 441639 705525 441673
rect 705581 441639 705649 441695
rect 705705 441639 705773 441695
rect 705829 441639 705897 441695
rect 705953 441639 706000 441695
rect 704353 441617 706000 441639
rect 702392 441571 706000 441617
rect 702392 441531 705525 441571
rect 702392 441475 702451 441531
rect 702507 441475 702593 441531
rect 702649 441475 702735 441531
rect 702791 441475 702877 441531
rect 702933 441475 703019 441531
rect 703075 441475 703161 441531
rect 703217 441475 703303 441531
rect 703359 441475 703445 441531
rect 703501 441475 703587 441531
rect 703643 441475 703729 441531
rect 703785 441475 703871 441531
rect 703927 441475 704013 441531
rect 704069 441475 704155 441531
rect 704211 441475 704297 441531
rect 704353 441515 705525 441531
rect 705581 441515 705649 441571
rect 705705 441515 705773 441571
rect 705829 441515 705897 441571
rect 705953 441515 706000 441571
rect 704353 441475 706000 441515
rect 702392 441447 706000 441475
rect 702392 441391 705525 441447
rect 705581 441391 705649 441447
rect 705705 441391 705773 441447
rect 705829 441391 705897 441447
rect 705953 441391 706000 441447
rect 702392 441389 706000 441391
rect 702392 441333 702451 441389
rect 702507 441333 702593 441389
rect 702649 441333 702735 441389
rect 702791 441333 702877 441389
rect 702933 441333 703019 441389
rect 703075 441333 703161 441389
rect 703217 441333 703303 441389
rect 703359 441333 703445 441389
rect 703501 441333 703587 441389
rect 703643 441333 703729 441389
rect 703785 441333 703871 441389
rect 703927 441333 704013 441389
rect 704069 441333 704155 441389
rect 704211 441333 704297 441389
rect 704353 441333 706000 441389
rect 702392 441323 706000 441333
rect 702392 441267 705525 441323
rect 705581 441267 705649 441323
rect 705705 441267 705773 441323
rect 705829 441267 705897 441323
rect 705953 441267 706000 441323
rect 702392 441247 706000 441267
rect 702392 441191 702451 441247
rect 702507 441191 702593 441247
rect 702649 441191 702735 441247
rect 702791 441191 702877 441247
rect 702933 441191 703019 441247
rect 703075 441191 703161 441247
rect 703217 441191 703303 441247
rect 703359 441191 703445 441247
rect 703501 441191 703587 441247
rect 703643 441191 703729 441247
rect 703785 441191 703871 441247
rect 703927 441191 704013 441247
rect 704069 441191 704155 441247
rect 704211 441191 704297 441247
rect 704353 441199 706000 441247
rect 704353 441191 705525 441199
rect 702392 441143 705525 441191
rect 705581 441143 705649 441199
rect 705705 441143 705773 441199
rect 705829 441143 705897 441199
rect 705953 441143 706000 441199
rect 702392 441105 706000 441143
rect 702392 441049 702451 441105
rect 702507 441049 702593 441105
rect 702649 441049 702735 441105
rect 702791 441049 702877 441105
rect 702933 441049 703019 441105
rect 703075 441049 703161 441105
rect 703217 441049 703303 441105
rect 703359 441049 703445 441105
rect 703501 441049 703587 441105
rect 703643 441049 703729 441105
rect 703785 441049 703871 441105
rect 703927 441049 704013 441105
rect 704069 441049 704155 441105
rect 704211 441049 704297 441105
rect 704353 441075 706000 441105
rect 704353 441049 705525 441075
rect 702392 441019 705525 441049
rect 705581 441019 705649 441075
rect 705705 441019 705773 441075
rect 705829 441019 705897 441075
rect 705953 441019 706000 441075
rect 702392 440963 706000 441019
rect 702392 440907 702451 440963
rect 702507 440907 702593 440963
rect 702649 440907 702735 440963
rect 702791 440907 702877 440963
rect 702933 440907 703019 440963
rect 703075 440907 703161 440963
rect 703217 440907 703303 440963
rect 703359 440907 703445 440963
rect 703501 440907 703587 440963
rect 703643 440907 703729 440963
rect 703785 440907 703871 440963
rect 703927 440907 704013 440963
rect 704069 440907 704155 440963
rect 704211 440907 704297 440963
rect 704353 440951 706000 440963
rect 704353 440907 705525 440951
rect 702392 440895 705525 440907
rect 705581 440895 705649 440951
rect 705705 440895 705773 440951
rect 705829 440895 705897 440951
rect 705953 440895 706000 440951
rect 702392 440828 706000 440895
rect 702392 440105 706000 440172
rect 702392 440103 705525 440105
rect 702392 440047 702451 440103
rect 702507 440047 702593 440103
rect 702649 440047 702735 440103
rect 702791 440047 702877 440103
rect 702933 440047 703019 440103
rect 703075 440047 703161 440103
rect 703217 440047 703303 440103
rect 703359 440047 703445 440103
rect 703501 440047 703587 440103
rect 703643 440047 703729 440103
rect 703785 440047 703871 440103
rect 703927 440047 704013 440103
rect 704069 440047 704155 440103
rect 704211 440047 704297 440103
rect 704353 440049 705525 440103
rect 705581 440049 705649 440105
rect 705705 440049 705773 440105
rect 705829 440049 705897 440105
rect 705953 440049 706000 440105
rect 704353 440047 706000 440049
rect 702392 439981 706000 440047
rect 702392 439961 705525 439981
rect 702392 439905 702451 439961
rect 702507 439905 702593 439961
rect 702649 439905 702735 439961
rect 702791 439905 702877 439961
rect 702933 439905 703019 439961
rect 703075 439905 703161 439961
rect 703217 439905 703303 439961
rect 703359 439905 703445 439961
rect 703501 439905 703587 439961
rect 703643 439905 703729 439961
rect 703785 439905 703871 439961
rect 703927 439905 704013 439961
rect 704069 439905 704155 439961
rect 704211 439905 704297 439961
rect 704353 439925 705525 439961
rect 705581 439925 705649 439981
rect 705705 439925 705773 439981
rect 705829 439925 705897 439981
rect 705953 439925 706000 439981
rect 704353 439905 706000 439925
rect 702392 439857 706000 439905
rect 702392 439819 705525 439857
rect 702392 439763 702451 439819
rect 702507 439763 702593 439819
rect 702649 439763 702735 439819
rect 702791 439763 702877 439819
rect 702933 439763 703019 439819
rect 703075 439763 703161 439819
rect 703217 439763 703303 439819
rect 703359 439763 703445 439819
rect 703501 439763 703587 439819
rect 703643 439763 703729 439819
rect 703785 439763 703871 439819
rect 703927 439763 704013 439819
rect 704069 439763 704155 439819
rect 704211 439763 704297 439819
rect 704353 439801 705525 439819
rect 705581 439801 705649 439857
rect 705705 439801 705773 439857
rect 705829 439801 705897 439857
rect 705953 439801 706000 439857
rect 704353 439763 706000 439801
rect 702392 439733 706000 439763
rect 702392 439677 705525 439733
rect 705581 439677 705649 439733
rect 705705 439677 705773 439733
rect 705829 439677 705897 439733
rect 705953 439677 706000 439733
rect 702392 439621 702451 439677
rect 702507 439621 702593 439677
rect 702649 439621 702735 439677
rect 702791 439621 702877 439677
rect 702933 439621 703019 439677
rect 703075 439621 703161 439677
rect 703217 439621 703303 439677
rect 703359 439621 703445 439677
rect 703501 439621 703587 439677
rect 703643 439621 703729 439677
rect 703785 439621 703871 439677
rect 703927 439621 704013 439677
rect 704069 439621 704155 439677
rect 704211 439621 704297 439677
rect 704353 439621 706000 439677
rect 702392 439609 706000 439621
rect 702392 439553 705525 439609
rect 705581 439553 705649 439609
rect 705705 439553 705773 439609
rect 705829 439553 705897 439609
rect 705953 439553 706000 439609
rect 702392 439535 706000 439553
rect 702392 439479 702451 439535
rect 702507 439479 702593 439535
rect 702649 439479 702735 439535
rect 702791 439479 702877 439535
rect 702933 439479 703019 439535
rect 703075 439479 703161 439535
rect 703217 439479 703303 439535
rect 703359 439479 703445 439535
rect 703501 439479 703587 439535
rect 703643 439479 703729 439535
rect 703785 439479 703871 439535
rect 703927 439479 704013 439535
rect 704069 439479 704155 439535
rect 704211 439479 704297 439535
rect 704353 439485 706000 439535
rect 704353 439479 705525 439485
rect 702392 439429 705525 439479
rect 705581 439429 705649 439485
rect 705705 439429 705773 439485
rect 705829 439429 705897 439485
rect 705953 439429 706000 439485
rect 702392 439393 706000 439429
rect 702392 439337 702451 439393
rect 702507 439337 702593 439393
rect 702649 439337 702735 439393
rect 702791 439337 702877 439393
rect 702933 439337 703019 439393
rect 703075 439337 703161 439393
rect 703217 439337 703303 439393
rect 703359 439337 703445 439393
rect 703501 439337 703587 439393
rect 703643 439337 703729 439393
rect 703785 439337 703871 439393
rect 703927 439337 704013 439393
rect 704069 439337 704155 439393
rect 704211 439337 704297 439393
rect 704353 439361 706000 439393
rect 704353 439337 705525 439361
rect 702392 439305 705525 439337
rect 705581 439305 705649 439361
rect 705705 439305 705773 439361
rect 705829 439305 705897 439361
rect 705953 439305 706000 439361
rect 702392 439251 706000 439305
rect 702392 439195 702451 439251
rect 702507 439195 702593 439251
rect 702649 439195 702735 439251
rect 702791 439195 702877 439251
rect 702933 439195 703019 439251
rect 703075 439195 703161 439251
rect 703217 439195 703303 439251
rect 703359 439195 703445 439251
rect 703501 439195 703587 439251
rect 703643 439195 703729 439251
rect 703785 439195 703871 439251
rect 703927 439195 704013 439251
rect 704069 439195 704155 439251
rect 704211 439195 704297 439251
rect 704353 439237 706000 439251
rect 704353 439195 705525 439237
rect 702392 439181 705525 439195
rect 705581 439181 705649 439237
rect 705705 439181 705773 439237
rect 705829 439181 705897 439237
rect 705953 439181 706000 439237
rect 702392 439113 706000 439181
rect 702392 439109 705525 439113
rect 702392 439053 702451 439109
rect 702507 439053 702593 439109
rect 702649 439053 702735 439109
rect 702791 439053 702877 439109
rect 702933 439053 703019 439109
rect 703075 439053 703161 439109
rect 703217 439053 703303 439109
rect 703359 439053 703445 439109
rect 703501 439053 703587 439109
rect 703643 439053 703729 439109
rect 703785 439053 703871 439109
rect 703927 439053 704013 439109
rect 704069 439053 704155 439109
rect 704211 439053 704297 439109
rect 704353 439057 705525 439109
rect 705581 439057 705649 439113
rect 705705 439057 705773 439113
rect 705829 439057 705897 439113
rect 705953 439057 706000 439113
rect 704353 439053 706000 439057
rect 702392 438989 706000 439053
rect 702392 438967 705525 438989
rect 702392 438911 702451 438967
rect 702507 438911 702593 438967
rect 702649 438911 702735 438967
rect 702791 438911 702877 438967
rect 702933 438911 703019 438967
rect 703075 438911 703161 438967
rect 703217 438911 703303 438967
rect 703359 438911 703445 438967
rect 703501 438911 703587 438967
rect 703643 438911 703729 438967
rect 703785 438911 703871 438967
rect 703927 438911 704013 438967
rect 704069 438911 704155 438967
rect 704211 438911 704297 438967
rect 704353 438933 705525 438967
rect 705581 438933 705649 438989
rect 705705 438933 705773 438989
rect 705829 438933 705897 438989
rect 705953 438933 706000 438989
rect 704353 438911 706000 438933
rect 702392 438865 706000 438911
rect 702392 438825 705525 438865
rect 702392 438769 702451 438825
rect 702507 438769 702593 438825
rect 702649 438769 702735 438825
rect 702791 438769 702877 438825
rect 702933 438769 703019 438825
rect 703075 438769 703161 438825
rect 703217 438769 703303 438825
rect 703359 438769 703445 438825
rect 703501 438769 703587 438825
rect 703643 438769 703729 438825
rect 703785 438769 703871 438825
rect 703927 438769 704013 438825
rect 704069 438769 704155 438825
rect 704211 438769 704297 438825
rect 704353 438809 705525 438825
rect 705581 438809 705649 438865
rect 705705 438809 705773 438865
rect 705829 438809 705897 438865
rect 705953 438809 706000 438865
rect 704353 438769 706000 438809
rect 702392 438741 706000 438769
rect 702392 438685 705525 438741
rect 705581 438685 705649 438741
rect 705705 438685 705773 438741
rect 705829 438685 705897 438741
rect 705953 438685 706000 438741
rect 702392 438683 706000 438685
rect 702392 438627 702451 438683
rect 702507 438627 702593 438683
rect 702649 438627 702735 438683
rect 702791 438627 702877 438683
rect 702933 438627 703019 438683
rect 703075 438627 703161 438683
rect 703217 438627 703303 438683
rect 703359 438627 703445 438683
rect 703501 438627 703587 438683
rect 703643 438627 703729 438683
rect 703785 438627 703871 438683
rect 703927 438627 704013 438683
rect 704069 438627 704155 438683
rect 704211 438627 704297 438683
rect 704353 438627 706000 438683
rect 702392 438617 706000 438627
rect 702392 438561 705525 438617
rect 705581 438561 705649 438617
rect 705705 438561 705773 438617
rect 705829 438561 705897 438617
rect 705953 438561 706000 438617
rect 702392 438541 706000 438561
rect 702392 438485 702451 438541
rect 702507 438485 702593 438541
rect 702649 438485 702735 438541
rect 702791 438485 702877 438541
rect 702933 438485 703019 438541
rect 703075 438485 703161 438541
rect 703217 438485 703303 438541
rect 703359 438485 703445 438541
rect 703501 438485 703587 438541
rect 703643 438485 703729 438541
rect 703785 438485 703871 438541
rect 703927 438485 704013 438541
rect 704069 438485 704155 438541
rect 704211 438485 704297 438541
rect 704353 438493 706000 438541
rect 704353 438485 705525 438493
rect 702392 438437 705525 438485
rect 705581 438437 705649 438493
rect 705705 438437 705773 438493
rect 705829 438437 705897 438493
rect 705953 438437 706000 438493
rect 702392 438399 706000 438437
rect 702392 438343 702451 438399
rect 702507 438343 702593 438399
rect 702649 438343 702735 438399
rect 702791 438343 702877 438399
rect 702933 438343 703019 438399
rect 703075 438343 703161 438399
rect 703217 438343 703303 438399
rect 703359 438343 703445 438399
rect 703501 438343 703587 438399
rect 703643 438343 703729 438399
rect 703785 438343 703871 438399
rect 703927 438343 704013 438399
rect 704069 438343 704155 438399
rect 704211 438343 704297 438399
rect 704353 438369 706000 438399
rect 704353 438343 705525 438369
rect 702392 438313 705525 438343
rect 705581 438313 705649 438369
rect 705705 438313 705773 438369
rect 705829 438313 705897 438369
rect 705953 438313 706000 438369
rect 702392 438257 706000 438313
rect 702392 438201 702451 438257
rect 702507 438201 702593 438257
rect 702649 438201 702735 438257
rect 702791 438201 702877 438257
rect 702933 438201 703019 438257
rect 703075 438201 703161 438257
rect 703217 438201 703303 438257
rect 703359 438201 703445 438257
rect 703501 438201 703587 438257
rect 703643 438201 703729 438257
rect 703785 438201 703871 438257
rect 703927 438201 704013 438257
rect 704069 438201 704155 438257
rect 704211 438201 704297 438257
rect 704353 438245 706000 438257
rect 704353 438201 705525 438245
rect 702392 438189 705525 438201
rect 705581 438189 705649 438245
rect 705705 438189 705773 438245
rect 705829 438189 705897 438245
rect 705953 438189 706000 438245
rect 702392 438122 706000 438189
rect 702392 437735 706000 437802
rect 702392 437733 705525 437735
rect 702392 437677 702451 437733
rect 702507 437677 702593 437733
rect 702649 437677 702735 437733
rect 702791 437677 702877 437733
rect 702933 437677 703019 437733
rect 703075 437677 703161 437733
rect 703217 437677 703303 437733
rect 703359 437677 703445 437733
rect 703501 437677 703587 437733
rect 703643 437677 703729 437733
rect 703785 437677 703871 437733
rect 703927 437677 704013 437733
rect 704069 437677 704155 437733
rect 704211 437677 704297 437733
rect 704353 437679 705525 437733
rect 705581 437679 705649 437735
rect 705705 437679 705773 437735
rect 705829 437679 705897 437735
rect 705953 437679 706000 437735
rect 704353 437677 706000 437679
rect 702392 437611 706000 437677
rect 702392 437591 705525 437611
rect 702392 437535 702451 437591
rect 702507 437535 702593 437591
rect 702649 437535 702735 437591
rect 702791 437535 702877 437591
rect 702933 437535 703019 437591
rect 703075 437535 703161 437591
rect 703217 437535 703303 437591
rect 703359 437535 703445 437591
rect 703501 437535 703587 437591
rect 703643 437535 703729 437591
rect 703785 437535 703871 437591
rect 703927 437535 704013 437591
rect 704069 437535 704155 437591
rect 704211 437535 704297 437591
rect 704353 437555 705525 437591
rect 705581 437555 705649 437611
rect 705705 437555 705773 437611
rect 705829 437555 705897 437611
rect 705953 437555 706000 437611
rect 704353 437535 706000 437555
rect 702392 437487 706000 437535
rect 702392 437449 705525 437487
rect 702392 437393 702451 437449
rect 702507 437393 702593 437449
rect 702649 437393 702735 437449
rect 702791 437393 702877 437449
rect 702933 437393 703019 437449
rect 703075 437393 703161 437449
rect 703217 437393 703303 437449
rect 703359 437393 703445 437449
rect 703501 437393 703587 437449
rect 703643 437393 703729 437449
rect 703785 437393 703871 437449
rect 703927 437393 704013 437449
rect 704069 437393 704155 437449
rect 704211 437393 704297 437449
rect 704353 437431 705525 437449
rect 705581 437431 705649 437487
rect 705705 437431 705773 437487
rect 705829 437431 705897 437487
rect 705953 437431 706000 437487
rect 704353 437393 706000 437431
rect 702392 437363 706000 437393
rect 702392 437307 705525 437363
rect 705581 437307 705649 437363
rect 705705 437307 705773 437363
rect 705829 437307 705897 437363
rect 705953 437307 706000 437363
rect 702392 437251 702451 437307
rect 702507 437251 702593 437307
rect 702649 437251 702735 437307
rect 702791 437251 702877 437307
rect 702933 437251 703019 437307
rect 703075 437251 703161 437307
rect 703217 437251 703303 437307
rect 703359 437251 703445 437307
rect 703501 437251 703587 437307
rect 703643 437251 703729 437307
rect 703785 437251 703871 437307
rect 703927 437251 704013 437307
rect 704069 437251 704155 437307
rect 704211 437251 704297 437307
rect 704353 437251 706000 437307
rect 702392 437239 706000 437251
rect 702392 437183 705525 437239
rect 705581 437183 705649 437239
rect 705705 437183 705773 437239
rect 705829 437183 705897 437239
rect 705953 437183 706000 437239
rect 702392 437165 706000 437183
rect 702392 437109 702451 437165
rect 702507 437109 702593 437165
rect 702649 437109 702735 437165
rect 702791 437109 702877 437165
rect 702933 437109 703019 437165
rect 703075 437109 703161 437165
rect 703217 437109 703303 437165
rect 703359 437109 703445 437165
rect 703501 437109 703587 437165
rect 703643 437109 703729 437165
rect 703785 437109 703871 437165
rect 703927 437109 704013 437165
rect 704069 437109 704155 437165
rect 704211 437109 704297 437165
rect 704353 437115 706000 437165
rect 704353 437109 705525 437115
rect 702392 437059 705525 437109
rect 705581 437059 705649 437115
rect 705705 437059 705773 437115
rect 705829 437059 705897 437115
rect 705953 437059 706000 437115
rect 702392 437023 706000 437059
rect 702392 436967 702451 437023
rect 702507 436967 702593 437023
rect 702649 436967 702735 437023
rect 702791 436967 702877 437023
rect 702933 436967 703019 437023
rect 703075 436967 703161 437023
rect 703217 436967 703303 437023
rect 703359 436967 703445 437023
rect 703501 436967 703587 437023
rect 703643 436967 703729 437023
rect 703785 436967 703871 437023
rect 703927 436967 704013 437023
rect 704069 436967 704155 437023
rect 704211 436967 704297 437023
rect 704353 436991 706000 437023
rect 704353 436967 705525 436991
rect 702392 436935 705525 436967
rect 705581 436935 705649 436991
rect 705705 436935 705773 436991
rect 705829 436935 705897 436991
rect 705953 436935 706000 436991
rect 702392 436881 706000 436935
rect 702392 436825 702451 436881
rect 702507 436825 702593 436881
rect 702649 436825 702735 436881
rect 702791 436825 702877 436881
rect 702933 436825 703019 436881
rect 703075 436825 703161 436881
rect 703217 436825 703303 436881
rect 703359 436825 703445 436881
rect 703501 436825 703587 436881
rect 703643 436825 703729 436881
rect 703785 436825 703871 436881
rect 703927 436825 704013 436881
rect 704069 436825 704155 436881
rect 704211 436825 704297 436881
rect 704353 436867 706000 436881
rect 704353 436825 705525 436867
rect 702392 436811 705525 436825
rect 705581 436811 705649 436867
rect 705705 436811 705773 436867
rect 705829 436811 705897 436867
rect 705953 436811 706000 436867
rect 702392 436743 706000 436811
rect 702392 436739 705525 436743
rect 702392 436683 702451 436739
rect 702507 436683 702593 436739
rect 702649 436683 702735 436739
rect 702791 436683 702877 436739
rect 702933 436683 703019 436739
rect 703075 436683 703161 436739
rect 703217 436683 703303 436739
rect 703359 436683 703445 436739
rect 703501 436683 703587 436739
rect 703643 436683 703729 436739
rect 703785 436683 703871 436739
rect 703927 436683 704013 436739
rect 704069 436683 704155 436739
rect 704211 436683 704297 436739
rect 704353 436687 705525 436739
rect 705581 436687 705649 436743
rect 705705 436687 705773 436743
rect 705829 436687 705897 436743
rect 705953 436687 706000 436743
rect 704353 436683 706000 436687
rect 702392 436619 706000 436683
rect 702392 436597 705525 436619
rect 702392 436541 702451 436597
rect 702507 436541 702593 436597
rect 702649 436541 702735 436597
rect 702791 436541 702877 436597
rect 702933 436541 703019 436597
rect 703075 436541 703161 436597
rect 703217 436541 703303 436597
rect 703359 436541 703445 436597
rect 703501 436541 703587 436597
rect 703643 436541 703729 436597
rect 703785 436541 703871 436597
rect 703927 436541 704013 436597
rect 704069 436541 704155 436597
rect 704211 436541 704297 436597
rect 704353 436563 705525 436597
rect 705581 436563 705649 436619
rect 705705 436563 705773 436619
rect 705829 436563 705897 436619
rect 705953 436563 706000 436619
rect 704353 436541 706000 436563
rect 702392 436495 706000 436541
rect 702392 436455 705525 436495
rect 702392 436399 702451 436455
rect 702507 436399 702593 436455
rect 702649 436399 702735 436455
rect 702791 436399 702877 436455
rect 702933 436399 703019 436455
rect 703075 436399 703161 436455
rect 703217 436399 703303 436455
rect 703359 436399 703445 436455
rect 703501 436399 703587 436455
rect 703643 436399 703729 436455
rect 703785 436399 703871 436455
rect 703927 436399 704013 436455
rect 704069 436399 704155 436455
rect 704211 436399 704297 436455
rect 704353 436439 705525 436455
rect 705581 436439 705649 436495
rect 705705 436439 705773 436495
rect 705829 436439 705897 436495
rect 705953 436439 706000 436495
rect 704353 436399 706000 436439
rect 702392 436371 706000 436399
rect 702392 436315 705525 436371
rect 705581 436315 705649 436371
rect 705705 436315 705773 436371
rect 705829 436315 705897 436371
rect 705953 436315 706000 436371
rect 702392 436313 706000 436315
rect 702392 436257 702451 436313
rect 702507 436257 702593 436313
rect 702649 436257 702735 436313
rect 702791 436257 702877 436313
rect 702933 436257 703019 436313
rect 703075 436257 703161 436313
rect 703217 436257 703303 436313
rect 703359 436257 703445 436313
rect 703501 436257 703587 436313
rect 703643 436257 703729 436313
rect 703785 436257 703871 436313
rect 703927 436257 704013 436313
rect 704069 436257 704155 436313
rect 704211 436257 704297 436313
rect 704353 436257 706000 436313
rect 702392 436247 706000 436257
rect 702392 436191 705525 436247
rect 705581 436191 705649 436247
rect 705705 436191 705773 436247
rect 705829 436191 705897 436247
rect 705953 436191 706000 436247
rect 702392 436171 706000 436191
rect 702392 436115 702451 436171
rect 702507 436115 702593 436171
rect 702649 436115 702735 436171
rect 702791 436115 702877 436171
rect 702933 436115 703019 436171
rect 703075 436115 703161 436171
rect 703217 436115 703303 436171
rect 703359 436115 703445 436171
rect 703501 436115 703587 436171
rect 703643 436115 703729 436171
rect 703785 436115 703871 436171
rect 703927 436115 704013 436171
rect 704069 436115 704155 436171
rect 704211 436115 704297 436171
rect 704353 436115 706000 436171
rect 702392 436080 706000 436115
rect 702392 435131 706000 435172
rect 702392 435110 705525 435131
rect 702392 435054 702440 435110
rect 702496 435054 702582 435110
rect 702638 435054 702724 435110
rect 702780 435054 702866 435110
rect 702922 435054 703008 435110
rect 703064 435054 703150 435110
rect 703206 435054 703292 435110
rect 703348 435054 703434 435110
rect 703490 435054 703576 435110
rect 703632 435054 703718 435110
rect 703774 435054 703860 435110
rect 703916 435054 704002 435110
rect 704058 435054 704144 435110
rect 704200 435054 704286 435110
rect 704342 435075 705525 435110
rect 705581 435075 705649 435131
rect 705705 435075 705773 435131
rect 705829 435075 705897 435131
rect 705953 435075 706000 435131
rect 704342 435054 706000 435075
rect 702392 435007 706000 435054
rect 702392 434968 705525 435007
rect 702392 434912 702440 434968
rect 702496 434912 702582 434968
rect 702638 434912 702724 434968
rect 702780 434912 702866 434968
rect 702922 434912 703008 434968
rect 703064 434912 703150 434968
rect 703206 434912 703292 434968
rect 703348 434912 703434 434968
rect 703490 434912 703576 434968
rect 703632 434912 703718 434968
rect 703774 434912 703860 434968
rect 703916 434912 704002 434968
rect 704058 434912 704144 434968
rect 704200 434912 704286 434968
rect 704342 434951 705525 434968
rect 705581 434951 705649 435007
rect 705705 434951 705773 435007
rect 705829 434951 705897 435007
rect 705953 434951 706000 435007
rect 704342 434912 706000 434951
rect 702392 434883 706000 434912
rect 702392 434827 705525 434883
rect 705581 434827 705649 434883
rect 705705 434827 705773 434883
rect 705829 434827 705897 434883
rect 705953 434827 706000 434883
rect 702392 434826 706000 434827
rect 702392 434770 702440 434826
rect 702496 434770 702582 434826
rect 702638 434770 702724 434826
rect 702780 434770 702866 434826
rect 702922 434770 703008 434826
rect 703064 434770 703150 434826
rect 703206 434770 703292 434826
rect 703348 434770 703434 434826
rect 703490 434770 703576 434826
rect 703632 434770 703718 434826
rect 703774 434770 703860 434826
rect 703916 434770 704002 434826
rect 704058 434770 704144 434826
rect 704200 434770 704286 434826
rect 704342 434770 706000 434826
rect 702392 434759 706000 434770
rect 702392 434703 705525 434759
rect 705581 434703 705649 434759
rect 705705 434703 705773 434759
rect 705829 434703 705897 434759
rect 705953 434703 706000 434759
rect 702392 434684 706000 434703
rect 702392 434628 702440 434684
rect 702496 434628 702582 434684
rect 702638 434628 702724 434684
rect 702780 434628 702866 434684
rect 702922 434628 703008 434684
rect 703064 434628 703150 434684
rect 703206 434628 703292 434684
rect 703348 434628 703434 434684
rect 703490 434628 703576 434684
rect 703632 434628 703718 434684
rect 703774 434628 703860 434684
rect 703916 434628 704002 434684
rect 704058 434628 704144 434684
rect 704200 434628 704286 434684
rect 704342 434635 706000 434684
rect 704342 434628 705525 434635
rect 702392 434579 705525 434628
rect 705581 434579 705649 434635
rect 705705 434579 705773 434635
rect 705829 434579 705897 434635
rect 705953 434579 706000 434635
rect 702392 434542 706000 434579
rect 702392 434486 702440 434542
rect 702496 434486 702582 434542
rect 702638 434486 702724 434542
rect 702780 434486 702866 434542
rect 702922 434486 703008 434542
rect 703064 434486 703150 434542
rect 703206 434486 703292 434542
rect 703348 434486 703434 434542
rect 703490 434486 703576 434542
rect 703632 434486 703718 434542
rect 703774 434486 703860 434542
rect 703916 434486 704002 434542
rect 704058 434486 704144 434542
rect 704200 434486 704286 434542
rect 704342 434511 706000 434542
rect 704342 434486 705525 434511
rect 702392 434455 705525 434486
rect 705581 434455 705649 434511
rect 705705 434455 705773 434511
rect 705829 434455 705897 434511
rect 705953 434455 706000 434511
rect 702392 434400 706000 434455
rect 702392 434344 702440 434400
rect 702496 434344 702582 434400
rect 702638 434344 702724 434400
rect 702780 434344 702866 434400
rect 702922 434344 703008 434400
rect 703064 434344 703150 434400
rect 703206 434344 703292 434400
rect 703348 434344 703434 434400
rect 703490 434344 703576 434400
rect 703632 434344 703718 434400
rect 703774 434344 703860 434400
rect 703916 434344 704002 434400
rect 704058 434344 704144 434400
rect 704200 434344 704286 434400
rect 704342 434387 706000 434400
rect 704342 434344 705525 434387
rect 702392 434331 705525 434344
rect 705581 434331 705649 434387
rect 705705 434331 705773 434387
rect 705829 434331 705897 434387
rect 705953 434331 706000 434387
rect 702392 434263 706000 434331
rect 702392 434258 705525 434263
rect 702392 434202 702440 434258
rect 702496 434202 702582 434258
rect 702638 434202 702724 434258
rect 702780 434202 702866 434258
rect 702922 434202 703008 434258
rect 703064 434202 703150 434258
rect 703206 434202 703292 434258
rect 703348 434202 703434 434258
rect 703490 434202 703576 434258
rect 703632 434202 703718 434258
rect 703774 434202 703860 434258
rect 703916 434202 704002 434258
rect 704058 434202 704144 434258
rect 704200 434202 704286 434258
rect 704342 434207 705525 434258
rect 705581 434207 705649 434263
rect 705705 434207 705773 434263
rect 705829 434207 705897 434263
rect 705953 434207 706000 434263
rect 704342 434202 706000 434207
rect 702392 434139 706000 434202
rect 702392 434116 705525 434139
rect 702392 434060 702440 434116
rect 702496 434060 702582 434116
rect 702638 434060 702724 434116
rect 702780 434060 702866 434116
rect 702922 434060 703008 434116
rect 703064 434060 703150 434116
rect 703206 434060 703292 434116
rect 703348 434060 703434 434116
rect 703490 434060 703576 434116
rect 703632 434060 703718 434116
rect 703774 434060 703860 434116
rect 703916 434060 704002 434116
rect 704058 434060 704144 434116
rect 704200 434060 704286 434116
rect 704342 434083 705525 434116
rect 705581 434083 705649 434139
rect 705705 434083 705773 434139
rect 705829 434083 705897 434139
rect 705953 434083 706000 434139
rect 704342 434060 706000 434083
rect 702392 434015 706000 434060
rect 702392 433974 705525 434015
rect 702392 433918 702440 433974
rect 702496 433918 702582 433974
rect 702638 433918 702724 433974
rect 702780 433918 702866 433974
rect 702922 433918 703008 433974
rect 703064 433918 703150 433974
rect 703206 433918 703292 433974
rect 703348 433918 703434 433974
rect 703490 433918 703576 433974
rect 703632 433918 703718 433974
rect 703774 433918 703860 433974
rect 703916 433918 704002 433974
rect 704058 433918 704144 433974
rect 704200 433918 704286 433974
rect 704342 433959 705525 433974
rect 705581 433959 705649 434015
rect 705705 433959 705773 434015
rect 705829 433959 705897 434015
rect 705953 433959 706000 434015
rect 704342 433918 706000 433959
rect 702392 433891 706000 433918
rect 702392 433835 705525 433891
rect 705581 433835 705649 433891
rect 705705 433835 705773 433891
rect 705829 433835 705897 433891
rect 705953 433835 706000 433891
rect 702392 433832 706000 433835
rect 702392 433776 702440 433832
rect 702496 433776 702582 433832
rect 702638 433776 702724 433832
rect 702780 433776 702866 433832
rect 702922 433776 703008 433832
rect 703064 433776 703150 433832
rect 703206 433776 703292 433832
rect 703348 433776 703434 433832
rect 703490 433776 703576 433832
rect 703632 433776 703718 433832
rect 703774 433776 703860 433832
rect 703916 433776 704002 433832
rect 704058 433776 704144 433832
rect 704200 433776 704286 433832
rect 704342 433776 706000 433832
rect 702392 433767 706000 433776
rect 702392 433711 705525 433767
rect 705581 433711 705649 433767
rect 705705 433711 705773 433767
rect 705829 433711 705897 433767
rect 705953 433711 706000 433767
rect 702392 433690 706000 433711
rect 702392 433634 702440 433690
rect 702496 433634 702582 433690
rect 702638 433634 702724 433690
rect 702780 433634 702866 433690
rect 702922 433634 703008 433690
rect 703064 433634 703150 433690
rect 703206 433634 703292 433690
rect 703348 433634 703434 433690
rect 703490 433634 703576 433690
rect 703632 433634 703718 433690
rect 703774 433634 703860 433690
rect 703916 433634 704002 433690
rect 704058 433634 704144 433690
rect 704200 433634 704286 433690
rect 704342 433643 706000 433690
rect 704342 433634 705525 433643
rect 702392 433587 705525 433634
rect 705581 433587 705649 433643
rect 705705 433587 705773 433643
rect 705829 433587 705897 433643
rect 705953 433587 706000 433643
rect 702392 433548 706000 433587
rect 702392 433492 702440 433548
rect 702496 433492 702582 433548
rect 702638 433492 702724 433548
rect 702780 433492 702866 433548
rect 702922 433492 703008 433548
rect 703064 433492 703150 433548
rect 703206 433492 703292 433548
rect 703348 433492 703434 433548
rect 703490 433492 703576 433548
rect 703632 433492 703718 433548
rect 703774 433492 703860 433548
rect 703916 433492 704002 433548
rect 704058 433492 704144 433548
rect 704200 433492 704286 433548
rect 704342 433519 706000 433548
rect 704342 433492 705525 433519
rect 702392 433463 705525 433492
rect 705581 433463 705649 433519
rect 705705 433463 705773 433519
rect 705829 433463 705897 433519
rect 705953 433463 706000 433519
rect 702392 433406 706000 433463
rect 702392 433350 702440 433406
rect 702496 433350 702582 433406
rect 702638 433350 702724 433406
rect 702780 433350 702866 433406
rect 702922 433350 703008 433406
rect 703064 433350 703150 433406
rect 703206 433350 703292 433406
rect 703348 433350 703434 433406
rect 703490 433350 703576 433406
rect 703632 433350 703718 433406
rect 703774 433350 703860 433406
rect 703916 433350 704002 433406
rect 704058 433350 704144 433406
rect 704200 433350 704286 433406
rect 704342 433395 706000 433406
rect 704342 433350 705525 433395
rect 702392 433339 705525 433350
rect 705581 433339 705649 433395
rect 705705 433339 705773 433395
rect 705829 433339 705897 433395
rect 705953 433339 706000 433395
rect 702392 433272 706000 433339
rect 70000 427661 73416 427728
rect 70000 427605 70047 427661
rect 70103 427605 70171 427661
rect 70227 427605 70295 427661
rect 70351 427605 70419 427661
rect 70475 427650 73416 427661
rect 70475 427605 71466 427650
rect 70000 427594 71466 427605
rect 71522 427594 71608 427650
rect 71664 427594 71750 427650
rect 71806 427594 71892 427650
rect 71948 427594 72034 427650
rect 72090 427594 72176 427650
rect 72232 427594 72318 427650
rect 72374 427594 72460 427650
rect 72516 427594 72602 427650
rect 72658 427594 72744 427650
rect 72800 427594 72886 427650
rect 72942 427594 73028 427650
rect 73084 427594 73170 427650
rect 73226 427594 73312 427650
rect 73368 427594 73416 427650
rect 70000 427537 73416 427594
rect 70000 427481 70047 427537
rect 70103 427481 70171 427537
rect 70227 427481 70295 427537
rect 70351 427481 70419 427537
rect 70475 427508 73416 427537
rect 70475 427481 71466 427508
rect 70000 427452 71466 427481
rect 71522 427452 71608 427508
rect 71664 427452 71750 427508
rect 71806 427452 71892 427508
rect 71948 427452 72034 427508
rect 72090 427452 72176 427508
rect 72232 427452 72318 427508
rect 72374 427452 72460 427508
rect 72516 427452 72602 427508
rect 72658 427452 72744 427508
rect 72800 427452 72886 427508
rect 72942 427452 73028 427508
rect 73084 427452 73170 427508
rect 73226 427452 73312 427508
rect 73368 427452 73416 427508
rect 70000 427413 73416 427452
rect 70000 427357 70047 427413
rect 70103 427357 70171 427413
rect 70227 427357 70295 427413
rect 70351 427357 70419 427413
rect 70475 427366 73416 427413
rect 70475 427357 71466 427366
rect 70000 427310 71466 427357
rect 71522 427310 71608 427366
rect 71664 427310 71750 427366
rect 71806 427310 71892 427366
rect 71948 427310 72034 427366
rect 72090 427310 72176 427366
rect 72232 427310 72318 427366
rect 72374 427310 72460 427366
rect 72516 427310 72602 427366
rect 72658 427310 72744 427366
rect 72800 427310 72886 427366
rect 72942 427310 73028 427366
rect 73084 427310 73170 427366
rect 73226 427310 73312 427366
rect 73368 427310 73416 427366
rect 70000 427289 73416 427310
rect 70000 427233 70047 427289
rect 70103 427233 70171 427289
rect 70227 427233 70295 427289
rect 70351 427233 70419 427289
rect 70475 427233 73416 427289
rect 70000 427224 73416 427233
rect 70000 427168 71466 427224
rect 71522 427168 71608 427224
rect 71664 427168 71750 427224
rect 71806 427168 71892 427224
rect 71948 427168 72034 427224
rect 72090 427168 72176 427224
rect 72232 427168 72318 427224
rect 72374 427168 72460 427224
rect 72516 427168 72602 427224
rect 72658 427168 72744 427224
rect 72800 427168 72886 427224
rect 72942 427168 73028 427224
rect 73084 427168 73170 427224
rect 73226 427168 73312 427224
rect 73368 427168 73416 427224
rect 70000 427165 73416 427168
rect 70000 427109 70047 427165
rect 70103 427109 70171 427165
rect 70227 427109 70295 427165
rect 70351 427109 70419 427165
rect 70475 427109 73416 427165
rect 70000 427082 73416 427109
rect 70000 427041 71466 427082
rect 70000 426985 70047 427041
rect 70103 426985 70171 427041
rect 70227 426985 70295 427041
rect 70351 426985 70419 427041
rect 70475 427026 71466 427041
rect 71522 427026 71608 427082
rect 71664 427026 71750 427082
rect 71806 427026 71892 427082
rect 71948 427026 72034 427082
rect 72090 427026 72176 427082
rect 72232 427026 72318 427082
rect 72374 427026 72460 427082
rect 72516 427026 72602 427082
rect 72658 427026 72744 427082
rect 72800 427026 72886 427082
rect 72942 427026 73028 427082
rect 73084 427026 73170 427082
rect 73226 427026 73312 427082
rect 73368 427026 73416 427082
rect 70475 426985 73416 427026
rect 70000 426940 73416 426985
rect 70000 426917 71466 426940
rect 70000 426861 70047 426917
rect 70103 426861 70171 426917
rect 70227 426861 70295 426917
rect 70351 426861 70419 426917
rect 70475 426884 71466 426917
rect 71522 426884 71608 426940
rect 71664 426884 71750 426940
rect 71806 426884 71892 426940
rect 71948 426884 72034 426940
rect 72090 426884 72176 426940
rect 72232 426884 72318 426940
rect 72374 426884 72460 426940
rect 72516 426884 72602 426940
rect 72658 426884 72744 426940
rect 72800 426884 72886 426940
rect 72942 426884 73028 426940
rect 73084 426884 73170 426940
rect 73226 426884 73312 426940
rect 73368 426884 73416 426940
rect 70475 426861 73416 426884
rect 70000 426798 73416 426861
rect 70000 426793 71466 426798
rect 70000 426737 70047 426793
rect 70103 426737 70171 426793
rect 70227 426737 70295 426793
rect 70351 426737 70419 426793
rect 70475 426742 71466 426793
rect 71522 426742 71608 426798
rect 71664 426742 71750 426798
rect 71806 426742 71892 426798
rect 71948 426742 72034 426798
rect 72090 426742 72176 426798
rect 72232 426742 72318 426798
rect 72374 426742 72460 426798
rect 72516 426742 72602 426798
rect 72658 426742 72744 426798
rect 72800 426742 72886 426798
rect 72942 426742 73028 426798
rect 73084 426742 73170 426798
rect 73226 426742 73312 426798
rect 73368 426742 73416 426798
rect 70475 426737 73416 426742
rect 70000 426669 73416 426737
rect 70000 426613 70047 426669
rect 70103 426613 70171 426669
rect 70227 426613 70295 426669
rect 70351 426613 70419 426669
rect 70475 426656 73416 426669
rect 70475 426613 71466 426656
rect 70000 426600 71466 426613
rect 71522 426600 71608 426656
rect 71664 426600 71750 426656
rect 71806 426600 71892 426656
rect 71948 426600 72034 426656
rect 72090 426600 72176 426656
rect 72232 426600 72318 426656
rect 72374 426600 72460 426656
rect 72516 426600 72602 426656
rect 72658 426600 72744 426656
rect 72800 426600 72886 426656
rect 72942 426600 73028 426656
rect 73084 426600 73170 426656
rect 73226 426600 73312 426656
rect 73368 426600 73416 426656
rect 70000 426545 73416 426600
rect 70000 426489 70047 426545
rect 70103 426489 70171 426545
rect 70227 426489 70295 426545
rect 70351 426489 70419 426545
rect 70475 426514 73416 426545
rect 70475 426489 71466 426514
rect 70000 426458 71466 426489
rect 71522 426458 71608 426514
rect 71664 426458 71750 426514
rect 71806 426458 71892 426514
rect 71948 426458 72034 426514
rect 72090 426458 72176 426514
rect 72232 426458 72318 426514
rect 72374 426458 72460 426514
rect 72516 426458 72602 426514
rect 72658 426458 72744 426514
rect 72800 426458 72886 426514
rect 72942 426458 73028 426514
rect 73084 426458 73170 426514
rect 73226 426458 73312 426514
rect 73368 426458 73416 426514
rect 70000 426421 73416 426458
rect 70000 426365 70047 426421
rect 70103 426365 70171 426421
rect 70227 426365 70295 426421
rect 70351 426365 70419 426421
rect 70475 426372 73416 426421
rect 70475 426365 71466 426372
rect 70000 426316 71466 426365
rect 71522 426316 71608 426372
rect 71664 426316 71750 426372
rect 71806 426316 71892 426372
rect 71948 426316 72034 426372
rect 72090 426316 72176 426372
rect 72232 426316 72318 426372
rect 72374 426316 72460 426372
rect 72516 426316 72602 426372
rect 72658 426316 72744 426372
rect 72800 426316 72886 426372
rect 72942 426316 73028 426372
rect 73084 426316 73170 426372
rect 73226 426316 73312 426372
rect 73368 426316 73416 426372
rect 70000 426297 73416 426316
rect 70000 426241 70047 426297
rect 70103 426241 70171 426297
rect 70227 426241 70295 426297
rect 70351 426241 70419 426297
rect 70475 426241 73416 426297
rect 70000 426230 73416 426241
rect 70000 426174 71466 426230
rect 71522 426174 71608 426230
rect 71664 426174 71750 426230
rect 71806 426174 71892 426230
rect 71948 426174 72034 426230
rect 72090 426174 72176 426230
rect 72232 426174 72318 426230
rect 72374 426174 72460 426230
rect 72516 426174 72602 426230
rect 72658 426174 72744 426230
rect 72800 426174 72886 426230
rect 72942 426174 73028 426230
rect 73084 426174 73170 426230
rect 73226 426174 73312 426230
rect 73368 426174 73416 426230
rect 70000 426173 73416 426174
rect 70000 426117 70047 426173
rect 70103 426117 70171 426173
rect 70227 426117 70295 426173
rect 70351 426117 70419 426173
rect 70475 426117 73416 426173
rect 70000 426088 73416 426117
rect 70000 426049 71466 426088
rect 70000 425993 70047 426049
rect 70103 425993 70171 426049
rect 70227 425993 70295 426049
rect 70351 425993 70419 426049
rect 70475 426032 71466 426049
rect 71522 426032 71608 426088
rect 71664 426032 71750 426088
rect 71806 426032 71892 426088
rect 71948 426032 72034 426088
rect 72090 426032 72176 426088
rect 72232 426032 72318 426088
rect 72374 426032 72460 426088
rect 72516 426032 72602 426088
rect 72658 426032 72744 426088
rect 72800 426032 72886 426088
rect 72942 426032 73028 426088
rect 73084 426032 73170 426088
rect 73226 426032 73312 426088
rect 73368 426032 73416 426088
rect 70475 425993 73416 426032
rect 70000 425946 73416 425993
rect 70000 425925 71466 425946
rect 70000 425869 70047 425925
rect 70103 425869 70171 425925
rect 70227 425869 70295 425925
rect 70351 425869 70419 425925
rect 70475 425890 71466 425925
rect 71522 425890 71608 425946
rect 71664 425890 71750 425946
rect 71806 425890 71892 425946
rect 71948 425890 72034 425946
rect 72090 425890 72176 425946
rect 72232 425890 72318 425946
rect 72374 425890 72460 425946
rect 72516 425890 72602 425946
rect 72658 425890 72744 425946
rect 72800 425890 72886 425946
rect 72942 425890 73028 425946
rect 73084 425890 73170 425946
rect 73226 425890 73312 425946
rect 73368 425890 73416 425946
rect 70475 425869 73416 425890
rect 70000 425828 73416 425869
rect 70000 425181 73416 425248
rect 70000 425125 70047 425181
rect 70103 425125 70171 425181
rect 70227 425125 70295 425181
rect 70351 425125 70419 425181
rect 70475 425169 73416 425181
rect 70475 425125 71455 425169
rect 70000 425113 71455 425125
rect 71511 425113 71597 425169
rect 71653 425113 71739 425169
rect 71795 425113 71881 425169
rect 71937 425113 72023 425169
rect 72079 425113 72165 425169
rect 72221 425113 72307 425169
rect 72363 425113 72449 425169
rect 72505 425113 72591 425169
rect 72647 425113 72733 425169
rect 72789 425113 72875 425169
rect 72931 425113 73017 425169
rect 73073 425113 73159 425169
rect 73215 425113 73301 425169
rect 73357 425113 73416 425169
rect 70000 425057 73416 425113
rect 70000 425001 70047 425057
rect 70103 425001 70171 425057
rect 70227 425001 70295 425057
rect 70351 425001 70419 425057
rect 70475 425027 73416 425057
rect 70475 425001 71455 425027
rect 70000 424971 71455 425001
rect 71511 424971 71597 425027
rect 71653 424971 71739 425027
rect 71795 424971 71881 425027
rect 71937 424971 72023 425027
rect 72079 424971 72165 425027
rect 72221 424971 72307 425027
rect 72363 424971 72449 425027
rect 72505 424971 72591 425027
rect 72647 424971 72733 425027
rect 72789 424971 72875 425027
rect 72931 424971 73017 425027
rect 73073 424971 73159 425027
rect 73215 424971 73301 425027
rect 73357 424971 73416 425027
rect 70000 424933 73416 424971
rect 70000 424877 70047 424933
rect 70103 424877 70171 424933
rect 70227 424877 70295 424933
rect 70351 424877 70419 424933
rect 70475 424885 73416 424933
rect 70475 424877 71455 424885
rect 70000 424829 71455 424877
rect 71511 424829 71597 424885
rect 71653 424829 71739 424885
rect 71795 424829 71881 424885
rect 71937 424829 72023 424885
rect 72079 424829 72165 424885
rect 72221 424829 72307 424885
rect 72363 424829 72449 424885
rect 72505 424829 72591 424885
rect 72647 424829 72733 424885
rect 72789 424829 72875 424885
rect 72931 424829 73017 424885
rect 73073 424829 73159 424885
rect 73215 424829 73301 424885
rect 73357 424829 73416 424885
rect 70000 424809 73416 424829
rect 70000 424753 70047 424809
rect 70103 424753 70171 424809
rect 70227 424753 70295 424809
rect 70351 424753 70419 424809
rect 70475 424753 73416 424809
rect 70000 424743 73416 424753
rect 70000 424687 71455 424743
rect 71511 424687 71597 424743
rect 71653 424687 71739 424743
rect 71795 424687 71881 424743
rect 71937 424687 72023 424743
rect 72079 424687 72165 424743
rect 72221 424687 72307 424743
rect 72363 424687 72449 424743
rect 72505 424687 72591 424743
rect 72647 424687 72733 424743
rect 72789 424687 72875 424743
rect 72931 424687 73017 424743
rect 73073 424687 73159 424743
rect 73215 424687 73301 424743
rect 73357 424687 73416 424743
rect 70000 424685 73416 424687
rect 70000 424629 70047 424685
rect 70103 424629 70171 424685
rect 70227 424629 70295 424685
rect 70351 424629 70419 424685
rect 70475 424629 73416 424685
rect 70000 424601 73416 424629
rect 70000 424561 71455 424601
rect 70000 424505 70047 424561
rect 70103 424505 70171 424561
rect 70227 424505 70295 424561
rect 70351 424505 70419 424561
rect 70475 424545 71455 424561
rect 71511 424545 71597 424601
rect 71653 424545 71739 424601
rect 71795 424545 71881 424601
rect 71937 424545 72023 424601
rect 72079 424545 72165 424601
rect 72221 424545 72307 424601
rect 72363 424545 72449 424601
rect 72505 424545 72591 424601
rect 72647 424545 72733 424601
rect 72789 424545 72875 424601
rect 72931 424545 73017 424601
rect 73073 424545 73159 424601
rect 73215 424545 73301 424601
rect 73357 424545 73416 424601
rect 70475 424505 73416 424545
rect 70000 424459 73416 424505
rect 70000 424437 71455 424459
rect 70000 424381 70047 424437
rect 70103 424381 70171 424437
rect 70227 424381 70295 424437
rect 70351 424381 70419 424437
rect 70475 424403 71455 424437
rect 71511 424403 71597 424459
rect 71653 424403 71739 424459
rect 71795 424403 71881 424459
rect 71937 424403 72023 424459
rect 72079 424403 72165 424459
rect 72221 424403 72307 424459
rect 72363 424403 72449 424459
rect 72505 424403 72591 424459
rect 72647 424403 72733 424459
rect 72789 424403 72875 424459
rect 72931 424403 73017 424459
rect 73073 424403 73159 424459
rect 73215 424403 73301 424459
rect 73357 424403 73416 424459
rect 70475 424381 73416 424403
rect 70000 424317 73416 424381
rect 70000 424313 71455 424317
rect 70000 424257 70047 424313
rect 70103 424257 70171 424313
rect 70227 424257 70295 424313
rect 70351 424257 70419 424313
rect 70475 424261 71455 424313
rect 71511 424261 71597 424317
rect 71653 424261 71739 424317
rect 71795 424261 71881 424317
rect 71937 424261 72023 424317
rect 72079 424261 72165 424317
rect 72221 424261 72307 424317
rect 72363 424261 72449 424317
rect 72505 424261 72591 424317
rect 72647 424261 72733 424317
rect 72789 424261 72875 424317
rect 72931 424261 73017 424317
rect 73073 424261 73159 424317
rect 73215 424261 73301 424317
rect 73357 424261 73416 424317
rect 70475 424257 73416 424261
rect 70000 424189 73416 424257
rect 70000 424133 70047 424189
rect 70103 424133 70171 424189
rect 70227 424133 70295 424189
rect 70351 424133 70419 424189
rect 70475 424175 73416 424189
rect 70475 424133 71455 424175
rect 70000 424119 71455 424133
rect 71511 424119 71597 424175
rect 71653 424119 71739 424175
rect 71795 424119 71881 424175
rect 71937 424119 72023 424175
rect 72079 424119 72165 424175
rect 72221 424119 72307 424175
rect 72363 424119 72449 424175
rect 72505 424119 72591 424175
rect 72647 424119 72733 424175
rect 72789 424119 72875 424175
rect 72931 424119 73017 424175
rect 73073 424119 73159 424175
rect 73215 424119 73301 424175
rect 73357 424119 73416 424175
rect 70000 424065 73416 424119
rect 70000 424009 70047 424065
rect 70103 424009 70171 424065
rect 70227 424009 70295 424065
rect 70351 424009 70419 424065
rect 70475 424033 73416 424065
rect 70475 424009 71455 424033
rect 70000 423977 71455 424009
rect 71511 423977 71597 424033
rect 71653 423977 71739 424033
rect 71795 423977 71881 424033
rect 71937 423977 72023 424033
rect 72079 423977 72165 424033
rect 72221 423977 72307 424033
rect 72363 423977 72449 424033
rect 72505 423977 72591 424033
rect 72647 423977 72733 424033
rect 72789 423977 72875 424033
rect 72931 423977 73017 424033
rect 73073 423977 73159 424033
rect 73215 423977 73301 424033
rect 73357 423977 73416 424033
rect 70000 423941 73416 423977
rect 70000 423885 70047 423941
rect 70103 423885 70171 423941
rect 70227 423885 70295 423941
rect 70351 423885 70419 423941
rect 70475 423891 73416 423941
rect 70475 423885 71455 423891
rect 70000 423835 71455 423885
rect 71511 423835 71597 423891
rect 71653 423835 71739 423891
rect 71795 423835 71881 423891
rect 71937 423835 72023 423891
rect 72079 423835 72165 423891
rect 72221 423835 72307 423891
rect 72363 423835 72449 423891
rect 72505 423835 72591 423891
rect 72647 423835 72733 423891
rect 72789 423835 72875 423891
rect 72931 423835 73017 423891
rect 73073 423835 73159 423891
rect 73215 423835 73301 423891
rect 73357 423835 73416 423891
rect 70000 423817 73416 423835
rect 70000 423761 70047 423817
rect 70103 423761 70171 423817
rect 70227 423761 70295 423817
rect 70351 423761 70419 423817
rect 70475 423761 73416 423817
rect 70000 423749 73416 423761
rect 70000 423693 71455 423749
rect 71511 423693 71597 423749
rect 71653 423693 71739 423749
rect 71795 423693 71881 423749
rect 71937 423693 72023 423749
rect 72079 423693 72165 423749
rect 72221 423693 72307 423749
rect 72363 423693 72449 423749
rect 72505 423693 72591 423749
rect 72647 423693 72733 423749
rect 72789 423693 72875 423749
rect 72931 423693 73017 423749
rect 73073 423693 73159 423749
rect 73215 423693 73301 423749
rect 73357 423693 73416 423749
rect 70000 423637 70047 423693
rect 70103 423637 70171 423693
rect 70227 423637 70295 423693
rect 70351 423637 70419 423693
rect 70475 423637 73416 423693
rect 70000 423607 73416 423637
rect 70000 423569 71455 423607
rect 70000 423513 70047 423569
rect 70103 423513 70171 423569
rect 70227 423513 70295 423569
rect 70351 423513 70419 423569
rect 70475 423551 71455 423569
rect 71511 423551 71597 423607
rect 71653 423551 71739 423607
rect 71795 423551 71881 423607
rect 71937 423551 72023 423607
rect 72079 423551 72165 423607
rect 72221 423551 72307 423607
rect 72363 423551 72449 423607
rect 72505 423551 72591 423607
rect 72647 423551 72733 423607
rect 72789 423551 72875 423607
rect 72931 423551 73017 423607
rect 73073 423551 73159 423607
rect 73215 423551 73301 423607
rect 73357 423551 73416 423607
rect 70475 423513 73416 423551
rect 70000 423465 73416 423513
rect 70000 423445 71455 423465
rect 70000 423389 70047 423445
rect 70103 423389 70171 423445
rect 70227 423389 70295 423445
rect 70351 423389 70419 423445
rect 70475 423409 71455 423445
rect 71511 423409 71597 423465
rect 71653 423409 71739 423465
rect 71795 423409 71881 423465
rect 71937 423409 72023 423465
rect 72079 423409 72165 423465
rect 72221 423409 72307 423465
rect 72363 423409 72449 423465
rect 72505 423409 72591 423465
rect 72647 423409 72733 423465
rect 72789 423409 72875 423465
rect 72931 423409 73017 423465
rect 73073 423409 73159 423465
rect 73215 423409 73301 423465
rect 73357 423409 73416 423465
rect 70475 423389 73416 423409
rect 70000 423323 73416 423389
rect 70000 423321 71455 423323
rect 70000 423265 70047 423321
rect 70103 423265 70171 423321
rect 70227 423265 70295 423321
rect 70351 423265 70419 423321
rect 70475 423267 71455 423321
rect 71511 423267 71597 423323
rect 71653 423267 71739 423323
rect 71795 423267 71881 423323
rect 71937 423267 72023 423323
rect 72079 423267 72165 423323
rect 72221 423267 72307 423323
rect 72363 423267 72449 423323
rect 72505 423267 72591 423323
rect 72647 423267 72733 423323
rect 72789 423267 72875 423323
rect 72931 423267 73017 423323
rect 73073 423267 73159 423323
rect 73215 423267 73301 423323
rect 73357 423267 73416 423323
rect 70475 423265 73416 423267
rect 70000 423198 73416 423265
rect 70000 422811 73416 422878
rect 70000 422755 70047 422811
rect 70103 422755 70171 422811
rect 70227 422755 70295 422811
rect 70351 422755 70419 422811
rect 70475 422799 73416 422811
rect 70475 422755 71455 422799
rect 70000 422743 71455 422755
rect 71511 422743 71597 422799
rect 71653 422743 71739 422799
rect 71795 422743 71881 422799
rect 71937 422743 72023 422799
rect 72079 422743 72165 422799
rect 72221 422743 72307 422799
rect 72363 422743 72449 422799
rect 72505 422743 72591 422799
rect 72647 422743 72733 422799
rect 72789 422743 72875 422799
rect 72931 422743 73017 422799
rect 73073 422743 73159 422799
rect 73215 422743 73301 422799
rect 73357 422743 73416 422799
rect 70000 422687 73416 422743
rect 70000 422631 70047 422687
rect 70103 422631 70171 422687
rect 70227 422631 70295 422687
rect 70351 422631 70419 422687
rect 70475 422657 73416 422687
rect 70475 422631 71455 422657
rect 70000 422601 71455 422631
rect 71511 422601 71597 422657
rect 71653 422601 71739 422657
rect 71795 422601 71881 422657
rect 71937 422601 72023 422657
rect 72079 422601 72165 422657
rect 72221 422601 72307 422657
rect 72363 422601 72449 422657
rect 72505 422601 72591 422657
rect 72647 422601 72733 422657
rect 72789 422601 72875 422657
rect 72931 422601 73017 422657
rect 73073 422601 73159 422657
rect 73215 422601 73301 422657
rect 73357 422601 73416 422657
rect 70000 422563 73416 422601
rect 70000 422507 70047 422563
rect 70103 422507 70171 422563
rect 70227 422507 70295 422563
rect 70351 422507 70419 422563
rect 70475 422515 73416 422563
rect 70475 422507 71455 422515
rect 70000 422459 71455 422507
rect 71511 422459 71597 422515
rect 71653 422459 71739 422515
rect 71795 422459 71881 422515
rect 71937 422459 72023 422515
rect 72079 422459 72165 422515
rect 72221 422459 72307 422515
rect 72363 422459 72449 422515
rect 72505 422459 72591 422515
rect 72647 422459 72733 422515
rect 72789 422459 72875 422515
rect 72931 422459 73017 422515
rect 73073 422459 73159 422515
rect 73215 422459 73301 422515
rect 73357 422459 73416 422515
rect 70000 422439 73416 422459
rect 70000 422383 70047 422439
rect 70103 422383 70171 422439
rect 70227 422383 70295 422439
rect 70351 422383 70419 422439
rect 70475 422383 73416 422439
rect 70000 422373 73416 422383
rect 70000 422317 71455 422373
rect 71511 422317 71597 422373
rect 71653 422317 71739 422373
rect 71795 422317 71881 422373
rect 71937 422317 72023 422373
rect 72079 422317 72165 422373
rect 72221 422317 72307 422373
rect 72363 422317 72449 422373
rect 72505 422317 72591 422373
rect 72647 422317 72733 422373
rect 72789 422317 72875 422373
rect 72931 422317 73017 422373
rect 73073 422317 73159 422373
rect 73215 422317 73301 422373
rect 73357 422317 73416 422373
rect 70000 422315 73416 422317
rect 70000 422259 70047 422315
rect 70103 422259 70171 422315
rect 70227 422259 70295 422315
rect 70351 422259 70419 422315
rect 70475 422259 73416 422315
rect 70000 422231 73416 422259
rect 70000 422191 71455 422231
rect 70000 422135 70047 422191
rect 70103 422135 70171 422191
rect 70227 422135 70295 422191
rect 70351 422135 70419 422191
rect 70475 422175 71455 422191
rect 71511 422175 71597 422231
rect 71653 422175 71739 422231
rect 71795 422175 71881 422231
rect 71937 422175 72023 422231
rect 72079 422175 72165 422231
rect 72221 422175 72307 422231
rect 72363 422175 72449 422231
rect 72505 422175 72591 422231
rect 72647 422175 72733 422231
rect 72789 422175 72875 422231
rect 72931 422175 73017 422231
rect 73073 422175 73159 422231
rect 73215 422175 73301 422231
rect 73357 422175 73416 422231
rect 70475 422135 73416 422175
rect 70000 422089 73416 422135
rect 70000 422067 71455 422089
rect 70000 422011 70047 422067
rect 70103 422011 70171 422067
rect 70227 422011 70295 422067
rect 70351 422011 70419 422067
rect 70475 422033 71455 422067
rect 71511 422033 71597 422089
rect 71653 422033 71739 422089
rect 71795 422033 71881 422089
rect 71937 422033 72023 422089
rect 72079 422033 72165 422089
rect 72221 422033 72307 422089
rect 72363 422033 72449 422089
rect 72505 422033 72591 422089
rect 72647 422033 72733 422089
rect 72789 422033 72875 422089
rect 72931 422033 73017 422089
rect 73073 422033 73159 422089
rect 73215 422033 73301 422089
rect 73357 422033 73416 422089
rect 70475 422011 73416 422033
rect 70000 421947 73416 422011
rect 70000 421943 71455 421947
rect 70000 421887 70047 421943
rect 70103 421887 70171 421943
rect 70227 421887 70295 421943
rect 70351 421887 70419 421943
rect 70475 421891 71455 421943
rect 71511 421891 71597 421947
rect 71653 421891 71739 421947
rect 71795 421891 71881 421947
rect 71937 421891 72023 421947
rect 72079 421891 72165 421947
rect 72221 421891 72307 421947
rect 72363 421891 72449 421947
rect 72505 421891 72591 421947
rect 72647 421891 72733 421947
rect 72789 421891 72875 421947
rect 72931 421891 73017 421947
rect 73073 421891 73159 421947
rect 73215 421891 73301 421947
rect 73357 421891 73416 421947
rect 70475 421887 73416 421891
rect 70000 421819 73416 421887
rect 70000 421763 70047 421819
rect 70103 421763 70171 421819
rect 70227 421763 70295 421819
rect 70351 421763 70419 421819
rect 70475 421805 73416 421819
rect 70475 421763 71455 421805
rect 70000 421749 71455 421763
rect 71511 421749 71597 421805
rect 71653 421749 71739 421805
rect 71795 421749 71881 421805
rect 71937 421749 72023 421805
rect 72079 421749 72165 421805
rect 72221 421749 72307 421805
rect 72363 421749 72449 421805
rect 72505 421749 72591 421805
rect 72647 421749 72733 421805
rect 72789 421749 72875 421805
rect 72931 421749 73017 421805
rect 73073 421749 73159 421805
rect 73215 421749 73301 421805
rect 73357 421749 73416 421805
rect 70000 421695 73416 421749
rect 70000 421639 70047 421695
rect 70103 421639 70171 421695
rect 70227 421639 70295 421695
rect 70351 421639 70419 421695
rect 70475 421663 73416 421695
rect 70475 421639 71455 421663
rect 70000 421607 71455 421639
rect 71511 421607 71597 421663
rect 71653 421607 71739 421663
rect 71795 421607 71881 421663
rect 71937 421607 72023 421663
rect 72079 421607 72165 421663
rect 72221 421607 72307 421663
rect 72363 421607 72449 421663
rect 72505 421607 72591 421663
rect 72647 421607 72733 421663
rect 72789 421607 72875 421663
rect 72931 421607 73017 421663
rect 73073 421607 73159 421663
rect 73215 421607 73301 421663
rect 73357 421607 73416 421663
rect 70000 421571 73416 421607
rect 70000 421515 70047 421571
rect 70103 421515 70171 421571
rect 70227 421515 70295 421571
rect 70351 421515 70419 421571
rect 70475 421521 73416 421571
rect 70475 421515 71455 421521
rect 70000 421465 71455 421515
rect 71511 421465 71597 421521
rect 71653 421465 71739 421521
rect 71795 421465 71881 421521
rect 71937 421465 72023 421521
rect 72079 421465 72165 421521
rect 72221 421465 72307 421521
rect 72363 421465 72449 421521
rect 72505 421465 72591 421521
rect 72647 421465 72733 421521
rect 72789 421465 72875 421521
rect 72931 421465 73017 421521
rect 73073 421465 73159 421521
rect 73215 421465 73301 421521
rect 73357 421465 73416 421521
rect 70000 421447 73416 421465
rect 70000 421391 70047 421447
rect 70103 421391 70171 421447
rect 70227 421391 70295 421447
rect 70351 421391 70419 421447
rect 70475 421391 73416 421447
rect 70000 421379 73416 421391
rect 70000 421323 71455 421379
rect 71511 421323 71597 421379
rect 71653 421323 71739 421379
rect 71795 421323 71881 421379
rect 71937 421323 72023 421379
rect 72079 421323 72165 421379
rect 72221 421323 72307 421379
rect 72363 421323 72449 421379
rect 72505 421323 72591 421379
rect 72647 421323 72733 421379
rect 72789 421323 72875 421379
rect 72931 421323 73017 421379
rect 73073 421323 73159 421379
rect 73215 421323 73301 421379
rect 73357 421323 73416 421379
rect 70000 421267 70047 421323
rect 70103 421267 70171 421323
rect 70227 421267 70295 421323
rect 70351 421267 70419 421323
rect 70475 421267 73416 421323
rect 70000 421237 73416 421267
rect 70000 421199 71455 421237
rect 70000 421143 70047 421199
rect 70103 421143 70171 421199
rect 70227 421143 70295 421199
rect 70351 421143 70419 421199
rect 70475 421181 71455 421199
rect 71511 421181 71597 421237
rect 71653 421181 71739 421237
rect 71795 421181 71881 421237
rect 71937 421181 72023 421237
rect 72079 421181 72165 421237
rect 72221 421181 72307 421237
rect 72363 421181 72449 421237
rect 72505 421181 72591 421237
rect 72647 421181 72733 421237
rect 72789 421181 72875 421237
rect 72931 421181 73017 421237
rect 73073 421181 73159 421237
rect 73215 421181 73301 421237
rect 73357 421181 73416 421237
rect 70475 421143 73416 421181
rect 70000 421095 73416 421143
rect 70000 421075 71455 421095
rect 70000 421019 70047 421075
rect 70103 421019 70171 421075
rect 70227 421019 70295 421075
rect 70351 421019 70419 421075
rect 70475 421039 71455 421075
rect 71511 421039 71597 421095
rect 71653 421039 71739 421095
rect 71795 421039 71881 421095
rect 71937 421039 72023 421095
rect 72079 421039 72165 421095
rect 72221 421039 72307 421095
rect 72363 421039 72449 421095
rect 72505 421039 72591 421095
rect 72647 421039 72733 421095
rect 72789 421039 72875 421095
rect 72931 421039 73017 421095
rect 73073 421039 73159 421095
rect 73215 421039 73301 421095
rect 73357 421039 73416 421095
rect 70475 421019 73416 421039
rect 70000 420953 73416 421019
rect 70000 420951 71455 420953
rect 70000 420895 70047 420951
rect 70103 420895 70171 420951
rect 70227 420895 70295 420951
rect 70351 420895 70419 420951
rect 70475 420897 71455 420951
rect 71511 420897 71597 420953
rect 71653 420897 71739 420953
rect 71795 420897 71881 420953
rect 71937 420897 72023 420953
rect 72079 420897 72165 420953
rect 72221 420897 72307 420953
rect 72363 420897 72449 420953
rect 72505 420897 72591 420953
rect 72647 420897 72733 420953
rect 72789 420897 72875 420953
rect 72931 420897 73017 420953
rect 73073 420897 73159 420953
rect 73215 420897 73301 420953
rect 73357 420897 73416 420953
rect 70475 420895 73416 420897
rect 70000 420828 73416 420895
rect 70000 420105 73416 420172
rect 70000 420049 70047 420105
rect 70103 420049 70171 420105
rect 70227 420049 70295 420105
rect 70351 420049 70419 420105
rect 70475 420093 73416 420105
rect 70475 420049 71455 420093
rect 70000 420037 71455 420049
rect 71511 420037 71597 420093
rect 71653 420037 71739 420093
rect 71795 420037 71881 420093
rect 71937 420037 72023 420093
rect 72079 420037 72165 420093
rect 72221 420037 72307 420093
rect 72363 420037 72449 420093
rect 72505 420037 72591 420093
rect 72647 420037 72733 420093
rect 72789 420037 72875 420093
rect 72931 420037 73017 420093
rect 73073 420037 73159 420093
rect 73215 420037 73301 420093
rect 73357 420037 73416 420093
rect 70000 419981 73416 420037
rect 70000 419925 70047 419981
rect 70103 419925 70171 419981
rect 70227 419925 70295 419981
rect 70351 419925 70419 419981
rect 70475 419951 73416 419981
rect 70475 419925 71455 419951
rect 70000 419895 71455 419925
rect 71511 419895 71597 419951
rect 71653 419895 71739 419951
rect 71795 419895 71881 419951
rect 71937 419895 72023 419951
rect 72079 419895 72165 419951
rect 72221 419895 72307 419951
rect 72363 419895 72449 419951
rect 72505 419895 72591 419951
rect 72647 419895 72733 419951
rect 72789 419895 72875 419951
rect 72931 419895 73017 419951
rect 73073 419895 73159 419951
rect 73215 419895 73301 419951
rect 73357 419895 73416 419951
rect 70000 419857 73416 419895
rect 70000 419801 70047 419857
rect 70103 419801 70171 419857
rect 70227 419801 70295 419857
rect 70351 419801 70419 419857
rect 70475 419809 73416 419857
rect 70475 419801 71455 419809
rect 70000 419753 71455 419801
rect 71511 419753 71597 419809
rect 71653 419753 71739 419809
rect 71795 419753 71881 419809
rect 71937 419753 72023 419809
rect 72079 419753 72165 419809
rect 72221 419753 72307 419809
rect 72363 419753 72449 419809
rect 72505 419753 72591 419809
rect 72647 419753 72733 419809
rect 72789 419753 72875 419809
rect 72931 419753 73017 419809
rect 73073 419753 73159 419809
rect 73215 419753 73301 419809
rect 73357 419753 73416 419809
rect 70000 419733 73416 419753
rect 70000 419677 70047 419733
rect 70103 419677 70171 419733
rect 70227 419677 70295 419733
rect 70351 419677 70419 419733
rect 70475 419677 73416 419733
rect 70000 419667 73416 419677
rect 70000 419611 71455 419667
rect 71511 419611 71597 419667
rect 71653 419611 71739 419667
rect 71795 419611 71881 419667
rect 71937 419611 72023 419667
rect 72079 419611 72165 419667
rect 72221 419611 72307 419667
rect 72363 419611 72449 419667
rect 72505 419611 72591 419667
rect 72647 419611 72733 419667
rect 72789 419611 72875 419667
rect 72931 419611 73017 419667
rect 73073 419611 73159 419667
rect 73215 419611 73301 419667
rect 73357 419611 73416 419667
rect 70000 419609 73416 419611
rect 70000 419553 70047 419609
rect 70103 419553 70171 419609
rect 70227 419553 70295 419609
rect 70351 419553 70419 419609
rect 70475 419553 73416 419609
rect 70000 419525 73416 419553
rect 70000 419485 71455 419525
rect 70000 419429 70047 419485
rect 70103 419429 70171 419485
rect 70227 419429 70295 419485
rect 70351 419429 70419 419485
rect 70475 419469 71455 419485
rect 71511 419469 71597 419525
rect 71653 419469 71739 419525
rect 71795 419469 71881 419525
rect 71937 419469 72023 419525
rect 72079 419469 72165 419525
rect 72221 419469 72307 419525
rect 72363 419469 72449 419525
rect 72505 419469 72591 419525
rect 72647 419469 72733 419525
rect 72789 419469 72875 419525
rect 72931 419469 73017 419525
rect 73073 419469 73159 419525
rect 73215 419469 73301 419525
rect 73357 419469 73416 419525
rect 70475 419429 73416 419469
rect 70000 419383 73416 419429
rect 70000 419361 71455 419383
rect 70000 419305 70047 419361
rect 70103 419305 70171 419361
rect 70227 419305 70295 419361
rect 70351 419305 70419 419361
rect 70475 419327 71455 419361
rect 71511 419327 71597 419383
rect 71653 419327 71739 419383
rect 71795 419327 71881 419383
rect 71937 419327 72023 419383
rect 72079 419327 72165 419383
rect 72221 419327 72307 419383
rect 72363 419327 72449 419383
rect 72505 419327 72591 419383
rect 72647 419327 72733 419383
rect 72789 419327 72875 419383
rect 72931 419327 73017 419383
rect 73073 419327 73159 419383
rect 73215 419327 73301 419383
rect 73357 419327 73416 419383
rect 70475 419305 73416 419327
rect 70000 419241 73416 419305
rect 70000 419237 71455 419241
rect 70000 419181 70047 419237
rect 70103 419181 70171 419237
rect 70227 419181 70295 419237
rect 70351 419181 70419 419237
rect 70475 419185 71455 419237
rect 71511 419185 71597 419241
rect 71653 419185 71739 419241
rect 71795 419185 71881 419241
rect 71937 419185 72023 419241
rect 72079 419185 72165 419241
rect 72221 419185 72307 419241
rect 72363 419185 72449 419241
rect 72505 419185 72591 419241
rect 72647 419185 72733 419241
rect 72789 419185 72875 419241
rect 72931 419185 73017 419241
rect 73073 419185 73159 419241
rect 73215 419185 73301 419241
rect 73357 419185 73416 419241
rect 70475 419181 73416 419185
rect 70000 419113 73416 419181
rect 70000 419057 70047 419113
rect 70103 419057 70171 419113
rect 70227 419057 70295 419113
rect 70351 419057 70419 419113
rect 70475 419099 73416 419113
rect 70475 419057 71455 419099
rect 70000 419043 71455 419057
rect 71511 419043 71597 419099
rect 71653 419043 71739 419099
rect 71795 419043 71881 419099
rect 71937 419043 72023 419099
rect 72079 419043 72165 419099
rect 72221 419043 72307 419099
rect 72363 419043 72449 419099
rect 72505 419043 72591 419099
rect 72647 419043 72733 419099
rect 72789 419043 72875 419099
rect 72931 419043 73017 419099
rect 73073 419043 73159 419099
rect 73215 419043 73301 419099
rect 73357 419043 73416 419099
rect 70000 418989 73416 419043
rect 70000 418933 70047 418989
rect 70103 418933 70171 418989
rect 70227 418933 70295 418989
rect 70351 418933 70419 418989
rect 70475 418957 73416 418989
rect 70475 418933 71455 418957
rect 70000 418901 71455 418933
rect 71511 418901 71597 418957
rect 71653 418901 71739 418957
rect 71795 418901 71881 418957
rect 71937 418901 72023 418957
rect 72079 418901 72165 418957
rect 72221 418901 72307 418957
rect 72363 418901 72449 418957
rect 72505 418901 72591 418957
rect 72647 418901 72733 418957
rect 72789 418901 72875 418957
rect 72931 418901 73017 418957
rect 73073 418901 73159 418957
rect 73215 418901 73301 418957
rect 73357 418901 73416 418957
rect 70000 418865 73416 418901
rect 70000 418809 70047 418865
rect 70103 418809 70171 418865
rect 70227 418809 70295 418865
rect 70351 418809 70419 418865
rect 70475 418815 73416 418865
rect 70475 418809 71455 418815
rect 70000 418759 71455 418809
rect 71511 418759 71597 418815
rect 71653 418759 71739 418815
rect 71795 418759 71881 418815
rect 71937 418759 72023 418815
rect 72079 418759 72165 418815
rect 72221 418759 72307 418815
rect 72363 418759 72449 418815
rect 72505 418759 72591 418815
rect 72647 418759 72733 418815
rect 72789 418759 72875 418815
rect 72931 418759 73017 418815
rect 73073 418759 73159 418815
rect 73215 418759 73301 418815
rect 73357 418759 73416 418815
rect 70000 418741 73416 418759
rect 70000 418685 70047 418741
rect 70103 418685 70171 418741
rect 70227 418685 70295 418741
rect 70351 418685 70419 418741
rect 70475 418685 73416 418741
rect 70000 418673 73416 418685
rect 70000 418617 71455 418673
rect 71511 418617 71597 418673
rect 71653 418617 71739 418673
rect 71795 418617 71881 418673
rect 71937 418617 72023 418673
rect 72079 418617 72165 418673
rect 72221 418617 72307 418673
rect 72363 418617 72449 418673
rect 72505 418617 72591 418673
rect 72647 418617 72733 418673
rect 72789 418617 72875 418673
rect 72931 418617 73017 418673
rect 73073 418617 73159 418673
rect 73215 418617 73301 418673
rect 73357 418617 73416 418673
rect 70000 418561 70047 418617
rect 70103 418561 70171 418617
rect 70227 418561 70295 418617
rect 70351 418561 70419 418617
rect 70475 418561 73416 418617
rect 70000 418531 73416 418561
rect 70000 418493 71455 418531
rect 70000 418437 70047 418493
rect 70103 418437 70171 418493
rect 70227 418437 70295 418493
rect 70351 418437 70419 418493
rect 70475 418475 71455 418493
rect 71511 418475 71597 418531
rect 71653 418475 71739 418531
rect 71795 418475 71881 418531
rect 71937 418475 72023 418531
rect 72079 418475 72165 418531
rect 72221 418475 72307 418531
rect 72363 418475 72449 418531
rect 72505 418475 72591 418531
rect 72647 418475 72733 418531
rect 72789 418475 72875 418531
rect 72931 418475 73017 418531
rect 73073 418475 73159 418531
rect 73215 418475 73301 418531
rect 73357 418475 73416 418531
rect 70475 418437 73416 418475
rect 70000 418389 73416 418437
rect 70000 418369 71455 418389
rect 70000 418313 70047 418369
rect 70103 418313 70171 418369
rect 70227 418313 70295 418369
rect 70351 418313 70419 418369
rect 70475 418333 71455 418369
rect 71511 418333 71597 418389
rect 71653 418333 71739 418389
rect 71795 418333 71881 418389
rect 71937 418333 72023 418389
rect 72079 418333 72165 418389
rect 72221 418333 72307 418389
rect 72363 418333 72449 418389
rect 72505 418333 72591 418389
rect 72647 418333 72733 418389
rect 72789 418333 72875 418389
rect 72931 418333 73017 418389
rect 73073 418333 73159 418389
rect 73215 418333 73301 418389
rect 73357 418333 73416 418389
rect 70475 418313 73416 418333
rect 70000 418247 73416 418313
rect 70000 418245 71455 418247
rect 70000 418189 70047 418245
rect 70103 418189 70171 418245
rect 70227 418189 70295 418245
rect 70351 418189 70419 418245
rect 70475 418191 71455 418245
rect 71511 418191 71597 418247
rect 71653 418191 71739 418247
rect 71795 418191 71881 418247
rect 71937 418191 72023 418247
rect 72079 418191 72165 418247
rect 72221 418191 72307 418247
rect 72363 418191 72449 418247
rect 72505 418191 72591 418247
rect 72647 418191 72733 418247
rect 72789 418191 72875 418247
rect 72931 418191 73017 418247
rect 73073 418191 73159 418247
rect 73215 418191 73301 418247
rect 73357 418191 73416 418247
rect 70475 418189 73416 418191
rect 70000 418122 73416 418189
rect 70000 417735 73416 417802
rect 70000 417679 70047 417735
rect 70103 417679 70171 417735
rect 70227 417679 70295 417735
rect 70351 417679 70419 417735
rect 70475 417723 73416 417735
rect 70475 417679 71455 417723
rect 70000 417667 71455 417679
rect 71511 417667 71597 417723
rect 71653 417667 71739 417723
rect 71795 417667 71881 417723
rect 71937 417667 72023 417723
rect 72079 417667 72165 417723
rect 72221 417667 72307 417723
rect 72363 417667 72449 417723
rect 72505 417667 72591 417723
rect 72647 417667 72733 417723
rect 72789 417667 72875 417723
rect 72931 417667 73017 417723
rect 73073 417667 73159 417723
rect 73215 417667 73301 417723
rect 73357 417667 73416 417723
rect 70000 417611 73416 417667
rect 70000 417555 70047 417611
rect 70103 417555 70171 417611
rect 70227 417555 70295 417611
rect 70351 417555 70419 417611
rect 70475 417581 73416 417611
rect 70475 417555 71455 417581
rect 70000 417525 71455 417555
rect 71511 417525 71597 417581
rect 71653 417525 71739 417581
rect 71795 417525 71881 417581
rect 71937 417525 72023 417581
rect 72079 417525 72165 417581
rect 72221 417525 72307 417581
rect 72363 417525 72449 417581
rect 72505 417525 72591 417581
rect 72647 417525 72733 417581
rect 72789 417525 72875 417581
rect 72931 417525 73017 417581
rect 73073 417525 73159 417581
rect 73215 417525 73301 417581
rect 73357 417525 73416 417581
rect 70000 417487 73416 417525
rect 70000 417431 70047 417487
rect 70103 417431 70171 417487
rect 70227 417431 70295 417487
rect 70351 417431 70419 417487
rect 70475 417439 73416 417487
rect 70475 417431 71455 417439
rect 70000 417383 71455 417431
rect 71511 417383 71597 417439
rect 71653 417383 71739 417439
rect 71795 417383 71881 417439
rect 71937 417383 72023 417439
rect 72079 417383 72165 417439
rect 72221 417383 72307 417439
rect 72363 417383 72449 417439
rect 72505 417383 72591 417439
rect 72647 417383 72733 417439
rect 72789 417383 72875 417439
rect 72931 417383 73017 417439
rect 73073 417383 73159 417439
rect 73215 417383 73301 417439
rect 73357 417383 73416 417439
rect 70000 417363 73416 417383
rect 70000 417307 70047 417363
rect 70103 417307 70171 417363
rect 70227 417307 70295 417363
rect 70351 417307 70419 417363
rect 70475 417307 73416 417363
rect 70000 417297 73416 417307
rect 70000 417241 71455 417297
rect 71511 417241 71597 417297
rect 71653 417241 71739 417297
rect 71795 417241 71881 417297
rect 71937 417241 72023 417297
rect 72079 417241 72165 417297
rect 72221 417241 72307 417297
rect 72363 417241 72449 417297
rect 72505 417241 72591 417297
rect 72647 417241 72733 417297
rect 72789 417241 72875 417297
rect 72931 417241 73017 417297
rect 73073 417241 73159 417297
rect 73215 417241 73301 417297
rect 73357 417241 73416 417297
rect 70000 417239 73416 417241
rect 70000 417183 70047 417239
rect 70103 417183 70171 417239
rect 70227 417183 70295 417239
rect 70351 417183 70419 417239
rect 70475 417183 73416 417239
rect 70000 417155 73416 417183
rect 70000 417115 71455 417155
rect 70000 417059 70047 417115
rect 70103 417059 70171 417115
rect 70227 417059 70295 417115
rect 70351 417059 70419 417115
rect 70475 417099 71455 417115
rect 71511 417099 71597 417155
rect 71653 417099 71739 417155
rect 71795 417099 71881 417155
rect 71937 417099 72023 417155
rect 72079 417099 72165 417155
rect 72221 417099 72307 417155
rect 72363 417099 72449 417155
rect 72505 417099 72591 417155
rect 72647 417099 72733 417155
rect 72789 417099 72875 417155
rect 72931 417099 73017 417155
rect 73073 417099 73159 417155
rect 73215 417099 73301 417155
rect 73357 417099 73416 417155
rect 70475 417059 73416 417099
rect 70000 417013 73416 417059
rect 70000 416991 71455 417013
rect 70000 416935 70047 416991
rect 70103 416935 70171 416991
rect 70227 416935 70295 416991
rect 70351 416935 70419 416991
rect 70475 416957 71455 416991
rect 71511 416957 71597 417013
rect 71653 416957 71739 417013
rect 71795 416957 71881 417013
rect 71937 416957 72023 417013
rect 72079 416957 72165 417013
rect 72221 416957 72307 417013
rect 72363 416957 72449 417013
rect 72505 416957 72591 417013
rect 72647 416957 72733 417013
rect 72789 416957 72875 417013
rect 72931 416957 73017 417013
rect 73073 416957 73159 417013
rect 73215 416957 73301 417013
rect 73357 416957 73416 417013
rect 70475 416935 73416 416957
rect 70000 416871 73416 416935
rect 70000 416867 71455 416871
rect 70000 416811 70047 416867
rect 70103 416811 70171 416867
rect 70227 416811 70295 416867
rect 70351 416811 70419 416867
rect 70475 416815 71455 416867
rect 71511 416815 71597 416871
rect 71653 416815 71739 416871
rect 71795 416815 71881 416871
rect 71937 416815 72023 416871
rect 72079 416815 72165 416871
rect 72221 416815 72307 416871
rect 72363 416815 72449 416871
rect 72505 416815 72591 416871
rect 72647 416815 72733 416871
rect 72789 416815 72875 416871
rect 72931 416815 73017 416871
rect 73073 416815 73159 416871
rect 73215 416815 73301 416871
rect 73357 416815 73416 416871
rect 70475 416811 73416 416815
rect 70000 416743 73416 416811
rect 70000 416687 70047 416743
rect 70103 416687 70171 416743
rect 70227 416687 70295 416743
rect 70351 416687 70419 416743
rect 70475 416729 73416 416743
rect 70475 416687 71455 416729
rect 70000 416673 71455 416687
rect 71511 416673 71597 416729
rect 71653 416673 71739 416729
rect 71795 416673 71881 416729
rect 71937 416673 72023 416729
rect 72079 416673 72165 416729
rect 72221 416673 72307 416729
rect 72363 416673 72449 416729
rect 72505 416673 72591 416729
rect 72647 416673 72733 416729
rect 72789 416673 72875 416729
rect 72931 416673 73017 416729
rect 73073 416673 73159 416729
rect 73215 416673 73301 416729
rect 73357 416673 73416 416729
rect 70000 416619 73416 416673
rect 70000 416563 70047 416619
rect 70103 416563 70171 416619
rect 70227 416563 70295 416619
rect 70351 416563 70419 416619
rect 70475 416587 73416 416619
rect 70475 416563 71455 416587
rect 70000 416531 71455 416563
rect 71511 416531 71597 416587
rect 71653 416531 71739 416587
rect 71795 416531 71881 416587
rect 71937 416531 72023 416587
rect 72079 416531 72165 416587
rect 72221 416531 72307 416587
rect 72363 416531 72449 416587
rect 72505 416531 72591 416587
rect 72647 416531 72733 416587
rect 72789 416531 72875 416587
rect 72931 416531 73017 416587
rect 73073 416531 73159 416587
rect 73215 416531 73301 416587
rect 73357 416531 73416 416587
rect 70000 416495 73416 416531
rect 70000 416439 70047 416495
rect 70103 416439 70171 416495
rect 70227 416439 70295 416495
rect 70351 416439 70419 416495
rect 70475 416445 73416 416495
rect 70475 416439 71455 416445
rect 70000 416389 71455 416439
rect 71511 416389 71597 416445
rect 71653 416389 71739 416445
rect 71795 416389 71881 416445
rect 71937 416389 72023 416445
rect 72079 416389 72165 416445
rect 72221 416389 72307 416445
rect 72363 416389 72449 416445
rect 72505 416389 72591 416445
rect 72647 416389 72733 416445
rect 72789 416389 72875 416445
rect 72931 416389 73017 416445
rect 73073 416389 73159 416445
rect 73215 416389 73301 416445
rect 73357 416389 73416 416445
rect 70000 416371 73416 416389
rect 70000 416315 70047 416371
rect 70103 416315 70171 416371
rect 70227 416315 70295 416371
rect 70351 416315 70419 416371
rect 70475 416315 73416 416371
rect 70000 416303 73416 416315
rect 70000 416247 71455 416303
rect 71511 416247 71597 416303
rect 71653 416247 71739 416303
rect 71795 416247 71881 416303
rect 71937 416247 72023 416303
rect 72079 416247 72165 416303
rect 72221 416247 72307 416303
rect 72363 416247 72449 416303
rect 72505 416247 72591 416303
rect 72647 416247 72733 416303
rect 72789 416247 72875 416303
rect 72931 416247 73017 416303
rect 73073 416247 73159 416303
rect 73215 416247 73301 416303
rect 73357 416247 73416 416303
rect 70000 416191 70047 416247
rect 70103 416191 70171 416247
rect 70227 416191 70295 416247
rect 70351 416191 70419 416247
rect 70475 416191 73416 416247
rect 70000 416161 73416 416191
rect 70000 416123 71455 416161
rect 70000 416067 70047 416123
rect 70103 416067 70171 416123
rect 70227 416067 70295 416123
rect 70351 416067 70419 416123
rect 70475 416105 71455 416123
rect 71511 416105 71597 416161
rect 71653 416105 71739 416161
rect 71795 416105 71881 416161
rect 71937 416105 72023 416161
rect 72079 416105 72165 416161
rect 72221 416105 72307 416161
rect 72363 416105 72449 416161
rect 72505 416105 72591 416161
rect 72647 416105 72733 416161
rect 72789 416105 72875 416161
rect 72931 416105 73017 416161
rect 73073 416105 73159 416161
rect 73215 416105 73301 416161
rect 73357 416105 73416 416161
rect 70475 416067 73416 416105
rect 70000 416019 73416 416067
rect 70000 415999 71455 416019
rect 70000 415943 70047 415999
rect 70103 415943 70171 415999
rect 70227 415943 70295 415999
rect 70351 415943 70419 415999
rect 70475 415963 71455 415999
rect 71511 415963 71597 416019
rect 71653 415963 71739 416019
rect 71795 415963 71881 416019
rect 71937 415963 72023 416019
rect 72079 415963 72165 416019
rect 72221 415963 72307 416019
rect 72363 415963 72449 416019
rect 72505 415963 72591 416019
rect 72647 415963 72733 416019
rect 72789 415963 72875 416019
rect 72931 415963 73017 416019
rect 73073 415963 73159 416019
rect 73215 415963 73301 416019
rect 73357 415963 73416 416019
rect 70475 415943 73416 415963
rect 70000 415877 73416 415943
rect 70000 415875 71455 415877
rect 70000 415819 70047 415875
rect 70103 415819 70171 415875
rect 70227 415819 70295 415875
rect 70351 415819 70419 415875
rect 70475 415821 71455 415875
rect 71511 415821 71597 415877
rect 71653 415821 71739 415877
rect 71795 415821 71881 415877
rect 71937 415821 72023 415877
rect 72079 415821 72165 415877
rect 72221 415821 72307 415877
rect 72363 415821 72449 415877
rect 72505 415821 72591 415877
rect 72647 415821 72733 415877
rect 72789 415821 72875 415877
rect 72931 415821 73017 415877
rect 73073 415821 73159 415877
rect 73215 415821 73301 415877
rect 73357 415821 73416 415877
rect 70475 415819 73416 415821
rect 70000 415752 73416 415819
rect 70000 415105 73416 415172
rect 70000 415049 70047 415105
rect 70103 415049 70171 415105
rect 70227 415049 70295 415105
rect 70351 415049 70419 415105
rect 70475 415094 73416 415105
rect 70475 415049 71466 415094
rect 70000 415038 71466 415049
rect 71522 415038 71608 415094
rect 71664 415038 71750 415094
rect 71806 415038 71892 415094
rect 71948 415038 72034 415094
rect 72090 415038 72176 415094
rect 72232 415038 72318 415094
rect 72374 415038 72460 415094
rect 72516 415038 72602 415094
rect 72658 415038 72744 415094
rect 72800 415038 72886 415094
rect 72942 415038 73028 415094
rect 73084 415038 73170 415094
rect 73226 415038 73312 415094
rect 73368 415038 73416 415094
rect 70000 414981 73416 415038
rect 70000 414925 70047 414981
rect 70103 414925 70171 414981
rect 70227 414925 70295 414981
rect 70351 414925 70419 414981
rect 70475 414952 73416 414981
rect 70475 414925 71466 414952
rect 70000 414896 71466 414925
rect 71522 414896 71608 414952
rect 71664 414896 71750 414952
rect 71806 414896 71892 414952
rect 71948 414896 72034 414952
rect 72090 414896 72176 414952
rect 72232 414896 72318 414952
rect 72374 414896 72460 414952
rect 72516 414896 72602 414952
rect 72658 414896 72744 414952
rect 72800 414896 72886 414952
rect 72942 414896 73028 414952
rect 73084 414896 73170 414952
rect 73226 414896 73312 414952
rect 73368 414896 73416 414952
rect 70000 414857 73416 414896
rect 70000 414801 70047 414857
rect 70103 414801 70171 414857
rect 70227 414801 70295 414857
rect 70351 414801 70419 414857
rect 70475 414810 73416 414857
rect 70475 414801 71466 414810
rect 70000 414754 71466 414801
rect 71522 414754 71608 414810
rect 71664 414754 71750 414810
rect 71806 414754 71892 414810
rect 71948 414754 72034 414810
rect 72090 414754 72176 414810
rect 72232 414754 72318 414810
rect 72374 414754 72460 414810
rect 72516 414754 72602 414810
rect 72658 414754 72744 414810
rect 72800 414754 72886 414810
rect 72942 414754 73028 414810
rect 73084 414754 73170 414810
rect 73226 414754 73312 414810
rect 73368 414754 73416 414810
rect 70000 414733 73416 414754
rect 70000 414677 70047 414733
rect 70103 414677 70171 414733
rect 70227 414677 70295 414733
rect 70351 414677 70419 414733
rect 70475 414677 73416 414733
rect 70000 414668 73416 414677
rect 70000 414612 71466 414668
rect 71522 414612 71608 414668
rect 71664 414612 71750 414668
rect 71806 414612 71892 414668
rect 71948 414612 72034 414668
rect 72090 414612 72176 414668
rect 72232 414612 72318 414668
rect 72374 414612 72460 414668
rect 72516 414612 72602 414668
rect 72658 414612 72744 414668
rect 72800 414612 72886 414668
rect 72942 414612 73028 414668
rect 73084 414612 73170 414668
rect 73226 414612 73312 414668
rect 73368 414612 73416 414668
rect 70000 414609 73416 414612
rect 70000 414553 70047 414609
rect 70103 414553 70171 414609
rect 70227 414553 70295 414609
rect 70351 414553 70419 414609
rect 70475 414553 73416 414609
rect 70000 414526 73416 414553
rect 70000 414485 71466 414526
rect 70000 414429 70047 414485
rect 70103 414429 70171 414485
rect 70227 414429 70295 414485
rect 70351 414429 70419 414485
rect 70475 414470 71466 414485
rect 71522 414470 71608 414526
rect 71664 414470 71750 414526
rect 71806 414470 71892 414526
rect 71948 414470 72034 414526
rect 72090 414470 72176 414526
rect 72232 414470 72318 414526
rect 72374 414470 72460 414526
rect 72516 414470 72602 414526
rect 72658 414470 72744 414526
rect 72800 414470 72886 414526
rect 72942 414470 73028 414526
rect 73084 414470 73170 414526
rect 73226 414470 73312 414526
rect 73368 414470 73416 414526
rect 70475 414429 73416 414470
rect 70000 414384 73416 414429
rect 70000 414361 71466 414384
rect 70000 414305 70047 414361
rect 70103 414305 70171 414361
rect 70227 414305 70295 414361
rect 70351 414305 70419 414361
rect 70475 414328 71466 414361
rect 71522 414328 71608 414384
rect 71664 414328 71750 414384
rect 71806 414328 71892 414384
rect 71948 414328 72034 414384
rect 72090 414328 72176 414384
rect 72232 414328 72318 414384
rect 72374 414328 72460 414384
rect 72516 414328 72602 414384
rect 72658 414328 72744 414384
rect 72800 414328 72886 414384
rect 72942 414328 73028 414384
rect 73084 414328 73170 414384
rect 73226 414328 73312 414384
rect 73368 414328 73416 414384
rect 70475 414305 73416 414328
rect 70000 414242 73416 414305
rect 70000 414237 71466 414242
rect 70000 414181 70047 414237
rect 70103 414181 70171 414237
rect 70227 414181 70295 414237
rect 70351 414181 70419 414237
rect 70475 414186 71466 414237
rect 71522 414186 71608 414242
rect 71664 414186 71750 414242
rect 71806 414186 71892 414242
rect 71948 414186 72034 414242
rect 72090 414186 72176 414242
rect 72232 414186 72318 414242
rect 72374 414186 72460 414242
rect 72516 414186 72602 414242
rect 72658 414186 72744 414242
rect 72800 414186 72886 414242
rect 72942 414186 73028 414242
rect 73084 414186 73170 414242
rect 73226 414186 73312 414242
rect 73368 414186 73416 414242
rect 70475 414181 73416 414186
rect 70000 414113 73416 414181
rect 70000 414057 70047 414113
rect 70103 414057 70171 414113
rect 70227 414057 70295 414113
rect 70351 414057 70419 414113
rect 70475 414100 73416 414113
rect 70475 414057 71466 414100
rect 70000 414044 71466 414057
rect 71522 414044 71608 414100
rect 71664 414044 71750 414100
rect 71806 414044 71892 414100
rect 71948 414044 72034 414100
rect 72090 414044 72176 414100
rect 72232 414044 72318 414100
rect 72374 414044 72460 414100
rect 72516 414044 72602 414100
rect 72658 414044 72744 414100
rect 72800 414044 72886 414100
rect 72942 414044 73028 414100
rect 73084 414044 73170 414100
rect 73226 414044 73312 414100
rect 73368 414044 73416 414100
rect 70000 413989 73416 414044
rect 70000 413933 70047 413989
rect 70103 413933 70171 413989
rect 70227 413933 70295 413989
rect 70351 413933 70419 413989
rect 70475 413958 73416 413989
rect 70475 413933 71466 413958
rect 70000 413902 71466 413933
rect 71522 413902 71608 413958
rect 71664 413902 71750 413958
rect 71806 413902 71892 413958
rect 71948 413902 72034 413958
rect 72090 413902 72176 413958
rect 72232 413902 72318 413958
rect 72374 413902 72460 413958
rect 72516 413902 72602 413958
rect 72658 413902 72744 413958
rect 72800 413902 72886 413958
rect 72942 413902 73028 413958
rect 73084 413902 73170 413958
rect 73226 413902 73312 413958
rect 73368 413902 73416 413958
rect 70000 413865 73416 413902
rect 70000 413809 70047 413865
rect 70103 413809 70171 413865
rect 70227 413809 70295 413865
rect 70351 413809 70419 413865
rect 70475 413816 73416 413865
rect 70475 413809 71466 413816
rect 70000 413760 71466 413809
rect 71522 413760 71608 413816
rect 71664 413760 71750 413816
rect 71806 413760 71892 413816
rect 71948 413760 72034 413816
rect 72090 413760 72176 413816
rect 72232 413760 72318 413816
rect 72374 413760 72460 413816
rect 72516 413760 72602 413816
rect 72658 413760 72744 413816
rect 72800 413760 72886 413816
rect 72942 413760 73028 413816
rect 73084 413760 73170 413816
rect 73226 413760 73312 413816
rect 73368 413760 73416 413816
rect 70000 413741 73416 413760
rect 70000 413685 70047 413741
rect 70103 413685 70171 413741
rect 70227 413685 70295 413741
rect 70351 413685 70419 413741
rect 70475 413685 73416 413741
rect 70000 413674 73416 413685
rect 70000 413618 71466 413674
rect 71522 413618 71608 413674
rect 71664 413618 71750 413674
rect 71806 413618 71892 413674
rect 71948 413618 72034 413674
rect 72090 413618 72176 413674
rect 72232 413618 72318 413674
rect 72374 413618 72460 413674
rect 72516 413618 72602 413674
rect 72658 413618 72744 413674
rect 72800 413618 72886 413674
rect 72942 413618 73028 413674
rect 73084 413618 73170 413674
rect 73226 413618 73312 413674
rect 73368 413618 73416 413674
rect 70000 413617 73416 413618
rect 70000 413561 70047 413617
rect 70103 413561 70171 413617
rect 70227 413561 70295 413617
rect 70351 413561 70419 413617
rect 70475 413561 73416 413617
rect 70000 413532 73416 413561
rect 70000 413493 71466 413532
rect 70000 413437 70047 413493
rect 70103 413437 70171 413493
rect 70227 413437 70295 413493
rect 70351 413437 70419 413493
rect 70475 413476 71466 413493
rect 71522 413476 71608 413532
rect 71664 413476 71750 413532
rect 71806 413476 71892 413532
rect 71948 413476 72034 413532
rect 72090 413476 72176 413532
rect 72232 413476 72318 413532
rect 72374 413476 72460 413532
rect 72516 413476 72602 413532
rect 72658 413476 72744 413532
rect 72800 413476 72886 413532
rect 72942 413476 73028 413532
rect 73084 413476 73170 413532
rect 73226 413476 73312 413532
rect 73368 413476 73416 413532
rect 70475 413437 73416 413476
rect 70000 413390 73416 413437
rect 70000 413369 71466 413390
rect 70000 413313 70047 413369
rect 70103 413313 70171 413369
rect 70227 413313 70295 413369
rect 70351 413313 70419 413369
rect 70475 413334 71466 413369
rect 71522 413334 71608 413390
rect 71664 413334 71750 413390
rect 71806 413334 71892 413390
rect 71948 413334 72034 413390
rect 72090 413334 72176 413390
rect 72232 413334 72318 413390
rect 72374 413334 72460 413390
rect 72516 413334 72602 413390
rect 72658 413334 72744 413390
rect 72800 413334 72886 413390
rect 72942 413334 73028 413390
rect 73084 413334 73170 413390
rect 73226 413334 73312 413390
rect 73368 413334 73416 413390
rect 70475 413313 73416 413334
rect 70000 413272 73416 413313
rect 702392 404687 706000 404728
rect 702392 404666 705525 404687
rect 702392 404610 702440 404666
rect 702496 404610 702582 404666
rect 702638 404610 702724 404666
rect 702780 404610 702866 404666
rect 702922 404610 703008 404666
rect 703064 404610 703150 404666
rect 703206 404610 703292 404666
rect 703348 404610 703434 404666
rect 703490 404610 703576 404666
rect 703632 404610 703718 404666
rect 703774 404610 703860 404666
rect 703916 404610 704002 404666
rect 704058 404610 704144 404666
rect 704200 404610 704286 404666
rect 704342 404631 705525 404666
rect 705581 404631 705649 404687
rect 705705 404631 705773 404687
rect 705829 404631 705897 404687
rect 705953 404631 706000 404687
rect 704342 404610 706000 404631
rect 702392 404563 706000 404610
rect 702392 404524 705525 404563
rect 702392 404468 702440 404524
rect 702496 404468 702582 404524
rect 702638 404468 702724 404524
rect 702780 404468 702866 404524
rect 702922 404468 703008 404524
rect 703064 404468 703150 404524
rect 703206 404468 703292 404524
rect 703348 404468 703434 404524
rect 703490 404468 703576 404524
rect 703632 404468 703718 404524
rect 703774 404468 703860 404524
rect 703916 404468 704002 404524
rect 704058 404468 704144 404524
rect 704200 404468 704286 404524
rect 704342 404507 705525 404524
rect 705581 404507 705649 404563
rect 705705 404507 705773 404563
rect 705829 404507 705897 404563
rect 705953 404507 706000 404563
rect 704342 404468 706000 404507
rect 702392 404439 706000 404468
rect 702392 404383 705525 404439
rect 705581 404383 705649 404439
rect 705705 404383 705773 404439
rect 705829 404383 705897 404439
rect 705953 404383 706000 404439
rect 702392 404382 706000 404383
rect 702392 404326 702440 404382
rect 702496 404326 702582 404382
rect 702638 404326 702724 404382
rect 702780 404326 702866 404382
rect 702922 404326 703008 404382
rect 703064 404326 703150 404382
rect 703206 404326 703292 404382
rect 703348 404326 703434 404382
rect 703490 404326 703576 404382
rect 703632 404326 703718 404382
rect 703774 404326 703860 404382
rect 703916 404326 704002 404382
rect 704058 404326 704144 404382
rect 704200 404326 704286 404382
rect 704342 404326 706000 404382
rect 702392 404315 706000 404326
rect 702392 404259 705525 404315
rect 705581 404259 705649 404315
rect 705705 404259 705773 404315
rect 705829 404259 705897 404315
rect 705953 404259 706000 404315
rect 702392 404240 706000 404259
rect 702392 404184 702440 404240
rect 702496 404184 702582 404240
rect 702638 404184 702724 404240
rect 702780 404184 702866 404240
rect 702922 404184 703008 404240
rect 703064 404184 703150 404240
rect 703206 404184 703292 404240
rect 703348 404184 703434 404240
rect 703490 404184 703576 404240
rect 703632 404184 703718 404240
rect 703774 404184 703860 404240
rect 703916 404184 704002 404240
rect 704058 404184 704144 404240
rect 704200 404184 704286 404240
rect 704342 404191 706000 404240
rect 704342 404184 705525 404191
rect 702392 404135 705525 404184
rect 705581 404135 705649 404191
rect 705705 404135 705773 404191
rect 705829 404135 705897 404191
rect 705953 404135 706000 404191
rect 702392 404098 706000 404135
rect 702392 404042 702440 404098
rect 702496 404042 702582 404098
rect 702638 404042 702724 404098
rect 702780 404042 702866 404098
rect 702922 404042 703008 404098
rect 703064 404042 703150 404098
rect 703206 404042 703292 404098
rect 703348 404042 703434 404098
rect 703490 404042 703576 404098
rect 703632 404042 703718 404098
rect 703774 404042 703860 404098
rect 703916 404042 704002 404098
rect 704058 404042 704144 404098
rect 704200 404042 704286 404098
rect 704342 404067 706000 404098
rect 704342 404042 705525 404067
rect 702392 404011 705525 404042
rect 705581 404011 705649 404067
rect 705705 404011 705773 404067
rect 705829 404011 705897 404067
rect 705953 404011 706000 404067
rect 702392 403956 706000 404011
rect 702392 403900 702440 403956
rect 702496 403900 702582 403956
rect 702638 403900 702724 403956
rect 702780 403900 702866 403956
rect 702922 403900 703008 403956
rect 703064 403900 703150 403956
rect 703206 403900 703292 403956
rect 703348 403900 703434 403956
rect 703490 403900 703576 403956
rect 703632 403900 703718 403956
rect 703774 403900 703860 403956
rect 703916 403900 704002 403956
rect 704058 403900 704144 403956
rect 704200 403900 704286 403956
rect 704342 403943 706000 403956
rect 704342 403900 705525 403943
rect 702392 403887 705525 403900
rect 705581 403887 705649 403943
rect 705705 403887 705773 403943
rect 705829 403887 705897 403943
rect 705953 403887 706000 403943
rect 702392 403819 706000 403887
rect 702392 403814 705525 403819
rect 702392 403758 702440 403814
rect 702496 403758 702582 403814
rect 702638 403758 702724 403814
rect 702780 403758 702866 403814
rect 702922 403758 703008 403814
rect 703064 403758 703150 403814
rect 703206 403758 703292 403814
rect 703348 403758 703434 403814
rect 703490 403758 703576 403814
rect 703632 403758 703718 403814
rect 703774 403758 703860 403814
rect 703916 403758 704002 403814
rect 704058 403758 704144 403814
rect 704200 403758 704286 403814
rect 704342 403763 705525 403814
rect 705581 403763 705649 403819
rect 705705 403763 705773 403819
rect 705829 403763 705897 403819
rect 705953 403763 706000 403819
rect 704342 403758 706000 403763
rect 702392 403695 706000 403758
rect 702392 403672 705525 403695
rect 702392 403616 702440 403672
rect 702496 403616 702582 403672
rect 702638 403616 702724 403672
rect 702780 403616 702866 403672
rect 702922 403616 703008 403672
rect 703064 403616 703150 403672
rect 703206 403616 703292 403672
rect 703348 403616 703434 403672
rect 703490 403616 703576 403672
rect 703632 403616 703718 403672
rect 703774 403616 703860 403672
rect 703916 403616 704002 403672
rect 704058 403616 704144 403672
rect 704200 403616 704286 403672
rect 704342 403639 705525 403672
rect 705581 403639 705649 403695
rect 705705 403639 705773 403695
rect 705829 403639 705897 403695
rect 705953 403639 706000 403695
rect 704342 403616 706000 403639
rect 702392 403571 706000 403616
rect 702392 403530 705525 403571
rect 702392 403474 702440 403530
rect 702496 403474 702582 403530
rect 702638 403474 702724 403530
rect 702780 403474 702866 403530
rect 702922 403474 703008 403530
rect 703064 403474 703150 403530
rect 703206 403474 703292 403530
rect 703348 403474 703434 403530
rect 703490 403474 703576 403530
rect 703632 403474 703718 403530
rect 703774 403474 703860 403530
rect 703916 403474 704002 403530
rect 704058 403474 704144 403530
rect 704200 403474 704286 403530
rect 704342 403515 705525 403530
rect 705581 403515 705649 403571
rect 705705 403515 705773 403571
rect 705829 403515 705897 403571
rect 705953 403515 706000 403571
rect 704342 403474 706000 403515
rect 702392 403447 706000 403474
rect 702392 403391 705525 403447
rect 705581 403391 705649 403447
rect 705705 403391 705773 403447
rect 705829 403391 705897 403447
rect 705953 403391 706000 403447
rect 702392 403388 706000 403391
rect 702392 403332 702440 403388
rect 702496 403332 702582 403388
rect 702638 403332 702724 403388
rect 702780 403332 702866 403388
rect 702922 403332 703008 403388
rect 703064 403332 703150 403388
rect 703206 403332 703292 403388
rect 703348 403332 703434 403388
rect 703490 403332 703576 403388
rect 703632 403332 703718 403388
rect 703774 403332 703860 403388
rect 703916 403332 704002 403388
rect 704058 403332 704144 403388
rect 704200 403332 704286 403388
rect 704342 403332 706000 403388
rect 702392 403323 706000 403332
rect 702392 403267 705525 403323
rect 705581 403267 705649 403323
rect 705705 403267 705773 403323
rect 705829 403267 705897 403323
rect 705953 403267 706000 403323
rect 702392 403246 706000 403267
rect 702392 403190 702440 403246
rect 702496 403190 702582 403246
rect 702638 403190 702724 403246
rect 702780 403190 702866 403246
rect 702922 403190 703008 403246
rect 703064 403190 703150 403246
rect 703206 403190 703292 403246
rect 703348 403190 703434 403246
rect 703490 403190 703576 403246
rect 703632 403190 703718 403246
rect 703774 403190 703860 403246
rect 703916 403190 704002 403246
rect 704058 403190 704144 403246
rect 704200 403190 704286 403246
rect 704342 403199 706000 403246
rect 704342 403190 705525 403199
rect 702392 403143 705525 403190
rect 705581 403143 705649 403199
rect 705705 403143 705773 403199
rect 705829 403143 705897 403199
rect 705953 403143 706000 403199
rect 702392 403104 706000 403143
rect 702392 403048 702440 403104
rect 702496 403048 702582 403104
rect 702638 403048 702724 403104
rect 702780 403048 702866 403104
rect 702922 403048 703008 403104
rect 703064 403048 703150 403104
rect 703206 403048 703292 403104
rect 703348 403048 703434 403104
rect 703490 403048 703576 403104
rect 703632 403048 703718 403104
rect 703774 403048 703860 403104
rect 703916 403048 704002 403104
rect 704058 403048 704144 403104
rect 704200 403048 704286 403104
rect 704342 403075 706000 403104
rect 704342 403048 705525 403075
rect 702392 403019 705525 403048
rect 705581 403019 705649 403075
rect 705705 403019 705773 403075
rect 705829 403019 705897 403075
rect 705953 403019 706000 403075
rect 702392 402962 706000 403019
rect 702392 402906 702440 402962
rect 702496 402906 702582 402962
rect 702638 402906 702724 402962
rect 702780 402906 702866 402962
rect 702922 402906 703008 402962
rect 703064 402906 703150 402962
rect 703206 402906 703292 402962
rect 703348 402906 703434 402962
rect 703490 402906 703576 402962
rect 703632 402906 703718 402962
rect 703774 402906 703860 402962
rect 703916 402906 704002 402962
rect 704058 402906 704144 402962
rect 704200 402906 704286 402962
rect 704342 402951 706000 402962
rect 704342 402906 705525 402951
rect 702392 402895 705525 402906
rect 705581 402895 705649 402951
rect 705705 402895 705773 402951
rect 705829 402895 705897 402951
rect 705953 402895 706000 402951
rect 702392 402828 706000 402895
rect 702392 402181 706000 402248
rect 702392 402179 705525 402181
rect 702392 402123 702451 402179
rect 702507 402123 702593 402179
rect 702649 402123 702735 402179
rect 702791 402123 702877 402179
rect 702933 402123 703019 402179
rect 703075 402123 703161 402179
rect 703217 402123 703303 402179
rect 703359 402123 703445 402179
rect 703501 402123 703587 402179
rect 703643 402123 703729 402179
rect 703785 402123 703871 402179
rect 703927 402123 704013 402179
rect 704069 402123 704155 402179
rect 704211 402123 704297 402179
rect 704353 402125 705525 402179
rect 705581 402125 705649 402181
rect 705705 402125 705773 402181
rect 705829 402125 705897 402181
rect 705953 402125 706000 402181
rect 704353 402123 706000 402125
rect 702392 402057 706000 402123
rect 702392 402037 705525 402057
rect 702392 401981 702451 402037
rect 702507 401981 702593 402037
rect 702649 401981 702735 402037
rect 702791 401981 702877 402037
rect 702933 401981 703019 402037
rect 703075 401981 703161 402037
rect 703217 401981 703303 402037
rect 703359 401981 703445 402037
rect 703501 401981 703587 402037
rect 703643 401981 703729 402037
rect 703785 401981 703871 402037
rect 703927 401981 704013 402037
rect 704069 401981 704155 402037
rect 704211 401981 704297 402037
rect 704353 402001 705525 402037
rect 705581 402001 705649 402057
rect 705705 402001 705773 402057
rect 705829 402001 705897 402057
rect 705953 402001 706000 402057
rect 704353 401981 706000 402001
rect 702392 401933 706000 401981
rect 702392 401895 705525 401933
rect 702392 401839 702451 401895
rect 702507 401839 702593 401895
rect 702649 401839 702735 401895
rect 702791 401839 702877 401895
rect 702933 401839 703019 401895
rect 703075 401839 703161 401895
rect 703217 401839 703303 401895
rect 703359 401839 703445 401895
rect 703501 401839 703587 401895
rect 703643 401839 703729 401895
rect 703785 401839 703871 401895
rect 703927 401839 704013 401895
rect 704069 401839 704155 401895
rect 704211 401839 704297 401895
rect 704353 401877 705525 401895
rect 705581 401877 705649 401933
rect 705705 401877 705773 401933
rect 705829 401877 705897 401933
rect 705953 401877 706000 401933
rect 704353 401839 706000 401877
rect 702392 401809 706000 401839
rect 702392 401753 705525 401809
rect 705581 401753 705649 401809
rect 705705 401753 705773 401809
rect 705829 401753 705897 401809
rect 705953 401753 706000 401809
rect 702392 401697 702451 401753
rect 702507 401697 702593 401753
rect 702649 401697 702735 401753
rect 702791 401697 702877 401753
rect 702933 401697 703019 401753
rect 703075 401697 703161 401753
rect 703217 401697 703303 401753
rect 703359 401697 703445 401753
rect 703501 401697 703587 401753
rect 703643 401697 703729 401753
rect 703785 401697 703871 401753
rect 703927 401697 704013 401753
rect 704069 401697 704155 401753
rect 704211 401697 704297 401753
rect 704353 401697 706000 401753
rect 702392 401685 706000 401697
rect 702392 401629 705525 401685
rect 705581 401629 705649 401685
rect 705705 401629 705773 401685
rect 705829 401629 705897 401685
rect 705953 401629 706000 401685
rect 702392 401611 706000 401629
rect 702392 401555 702451 401611
rect 702507 401555 702593 401611
rect 702649 401555 702735 401611
rect 702791 401555 702877 401611
rect 702933 401555 703019 401611
rect 703075 401555 703161 401611
rect 703217 401555 703303 401611
rect 703359 401555 703445 401611
rect 703501 401555 703587 401611
rect 703643 401555 703729 401611
rect 703785 401555 703871 401611
rect 703927 401555 704013 401611
rect 704069 401555 704155 401611
rect 704211 401555 704297 401611
rect 704353 401561 706000 401611
rect 704353 401555 705525 401561
rect 702392 401505 705525 401555
rect 705581 401505 705649 401561
rect 705705 401505 705773 401561
rect 705829 401505 705897 401561
rect 705953 401505 706000 401561
rect 702392 401469 706000 401505
rect 702392 401413 702451 401469
rect 702507 401413 702593 401469
rect 702649 401413 702735 401469
rect 702791 401413 702877 401469
rect 702933 401413 703019 401469
rect 703075 401413 703161 401469
rect 703217 401413 703303 401469
rect 703359 401413 703445 401469
rect 703501 401413 703587 401469
rect 703643 401413 703729 401469
rect 703785 401413 703871 401469
rect 703927 401413 704013 401469
rect 704069 401413 704155 401469
rect 704211 401413 704297 401469
rect 704353 401437 706000 401469
rect 704353 401413 705525 401437
rect 702392 401381 705525 401413
rect 705581 401381 705649 401437
rect 705705 401381 705773 401437
rect 705829 401381 705897 401437
rect 705953 401381 706000 401437
rect 702392 401327 706000 401381
rect 702392 401271 702451 401327
rect 702507 401271 702593 401327
rect 702649 401271 702735 401327
rect 702791 401271 702877 401327
rect 702933 401271 703019 401327
rect 703075 401271 703161 401327
rect 703217 401271 703303 401327
rect 703359 401271 703445 401327
rect 703501 401271 703587 401327
rect 703643 401271 703729 401327
rect 703785 401271 703871 401327
rect 703927 401271 704013 401327
rect 704069 401271 704155 401327
rect 704211 401271 704297 401327
rect 704353 401313 706000 401327
rect 704353 401271 705525 401313
rect 702392 401257 705525 401271
rect 705581 401257 705649 401313
rect 705705 401257 705773 401313
rect 705829 401257 705897 401313
rect 705953 401257 706000 401313
rect 702392 401189 706000 401257
rect 702392 401185 705525 401189
rect 702392 401129 702451 401185
rect 702507 401129 702593 401185
rect 702649 401129 702735 401185
rect 702791 401129 702877 401185
rect 702933 401129 703019 401185
rect 703075 401129 703161 401185
rect 703217 401129 703303 401185
rect 703359 401129 703445 401185
rect 703501 401129 703587 401185
rect 703643 401129 703729 401185
rect 703785 401129 703871 401185
rect 703927 401129 704013 401185
rect 704069 401129 704155 401185
rect 704211 401129 704297 401185
rect 704353 401133 705525 401185
rect 705581 401133 705649 401189
rect 705705 401133 705773 401189
rect 705829 401133 705897 401189
rect 705953 401133 706000 401189
rect 704353 401129 706000 401133
rect 702392 401065 706000 401129
rect 702392 401043 705525 401065
rect 702392 400987 702451 401043
rect 702507 400987 702593 401043
rect 702649 400987 702735 401043
rect 702791 400987 702877 401043
rect 702933 400987 703019 401043
rect 703075 400987 703161 401043
rect 703217 400987 703303 401043
rect 703359 400987 703445 401043
rect 703501 400987 703587 401043
rect 703643 400987 703729 401043
rect 703785 400987 703871 401043
rect 703927 400987 704013 401043
rect 704069 400987 704155 401043
rect 704211 400987 704297 401043
rect 704353 401009 705525 401043
rect 705581 401009 705649 401065
rect 705705 401009 705773 401065
rect 705829 401009 705897 401065
rect 705953 401009 706000 401065
rect 704353 400987 706000 401009
rect 702392 400941 706000 400987
rect 702392 400901 705525 400941
rect 702392 400845 702451 400901
rect 702507 400845 702593 400901
rect 702649 400845 702735 400901
rect 702791 400845 702877 400901
rect 702933 400845 703019 400901
rect 703075 400845 703161 400901
rect 703217 400845 703303 400901
rect 703359 400845 703445 400901
rect 703501 400845 703587 400901
rect 703643 400845 703729 400901
rect 703785 400845 703871 400901
rect 703927 400845 704013 400901
rect 704069 400845 704155 400901
rect 704211 400845 704297 400901
rect 704353 400885 705525 400901
rect 705581 400885 705649 400941
rect 705705 400885 705773 400941
rect 705829 400885 705897 400941
rect 705953 400885 706000 400941
rect 704353 400845 706000 400885
rect 702392 400817 706000 400845
rect 702392 400761 705525 400817
rect 705581 400761 705649 400817
rect 705705 400761 705773 400817
rect 705829 400761 705897 400817
rect 705953 400761 706000 400817
rect 702392 400759 706000 400761
rect 702392 400703 702451 400759
rect 702507 400703 702593 400759
rect 702649 400703 702735 400759
rect 702791 400703 702877 400759
rect 702933 400703 703019 400759
rect 703075 400703 703161 400759
rect 703217 400703 703303 400759
rect 703359 400703 703445 400759
rect 703501 400703 703587 400759
rect 703643 400703 703729 400759
rect 703785 400703 703871 400759
rect 703927 400703 704013 400759
rect 704069 400703 704155 400759
rect 704211 400703 704297 400759
rect 704353 400703 706000 400759
rect 702392 400693 706000 400703
rect 702392 400637 705525 400693
rect 705581 400637 705649 400693
rect 705705 400637 705773 400693
rect 705829 400637 705897 400693
rect 705953 400637 706000 400693
rect 702392 400617 706000 400637
rect 702392 400561 702451 400617
rect 702507 400561 702593 400617
rect 702649 400561 702735 400617
rect 702791 400561 702877 400617
rect 702933 400561 703019 400617
rect 703075 400561 703161 400617
rect 703217 400561 703303 400617
rect 703359 400561 703445 400617
rect 703501 400561 703587 400617
rect 703643 400561 703729 400617
rect 703785 400561 703871 400617
rect 703927 400561 704013 400617
rect 704069 400561 704155 400617
rect 704211 400561 704297 400617
rect 704353 400569 706000 400617
rect 704353 400561 705525 400569
rect 702392 400513 705525 400561
rect 705581 400513 705649 400569
rect 705705 400513 705773 400569
rect 705829 400513 705897 400569
rect 705953 400513 706000 400569
rect 702392 400475 706000 400513
rect 702392 400419 702451 400475
rect 702507 400419 702593 400475
rect 702649 400419 702735 400475
rect 702791 400419 702877 400475
rect 702933 400419 703019 400475
rect 703075 400419 703161 400475
rect 703217 400419 703303 400475
rect 703359 400419 703445 400475
rect 703501 400419 703587 400475
rect 703643 400419 703729 400475
rect 703785 400419 703871 400475
rect 703927 400419 704013 400475
rect 704069 400419 704155 400475
rect 704211 400419 704297 400475
rect 704353 400445 706000 400475
rect 704353 400419 705525 400445
rect 702392 400389 705525 400419
rect 705581 400389 705649 400445
rect 705705 400389 705773 400445
rect 705829 400389 705897 400445
rect 705953 400389 706000 400445
rect 702392 400333 706000 400389
rect 702392 400277 702451 400333
rect 702507 400277 702593 400333
rect 702649 400277 702735 400333
rect 702791 400277 702877 400333
rect 702933 400277 703019 400333
rect 703075 400277 703161 400333
rect 703217 400277 703303 400333
rect 703359 400277 703445 400333
rect 703501 400277 703587 400333
rect 703643 400277 703729 400333
rect 703785 400277 703871 400333
rect 703927 400277 704013 400333
rect 704069 400277 704155 400333
rect 704211 400277 704297 400333
rect 704353 400321 706000 400333
rect 704353 400277 705525 400321
rect 702392 400265 705525 400277
rect 705581 400265 705649 400321
rect 705705 400265 705773 400321
rect 705829 400265 705897 400321
rect 705953 400265 706000 400321
rect 702392 400198 706000 400265
rect 702392 399811 706000 399878
rect 702392 399809 705525 399811
rect 702392 399753 702451 399809
rect 702507 399753 702593 399809
rect 702649 399753 702735 399809
rect 702791 399753 702877 399809
rect 702933 399753 703019 399809
rect 703075 399753 703161 399809
rect 703217 399753 703303 399809
rect 703359 399753 703445 399809
rect 703501 399753 703587 399809
rect 703643 399753 703729 399809
rect 703785 399753 703871 399809
rect 703927 399753 704013 399809
rect 704069 399753 704155 399809
rect 704211 399753 704297 399809
rect 704353 399755 705525 399809
rect 705581 399755 705649 399811
rect 705705 399755 705773 399811
rect 705829 399755 705897 399811
rect 705953 399755 706000 399811
rect 704353 399753 706000 399755
rect 702392 399687 706000 399753
rect 702392 399667 705525 399687
rect 702392 399611 702451 399667
rect 702507 399611 702593 399667
rect 702649 399611 702735 399667
rect 702791 399611 702877 399667
rect 702933 399611 703019 399667
rect 703075 399611 703161 399667
rect 703217 399611 703303 399667
rect 703359 399611 703445 399667
rect 703501 399611 703587 399667
rect 703643 399611 703729 399667
rect 703785 399611 703871 399667
rect 703927 399611 704013 399667
rect 704069 399611 704155 399667
rect 704211 399611 704297 399667
rect 704353 399631 705525 399667
rect 705581 399631 705649 399687
rect 705705 399631 705773 399687
rect 705829 399631 705897 399687
rect 705953 399631 706000 399687
rect 704353 399611 706000 399631
rect 702392 399563 706000 399611
rect 702392 399525 705525 399563
rect 702392 399469 702451 399525
rect 702507 399469 702593 399525
rect 702649 399469 702735 399525
rect 702791 399469 702877 399525
rect 702933 399469 703019 399525
rect 703075 399469 703161 399525
rect 703217 399469 703303 399525
rect 703359 399469 703445 399525
rect 703501 399469 703587 399525
rect 703643 399469 703729 399525
rect 703785 399469 703871 399525
rect 703927 399469 704013 399525
rect 704069 399469 704155 399525
rect 704211 399469 704297 399525
rect 704353 399507 705525 399525
rect 705581 399507 705649 399563
rect 705705 399507 705773 399563
rect 705829 399507 705897 399563
rect 705953 399507 706000 399563
rect 704353 399469 706000 399507
rect 702392 399439 706000 399469
rect 702392 399383 705525 399439
rect 705581 399383 705649 399439
rect 705705 399383 705773 399439
rect 705829 399383 705897 399439
rect 705953 399383 706000 399439
rect 702392 399327 702451 399383
rect 702507 399327 702593 399383
rect 702649 399327 702735 399383
rect 702791 399327 702877 399383
rect 702933 399327 703019 399383
rect 703075 399327 703161 399383
rect 703217 399327 703303 399383
rect 703359 399327 703445 399383
rect 703501 399327 703587 399383
rect 703643 399327 703729 399383
rect 703785 399327 703871 399383
rect 703927 399327 704013 399383
rect 704069 399327 704155 399383
rect 704211 399327 704297 399383
rect 704353 399327 706000 399383
rect 702392 399315 706000 399327
rect 702392 399259 705525 399315
rect 705581 399259 705649 399315
rect 705705 399259 705773 399315
rect 705829 399259 705897 399315
rect 705953 399259 706000 399315
rect 702392 399241 706000 399259
rect 702392 399185 702451 399241
rect 702507 399185 702593 399241
rect 702649 399185 702735 399241
rect 702791 399185 702877 399241
rect 702933 399185 703019 399241
rect 703075 399185 703161 399241
rect 703217 399185 703303 399241
rect 703359 399185 703445 399241
rect 703501 399185 703587 399241
rect 703643 399185 703729 399241
rect 703785 399185 703871 399241
rect 703927 399185 704013 399241
rect 704069 399185 704155 399241
rect 704211 399185 704297 399241
rect 704353 399191 706000 399241
rect 704353 399185 705525 399191
rect 702392 399135 705525 399185
rect 705581 399135 705649 399191
rect 705705 399135 705773 399191
rect 705829 399135 705897 399191
rect 705953 399135 706000 399191
rect 702392 399099 706000 399135
rect 702392 399043 702451 399099
rect 702507 399043 702593 399099
rect 702649 399043 702735 399099
rect 702791 399043 702877 399099
rect 702933 399043 703019 399099
rect 703075 399043 703161 399099
rect 703217 399043 703303 399099
rect 703359 399043 703445 399099
rect 703501 399043 703587 399099
rect 703643 399043 703729 399099
rect 703785 399043 703871 399099
rect 703927 399043 704013 399099
rect 704069 399043 704155 399099
rect 704211 399043 704297 399099
rect 704353 399067 706000 399099
rect 704353 399043 705525 399067
rect 702392 399011 705525 399043
rect 705581 399011 705649 399067
rect 705705 399011 705773 399067
rect 705829 399011 705897 399067
rect 705953 399011 706000 399067
rect 702392 398957 706000 399011
rect 702392 398901 702451 398957
rect 702507 398901 702593 398957
rect 702649 398901 702735 398957
rect 702791 398901 702877 398957
rect 702933 398901 703019 398957
rect 703075 398901 703161 398957
rect 703217 398901 703303 398957
rect 703359 398901 703445 398957
rect 703501 398901 703587 398957
rect 703643 398901 703729 398957
rect 703785 398901 703871 398957
rect 703927 398901 704013 398957
rect 704069 398901 704155 398957
rect 704211 398901 704297 398957
rect 704353 398943 706000 398957
rect 704353 398901 705525 398943
rect 702392 398887 705525 398901
rect 705581 398887 705649 398943
rect 705705 398887 705773 398943
rect 705829 398887 705897 398943
rect 705953 398887 706000 398943
rect 702392 398819 706000 398887
rect 702392 398815 705525 398819
rect 702392 398759 702451 398815
rect 702507 398759 702593 398815
rect 702649 398759 702735 398815
rect 702791 398759 702877 398815
rect 702933 398759 703019 398815
rect 703075 398759 703161 398815
rect 703217 398759 703303 398815
rect 703359 398759 703445 398815
rect 703501 398759 703587 398815
rect 703643 398759 703729 398815
rect 703785 398759 703871 398815
rect 703927 398759 704013 398815
rect 704069 398759 704155 398815
rect 704211 398759 704297 398815
rect 704353 398763 705525 398815
rect 705581 398763 705649 398819
rect 705705 398763 705773 398819
rect 705829 398763 705897 398819
rect 705953 398763 706000 398819
rect 704353 398759 706000 398763
rect 702392 398695 706000 398759
rect 702392 398673 705525 398695
rect 702392 398617 702451 398673
rect 702507 398617 702593 398673
rect 702649 398617 702735 398673
rect 702791 398617 702877 398673
rect 702933 398617 703019 398673
rect 703075 398617 703161 398673
rect 703217 398617 703303 398673
rect 703359 398617 703445 398673
rect 703501 398617 703587 398673
rect 703643 398617 703729 398673
rect 703785 398617 703871 398673
rect 703927 398617 704013 398673
rect 704069 398617 704155 398673
rect 704211 398617 704297 398673
rect 704353 398639 705525 398673
rect 705581 398639 705649 398695
rect 705705 398639 705773 398695
rect 705829 398639 705897 398695
rect 705953 398639 706000 398695
rect 704353 398617 706000 398639
rect 702392 398571 706000 398617
rect 702392 398531 705525 398571
rect 702392 398475 702451 398531
rect 702507 398475 702593 398531
rect 702649 398475 702735 398531
rect 702791 398475 702877 398531
rect 702933 398475 703019 398531
rect 703075 398475 703161 398531
rect 703217 398475 703303 398531
rect 703359 398475 703445 398531
rect 703501 398475 703587 398531
rect 703643 398475 703729 398531
rect 703785 398475 703871 398531
rect 703927 398475 704013 398531
rect 704069 398475 704155 398531
rect 704211 398475 704297 398531
rect 704353 398515 705525 398531
rect 705581 398515 705649 398571
rect 705705 398515 705773 398571
rect 705829 398515 705897 398571
rect 705953 398515 706000 398571
rect 704353 398475 706000 398515
rect 702392 398447 706000 398475
rect 702392 398391 705525 398447
rect 705581 398391 705649 398447
rect 705705 398391 705773 398447
rect 705829 398391 705897 398447
rect 705953 398391 706000 398447
rect 702392 398389 706000 398391
rect 702392 398333 702451 398389
rect 702507 398333 702593 398389
rect 702649 398333 702735 398389
rect 702791 398333 702877 398389
rect 702933 398333 703019 398389
rect 703075 398333 703161 398389
rect 703217 398333 703303 398389
rect 703359 398333 703445 398389
rect 703501 398333 703587 398389
rect 703643 398333 703729 398389
rect 703785 398333 703871 398389
rect 703927 398333 704013 398389
rect 704069 398333 704155 398389
rect 704211 398333 704297 398389
rect 704353 398333 706000 398389
rect 702392 398323 706000 398333
rect 702392 398267 705525 398323
rect 705581 398267 705649 398323
rect 705705 398267 705773 398323
rect 705829 398267 705897 398323
rect 705953 398267 706000 398323
rect 702392 398247 706000 398267
rect 702392 398191 702451 398247
rect 702507 398191 702593 398247
rect 702649 398191 702735 398247
rect 702791 398191 702877 398247
rect 702933 398191 703019 398247
rect 703075 398191 703161 398247
rect 703217 398191 703303 398247
rect 703359 398191 703445 398247
rect 703501 398191 703587 398247
rect 703643 398191 703729 398247
rect 703785 398191 703871 398247
rect 703927 398191 704013 398247
rect 704069 398191 704155 398247
rect 704211 398191 704297 398247
rect 704353 398199 706000 398247
rect 704353 398191 705525 398199
rect 702392 398143 705525 398191
rect 705581 398143 705649 398199
rect 705705 398143 705773 398199
rect 705829 398143 705897 398199
rect 705953 398143 706000 398199
rect 702392 398105 706000 398143
rect 702392 398049 702451 398105
rect 702507 398049 702593 398105
rect 702649 398049 702735 398105
rect 702791 398049 702877 398105
rect 702933 398049 703019 398105
rect 703075 398049 703161 398105
rect 703217 398049 703303 398105
rect 703359 398049 703445 398105
rect 703501 398049 703587 398105
rect 703643 398049 703729 398105
rect 703785 398049 703871 398105
rect 703927 398049 704013 398105
rect 704069 398049 704155 398105
rect 704211 398049 704297 398105
rect 704353 398075 706000 398105
rect 704353 398049 705525 398075
rect 702392 398019 705525 398049
rect 705581 398019 705649 398075
rect 705705 398019 705773 398075
rect 705829 398019 705897 398075
rect 705953 398019 706000 398075
rect 702392 397963 706000 398019
rect 702392 397907 702451 397963
rect 702507 397907 702593 397963
rect 702649 397907 702735 397963
rect 702791 397907 702877 397963
rect 702933 397907 703019 397963
rect 703075 397907 703161 397963
rect 703217 397907 703303 397963
rect 703359 397907 703445 397963
rect 703501 397907 703587 397963
rect 703643 397907 703729 397963
rect 703785 397907 703871 397963
rect 703927 397907 704013 397963
rect 704069 397907 704155 397963
rect 704211 397907 704297 397963
rect 704353 397951 706000 397963
rect 704353 397907 705525 397951
rect 702392 397895 705525 397907
rect 705581 397895 705649 397951
rect 705705 397895 705773 397951
rect 705829 397895 705897 397951
rect 705953 397895 706000 397951
rect 702392 397828 706000 397895
rect 702392 397105 706000 397172
rect 702392 397103 705525 397105
rect 702392 397047 702451 397103
rect 702507 397047 702593 397103
rect 702649 397047 702735 397103
rect 702791 397047 702877 397103
rect 702933 397047 703019 397103
rect 703075 397047 703161 397103
rect 703217 397047 703303 397103
rect 703359 397047 703445 397103
rect 703501 397047 703587 397103
rect 703643 397047 703729 397103
rect 703785 397047 703871 397103
rect 703927 397047 704013 397103
rect 704069 397047 704155 397103
rect 704211 397047 704297 397103
rect 704353 397049 705525 397103
rect 705581 397049 705649 397105
rect 705705 397049 705773 397105
rect 705829 397049 705897 397105
rect 705953 397049 706000 397105
rect 704353 397047 706000 397049
rect 702392 396981 706000 397047
rect 702392 396961 705525 396981
rect 702392 396905 702451 396961
rect 702507 396905 702593 396961
rect 702649 396905 702735 396961
rect 702791 396905 702877 396961
rect 702933 396905 703019 396961
rect 703075 396905 703161 396961
rect 703217 396905 703303 396961
rect 703359 396905 703445 396961
rect 703501 396905 703587 396961
rect 703643 396905 703729 396961
rect 703785 396905 703871 396961
rect 703927 396905 704013 396961
rect 704069 396905 704155 396961
rect 704211 396905 704297 396961
rect 704353 396925 705525 396961
rect 705581 396925 705649 396981
rect 705705 396925 705773 396981
rect 705829 396925 705897 396981
rect 705953 396925 706000 396981
rect 704353 396905 706000 396925
rect 702392 396857 706000 396905
rect 702392 396819 705525 396857
rect 702392 396763 702451 396819
rect 702507 396763 702593 396819
rect 702649 396763 702735 396819
rect 702791 396763 702877 396819
rect 702933 396763 703019 396819
rect 703075 396763 703161 396819
rect 703217 396763 703303 396819
rect 703359 396763 703445 396819
rect 703501 396763 703587 396819
rect 703643 396763 703729 396819
rect 703785 396763 703871 396819
rect 703927 396763 704013 396819
rect 704069 396763 704155 396819
rect 704211 396763 704297 396819
rect 704353 396801 705525 396819
rect 705581 396801 705649 396857
rect 705705 396801 705773 396857
rect 705829 396801 705897 396857
rect 705953 396801 706000 396857
rect 704353 396763 706000 396801
rect 702392 396733 706000 396763
rect 702392 396677 705525 396733
rect 705581 396677 705649 396733
rect 705705 396677 705773 396733
rect 705829 396677 705897 396733
rect 705953 396677 706000 396733
rect 702392 396621 702451 396677
rect 702507 396621 702593 396677
rect 702649 396621 702735 396677
rect 702791 396621 702877 396677
rect 702933 396621 703019 396677
rect 703075 396621 703161 396677
rect 703217 396621 703303 396677
rect 703359 396621 703445 396677
rect 703501 396621 703587 396677
rect 703643 396621 703729 396677
rect 703785 396621 703871 396677
rect 703927 396621 704013 396677
rect 704069 396621 704155 396677
rect 704211 396621 704297 396677
rect 704353 396621 706000 396677
rect 702392 396609 706000 396621
rect 702392 396553 705525 396609
rect 705581 396553 705649 396609
rect 705705 396553 705773 396609
rect 705829 396553 705897 396609
rect 705953 396553 706000 396609
rect 702392 396535 706000 396553
rect 702392 396479 702451 396535
rect 702507 396479 702593 396535
rect 702649 396479 702735 396535
rect 702791 396479 702877 396535
rect 702933 396479 703019 396535
rect 703075 396479 703161 396535
rect 703217 396479 703303 396535
rect 703359 396479 703445 396535
rect 703501 396479 703587 396535
rect 703643 396479 703729 396535
rect 703785 396479 703871 396535
rect 703927 396479 704013 396535
rect 704069 396479 704155 396535
rect 704211 396479 704297 396535
rect 704353 396485 706000 396535
rect 704353 396479 705525 396485
rect 702392 396429 705525 396479
rect 705581 396429 705649 396485
rect 705705 396429 705773 396485
rect 705829 396429 705897 396485
rect 705953 396429 706000 396485
rect 702392 396393 706000 396429
rect 702392 396337 702451 396393
rect 702507 396337 702593 396393
rect 702649 396337 702735 396393
rect 702791 396337 702877 396393
rect 702933 396337 703019 396393
rect 703075 396337 703161 396393
rect 703217 396337 703303 396393
rect 703359 396337 703445 396393
rect 703501 396337 703587 396393
rect 703643 396337 703729 396393
rect 703785 396337 703871 396393
rect 703927 396337 704013 396393
rect 704069 396337 704155 396393
rect 704211 396337 704297 396393
rect 704353 396361 706000 396393
rect 704353 396337 705525 396361
rect 702392 396305 705525 396337
rect 705581 396305 705649 396361
rect 705705 396305 705773 396361
rect 705829 396305 705897 396361
rect 705953 396305 706000 396361
rect 702392 396251 706000 396305
rect 702392 396195 702451 396251
rect 702507 396195 702593 396251
rect 702649 396195 702735 396251
rect 702791 396195 702877 396251
rect 702933 396195 703019 396251
rect 703075 396195 703161 396251
rect 703217 396195 703303 396251
rect 703359 396195 703445 396251
rect 703501 396195 703587 396251
rect 703643 396195 703729 396251
rect 703785 396195 703871 396251
rect 703927 396195 704013 396251
rect 704069 396195 704155 396251
rect 704211 396195 704297 396251
rect 704353 396237 706000 396251
rect 704353 396195 705525 396237
rect 702392 396181 705525 396195
rect 705581 396181 705649 396237
rect 705705 396181 705773 396237
rect 705829 396181 705897 396237
rect 705953 396181 706000 396237
rect 702392 396113 706000 396181
rect 702392 396109 705525 396113
rect 702392 396053 702451 396109
rect 702507 396053 702593 396109
rect 702649 396053 702735 396109
rect 702791 396053 702877 396109
rect 702933 396053 703019 396109
rect 703075 396053 703161 396109
rect 703217 396053 703303 396109
rect 703359 396053 703445 396109
rect 703501 396053 703587 396109
rect 703643 396053 703729 396109
rect 703785 396053 703871 396109
rect 703927 396053 704013 396109
rect 704069 396053 704155 396109
rect 704211 396053 704297 396109
rect 704353 396057 705525 396109
rect 705581 396057 705649 396113
rect 705705 396057 705773 396113
rect 705829 396057 705897 396113
rect 705953 396057 706000 396113
rect 704353 396053 706000 396057
rect 702392 395989 706000 396053
rect 702392 395967 705525 395989
rect 702392 395911 702451 395967
rect 702507 395911 702593 395967
rect 702649 395911 702735 395967
rect 702791 395911 702877 395967
rect 702933 395911 703019 395967
rect 703075 395911 703161 395967
rect 703217 395911 703303 395967
rect 703359 395911 703445 395967
rect 703501 395911 703587 395967
rect 703643 395911 703729 395967
rect 703785 395911 703871 395967
rect 703927 395911 704013 395967
rect 704069 395911 704155 395967
rect 704211 395911 704297 395967
rect 704353 395933 705525 395967
rect 705581 395933 705649 395989
rect 705705 395933 705773 395989
rect 705829 395933 705897 395989
rect 705953 395933 706000 395989
rect 704353 395911 706000 395933
rect 702392 395865 706000 395911
rect 702392 395825 705525 395865
rect 702392 395769 702451 395825
rect 702507 395769 702593 395825
rect 702649 395769 702735 395825
rect 702791 395769 702877 395825
rect 702933 395769 703019 395825
rect 703075 395769 703161 395825
rect 703217 395769 703303 395825
rect 703359 395769 703445 395825
rect 703501 395769 703587 395825
rect 703643 395769 703729 395825
rect 703785 395769 703871 395825
rect 703927 395769 704013 395825
rect 704069 395769 704155 395825
rect 704211 395769 704297 395825
rect 704353 395809 705525 395825
rect 705581 395809 705649 395865
rect 705705 395809 705773 395865
rect 705829 395809 705897 395865
rect 705953 395809 706000 395865
rect 704353 395769 706000 395809
rect 702392 395741 706000 395769
rect 702392 395685 705525 395741
rect 705581 395685 705649 395741
rect 705705 395685 705773 395741
rect 705829 395685 705897 395741
rect 705953 395685 706000 395741
rect 702392 395683 706000 395685
rect 702392 395627 702451 395683
rect 702507 395627 702593 395683
rect 702649 395627 702735 395683
rect 702791 395627 702877 395683
rect 702933 395627 703019 395683
rect 703075 395627 703161 395683
rect 703217 395627 703303 395683
rect 703359 395627 703445 395683
rect 703501 395627 703587 395683
rect 703643 395627 703729 395683
rect 703785 395627 703871 395683
rect 703927 395627 704013 395683
rect 704069 395627 704155 395683
rect 704211 395627 704297 395683
rect 704353 395627 706000 395683
rect 702392 395617 706000 395627
rect 702392 395561 705525 395617
rect 705581 395561 705649 395617
rect 705705 395561 705773 395617
rect 705829 395561 705897 395617
rect 705953 395561 706000 395617
rect 702392 395541 706000 395561
rect 702392 395485 702451 395541
rect 702507 395485 702593 395541
rect 702649 395485 702735 395541
rect 702791 395485 702877 395541
rect 702933 395485 703019 395541
rect 703075 395485 703161 395541
rect 703217 395485 703303 395541
rect 703359 395485 703445 395541
rect 703501 395485 703587 395541
rect 703643 395485 703729 395541
rect 703785 395485 703871 395541
rect 703927 395485 704013 395541
rect 704069 395485 704155 395541
rect 704211 395485 704297 395541
rect 704353 395493 706000 395541
rect 704353 395485 705525 395493
rect 702392 395437 705525 395485
rect 705581 395437 705649 395493
rect 705705 395437 705773 395493
rect 705829 395437 705897 395493
rect 705953 395437 706000 395493
rect 702392 395399 706000 395437
rect 702392 395343 702451 395399
rect 702507 395343 702593 395399
rect 702649 395343 702735 395399
rect 702791 395343 702877 395399
rect 702933 395343 703019 395399
rect 703075 395343 703161 395399
rect 703217 395343 703303 395399
rect 703359 395343 703445 395399
rect 703501 395343 703587 395399
rect 703643 395343 703729 395399
rect 703785 395343 703871 395399
rect 703927 395343 704013 395399
rect 704069 395343 704155 395399
rect 704211 395343 704297 395399
rect 704353 395369 706000 395399
rect 704353 395343 705525 395369
rect 702392 395313 705525 395343
rect 705581 395313 705649 395369
rect 705705 395313 705773 395369
rect 705829 395313 705897 395369
rect 705953 395313 706000 395369
rect 702392 395257 706000 395313
rect 702392 395201 702451 395257
rect 702507 395201 702593 395257
rect 702649 395201 702735 395257
rect 702791 395201 702877 395257
rect 702933 395201 703019 395257
rect 703075 395201 703161 395257
rect 703217 395201 703303 395257
rect 703359 395201 703445 395257
rect 703501 395201 703587 395257
rect 703643 395201 703729 395257
rect 703785 395201 703871 395257
rect 703927 395201 704013 395257
rect 704069 395201 704155 395257
rect 704211 395201 704297 395257
rect 704353 395245 706000 395257
rect 704353 395201 705525 395245
rect 702392 395189 705525 395201
rect 705581 395189 705649 395245
rect 705705 395189 705773 395245
rect 705829 395189 705897 395245
rect 705953 395189 706000 395245
rect 702392 395122 706000 395189
rect 702392 394735 706000 394802
rect 702392 394733 705525 394735
rect 702392 394677 702451 394733
rect 702507 394677 702593 394733
rect 702649 394677 702735 394733
rect 702791 394677 702877 394733
rect 702933 394677 703019 394733
rect 703075 394677 703161 394733
rect 703217 394677 703303 394733
rect 703359 394677 703445 394733
rect 703501 394677 703587 394733
rect 703643 394677 703729 394733
rect 703785 394677 703871 394733
rect 703927 394677 704013 394733
rect 704069 394677 704155 394733
rect 704211 394677 704297 394733
rect 704353 394679 705525 394733
rect 705581 394679 705649 394735
rect 705705 394679 705773 394735
rect 705829 394679 705897 394735
rect 705953 394679 706000 394735
rect 704353 394677 706000 394679
rect 702392 394611 706000 394677
rect 702392 394591 705525 394611
rect 702392 394535 702451 394591
rect 702507 394535 702593 394591
rect 702649 394535 702735 394591
rect 702791 394535 702877 394591
rect 702933 394535 703019 394591
rect 703075 394535 703161 394591
rect 703217 394535 703303 394591
rect 703359 394535 703445 394591
rect 703501 394535 703587 394591
rect 703643 394535 703729 394591
rect 703785 394535 703871 394591
rect 703927 394535 704013 394591
rect 704069 394535 704155 394591
rect 704211 394535 704297 394591
rect 704353 394555 705525 394591
rect 705581 394555 705649 394611
rect 705705 394555 705773 394611
rect 705829 394555 705897 394611
rect 705953 394555 706000 394611
rect 704353 394535 706000 394555
rect 702392 394487 706000 394535
rect 702392 394449 705525 394487
rect 702392 394393 702451 394449
rect 702507 394393 702593 394449
rect 702649 394393 702735 394449
rect 702791 394393 702877 394449
rect 702933 394393 703019 394449
rect 703075 394393 703161 394449
rect 703217 394393 703303 394449
rect 703359 394393 703445 394449
rect 703501 394393 703587 394449
rect 703643 394393 703729 394449
rect 703785 394393 703871 394449
rect 703927 394393 704013 394449
rect 704069 394393 704155 394449
rect 704211 394393 704297 394449
rect 704353 394431 705525 394449
rect 705581 394431 705649 394487
rect 705705 394431 705773 394487
rect 705829 394431 705897 394487
rect 705953 394431 706000 394487
rect 704353 394393 706000 394431
rect 702392 394363 706000 394393
rect 702392 394307 705525 394363
rect 705581 394307 705649 394363
rect 705705 394307 705773 394363
rect 705829 394307 705897 394363
rect 705953 394307 706000 394363
rect 702392 394251 702451 394307
rect 702507 394251 702593 394307
rect 702649 394251 702735 394307
rect 702791 394251 702877 394307
rect 702933 394251 703019 394307
rect 703075 394251 703161 394307
rect 703217 394251 703303 394307
rect 703359 394251 703445 394307
rect 703501 394251 703587 394307
rect 703643 394251 703729 394307
rect 703785 394251 703871 394307
rect 703927 394251 704013 394307
rect 704069 394251 704155 394307
rect 704211 394251 704297 394307
rect 704353 394251 706000 394307
rect 702392 394239 706000 394251
rect 702392 394183 705525 394239
rect 705581 394183 705649 394239
rect 705705 394183 705773 394239
rect 705829 394183 705897 394239
rect 705953 394183 706000 394239
rect 702392 394165 706000 394183
rect 702392 394109 702451 394165
rect 702507 394109 702593 394165
rect 702649 394109 702735 394165
rect 702791 394109 702877 394165
rect 702933 394109 703019 394165
rect 703075 394109 703161 394165
rect 703217 394109 703303 394165
rect 703359 394109 703445 394165
rect 703501 394109 703587 394165
rect 703643 394109 703729 394165
rect 703785 394109 703871 394165
rect 703927 394109 704013 394165
rect 704069 394109 704155 394165
rect 704211 394109 704297 394165
rect 704353 394115 706000 394165
rect 704353 394109 705525 394115
rect 702392 394059 705525 394109
rect 705581 394059 705649 394115
rect 705705 394059 705773 394115
rect 705829 394059 705897 394115
rect 705953 394059 706000 394115
rect 702392 394023 706000 394059
rect 702392 393967 702451 394023
rect 702507 393967 702593 394023
rect 702649 393967 702735 394023
rect 702791 393967 702877 394023
rect 702933 393967 703019 394023
rect 703075 393967 703161 394023
rect 703217 393967 703303 394023
rect 703359 393967 703445 394023
rect 703501 393967 703587 394023
rect 703643 393967 703729 394023
rect 703785 393967 703871 394023
rect 703927 393967 704013 394023
rect 704069 393967 704155 394023
rect 704211 393967 704297 394023
rect 704353 393991 706000 394023
rect 704353 393967 705525 393991
rect 702392 393935 705525 393967
rect 705581 393935 705649 393991
rect 705705 393935 705773 393991
rect 705829 393935 705897 393991
rect 705953 393935 706000 393991
rect 702392 393881 706000 393935
rect 702392 393825 702451 393881
rect 702507 393825 702593 393881
rect 702649 393825 702735 393881
rect 702791 393825 702877 393881
rect 702933 393825 703019 393881
rect 703075 393825 703161 393881
rect 703217 393825 703303 393881
rect 703359 393825 703445 393881
rect 703501 393825 703587 393881
rect 703643 393825 703729 393881
rect 703785 393825 703871 393881
rect 703927 393825 704013 393881
rect 704069 393825 704155 393881
rect 704211 393825 704297 393881
rect 704353 393867 706000 393881
rect 704353 393825 705525 393867
rect 702392 393811 705525 393825
rect 705581 393811 705649 393867
rect 705705 393811 705773 393867
rect 705829 393811 705897 393867
rect 705953 393811 706000 393867
rect 702392 393743 706000 393811
rect 702392 393739 705525 393743
rect 702392 393683 702451 393739
rect 702507 393683 702593 393739
rect 702649 393683 702735 393739
rect 702791 393683 702877 393739
rect 702933 393683 703019 393739
rect 703075 393683 703161 393739
rect 703217 393683 703303 393739
rect 703359 393683 703445 393739
rect 703501 393683 703587 393739
rect 703643 393683 703729 393739
rect 703785 393683 703871 393739
rect 703927 393683 704013 393739
rect 704069 393683 704155 393739
rect 704211 393683 704297 393739
rect 704353 393687 705525 393739
rect 705581 393687 705649 393743
rect 705705 393687 705773 393743
rect 705829 393687 705897 393743
rect 705953 393687 706000 393743
rect 704353 393683 706000 393687
rect 702392 393619 706000 393683
rect 702392 393597 705525 393619
rect 702392 393541 702451 393597
rect 702507 393541 702593 393597
rect 702649 393541 702735 393597
rect 702791 393541 702877 393597
rect 702933 393541 703019 393597
rect 703075 393541 703161 393597
rect 703217 393541 703303 393597
rect 703359 393541 703445 393597
rect 703501 393541 703587 393597
rect 703643 393541 703729 393597
rect 703785 393541 703871 393597
rect 703927 393541 704013 393597
rect 704069 393541 704155 393597
rect 704211 393541 704297 393597
rect 704353 393563 705525 393597
rect 705581 393563 705649 393619
rect 705705 393563 705773 393619
rect 705829 393563 705897 393619
rect 705953 393563 706000 393619
rect 704353 393541 706000 393563
rect 702392 393495 706000 393541
rect 702392 393455 705525 393495
rect 702392 393399 702451 393455
rect 702507 393399 702593 393455
rect 702649 393399 702735 393455
rect 702791 393399 702877 393455
rect 702933 393399 703019 393455
rect 703075 393399 703161 393455
rect 703217 393399 703303 393455
rect 703359 393399 703445 393455
rect 703501 393399 703587 393455
rect 703643 393399 703729 393455
rect 703785 393399 703871 393455
rect 703927 393399 704013 393455
rect 704069 393399 704155 393455
rect 704211 393399 704297 393455
rect 704353 393439 705525 393455
rect 705581 393439 705649 393495
rect 705705 393439 705773 393495
rect 705829 393439 705897 393495
rect 705953 393439 706000 393495
rect 704353 393399 706000 393439
rect 702392 393371 706000 393399
rect 702392 393315 705525 393371
rect 705581 393315 705649 393371
rect 705705 393315 705773 393371
rect 705829 393315 705897 393371
rect 705953 393315 706000 393371
rect 702392 393313 706000 393315
rect 702392 393257 702451 393313
rect 702507 393257 702593 393313
rect 702649 393257 702735 393313
rect 702791 393257 702877 393313
rect 702933 393257 703019 393313
rect 703075 393257 703161 393313
rect 703217 393257 703303 393313
rect 703359 393257 703445 393313
rect 703501 393257 703587 393313
rect 703643 393257 703729 393313
rect 703785 393257 703871 393313
rect 703927 393257 704013 393313
rect 704069 393257 704155 393313
rect 704211 393257 704297 393313
rect 704353 393257 706000 393313
rect 702392 393247 706000 393257
rect 702392 393191 705525 393247
rect 705581 393191 705649 393247
rect 705705 393191 705773 393247
rect 705829 393191 705897 393247
rect 705953 393191 706000 393247
rect 702392 393171 706000 393191
rect 702392 393115 702451 393171
rect 702507 393115 702593 393171
rect 702649 393115 702735 393171
rect 702791 393115 702877 393171
rect 702933 393115 703019 393171
rect 703075 393115 703161 393171
rect 703217 393115 703303 393171
rect 703359 393115 703445 393171
rect 703501 393115 703587 393171
rect 703643 393115 703729 393171
rect 703785 393115 703871 393171
rect 703927 393115 704013 393171
rect 704069 393115 704155 393171
rect 704211 393115 704297 393171
rect 704353 393123 706000 393171
rect 704353 393115 705525 393123
rect 702392 393067 705525 393115
rect 705581 393067 705649 393123
rect 705705 393067 705773 393123
rect 705829 393067 705897 393123
rect 705953 393067 706000 393123
rect 702392 393029 706000 393067
rect 702392 392973 702451 393029
rect 702507 392973 702593 393029
rect 702649 392973 702735 393029
rect 702791 392973 702877 393029
rect 702933 392973 703019 393029
rect 703075 392973 703161 393029
rect 703217 392973 703303 393029
rect 703359 392973 703445 393029
rect 703501 392973 703587 393029
rect 703643 392973 703729 393029
rect 703785 392973 703871 393029
rect 703927 392973 704013 393029
rect 704069 392973 704155 393029
rect 704211 392973 704297 393029
rect 704353 392999 706000 393029
rect 704353 392973 705525 392999
rect 702392 392943 705525 392973
rect 705581 392943 705649 392999
rect 705705 392943 705773 392999
rect 705829 392943 705897 392999
rect 705953 392943 706000 392999
rect 702392 392887 706000 392943
rect 702392 392831 702451 392887
rect 702507 392831 702593 392887
rect 702649 392831 702735 392887
rect 702791 392831 702877 392887
rect 702933 392831 703019 392887
rect 703075 392831 703161 392887
rect 703217 392831 703303 392887
rect 703359 392831 703445 392887
rect 703501 392831 703587 392887
rect 703643 392831 703729 392887
rect 703785 392831 703871 392887
rect 703927 392831 704013 392887
rect 704069 392831 704155 392887
rect 704211 392831 704297 392887
rect 704353 392875 706000 392887
rect 704353 392831 705525 392875
rect 702392 392819 705525 392831
rect 705581 392819 705649 392875
rect 705705 392819 705773 392875
rect 705829 392819 705897 392875
rect 705953 392819 706000 392875
rect 702392 392752 706000 392819
rect 702392 392131 706000 392172
rect 702392 392110 705525 392131
rect 702392 392054 702440 392110
rect 702496 392054 702582 392110
rect 702638 392054 702724 392110
rect 702780 392054 702866 392110
rect 702922 392054 703008 392110
rect 703064 392054 703150 392110
rect 703206 392054 703292 392110
rect 703348 392054 703434 392110
rect 703490 392054 703576 392110
rect 703632 392054 703718 392110
rect 703774 392054 703860 392110
rect 703916 392054 704002 392110
rect 704058 392054 704144 392110
rect 704200 392054 704286 392110
rect 704342 392075 705525 392110
rect 705581 392075 705649 392131
rect 705705 392075 705773 392131
rect 705829 392075 705897 392131
rect 705953 392075 706000 392131
rect 704342 392054 706000 392075
rect 702392 392007 706000 392054
rect 702392 391968 705525 392007
rect 702392 391912 702440 391968
rect 702496 391912 702582 391968
rect 702638 391912 702724 391968
rect 702780 391912 702866 391968
rect 702922 391912 703008 391968
rect 703064 391912 703150 391968
rect 703206 391912 703292 391968
rect 703348 391912 703434 391968
rect 703490 391912 703576 391968
rect 703632 391912 703718 391968
rect 703774 391912 703860 391968
rect 703916 391912 704002 391968
rect 704058 391912 704144 391968
rect 704200 391912 704286 391968
rect 704342 391951 705525 391968
rect 705581 391951 705649 392007
rect 705705 391951 705773 392007
rect 705829 391951 705897 392007
rect 705953 391951 706000 392007
rect 704342 391912 706000 391951
rect 702392 391883 706000 391912
rect 702392 391827 705525 391883
rect 705581 391827 705649 391883
rect 705705 391827 705773 391883
rect 705829 391827 705897 391883
rect 705953 391827 706000 391883
rect 702392 391826 706000 391827
rect 702392 391770 702440 391826
rect 702496 391770 702582 391826
rect 702638 391770 702724 391826
rect 702780 391770 702866 391826
rect 702922 391770 703008 391826
rect 703064 391770 703150 391826
rect 703206 391770 703292 391826
rect 703348 391770 703434 391826
rect 703490 391770 703576 391826
rect 703632 391770 703718 391826
rect 703774 391770 703860 391826
rect 703916 391770 704002 391826
rect 704058 391770 704144 391826
rect 704200 391770 704286 391826
rect 704342 391770 706000 391826
rect 702392 391759 706000 391770
rect 702392 391703 705525 391759
rect 705581 391703 705649 391759
rect 705705 391703 705773 391759
rect 705829 391703 705897 391759
rect 705953 391703 706000 391759
rect 702392 391684 706000 391703
rect 702392 391628 702440 391684
rect 702496 391628 702582 391684
rect 702638 391628 702724 391684
rect 702780 391628 702866 391684
rect 702922 391628 703008 391684
rect 703064 391628 703150 391684
rect 703206 391628 703292 391684
rect 703348 391628 703434 391684
rect 703490 391628 703576 391684
rect 703632 391628 703718 391684
rect 703774 391628 703860 391684
rect 703916 391628 704002 391684
rect 704058 391628 704144 391684
rect 704200 391628 704286 391684
rect 704342 391635 706000 391684
rect 704342 391628 705525 391635
rect 702392 391579 705525 391628
rect 705581 391579 705649 391635
rect 705705 391579 705773 391635
rect 705829 391579 705897 391635
rect 705953 391579 706000 391635
rect 702392 391542 706000 391579
rect 702392 391486 702440 391542
rect 702496 391486 702582 391542
rect 702638 391486 702724 391542
rect 702780 391486 702866 391542
rect 702922 391486 703008 391542
rect 703064 391486 703150 391542
rect 703206 391486 703292 391542
rect 703348 391486 703434 391542
rect 703490 391486 703576 391542
rect 703632 391486 703718 391542
rect 703774 391486 703860 391542
rect 703916 391486 704002 391542
rect 704058 391486 704144 391542
rect 704200 391486 704286 391542
rect 704342 391511 706000 391542
rect 704342 391486 705525 391511
rect 702392 391455 705525 391486
rect 705581 391455 705649 391511
rect 705705 391455 705773 391511
rect 705829 391455 705897 391511
rect 705953 391455 706000 391511
rect 702392 391400 706000 391455
rect 702392 391344 702440 391400
rect 702496 391344 702582 391400
rect 702638 391344 702724 391400
rect 702780 391344 702866 391400
rect 702922 391344 703008 391400
rect 703064 391344 703150 391400
rect 703206 391344 703292 391400
rect 703348 391344 703434 391400
rect 703490 391344 703576 391400
rect 703632 391344 703718 391400
rect 703774 391344 703860 391400
rect 703916 391344 704002 391400
rect 704058 391344 704144 391400
rect 704200 391344 704286 391400
rect 704342 391387 706000 391400
rect 704342 391344 705525 391387
rect 702392 391331 705525 391344
rect 705581 391331 705649 391387
rect 705705 391331 705773 391387
rect 705829 391331 705897 391387
rect 705953 391331 706000 391387
rect 702392 391263 706000 391331
rect 702392 391258 705525 391263
rect 702392 391202 702440 391258
rect 702496 391202 702582 391258
rect 702638 391202 702724 391258
rect 702780 391202 702866 391258
rect 702922 391202 703008 391258
rect 703064 391202 703150 391258
rect 703206 391202 703292 391258
rect 703348 391202 703434 391258
rect 703490 391202 703576 391258
rect 703632 391202 703718 391258
rect 703774 391202 703860 391258
rect 703916 391202 704002 391258
rect 704058 391202 704144 391258
rect 704200 391202 704286 391258
rect 704342 391207 705525 391258
rect 705581 391207 705649 391263
rect 705705 391207 705773 391263
rect 705829 391207 705897 391263
rect 705953 391207 706000 391263
rect 704342 391202 706000 391207
rect 702392 391139 706000 391202
rect 702392 391116 705525 391139
rect 702392 391060 702440 391116
rect 702496 391060 702582 391116
rect 702638 391060 702724 391116
rect 702780 391060 702866 391116
rect 702922 391060 703008 391116
rect 703064 391060 703150 391116
rect 703206 391060 703292 391116
rect 703348 391060 703434 391116
rect 703490 391060 703576 391116
rect 703632 391060 703718 391116
rect 703774 391060 703860 391116
rect 703916 391060 704002 391116
rect 704058 391060 704144 391116
rect 704200 391060 704286 391116
rect 704342 391083 705525 391116
rect 705581 391083 705649 391139
rect 705705 391083 705773 391139
rect 705829 391083 705897 391139
rect 705953 391083 706000 391139
rect 704342 391060 706000 391083
rect 702392 391015 706000 391060
rect 702392 390974 705525 391015
rect 702392 390918 702440 390974
rect 702496 390918 702582 390974
rect 702638 390918 702724 390974
rect 702780 390918 702866 390974
rect 702922 390918 703008 390974
rect 703064 390918 703150 390974
rect 703206 390918 703292 390974
rect 703348 390918 703434 390974
rect 703490 390918 703576 390974
rect 703632 390918 703718 390974
rect 703774 390918 703860 390974
rect 703916 390918 704002 390974
rect 704058 390918 704144 390974
rect 704200 390918 704286 390974
rect 704342 390959 705525 390974
rect 705581 390959 705649 391015
rect 705705 390959 705773 391015
rect 705829 390959 705897 391015
rect 705953 390959 706000 391015
rect 704342 390918 706000 390959
rect 702392 390891 706000 390918
rect 702392 390835 705525 390891
rect 705581 390835 705649 390891
rect 705705 390835 705773 390891
rect 705829 390835 705897 390891
rect 705953 390835 706000 390891
rect 702392 390832 706000 390835
rect 702392 390776 702440 390832
rect 702496 390776 702582 390832
rect 702638 390776 702724 390832
rect 702780 390776 702866 390832
rect 702922 390776 703008 390832
rect 703064 390776 703150 390832
rect 703206 390776 703292 390832
rect 703348 390776 703434 390832
rect 703490 390776 703576 390832
rect 703632 390776 703718 390832
rect 703774 390776 703860 390832
rect 703916 390776 704002 390832
rect 704058 390776 704144 390832
rect 704200 390776 704286 390832
rect 704342 390776 706000 390832
rect 702392 390767 706000 390776
rect 702392 390711 705525 390767
rect 705581 390711 705649 390767
rect 705705 390711 705773 390767
rect 705829 390711 705897 390767
rect 705953 390711 706000 390767
rect 702392 390690 706000 390711
rect 702392 390634 702440 390690
rect 702496 390634 702582 390690
rect 702638 390634 702724 390690
rect 702780 390634 702866 390690
rect 702922 390634 703008 390690
rect 703064 390634 703150 390690
rect 703206 390634 703292 390690
rect 703348 390634 703434 390690
rect 703490 390634 703576 390690
rect 703632 390634 703718 390690
rect 703774 390634 703860 390690
rect 703916 390634 704002 390690
rect 704058 390634 704144 390690
rect 704200 390634 704286 390690
rect 704342 390643 706000 390690
rect 704342 390634 705525 390643
rect 702392 390587 705525 390634
rect 705581 390587 705649 390643
rect 705705 390587 705773 390643
rect 705829 390587 705897 390643
rect 705953 390587 706000 390643
rect 702392 390548 706000 390587
rect 702392 390492 702440 390548
rect 702496 390492 702582 390548
rect 702638 390492 702724 390548
rect 702780 390492 702866 390548
rect 702922 390492 703008 390548
rect 703064 390492 703150 390548
rect 703206 390492 703292 390548
rect 703348 390492 703434 390548
rect 703490 390492 703576 390548
rect 703632 390492 703718 390548
rect 703774 390492 703860 390548
rect 703916 390492 704002 390548
rect 704058 390492 704144 390548
rect 704200 390492 704286 390548
rect 704342 390519 706000 390548
rect 704342 390492 705525 390519
rect 702392 390463 705525 390492
rect 705581 390463 705649 390519
rect 705705 390463 705773 390519
rect 705829 390463 705897 390519
rect 705953 390463 706000 390519
rect 702392 390406 706000 390463
rect 702392 390350 702440 390406
rect 702496 390350 702582 390406
rect 702638 390350 702724 390406
rect 702780 390350 702866 390406
rect 702922 390350 703008 390406
rect 703064 390350 703150 390406
rect 703206 390350 703292 390406
rect 703348 390350 703434 390406
rect 703490 390350 703576 390406
rect 703632 390350 703718 390406
rect 703774 390350 703860 390406
rect 703916 390350 704002 390406
rect 704058 390350 704144 390406
rect 704200 390350 704286 390406
rect 704342 390395 706000 390406
rect 704342 390350 705525 390395
rect 702392 390339 705525 390350
rect 705581 390339 705649 390395
rect 705705 390339 705773 390395
rect 705829 390339 705897 390395
rect 705953 390339 706000 390395
rect 702392 390272 706000 390339
rect 70000 140661 75416 140728
rect 70000 140605 70047 140661
rect 70103 140605 70171 140661
rect 70227 140605 70295 140661
rect 70351 140605 70419 140661
rect 70475 140650 75416 140661
rect 70475 140605 73866 140650
rect 70000 140594 73866 140605
rect 73922 140594 74008 140650
rect 74064 140594 74150 140650
rect 74206 140594 74292 140650
rect 74348 140594 74434 140650
rect 74490 140594 74576 140650
rect 74632 140594 74718 140650
rect 74774 140594 74860 140650
rect 74916 140594 75002 140650
rect 75058 140594 75144 140650
rect 75200 140594 75286 140650
rect 75342 140594 75416 140650
rect 70000 140537 75416 140594
rect 70000 140481 70047 140537
rect 70103 140481 70171 140537
rect 70227 140481 70295 140537
rect 70351 140481 70419 140537
rect 70475 140508 75416 140537
rect 70475 140481 73866 140508
rect 70000 140452 73866 140481
rect 73922 140452 74008 140508
rect 74064 140452 74150 140508
rect 74206 140452 74292 140508
rect 74348 140452 74434 140508
rect 74490 140452 74576 140508
rect 74632 140452 74718 140508
rect 74774 140452 74860 140508
rect 74916 140452 75002 140508
rect 75058 140452 75144 140508
rect 75200 140452 75286 140508
rect 75342 140452 75416 140508
rect 70000 140413 75416 140452
rect 70000 140357 70047 140413
rect 70103 140357 70171 140413
rect 70227 140357 70295 140413
rect 70351 140357 70419 140413
rect 70475 140366 75416 140413
rect 70475 140357 73866 140366
rect 70000 140310 73866 140357
rect 73922 140310 74008 140366
rect 74064 140310 74150 140366
rect 74206 140310 74292 140366
rect 74348 140310 74434 140366
rect 74490 140310 74576 140366
rect 74632 140310 74718 140366
rect 74774 140310 74860 140366
rect 74916 140310 75002 140366
rect 75058 140310 75144 140366
rect 75200 140310 75286 140366
rect 75342 140310 75416 140366
rect 70000 140289 75416 140310
rect 70000 140233 70047 140289
rect 70103 140233 70171 140289
rect 70227 140233 70295 140289
rect 70351 140233 70419 140289
rect 70475 140233 75416 140289
rect 70000 140224 75416 140233
rect 70000 140168 73866 140224
rect 73922 140168 74008 140224
rect 74064 140168 74150 140224
rect 74206 140168 74292 140224
rect 74348 140168 74434 140224
rect 74490 140168 74576 140224
rect 74632 140168 74718 140224
rect 74774 140168 74860 140224
rect 74916 140168 75002 140224
rect 75058 140168 75144 140224
rect 75200 140168 75286 140224
rect 75342 140168 75416 140224
rect 70000 140165 75416 140168
rect 70000 140109 70047 140165
rect 70103 140109 70171 140165
rect 70227 140109 70295 140165
rect 70351 140109 70419 140165
rect 70475 140109 75416 140165
rect 70000 140082 75416 140109
rect 70000 140041 73866 140082
rect 70000 139985 70047 140041
rect 70103 139985 70171 140041
rect 70227 139985 70295 140041
rect 70351 139985 70419 140041
rect 70475 140026 73866 140041
rect 73922 140026 74008 140082
rect 74064 140026 74150 140082
rect 74206 140026 74292 140082
rect 74348 140026 74434 140082
rect 74490 140026 74576 140082
rect 74632 140026 74718 140082
rect 74774 140026 74860 140082
rect 74916 140026 75002 140082
rect 75058 140026 75144 140082
rect 75200 140026 75286 140082
rect 75342 140026 75416 140082
rect 70475 139985 75416 140026
rect 70000 139940 75416 139985
rect 70000 139917 73866 139940
rect 70000 139861 70047 139917
rect 70103 139861 70171 139917
rect 70227 139861 70295 139917
rect 70351 139861 70419 139917
rect 70475 139884 73866 139917
rect 73922 139884 74008 139940
rect 74064 139884 74150 139940
rect 74206 139884 74292 139940
rect 74348 139884 74434 139940
rect 74490 139884 74576 139940
rect 74632 139884 74718 139940
rect 74774 139884 74860 139940
rect 74916 139884 75002 139940
rect 75058 139884 75144 139940
rect 75200 139884 75286 139940
rect 75342 139884 75416 139940
rect 70475 139861 75416 139884
rect 70000 139798 75416 139861
rect 70000 139793 73866 139798
rect 70000 139737 70047 139793
rect 70103 139737 70171 139793
rect 70227 139737 70295 139793
rect 70351 139737 70419 139793
rect 70475 139742 73866 139793
rect 73922 139742 74008 139798
rect 74064 139742 74150 139798
rect 74206 139742 74292 139798
rect 74348 139742 74434 139798
rect 74490 139742 74576 139798
rect 74632 139742 74718 139798
rect 74774 139742 74860 139798
rect 74916 139742 75002 139798
rect 75058 139742 75144 139798
rect 75200 139742 75286 139798
rect 75342 139742 75416 139798
rect 70475 139737 75416 139742
rect 70000 139669 75416 139737
rect 70000 139613 70047 139669
rect 70103 139613 70171 139669
rect 70227 139613 70295 139669
rect 70351 139613 70419 139669
rect 70475 139656 75416 139669
rect 70475 139613 73866 139656
rect 70000 139600 73866 139613
rect 73922 139600 74008 139656
rect 74064 139600 74150 139656
rect 74206 139600 74292 139656
rect 74348 139600 74434 139656
rect 74490 139600 74576 139656
rect 74632 139600 74718 139656
rect 74774 139600 74860 139656
rect 74916 139600 75002 139656
rect 75058 139600 75144 139656
rect 75200 139600 75286 139656
rect 75342 139600 75416 139656
rect 70000 139545 75416 139600
rect 70000 139489 70047 139545
rect 70103 139489 70171 139545
rect 70227 139489 70295 139545
rect 70351 139489 70419 139545
rect 70475 139514 75416 139545
rect 70475 139489 73866 139514
rect 70000 139458 73866 139489
rect 73922 139458 74008 139514
rect 74064 139458 74150 139514
rect 74206 139458 74292 139514
rect 74348 139458 74434 139514
rect 74490 139458 74576 139514
rect 74632 139458 74718 139514
rect 74774 139458 74860 139514
rect 74916 139458 75002 139514
rect 75058 139458 75144 139514
rect 75200 139458 75286 139514
rect 75342 139458 75416 139514
rect 70000 139421 75416 139458
rect 70000 139365 70047 139421
rect 70103 139365 70171 139421
rect 70227 139365 70295 139421
rect 70351 139365 70419 139421
rect 70475 139372 75416 139421
rect 70475 139365 73866 139372
rect 70000 139316 73866 139365
rect 73922 139316 74008 139372
rect 74064 139316 74150 139372
rect 74206 139316 74292 139372
rect 74348 139316 74434 139372
rect 74490 139316 74576 139372
rect 74632 139316 74718 139372
rect 74774 139316 74860 139372
rect 74916 139316 75002 139372
rect 75058 139316 75144 139372
rect 75200 139316 75286 139372
rect 75342 139316 75416 139372
rect 70000 139297 75416 139316
rect 70000 139241 70047 139297
rect 70103 139241 70171 139297
rect 70227 139241 70295 139297
rect 70351 139241 70419 139297
rect 70475 139241 75416 139297
rect 70000 139230 75416 139241
rect 70000 139174 73866 139230
rect 73922 139174 74008 139230
rect 74064 139174 74150 139230
rect 74206 139174 74292 139230
rect 74348 139174 74434 139230
rect 74490 139174 74576 139230
rect 74632 139174 74718 139230
rect 74774 139174 74860 139230
rect 74916 139174 75002 139230
rect 75058 139174 75144 139230
rect 75200 139174 75286 139230
rect 75342 139174 75416 139230
rect 70000 139173 75416 139174
rect 70000 139117 70047 139173
rect 70103 139117 70171 139173
rect 70227 139117 70295 139173
rect 70351 139117 70419 139173
rect 70475 139117 75416 139173
rect 70000 139088 75416 139117
rect 70000 139049 73866 139088
rect 70000 138993 70047 139049
rect 70103 138993 70171 139049
rect 70227 138993 70295 139049
rect 70351 138993 70419 139049
rect 70475 139032 73866 139049
rect 73922 139032 74008 139088
rect 74064 139032 74150 139088
rect 74206 139032 74292 139088
rect 74348 139032 74434 139088
rect 74490 139032 74576 139088
rect 74632 139032 74718 139088
rect 74774 139032 74860 139088
rect 74916 139032 75002 139088
rect 75058 139032 75144 139088
rect 75200 139032 75286 139088
rect 75342 139032 75416 139088
rect 70475 138993 75416 139032
rect 70000 138946 75416 138993
rect 70000 138925 73866 138946
rect 70000 138869 70047 138925
rect 70103 138869 70171 138925
rect 70227 138869 70295 138925
rect 70351 138869 70419 138925
rect 70475 138890 73866 138925
rect 73922 138890 74008 138946
rect 74064 138890 74150 138946
rect 74206 138890 74292 138946
rect 74348 138890 74434 138946
rect 74490 138890 74576 138946
rect 74632 138890 74718 138946
rect 74774 138890 74860 138946
rect 74916 138890 75002 138946
rect 75058 138890 75144 138946
rect 75200 138890 75286 138946
rect 75342 138890 75416 138946
rect 70475 138869 75416 138890
rect 70000 138828 75416 138869
rect 70000 138181 75416 138248
rect 70000 138125 70047 138181
rect 70103 138125 70171 138181
rect 70227 138125 70295 138181
rect 70351 138125 70419 138181
rect 70475 138169 75416 138181
rect 70475 138125 73855 138169
rect 70000 138113 73855 138125
rect 73911 138113 73997 138169
rect 74053 138113 74139 138169
rect 74195 138113 74281 138169
rect 74337 138113 74423 138169
rect 74479 138113 74565 138169
rect 74621 138113 74707 138169
rect 74763 138113 74849 138169
rect 74905 138113 74991 138169
rect 75047 138113 75133 138169
rect 75189 138113 75275 138169
rect 75331 138113 75416 138169
rect 70000 138057 75416 138113
rect 70000 138001 70047 138057
rect 70103 138001 70171 138057
rect 70227 138001 70295 138057
rect 70351 138001 70419 138057
rect 70475 138027 75416 138057
rect 70475 138001 73855 138027
rect 70000 137971 73855 138001
rect 73911 137971 73997 138027
rect 74053 137971 74139 138027
rect 74195 137971 74281 138027
rect 74337 137971 74423 138027
rect 74479 137971 74565 138027
rect 74621 137971 74707 138027
rect 74763 137971 74849 138027
rect 74905 137971 74991 138027
rect 75047 137971 75133 138027
rect 75189 137971 75275 138027
rect 75331 137971 75416 138027
rect 70000 137933 75416 137971
rect 70000 137877 70047 137933
rect 70103 137877 70171 137933
rect 70227 137877 70295 137933
rect 70351 137877 70419 137933
rect 70475 137885 75416 137933
rect 70475 137877 73855 137885
rect 70000 137829 73855 137877
rect 73911 137829 73997 137885
rect 74053 137829 74139 137885
rect 74195 137829 74281 137885
rect 74337 137829 74423 137885
rect 74479 137829 74565 137885
rect 74621 137829 74707 137885
rect 74763 137829 74849 137885
rect 74905 137829 74991 137885
rect 75047 137829 75133 137885
rect 75189 137829 75275 137885
rect 75331 137829 75416 137885
rect 70000 137809 75416 137829
rect 70000 137753 70047 137809
rect 70103 137753 70171 137809
rect 70227 137753 70295 137809
rect 70351 137753 70419 137809
rect 70475 137753 75416 137809
rect 70000 137743 75416 137753
rect 70000 137687 73855 137743
rect 73911 137687 73997 137743
rect 74053 137687 74139 137743
rect 74195 137687 74281 137743
rect 74337 137687 74423 137743
rect 74479 137687 74565 137743
rect 74621 137687 74707 137743
rect 74763 137687 74849 137743
rect 74905 137687 74991 137743
rect 75047 137687 75133 137743
rect 75189 137687 75275 137743
rect 75331 137687 75416 137743
rect 70000 137685 75416 137687
rect 70000 137629 70047 137685
rect 70103 137629 70171 137685
rect 70227 137629 70295 137685
rect 70351 137629 70419 137685
rect 70475 137629 75416 137685
rect 70000 137601 75416 137629
rect 70000 137561 73855 137601
rect 70000 137505 70047 137561
rect 70103 137505 70171 137561
rect 70227 137505 70295 137561
rect 70351 137505 70419 137561
rect 70475 137545 73855 137561
rect 73911 137545 73997 137601
rect 74053 137545 74139 137601
rect 74195 137545 74281 137601
rect 74337 137545 74423 137601
rect 74479 137545 74565 137601
rect 74621 137545 74707 137601
rect 74763 137545 74849 137601
rect 74905 137545 74991 137601
rect 75047 137545 75133 137601
rect 75189 137545 75275 137601
rect 75331 137545 75416 137601
rect 70475 137505 75416 137545
rect 70000 137459 75416 137505
rect 70000 137437 73855 137459
rect 70000 137381 70047 137437
rect 70103 137381 70171 137437
rect 70227 137381 70295 137437
rect 70351 137381 70419 137437
rect 70475 137403 73855 137437
rect 73911 137403 73997 137459
rect 74053 137403 74139 137459
rect 74195 137403 74281 137459
rect 74337 137403 74423 137459
rect 74479 137403 74565 137459
rect 74621 137403 74707 137459
rect 74763 137403 74849 137459
rect 74905 137403 74991 137459
rect 75047 137403 75133 137459
rect 75189 137403 75275 137459
rect 75331 137403 75416 137459
rect 70475 137381 75416 137403
rect 70000 137317 75416 137381
rect 70000 137313 73855 137317
rect 70000 137257 70047 137313
rect 70103 137257 70171 137313
rect 70227 137257 70295 137313
rect 70351 137257 70419 137313
rect 70475 137261 73855 137313
rect 73911 137261 73997 137317
rect 74053 137261 74139 137317
rect 74195 137261 74281 137317
rect 74337 137261 74423 137317
rect 74479 137261 74565 137317
rect 74621 137261 74707 137317
rect 74763 137261 74849 137317
rect 74905 137261 74991 137317
rect 75047 137261 75133 137317
rect 75189 137261 75275 137317
rect 75331 137261 75416 137317
rect 70475 137257 75416 137261
rect 70000 137189 75416 137257
rect 70000 137133 70047 137189
rect 70103 137133 70171 137189
rect 70227 137133 70295 137189
rect 70351 137133 70419 137189
rect 70475 137175 75416 137189
rect 70475 137133 73855 137175
rect 70000 137119 73855 137133
rect 73911 137119 73997 137175
rect 74053 137119 74139 137175
rect 74195 137119 74281 137175
rect 74337 137119 74423 137175
rect 74479 137119 74565 137175
rect 74621 137119 74707 137175
rect 74763 137119 74849 137175
rect 74905 137119 74991 137175
rect 75047 137119 75133 137175
rect 75189 137119 75275 137175
rect 75331 137119 75416 137175
rect 70000 137065 75416 137119
rect 70000 137009 70047 137065
rect 70103 137009 70171 137065
rect 70227 137009 70295 137065
rect 70351 137009 70419 137065
rect 70475 137033 75416 137065
rect 70475 137009 73855 137033
rect 70000 136977 73855 137009
rect 73911 136977 73997 137033
rect 74053 136977 74139 137033
rect 74195 136977 74281 137033
rect 74337 136977 74423 137033
rect 74479 136977 74565 137033
rect 74621 136977 74707 137033
rect 74763 136977 74849 137033
rect 74905 136977 74991 137033
rect 75047 136977 75133 137033
rect 75189 136977 75275 137033
rect 75331 136977 75416 137033
rect 70000 136941 75416 136977
rect 70000 136885 70047 136941
rect 70103 136885 70171 136941
rect 70227 136885 70295 136941
rect 70351 136885 70419 136941
rect 70475 136891 75416 136941
rect 70475 136885 73855 136891
rect 70000 136835 73855 136885
rect 73911 136835 73997 136891
rect 74053 136835 74139 136891
rect 74195 136835 74281 136891
rect 74337 136835 74423 136891
rect 74479 136835 74565 136891
rect 74621 136835 74707 136891
rect 74763 136835 74849 136891
rect 74905 136835 74991 136891
rect 75047 136835 75133 136891
rect 75189 136835 75275 136891
rect 75331 136835 75416 136891
rect 70000 136817 75416 136835
rect 70000 136761 70047 136817
rect 70103 136761 70171 136817
rect 70227 136761 70295 136817
rect 70351 136761 70419 136817
rect 70475 136761 75416 136817
rect 70000 136749 75416 136761
rect 70000 136693 73855 136749
rect 73911 136693 73997 136749
rect 74053 136693 74139 136749
rect 74195 136693 74281 136749
rect 74337 136693 74423 136749
rect 74479 136693 74565 136749
rect 74621 136693 74707 136749
rect 74763 136693 74849 136749
rect 74905 136693 74991 136749
rect 75047 136693 75133 136749
rect 75189 136693 75275 136749
rect 75331 136693 75416 136749
rect 70000 136637 70047 136693
rect 70103 136637 70171 136693
rect 70227 136637 70295 136693
rect 70351 136637 70419 136693
rect 70475 136637 75416 136693
rect 70000 136607 75416 136637
rect 70000 136569 73855 136607
rect 70000 136513 70047 136569
rect 70103 136513 70171 136569
rect 70227 136513 70295 136569
rect 70351 136513 70419 136569
rect 70475 136551 73855 136569
rect 73911 136551 73997 136607
rect 74053 136551 74139 136607
rect 74195 136551 74281 136607
rect 74337 136551 74423 136607
rect 74479 136551 74565 136607
rect 74621 136551 74707 136607
rect 74763 136551 74849 136607
rect 74905 136551 74991 136607
rect 75047 136551 75133 136607
rect 75189 136551 75275 136607
rect 75331 136551 75416 136607
rect 70475 136513 75416 136551
rect 70000 136465 75416 136513
rect 70000 136445 73855 136465
rect 70000 136389 70047 136445
rect 70103 136389 70171 136445
rect 70227 136389 70295 136445
rect 70351 136389 70419 136445
rect 70475 136409 73855 136445
rect 73911 136409 73997 136465
rect 74053 136409 74139 136465
rect 74195 136409 74281 136465
rect 74337 136409 74423 136465
rect 74479 136409 74565 136465
rect 74621 136409 74707 136465
rect 74763 136409 74849 136465
rect 74905 136409 74991 136465
rect 75047 136409 75133 136465
rect 75189 136409 75275 136465
rect 75331 136409 75416 136465
rect 70475 136389 75416 136409
rect 70000 136323 75416 136389
rect 70000 136321 73855 136323
rect 70000 136265 70047 136321
rect 70103 136265 70171 136321
rect 70227 136265 70295 136321
rect 70351 136265 70419 136321
rect 70475 136267 73855 136321
rect 73911 136267 73997 136323
rect 74053 136267 74139 136323
rect 74195 136267 74281 136323
rect 74337 136267 74423 136323
rect 74479 136267 74565 136323
rect 74621 136267 74707 136323
rect 74763 136267 74849 136323
rect 74905 136267 74991 136323
rect 75047 136267 75133 136323
rect 75189 136267 75275 136323
rect 75331 136267 75416 136323
rect 70475 136265 75416 136267
rect 70000 136198 75416 136265
rect 70000 135811 75416 135878
rect 70000 135755 70047 135811
rect 70103 135755 70171 135811
rect 70227 135755 70295 135811
rect 70351 135755 70419 135811
rect 70475 135799 75416 135811
rect 70475 135755 73855 135799
rect 70000 135743 73855 135755
rect 73911 135743 73997 135799
rect 74053 135743 74139 135799
rect 74195 135743 74281 135799
rect 74337 135743 74423 135799
rect 74479 135743 74565 135799
rect 74621 135743 74707 135799
rect 74763 135743 74849 135799
rect 74905 135743 74991 135799
rect 75047 135743 75133 135799
rect 75189 135743 75275 135799
rect 75331 135743 75416 135799
rect 70000 135687 75416 135743
rect 70000 135631 70047 135687
rect 70103 135631 70171 135687
rect 70227 135631 70295 135687
rect 70351 135631 70419 135687
rect 70475 135657 75416 135687
rect 70475 135631 73855 135657
rect 70000 135601 73855 135631
rect 73911 135601 73997 135657
rect 74053 135601 74139 135657
rect 74195 135601 74281 135657
rect 74337 135601 74423 135657
rect 74479 135601 74565 135657
rect 74621 135601 74707 135657
rect 74763 135601 74849 135657
rect 74905 135601 74991 135657
rect 75047 135601 75133 135657
rect 75189 135601 75275 135657
rect 75331 135601 75416 135657
rect 70000 135563 75416 135601
rect 70000 135507 70047 135563
rect 70103 135507 70171 135563
rect 70227 135507 70295 135563
rect 70351 135507 70419 135563
rect 70475 135515 75416 135563
rect 70475 135507 73855 135515
rect 70000 135459 73855 135507
rect 73911 135459 73997 135515
rect 74053 135459 74139 135515
rect 74195 135459 74281 135515
rect 74337 135459 74423 135515
rect 74479 135459 74565 135515
rect 74621 135459 74707 135515
rect 74763 135459 74849 135515
rect 74905 135459 74991 135515
rect 75047 135459 75133 135515
rect 75189 135459 75275 135515
rect 75331 135459 75416 135515
rect 70000 135439 75416 135459
rect 70000 135383 70047 135439
rect 70103 135383 70171 135439
rect 70227 135383 70295 135439
rect 70351 135383 70419 135439
rect 70475 135383 75416 135439
rect 70000 135373 75416 135383
rect 70000 135317 73855 135373
rect 73911 135317 73997 135373
rect 74053 135317 74139 135373
rect 74195 135317 74281 135373
rect 74337 135317 74423 135373
rect 74479 135317 74565 135373
rect 74621 135317 74707 135373
rect 74763 135317 74849 135373
rect 74905 135317 74991 135373
rect 75047 135317 75133 135373
rect 75189 135317 75275 135373
rect 75331 135317 75416 135373
rect 70000 135315 75416 135317
rect 70000 135259 70047 135315
rect 70103 135259 70171 135315
rect 70227 135259 70295 135315
rect 70351 135259 70419 135315
rect 70475 135259 75416 135315
rect 70000 135231 75416 135259
rect 70000 135191 73855 135231
rect 70000 135135 70047 135191
rect 70103 135135 70171 135191
rect 70227 135135 70295 135191
rect 70351 135135 70419 135191
rect 70475 135175 73855 135191
rect 73911 135175 73997 135231
rect 74053 135175 74139 135231
rect 74195 135175 74281 135231
rect 74337 135175 74423 135231
rect 74479 135175 74565 135231
rect 74621 135175 74707 135231
rect 74763 135175 74849 135231
rect 74905 135175 74991 135231
rect 75047 135175 75133 135231
rect 75189 135175 75275 135231
rect 75331 135175 75416 135231
rect 70475 135135 75416 135175
rect 70000 135089 75416 135135
rect 70000 135067 73855 135089
rect 70000 135011 70047 135067
rect 70103 135011 70171 135067
rect 70227 135011 70295 135067
rect 70351 135011 70419 135067
rect 70475 135033 73855 135067
rect 73911 135033 73997 135089
rect 74053 135033 74139 135089
rect 74195 135033 74281 135089
rect 74337 135033 74423 135089
rect 74479 135033 74565 135089
rect 74621 135033 74707 135089
rect 74763 135033 74849 135089
rect 74905 135033 74991 135089
rect 75047 135033 75133 135089
rect 75189 135033 75275 135089
rect 75331 135033 75416 135089
rect 70475 135011 75416 135033
rect 70000 134947 75416 135011
rect 70000 134943 73855 134947
rect 70000 134887 70047 134943
rect 70103 134887 70171 134943
rect 70227 134887 70295 134943
rect 70351 134887 70419 134943
rect 70475 134891 73855 134943
rect 73911 134891 73997 134947
rect 74053 134891 74139 134947
rect 74195 134891 74281 134947
rect 74337 134891 74423 134947
rect 74479 134891 74565 134947
rect 74621 134891 74707 134947
rect 74763 134891 74849 134947
rect 74905 134891 74991 134947
rect 75047 134891 75133 134947
rect 75189 134891 75275 134947
rect 75331 134891 75416 134947
rect 70475 134887 75416 134891
rect 70000 134819 75416 134887
rect 70000 134763 70047 134819
rect 70103 134763 70171 134819
rect 70227 134763 70295 134819
rect 70351 134763 70419 134819
rect 70475 134805 75416 134819
rect 70475 134763 73855 134805
rect 70000 134749 73855 134763
rect 73911 134749 73997 134805
rect 74053 134749 74139 134805
rect 74195 134749 74281 134805
rect 74337 134749 74423 134805
rect 74479 134749 74565 134805
rect 74621 134749 74707 134805
rect 74763 134749 74849 134805
rect 74905 134749 74991 134805
rect 75047 134749 75133 134805
rect 75189 134749 75275 134805
rect 75331 134749 75416 134805
rect 70000 134695 75416 134749
rect 70000 134639 70047 134695
rect 70103 134639 70171 134695
rect 70227 134639 70295 134695
rect 70351 134639 70419 134695
rect 70475 134663 75416 134695
rect 70475 134639 73855 134663
rect 70000 134607 73855 134639
rect 73911 134607 73997 134663
rect 74053 134607 74139 134663
rect 74195 134607 74281 134663
rect 74337 134607 74423 134663
rect 74479 134607 74565 134663
rect 74621 134607 74707 134663
rect 74763 134607 74849 134663
rect 74905 134607 74991 134663
rect 75047 134607 75133 134663
rect 75189 134607 75275 134663
rect 75331 134607 75416 134663
rect 70000 134571 75416 134607
rect 70000 134515 70047 134571
rect 70103 134515 70171 134571
rect 70227 134515 70295 134571
rect 70351 134515 70419 134571
rect 70475 134521 75416 134571
rect 70475 134515 73855 134521
rect 70000 134465 73855 134515
rect 73911 134465 73997 134521
rect 74053 134465 74139 134521
rect 74195 134465 74281 134521
rect 74337 134465 74423 134521
rect 74479 134465 74565 134521
rect 74621 134465 74707 134521
rect 74763 134465 74849 134521
rect 74905 134465 74991 134521
rect 75047 134465 75133 134521
rect 75189 134465 75275 134521
rect 75331 134465 75416 134521
rect 70000 134447 75416 134465
rect 70000 134391 70047 134447
rect 70103 134391 70171 134447
rect 70227 134391 70295 134447
rect 70351 134391 70419 134447
rect 70475 134391 75416 134447
rect 70000 134379 75416 134391
rect 70000 134323 73855 134379
rect 73911 134323 73997 134379
rect 74053 134323 74139 134379
rect 74195 134323 74281 134379
rect 74337 134323 74423 134379
rect 74479 134323 74565 134379
rect 74621 134323 74707 134379
rect 74763 134323 74849 134379
rect 74905 134323 74991 134379
rect 75047 134323 75133 134379
rect 75189 134323 75275 134379
rect 75331 134323 75416 134379
rect 70000 134267 70047 134323
rect 70103 134267 70171 134323
rect 70227 134267 70295 134323
rect 70351 134267 70419 134323
rect 70475 134267 75416 134323
rect 70000 134237 75416 134267
rect 70000 134199 73855 134237
rect 70000 134143 70047 134199
rect 70103 134143 70171 134199
rect 70227 134143 70295 134199
rect 70351 134143 70419 134199
rect 70475 134181 73855 134199
rect 73911 134181 73997 134237
rect 74053 134181 74139 134237
rect 74195 134181 74281 134237
rect 74337 134181 74423 134237
rect 74479 134181 74565 134237
rect 74621 134181 74707 134237
rect 74763 134181 74849 134237
rect 74905 134181 74991 134237
rect 75047 134181 75133 134237
rect 75189 134181 75275 134237
rect 75331 134181 75416 134237
rect 70475 134143 75416 134181
rect 70000 134095 75416 134143
rect 70000 134075 73855 134095
rect 70000 134019 70047 134075
rect 70103 134019 70171 134075
rect 70227 134019 70295 134075
rect 70351 134019 70419 134075
rect 70475 134039 73855 134075
rect 73911 134039 73997 134095
rect 74053 134039 74139 134095
rect 74195 134039 74281 134095
rect 74337 134039 74423 134095
rect 74479 134039 74565 134095
rect 74621 134039 74707 134095
rect 74763 134039 74849 134095
rect 74905 134039 74991 134095
rect 75047 134039 75133 134095
rect 75189 134039 75275 134095
rect 75331 134039 75416 134095
rect 70475 134019 75416 134039
rect 70000 133953 75416 134019
rect 70000 133951 73855 133953
rect 70000 133895 70047 133951
rect 70103 133895 70171 133951
rect 70227 133895 70295 133951
rect 70351 133895 70419 133951
rect 70475 133897 73855 133951
rect 73911 133897 73997 133953
rect 74053 133897 74139 133953
rect 74195 133897 74281 133953
rect 74337 133897 74423 133953
rect 74479 133897 74565 133953
rect 74621 133897 74707 133953
rect 74763 133897 74849 133953
rect 74905 133897 74991 133953
rect 75047 133897 75133 133953
rect 75189 133897 75275 133953
rect 75331 133897 75416 133953
rect 70475 133895 75416 133897
rect 70000 133828 75416 133895
rect 70000 133105 75416 133172
rect 70000 133049 70047 133105
rect 70103 133049 70171 133105
rect 70227 133049 70295 133105
rect 70351 133049 70419 133105
rect 70475 133093 75416 133105
rect 70475 133049 73855 133093
rect 70000 133037 73855 133049
rect 73911 133037 73997 133093
rect 74053 133037 74139 133093
rect 74195 133037 74281 133093
rect 74337 133037 74423 133093
rect 74479 133037 74565 133093
rect 74621 133037 74707 133093
rect 74763 133037 74849 133093
rect 74905 133037 74991 133093
rect 75047 133037 75133 133093
rect 75189 133037 75275 133093
rect 75331 133037 75416 133093
rect 70000 132981 75416 133037
rect 70000 132925 70047 132981
rect 70103 132925 70171 132981
rect 70227 132925 70295 132981
rect 70351 132925 70419 132981
rect 70475 132951 75416 132981
rect 70475 132925 73855 132951
rect 70000 132895 73855 132925
rect 73911 132895 73997 132951
rect 74053 132895 74139 132951
rect 74195 132895 74281 132951
rect 74337 132895 74423 132951
rect 74479 132895 74565 132951
rect 74621 132895 74707 132951
rect 74763 132895 74849 132951
rect 74905 132895 74991 132951
rect 75047 132895 75133 132951
rect 75189 132895 75275 132951
rect 75331 132895 75416 132951
rect 70000 132857 75416 132895
rect 70000 132801 70047 132857
rect 70103 132801 70171 132857
rect 70227 132801 70295 132857
rect 70351 132801 70419 132857
rect 70475 132809 75416 132857
rect 70475 132801 73855 132809
rect 70000 132753 73855 132801
rect 73911 132753 73997 132809
rect 74053 132753 74139 132809
rect 74195 132753 74281 132809
rect 74337 132753 74423 132809
rect 74479 132753 74565 132809
rect 74621 132753 74707 132809
rect 74763 132753 74849 132809
rect 74905 132753 74991 132809
rect 75047 132753 75133 132809
rect 75189 132753 75275 132809
rect 75331 132753 75416 132809
rect 70000 132733 75416 132753
rect 70000 132677 70047 132733
rect 70103 132677 70171 132733
rect 70227 132677 70295 132733
rect 70351 132677 70419 132733
rect 70475 132677 75416 132733
rect 70000 132667 75416 132677
rect 70000 132611 73855 132667
rect 73911 132611 73997 132667
rect 74053 132611 74139 132667
rect 74195 132611 74281 132667
rect 74337 132611 74423 132667
rect 74479 132611 74565 132667
rect 74621 132611 74707 132667
rect 74763 132611 74849 132667
rect 74905 132611 74991 132667
rect 75047 132611 75133 132667
rect 75189 132611 75275 132667
rect 75331 132611 75416 132667
rect 70000 132609 75416 132611
rect 70000 132553 70047 132609
rect 70103 132553 70171 132609
rect 70227 132553 70295 132609
rect 70351 132553 70419 132609
rect 70475 132553 75416 132609
rect 70000 132525 75416 132553
rect 70000 132485 73855 132525
rect 70000 132429 70047 132485
rect 70103 132429 70171 132485
rect 70227 132429 70295 132485
rect 70351 132429 70419 132485
rect 70475 132469 73855 132485
rect 73911 132469 73997 132525
rect 74053 132469 74139 132525
rect 74195 132469 74281 132525
rect 74337 132469 74423 132525
rect 74479 132469 74565 132525
rect 74621 132469 74707 132525
rect 74763 132469 74849 132525
rect 74905 132469 74991 132525
rect 75047 132469 75133 132525
rect 75189 132469 75275 132525
rect 75331 132469 75416 132525
rect 70475 132429 75416 132469
rect 70000 132383 75416 132429
rect 70000 132361 73855 132383
rect 70000 132305 70047 132361
rect 70103 132305 70171 132361
rect 70227 132305 70295 132361
rect 70351 132305 70419 132361
rect 70475 132327 73855 132361
rect 73911 132327 73997 132383
rect 74053 132327 74139 132383
rect 74195 132327 74281 132383
rect 74337 132327 74423 132383
rect 74479 132327 74565 132383
rect 74621 132327 74707 132383
rect 74763 132327 74849 132383
rect 74905 132327 74991 132383
rect 75047 132327 75133 132383
rect 75189 132327 75275 132383
rect 75331 132327 75416 132383
rect 70475 132305 75416 132327
rect 70000 132241 75416 132305
rect 70000 132237 73855 132241
rect 70000 132181 70047 132237
rect 70103 132181 70171 132237
rect 70227 132181 70295 132237
rect 70351 132181 70419 132237
rect 70475 132185 73855 132237
rect 73911 132185 73997 132241
rect 74053 132185 74139 132241
rect 74195 132185 74281 132241
rect 74337 132185 74423 132241
rect 74479 132185 74565 132241
rect 74621 132185 74707 132241
rect 74763 132185 74849 132241
rect 74905 132185 74991 132241
rect 75047 132185 75133 132241
rect 75189 132185 75275 132241
rect 75331 132185 75416 132241
rect 70475 132181 75416 132185
rect 70000 132113 75416 132181
rect 70000 132057 70047 132113
rect 70103 132057 70171 132113
rect 70227 132057 70295 132113
rect 70351 132057 70419 132113
rect 70475 132099 75416 132113
rect 70475 132057 73855 132099
rect 70000 132043 73855 132057
rect 73911 132043 73997 132099
rect 74053 132043 74139 132099
rect 74195 132043 74281 132099
rect 74337 132043 74423 132099
rect 74479 132043 74565 132099
rect 74621 132043 74707 132099
rect 74763 132043 74849 132099
rect 74905 132043 74991 132099
rect 75047 132043 75133 132099
rect 75189 132043 75275 132099
rect 75331 132043 75416 132099
rect 70000 131989 75416 132043
rect 70000 131933 70047 131989
rect 70103 131933 70171 131989
rect 70227 131933 70295 131989
rect 70351 131933 70419 131989
rect 70475 131957 75416 131989
rect 70475 131933 73855 131957
rect 70000 131901 73855 131933
rect 73911 131901 73997 131957
rect 74053 131901 74139 131957
rect 74195 131901 74281 131957
rect 74337 131901 74423 131957
rect 74479 131901 74565 131957
rect 74621 131901 74707 131957
rect 74763 131901 74849 131957
rect 74905 131901 74991 131957
rect 75047 131901 75133 131957
rect 75189 131901 75275 131957
rect 75331 131901 75416 131957
rect 70000 131865 75416 131901
rect 70000 131809 70047 131865
rect 70103 131809 70171 131865
rect 70227 131809 70295 131865
rect 70351 131809 70419 131865
rect 70475 131815 75416 131865
rect 70475 131809 73855 131815
rect 70000 131759 73855 131809
rect 73911 131759 73997 131815
rect 74053 131759 74139 131815
rect 74195 131759 74281 131815
rect 74337 131759 74423 131815
rect 74479 131759 74565 131815
rect 74621 131759 74707 131815
rect 74763 131759 74849 131815
rect 74905 131759 74991 131815
rect 75047 131759 75133 131815
rect 75189 131759 75275 131815
rect 75331 131759 75416 131815
rect 70000 131741 75416 131759
rect 70000 131685 70047 131741
rect 70103 131685 70171 131741
rect 70227 131685 70295 131741
rect 70351 131685 70419 131741
rect 70475 131685 75416 131741
rect 70000 131673 75416 131685
rect 70000 131617 73855 131673
rect 73911 131617 73997 131673
rect 74053 131617 74139 131673
rect 74195 131617 74281 131673
rect 74337 131617 74423 131673
rect 74479 131617 74565 131673
rect 74621 131617 74707 131673
rect 74763 131617 74849 131673
rect 74905 131617 74991 131673
rect 75047 131617 75133 131673
rect 75189 131617 75275 131673
rect 75331 131617 75416 131673
rect 70000 131561 70047 131617
rect 70103 131561 70171 131617
rect 70227 131561 70295 131617
rect 70351 131561 70419 131617
rect 70475 131561 75416 131617
rect 70000 131531 75416 131561
rect 70000 131493 73855 131531
rect 70000 131437 70047 131493
rect 70103 131437 70171 131493
rect 70227 131437 70295 131493
rect 70351 131437 70419 131493
rect 70475 131475 73855 131493
rect 73911 131475 73997 131531
rect 74053 131475 74139 131531
rect 74195 131475 74281 131531
rect 74337 131475 74423 131531
rect 74479 131475 74565 131531
rect 74621 131475 74707 131531
rect 74763 131475 74849 131531
rect 74905 131475 74991 131531
rect 75047 131475 75133 131531
rect 75189 131475 75275 131531
rect 75331 131475 75416 131531
rect 70475 131437 75416 131475
rect 70000 131389 75416 131437
rect 70000 131369 73855 131389
rect 70000 131313 70047 131369
rect 70103 131313 70171 131369
rect 70227 131313 70295 131369
rect 70351 131313 70419 131369
rect 70475 131333 73855 131369
rect 73911 131333 73997 131389
rect 74053 131333 74139 131389
rect 74195 131333 74281 131389
rect 74337 131333 74423 131389
rect 74479 131333 74565 131389
rect 74621 131333 74707 131389
rect 74763 131333 74849 131389
rect 74905 131333 74991 131389
rect 75047 131333 75133 131389
rect 75189 131333 75275 131389
rect 75331 131333 75416 131389
rect 70475 131313 75416 131333
rect 70000 131247 75416 131313
rect 70000 131245 73855 131247
rect 70000 131189 70047 131245
rect 70103 131189 70171 131245
rect 70227 131189 70295 131245
rect 70351 131189 70419 131245
rect 70475 131191 73855 131245
rect 73911 131191 73997 131247
rect 74053 131191 74139 131247
rect 74195 131191 74281 131247
rect 74337 131191 74423 131247
rect 74479 131191 74565 131247
rect 74621 131191 74707 131247
rect 74763 131191 74849 131247
rect 74905 131191 74991 131247
rect 75047 131191 75133 131247
rect 75189 131191 75275 131247
rect 75331 131191 75416 131247
rect 70475 131189 75416 131191
rect 70000 131122 75416 131189
rect 70000 130735 75416 130802
rect 70000 130679 70047 130735
rect 70103 130679 70171 130735
rect 70227 130679 70295 130735
rect 70351 130679 70419 130735
rect 70475 130723 75416 130735
rect 70475 130679 73855 130723
rect 70000 130667 73855 130679
rect 73911 130667 73997 130723
rect 74053 130667 74139 130723
rect 74195 130667 74281 130723
rect 74337 130667 74423 130723
rect 74479 130667 74565 130723
rect 74621 130667 74707 130723
rect 74763 130667 74849 130723
rect 74905 130667 74991 130723
rect 75047 130667 75133 130723
rect 75189 130667 75275 130723
rect 75331 130667 75416 130723
rect 70000 130611 75416 130667
rect 70000 130555 70047 130611
rect 70103 130555 70171 130611
rect 70227 130555 70295 130611
rect 70351 130555 70419 130611
rect 70475 130581 75416 130611
rect 70475 130555 73855 130581
rect 70000 130525 73855 130555
rect 73911 130525 73997 130581
rect 74053 130525 74139 130581
rect 74195 130525 74281 130581
rect 74337 130525 74423 130581
rect 74479 130525 74565 130581
rect 74621 130525 74707 130581
rect 74763 130525 74849 130581
rect 74905 130525 74991 130581
rect 75047 130525 75133 130581
rect 75189 130525 75275 130581
rect 75331 130525 75416 130581
rect 70000 130487 75416 130525
rect 70000 130431 70047 130487
rect 70103 130431 70171 130487
rect 70227 130431 70295 130487
rect 70351 130431 70419 130487
rect 70475 130439 75416 130487
rect 70475 130431 73855 130439
rect 70000 130383 73855 130431
rect 73911 130383 73997 130439
rect 74053 130383 74139 130439
rect 74195 130383 74281 130439
rect 74337 130383 74423 130439
rect 74479 130383 74565 130439
rect 74621 130383 74707 130439
rect 74763 130383 74849 130439
rect 74905 130383 74991 130439
rect 75047 130383 75133 130439
rect 75189 130383 75275 130439
rect 75331 130383 75416 130439
rect 70000 130363 75416 130383
rect 70000 130307 70047 130363
rect 70103 130307 70171 130363
rect 70227 130307 70295 130363
rect 70351 130307 70419 130363
rect 70475 130307 75416 130363
rect 70000 130297 75416 130307
rect 70000 130241 73855 130297
rect 73911 130241 73997 130297
rect 74053 130241 74139 130297
rect 74195 130241 74281 130297
rect 74337 130241 74423 130297
rect 74479 130241 74565 130297
rect 74621 130241 74707 130297
rect 74763 130241 74849 130297
rect 74905 130241 74991 130297
rect 75047 130241 75133 130297
rect 75189 130241 75275 130297
rect 75331 130241 75416 130297
rect 70000 130239 75416 130241
rect 70000 130183 70047 130239
rect 70103 130183 70171 130239
rect 70227 130183 70295 130239
rect 70351 130183 70419 130239
rect 70475 130183 75416 130239
rect 70000 130155 75416 130183
rect 70000 130115 73855 130155
rect 70000 130059 70047 130115
rect 70103 130059 70171 130115
rect 70227 130059 70295 130115
rect 70351 130059 70419 130115
rect 70475 130099 73855 130115
rect 73911 130099 73997 130155
rect 74053 130099 74139 130155
rect 74195 130099 74281 130155
rect 74337 130099 74423 130155
rect 74479 130099 74565 130155
rect 74621 130099 74707 130155
rect 74763 130099 74849 130155
rect 74905 130099 74991 130155
rect 75047 130099 75133 130155
rect 75189 130099 75275 130155
rect 75331 130099 75416 130155
rect 70475 130059 75416 130099
rect 70000 130013 75416 130059
rect 70000 129991 73855 130013
rect 70000 129935 70047 129991
rect 70103 129935 70171 129991
rect 70227 129935 70295 129991
rect 70351 129935 70419 129991
rect 70475 129957 73855 129991
rect 73911 129957 73997 130013
rect 74053 129957 74139 130013
rect 74195 129957 74281 130013
rect 74337 129957 74423 130013
rect 74479 129957 74565 130013
rect 74621 129957 74707 130013
rect 74763 129957 74849 130013
rect 74905 129957 74991 130013
rect 75047 129957 75133 130013
rect 75189 129957 75275 130013
rect 75331 129957 75416 130013
rect 70475 129935 75416 129957
rect 70000 129871 75416 129935
rect 70000 129867 73855 129871
rect 70000 129811 70047 129867
rect 70103 129811 70171 129867
rect 70227 129811 70295 129867
rect 70351 129811 70419 129867
rect 70475 129815 73855 129867
rect 73911 129815 73997 129871
rect 74053 129815 74139 129871
rect 74195 129815 74281 129871
rect 74337 129815 74423 129871
rect 74479 129815 74565 129871
rect 74621 129815 74707 129871
rect 74763 129815 74849 129871
rect 74905 129815 74991 129871
rect 75047 129815 75133 129871
rect 75189 129815 75275 129871
rect 75331 129815 75416 129871
rect 70475 129811 75416 129815
rect 70000 129743 75416 129811
rect 70000 129687 70047 129743
rect 70103 129687 70171 129743
rect 70227 129687 70295 129743
rect 70351 129687 70419 129743
rect 70475 129729 75416 129743
rect 70475 129687 73855 129729
rect 70000 129673 73855 129687
rect 73911 129673 73997 129729
rect 74053 129673 74139 129729
rect 74195 129673 74281 129729
rect 74337 129673 74423 129729
rect 74479 129673 74565 129729
rect 74621 129673 74707 129729
rect 74763 129673 74849 129729
rect 74905 129673 74991 129729
rect 75047 129673 75133 129729
rect 75189 129673 75275 129729
rect 75331 129673 75416 129729
rect 70000 129619 75416 129673
rect 70000 129563 70047 129619
rect 70103 129563 70171 129619
rect 70227 129563 70295 129619
rect 70351 129563 70419 129619
rect 70475 129587 75416 129619
rect 70475 129563 73855 129587
rect 70000 129531 73855 129563
rect 73911 129531 73997 129587
rect 74053 129531 74139 129587
rect 74195 129531 74281 129587
rect 74337 129531 74423 129587
rect 74479 129531 74565 129587
rect 74621 129531 74707 129587
rect 74763 129531 74849 129587
rect 74905 129531 74991 129587
rect 75047 129531 75133 129587
rect 75189 129531 75275 129587
rect 75331 129531 75416 129587
rect 70000 129495 75416 129531
rect 70000 129439 70047 129495
rect 70103 129439 70171 129495
rect 70227 129439 70295 129495
rect 70351 129439 70419 129495
rect 70475 129445 75416 129495
rect 70475 129439 73855 129445
rect 70000 129389 73855 129439
rect 73911 129389 73997 129445
rect 74053 129389 74139 129445
rect 74195 129389 74281 129445
rect 74337 129389 74423 129445
rect 74479 129389 74565 129445
rect 74621 129389 74707 129445
rect 74763 129389 74849 129445
rect 74905 129389 74991 129445
rect 75047 129389 75133 129445
rect 75189 129389 75275 129445
rect 75331 129389 75416 129445
rect 70000 129371 75416 129389
rect 70000 129315 70047 129371
rect 70103 129315 70171 129371
rect 70227 129315 70295 129371
rect 70351 129315 70419 129371
rect 70475 129315 75416 129371
rect 70000 129303 75416 129315
rect 70000 129247 73855 129303
rect 73911 129247 73997 129303
rect 74053 129247 74139 129303
rect 74195 129247 74281 129303
rect 74337 129247 74423 129303
rect 74479 129247 74565 129303
rect 74621 129247 74707 129303
rect 74763 129247 74849 129303
rect 74905 129247 74991 129303
rect 75047 129247 75133 129303
rect 75189 129247 75275 129303
rect 75331 129247 75416 129303
rect 70000 129191 70047 129247
rect 70103 129191 70171 129247
rect 70227 129191 70295 129247
rect 70351 129191 70419 129247
rect 70475 129191 75416 129247
rect 70000 129161 75416 129191
rect 70000 129123 73855 129161
rect 70000 129067 70047 129123
rect 70103 129067 70171 129123
rect 70227 129067 70295 129123
rect 70351 129067 70419 129123
rect 70475 129105 73855 129123
rect 73911 129105 73997 129161
rect 74053 129105 74139 129161
rect 74195 129105 74281 129161
rect 74337 129105 74423 129161
rect 74479 129105 74565 129161
rect 74621 129105 74707 129161
rect 74763 129105 74849 129161
rect 74905 129105 74991 129161
rect 75047 129105 75133 129161
rect 75189 129105 75275 129161
rect 75331 129105 75416 129161
rect 70475 129067 75416 129105
rect 70000 129019 75416 129067
rect 70000 128999 73855 129019
rect 70000 128943 70047 128999
rect 70103 128943 70171 128999
rect 70227 128943 70295 128999
rect 70351 128943 70419 128999
rect 70475 128963 73855 128999
rect 73911 128963 73997 129019
rect 74053 128963 74139 129019
rect 74195 128963 74281 129019
rect 74337 128963 74423 129019
rect 74479 128963 74565 129019
rect 74621 128963 74707 129019
rect 74763 128963 74849 129019
rect 74905 128963 74991 129019
rect 75047 128963 75133 129019
rect 75189 128963 75275 129019
rect 75331 128963 75416 129019
rect 70475 128943 75416 128963
rect 70000 128877 75416 128943
rect 70000 128875 73855 128877
rect 70000 128819 70047 128875
rect 70103 128819 70171 128875
rect 70227 128819 70295 128875
rect 70351 128819 70419 128875
rect 70475 128821 73855 128875
rect 73911 128821 73997 128877
rect 74053 128821 74139 128877
rect 74195 128821 74281 128877
rect 74337 128821 74423 128877
rect 74479 128821 74565 128877
rect 74621 128821 74707 128877
rect 74763 128821 74849 128877
rect 74905 128821 74991 128877
rect 75047 128821 75133 128877
rect 75189 128821 75275 128877
rect 75331 128821 75416 128877
rect 70475 128819 75416 128821
rect 70000 128752 75416 128819
rect 70000 128105 75416 128172
rect 70000 128049 70047 128105
rect 70103 128049 70171 128105
rect 70227 128049 70295 128105
rect 70351 128049 70419 128105
rect 70475 128094 75416 128105
rect 70475 128049 73866 128094
rect 70000 128038 73866 128049
rect 73922 128038 74008 128094
rect 74064 128038 74150 128094
rect 74206 128038 74292 128094
rect 74348 128038 74434 128094
rect 74490 128038 74576 128094
rect 74632 128038 74718 128094
rect 74774 128038 74860 128094
rect 74916 128038 75002 128094
rect 75058 128038 75144 128094
rect 75200 128038 75286 128094
rect 75342 128038 75416 128094
rect 70000 127981 75416 128038
rect 70000 127925 70047 127981
rect 70103 127925 70171 127981
rect 70227 127925 70295 127981
rect 70351 127925 70419 127981
rect 70475 127952 75416 127981
rect 70475 127925 73866 127952
rect 70000 127896 73866 127925
rect 73922 127896 74008 127952
rect 74064 127896 74150 127952
rect 74206 127896 74292 127952
rect 74348 127896 74434 127952
rect 74490 127896 74576 127952
rect 74632 127896 74718 127952
rect 74774 127896 74860 127952
rect 74916 127896 75002 127952
rect 75058 127896 75144 127952
rect 75200 127896 75286 127952
rect 75342 127896 75416 127952
rect 70000 127857 75416 127896
rect 70000 127801 70047 127857
rect 70103 127801 70171 127857
rect 70227 127801 70295 127857
rect 70351 127801 70419 127857
rect 70475 127810 75416 127857
rect 70475 127801 73866 127810
rect 70000 127754 73866 127801
rect 73922 127754 74008 127810
rect 74064 127754 74150 127810
rect 74206 127754 74292 127810
rect 74348 127754 74434 127810
rect 74490 127754 74576 127810
rect 74632 127754 74718 127810
rect 74774 127754 74860 127810
rect 74916 127754 75002 127810
rect 75058 127754 75144 127810
rect 75200 127754 75286 127810
rect 75342 127754 75416 127810
rect 70000 127733 75416 127754
rect 70000 127677 70047 127733
rect 70103 127677 70171 127733
rect 70227 127677 70295 127733
rect 70351 127677 70419 127733
rect 70475 127677 75416 127733
rect 70000 127668 75416 127677
rect 70000 127612 73866 127668
rect 73922 127612 74008 127668
rect 74064 127612 74150 127668
rect 74206 127612 74292 127668
rect 74348 127612 74434 127668
rect 74490 127612 74576 127668
rect 74632 127612 74718 127668
rect 74774 127612 74860 127668
rect 74916 127612 75002 127668
rect 75058 127612 75144 127668
rect 75200 127612 75286 127668
rect 75342 127612 75416 127668
rect 70000 127609 75416 127612
rect 70000 127553 70047 127609
rect 70103 127553 70171 127609
rect 70227 127553 70295 127609
rect 70351 127553 70419 127609
rect 70475 127553 75416 127609
rect 70000 127526 75416 127553
rect 70000 127485 73866 127526
rect 70000 127429 70047 127485
rect 70103 127429 70171 127485
rect 70227 127429 70295 127485
rect 70351 127429 70419 127485
rect 70475 127470 73866 127485
rect 73922 127470 74008 127526
rect 74064 127470 74150 127526
rect 74206 127470 74292 127526
rect 74348 127470 74434 127526
rect 74490 127470 74576 127526
rect 74632 127470 74718 127526
rect 74774 127470 74860 127526
rect 74916 127470 75002 127526
rect 75058 127470 75144 127526
rect 75200 127470 75286 127526
rect 75342 127470 75416 127526
rect 70475 127429 75416 127470
rect 70000 127384 75416 127429
rect 70000 127361 73866 127384
rect 70000 127305 70047 127361
rect 70103 127305 70171 127361
rect 70227 127305 70295 127361
rect 70351 127305 70419 127361
rect 70475 127328 73866 127361
rect 73922 127328 74008 127384
rect 74064 127328 74150 127384
rect 74206 127328 74292 127384
rect 74348 127328 74434 127384
rect 74490 127328 74576 127384
rect 74632 127328 74718 127384
rect 74774 127328 74860 127384
rect 74916 127328 75002 127384
rect 75058 127328 75144 127384
rect 75200 127328 75286 127384
rect 75342 127328 75416 127384
rect 70475 127305 75416 127328
rect 70000 127242 75416 127305
rect 70000 127237 73866 127242
rect 70000 127181 70047 127237
rect 70103 127181 70171 127237
rect 70227 127181 70295 127237
rect 70351 127181 70419 127237
rect 70475 127186 73866 127237
rect 73922 127186 74008 127242
rect 74064 127186 74150 127242
rect 74206 127186 74292 127242
rect 74348 127186 74434 127242
rect 74490 127186 74576 127242
rect 74632 127186 74718 127242
rect 74774 127186 74860 127242
rect 74916 127186 75002 127242
rect 75058 127186 75144 127242
rect 75200 127186 75286 127242
rect 75342 127186 75416 127242
rect 70475 127181 75416 127186
rect 70000 127113 75416 127181
rect 70000 127057 70047 127113
rect 70103 127057 70171 127113
rect 70227 127057 70295 127113
rect 70351 127057 70419 127113
rect 70475 127100 75416 127113
rect 70475 127057 73866 127100
rect 70000 127044 73866 127057
rect 73922 127044 74008 127100
rect 74064 127044 74150 127100
rect 74206 127044 74292 127100
rect 74348 127044 74434 127100
rect 74490 127044 74576 127100
rect 74632 127044 74718 127100
rect 74774 127044 74860 127100
rect 74916 127044 75002 127100
rect 75058 127044 75144 127100
rect 75200 127044 75286 127100
rect 75342 127044 75416 127100
rect 70000 126989 75416 127044
rect 70000 126933 70047 126989
rect 70103 126933 70171 126989
rect 70227 126933 70295 126989
rect 70351 126933 70419 126989
rect 70475 126958 75416 126989
rect 70475 126933 73866 126958
rect 70000 126902 73866 126933
rect 73922 126902 74008 126958
rect 74064 126902 74150 126958
rect 74206 126902 74292 126958
rect 74348 126902 74434 126958
rect 74490 126902 74576 126958
rect 74632 126902 74718 126958
rect 74774 126902 74860 126958
rect 74916 126902 75002 126958
rect 75058 126902 75144 126958
rect 75200 126902 75286 126958
rect 75342 126902 75416 126958
rect 70000 126865 75416 126902
rect 70000 126809 70047 126865
rect 70103 126809 70171 126865
rect 70227 126809 70295 126865
rect 70351 126809 70419 126865
rect 70475 126816 75416 126865
rect 70475 126809 73866 126816
rect 70000 126760 73866 126809
rect 73922 126760 74008 126816
rect 74064 126760 74150 126816
rect 74206 126760 74292 126816
rect 74348 126760 74434 126816
rect 74490 126760 74576 126816
rect 74632 126760 74718 126816
rect 74774 126760 74860 126816
rect 74916 126760 75002 126816
rect 75058 126760 75144 126816
rect 75200 126760 75286 126816
rect 75342 126760 75416 126816
rect 70000 126741 75416 126760
rect 70000 126685 70047 126741
rect 70103 126685 70171 126741
rect 70227 126685 70295 126741
rect 70351 126685 70419 126741
rect 70475 126685 75416 126741
rect 70000 126674 75416 126685
rect 70000 126618 73866 126674
rect 73922 126618 74008 126674
rect 74064 126618 74150 126674
rect 74206 126618 74292 126674
rect 74348 126618 74434 126674
rect 74490 126618 74576 126674
rect 74632 126618 74718 126674
rect 74774 126618 74860 126674
rect 74916 126618 75002 126674
rect 75058 126618 75144 126674
rect 75200 126618 75286 126674
rect 75342 126618 75416 126674
rect 70000 126617 75416 126618
rect 70000 126561 70047 126617
rect 70103 126561 70171 126617
rect 70227 126561 70295 126617
rect 70351 126561 70419 126617
rect 70475 126561 75416 126617
rect 70000 126532 75416 126561
rect 70000 126493 73866 126532
rect 70000 126437 70047 126493
rect 70103 126437 70171 126493
rect 70227 126437 70295 126493
rect 70351 126437 70419 126493
rect 70475 126476 73866 126493
rect 73922 126476 74008 126532
rect 74064 126476 74150 126532
rect 74206 126476 74292 126532
rect 74348 126476 74434 126532
rect 74490 126476 74576 126532
rect 74632 126476 74718 126532
rect 74774 126476 74860 126532
rect 74916 126476 75002 126532
rect 75058 126476 75144 126532
rect 75200 126476 75286 126532
rect 75342 126476 75416 126532
rect 70475 126437 75416 126476
rect 70000 126390 75416 126437
rect 70000 126369 73866 126390
rect 70000 126313 70047 126369
rect 70103 126313 70171 126369
rect 70227 126313 70295 126369
rect 70351 126313 70419 126369
rect 70475 126334 73866 126369
rect 73922 126334 74008 126390
rect 74064 126334 74150 126390
rect 74206 126334 74292 126390
rect 74348 126334 74434 126390
rect 74490 126334 74576 126390
rect 74632 126334 74718 126390
rect 74774 126334 74860 126390
rect 74916 126334 75002 126390
rect 75058 126334 75144 126390
rect 75200 126334 75286 126390
rect 75342 126334 75416 126390
rect 70475 126313 75416 126334
rect 70000 126272 75416 126313
rect 70000 99661 75416 99728
rect 70000 99605 70047 99661
rect 70103 99605 70171 99661
rect 70227 99605 70295 99661
rect 70351 99605 70419 99661
rect 70475 99650 75416 99661
rect 70475 99605 73866 99650
rect 70000 99594 73866 99605
rect 73922 99594 74008 99650
rect 74064 99594 74150 99650
rect 74206 99594 74292 99650
rect 74348 99594 74434 99650
rect 74490 99594 74576 99650
rect 74632 99594 74718 99650
rect 74774 99594 74860 99650
rect 74916 99594 75002 99650
rect 75058 99594 75144 99650
rect 75200 99594 75286 99650
rect 75342 99594 75416 99650
rect 70000 99537 75416 99594
rect 70000 99481 70047 99537
rect 70103 99481 70171 99537
rect 70227 99481 70295 99537
rect 70351 99481 70419 99537
rect 70475 99508 75416 99537
rect 70475 99481 73866 99508
rect 70000 99452 73866 99481
rect 73922 99452 74008 99508
rect 74064 99452 74150 99508
rect 74206 99452 74292 99508
rect 74348 99452 74434 99508
rect 74490 99452 74576 99508
rect 74632 99452 74718 99508
rect 74774 99452 74860 99508
rect 74916 99452 75002 99508
rect 75058 99452 75144 99508
rect 75200 99452 75286 99508
rect 75342 99452 75416 99508
rect 70000 99413 75416 99452
rect 70000 99357 70047 99413
rect 70103 99357 70171 99413
rect 70227 99357 70295 99413
rect 70351 99357 70419 99413
rect 70475 99366 75416 99413
rect 70475 99357 73866 99366
rect 70000 99310 73866 99357
rect 73922 99310 74008 99366
rect 74064 99310 74150 99366
rect 74206 99310 74292 99366
rect 74348 99310 74434 99366
rect 74490 99310 74576 99366
rect 74632 99310 74718 99366
rect 74774 99310 74860 99366
rect 74916 99310 75002 99366
rect 75058 99310 75144 99366
rect 75200 99310 75286 99366
rect 75342 99310 75416 99366
rect 70000 99289 75416 99310
rect 70000 99233 70047 99289
rect 70103 99233 70171 99289
rect 70227 99233 70295 99289
rect 70351 99233 70419 99289
rect 70475 99233 75416 99289
rect 70000 99224 75416 99233
rect 70000 99168 73866 99224
rect 73922 99168 74008 99224
rect 74064 99168 74150 99224
rect 74206 99168 74292 99224
rect 74348 99168 74434 99224
rect 74490 99168 74576 99224
rect 74632 99168 74718 99224
rect 74774 99168 74860 99224
rect 74916 99168 75002 99224
rect 75058 99168 75144 99224
rect 75200 99168 75286 99224
rect 75342 99168 75416 99224
rect 70000 99165 75416 99168
rect 70000 99109 70047 99165
rect 70103 99109 70171 99165
rect 70227 99109 70295 99165
rect 70351 99109 70419 99165
rect 70475 99109 75416 99165
rect 70000 99082 75416 99109
rect 70000 99041 73866 99082
rect 70000 98985 70047 99041
rect 70103 98985 70171 99041
rect 70227 98985 70295 99041
rect 70351 98985 70419 99041
rect 70475 99026 73866 99041
rect 73922 99026 74008 99082
rect 74064 99026 74150 99082
rect 74206 99026 74292 99082
rect 74348 99026 74434 99082
rect 74490 99026 74576 99082
rect 74632 99026 74718 99082
rect 74774 99026 74860 99082
rect 74916 99026 75002 99082
rect 75058 99026 75144 99082
rect 75200 99026 75286 99082
rect 75342 99026 75416 99082
rect 70475 98985 75416 99026
rect 70000 98940 75416 98985
rect 70000 98917 73866 98940
rect 70000 98861 70047 98917
rect 70103 98861 70171 98917
rect 70227 98861 70295 98917
rect 70351 98861 70419 98917
rect 70475 98884 73866 98917
rect 73922 98884 74008 98940
rect 74064 98884 74150 98940
rect 74206 98884 74292 98940
rect 74348 98884 74434 98940
rect 74490 98884 74576 98940
rect 74632 98884 74718 98940
rect 74774 98884 74860 98940
rect 74916 98884 75002 98940
rect 75058 98884 75144 98940
rect 75200 98884 75286 98940
rect 75342 98884 75416 98940
rect 70475 98861 75416 98884
rect 70000 98798 75416 98861
rect 70000 98793 73866 98798
rect 70000 98737 70047 98793
rect 70103 98737 70171 98793
rect 70227 98737 70295 98793
rect 70351 98737 70419 98793
rect 70475 98742 73866 98793
rect 73922 98742 74008 98798
rect 74064 98742 74150 98798
rect 74206 98742 74292 98798
rect 74348 98742 74434 98798
rect 74490 98742 74576 98798
rect 74632 98742 74718 98798
rect 74774 98742 74860 98798
rect 74916 98742 75002 98798
rect 75058 98742 75144 98798
rect 75200 98742 75286 98798
rect 75342 98742 75416 98798
rect 70475 98737 75416 98742
rect 70000 98669 75416 98737
rect 70000 98613 70047 98669
rect 70103 98613 70171 98669
rect 70227 98613 70295 98669
rect 70351 98613 70419 98669
rect 70475 98656 75416 98669
rect 70475 98613 73866 98656
rect 70000 98600 73866 98613
rect 73922 98600 74008 98656
rect 74064 98600 74150 98656
rect 74206 98600 74292 98656
rect 74348 98600 74434 98656
rect 74490 98600 74576 98656
rect 74632 98600 74718 98656
rect 74774 98600 74860 98656
rect 74916 98600 75002 98656
rect 75058 98600 75144 98656
rect 75200 98600 75286 98656
rect 75342 98600 75416 98656
rect 70000 98545 75416 98600
rect 70000 98489 70047 98545
rect 70103 98489 70171 98545
rect 70227 98489 70295 98545
rect 70351 98489 70419 98545
rect 70475 98514 75416 98545
rect 70475 98489 73866 98514
rect 70000 98458 73866 98489
rect 73922 98458 74008 98514
rect 74064 98458 74150 98514
rect 74206 98458 74292 98514
rect 74348 98458 74434 98514
rect 74490 98458 74576 98514
rect 74632 98458 74718 98514
rect 74774 98458 74860 98514
rect 74916 98458 75002 98514
rect 75058 98458 75144 98514
rect 75200 98458 75286 98514
rect 75342 98458 75416 98514
rect 70000 98421 75416 98458
rect 70000 98365 70047 98421
rect 70103 98365 70171 98421
rect 70227 98365 70295 98421
rect 70351 98365 70419 98421
rect 70475 98372 75416 98421
rect 70475 98365 73866 98372
rect 70000 98316 73866 98365
rect 73922 98316 74008 98372
rect 74064 98316 74150 98372
rect 74206 98316 74292 98372
rect 74348 98316 74434 98372
rect 74490 98316 74576 98372
rect 74632 98316 74718 98372
rect 74774 98316 74860 98372
rect 74916 98316 75002 98372
rect 75058 98316 75144 98372
rect 75200 98316 75286 98372
rect 75342 98316 75416 98372
rect 70000 98297 75416 98316
rect 70000 98241 70047 98297
rect 70103 98241 70171 98297
rect 70227 98241 70295 98297
rect 70351 98241 70419 98297
rect 70475 98241 75416 98297
rect 70000 98230 75416 98241
rect 70000 98174 73866 98230
rect 73922 98174 74008 98230
rect 74064 98174 74150 98230
rect 74206 98174 74292 98230
rect 74348 98174 74434 98230
rect 74490 98174 74576 98230
rect 74632 98174 74718 98230
rect 74774 98174 74860 98230
rect 74916 98174 75002 98230
rect 75058 98174 75144 98230
rect 75200 98174 75286 98230
rect 75342 98174 75416 98230
rect 70000 98173 75416 98174
rect 70000 98117 70047 98173
rect 70103 98117 70171 98173
rect 70227 98117 70295 98173
rect 70351 98117 70419 98173
rect 70475 98117 75416 98173
rect 70000 98088 75416 98117
rect 70000 98049 73866 98088
rect 70000 97993 70047 98049
rect 70103 97993 70171 98049
rect 70227 97993 70295 98049
rect 70351 97993 70419 98049
rect 70475 98032 73866 98049
rect 73922 98032 74008 98088
rect 74064 98032 74150 98088
rect 74206 98032 74292 98088
rect 74348 98032 74434 98088
rect 74490 98032 74576 98088
rect 74632 98032 74718 98088
rect 74774 98032 74860 98088
rect 74916 98032 75002 98088
rect 75058 98032 75144 98088
rect 75200 98032 75286 98088
rect 75342 98032 75416 98088
rect 70475 97993 75416 98032
rect 70000 97946 75416 97993
rect 70000 97925 73866 97946
rect 70000 97869 70047 97925
rect 70103 97869 70171 97925
rect 70227 97869 70295 97925
rect 70351 97869 70419 97925
rect 70475 97890 73866 97925
rect 73922 97890 74008 97946
rect 74064 97890 74150 97946
rect 74206 97890 74292 97946
rect 74348 97890 74434 97946
rect 74490 97890 74576 97946
rect 74632 97890 74718 97946
rect 74774 97890 74860 97946
rect 74916 97890 75002 97946
rect 75058 97890 75144 97946
rect 75200 97890 75286 97946
rect 75342 97890 75416 97946
rect 70475 97869 75416 97890
rect 70000 97828 75416 97869
rect 70000 97181 75416 97248
rect 70000 97125 70047 97181
rect 70103 97125 70171 97181
rect 70227 97125 70295 97181
rect 70351 97125 70419 97181
rect 70475 97169 75416 97181
rect 70475 97125 73855 97169
rect 70000 97113 73855 97125
rect 73911 97113 73997 97169
rect 74053 97113 74139 97169
rect 74195 97113 74281 97169
rect 74337 97113 74423 97169
rect 74479 97113 74565 97169
rect 74621 97113 74707 97169
rect 74763 97113 74849 97169
rect 74905 97113 74991 97169
rect 75047 97113 75133 97169
rect 75189 97113 75275 97169
rect 75331 97113 75416 97169
rect 70000 97057 75416 97113
rect 70000 97001 70047 97057
rect 70103 97001 70171 97057
rect 70227 97001 70295 97057
rect 70351 97001 70419 97057
rect 70475 97027 75416 97057
rect 70475 97001 73855 97027
rect 70000 96971 73855 97001
rect 73911 96971 73997 97027
rect 74053 96971 74139 97027
rect 74195 96971 74281 97027
rect 74337 96971 74423 97027
rect 74479 96971 74565 97027
rect 74621 96971 74707 97027
rect 74763 96971 74849 97027
rect 74905 96971 74991 97027
rect 75047 96971 75133 97027
rect 75189 96971 75275 97027
rect 75331 96971 75416 97027
rect 70000 96933 75416 96971
rect 70000 96877 70047 96933
rect 70103 96877 70171 96933
rect 70227 96877 70295 96933
rect 70351 96877 70419 96933
rect 70475 96885 75416 96933
rect 70475 96877 73855 96885
rect 70000 96829 73855 96877
rect 73911 96829 73997 96885
rect 74053 96829 74139 96885
rect 74195 96829 74281 96885
rect 74337 96829 74423 96885
rect 74479 96829 74565 96885
rect 74621 96829 74707 96885
rect 74763 96829 74849 96885
rect 74905 96829 74991 96885
rect 75047 96829 75133 96885
rect 75189 96829 75275 96885
rect 75331 96829 75416 96885
rect 70000 96809 75416 96829
rect 70000 96753 70047 96809
rect 70103 96753 70171 96809
rect 70227 96753 70295 96809
rect 70351 96753 70419 96809
rect 70475 96753 75416 96809
rect 70000 96743 75416 96753
rect 70000 96687 73855 96743
rect 73911 96687 73997 96743
rect 74053 96687 74139 96743
rect 74195 96687 74281 96743
rect 74337 96687 74423 96743
rect 74479 96687 74565 96743
rect 74621 96687 74707 96743
rect 74763 96687 74849 96743
rect 74905 96687 74991 96743
rect 75047 96687 75133 96743
rect 75189 96687 75275 96743
rect 75331 96687 75416 96743
rect 70000 96685 75416 96687
rect 70000 96629 70047 96685
rect 70103 96629 70171 96685
rect 70227 96629 70295 96685
rect 70351 96629 70419 96685
rect 70475 96629 75416 96685
rect 70000 96601 75416 96629
rect 70000 96561 73855 96601
rect 70000 96505 70047 96561
rect 70103 96505 70171 96561
rect 70227 96505 70295 96561
rect 70351 96505 70419 96561
rect 70475 96545 73855 96561
rect 73911 96545 73997 96601
rect 74053 96545 74139 96601
rect 74195 96545 74281 96601
rect 74337 96545 74423 96601
rect 74479 96545 74565 96601
rect 74621 96545 74707 96601
rect 74763 96545 74849 96601
rect 74905 96545 74991 96601
rect 75047 96545 75133 96601
rect 75189 96545 75275 96601
rect 75331 96545 75416 96601
rect 70475 96505 75416 96545
rect 70000 96459 75416 96505
rect 70000 96437 73855 96459
rect 70000 96381 70047 96437
rect 70103 96381 70171 96437
rect 70227 96381 70295 96437
rect 70351 96381 70419 96437
rect 70475 96403 73855 96437
rect 73911 96403 73997 96459
rect 74053 96403 74139 96459
rect 74195 96403 74281 96459
rect 74337 96403 74423 96459
rect 74479 96403 74565 96459
rect 74621 96403 74707 96459
rect 74763 96403 74849 96459
rect 74905 96403 74991 96459
rect 75047 96403 75133 96459
rect 75189 96403 75275 96459
rect 75331 96403 75416 96459
rect 70475 96381 75416 96403
rect 70000 96317 75416 96381
rect 70000 96313 73855 96317
rect 70000 96257 70047 96313
rect 70103 96257 70171 96313
rect 70227 96257 70295 96313
rect 70351 96257 70419 96313
rect 70475 96261 73855 96313
rect 73911 96261 73997 96317
rect 74053 96261 74139 96317
rect 74195 96261 74281 96317
rect 74337 96261 74423 96317
rect 74479 96261 74565 96317
rect 74621 96261 74707 96317
rect 74763 96261 74849 96317
rect 74905 96261 74991 96317
rect 75047 96261 75133 96317
rect 75189 96261 75275 96317
rect 75331 96261 75416 96317
rect 70475 96257 75416 96261
rect 70000 96189 75416 96257
rect 70000 96133 70047 96189
rect 70103 96133 70171 96189
rect 70227 96133 70295 96189
rect 70351 96133 70419 96189
rect 70475 96175 75416 96189
rect 70475 96133 73855 96175
rect 70000 96119 73855 96133
rect 73911 96119 73997 96175
rect 74053 96119 74139 96175
rect 74195 96119 74281 96175
rect 74337 96119 74423 96175
rect 74479 96119 74565 96175
rect 74621 96119 74707 96175
rect 74763 96119 74849 96175
rect 74905 96119 74991 96175
rect 75047 96119 75133 96175
rect 75189 96119 75275 96175
rect 75331 96119 75416 96175
rect 70000 96065 75416 96119
rect 70000 96009 70047 96065
rect 70103 96009 70171 96065
rect 70227 96009 70295 96065
rect 70351 96009 70419 96065
rect 70475 96033 75416 96065
rect 70475 96009 73855 96033
rect 70000 95977 73855 96009
rect 73911 95977 73997 96033
rect 74053 95977 74139 96033
rect 74195 95977 74281 96033
rect 74337 95977 74423 96033
rect 74479 95977 74565 96033
rect 74621 95977 74707 96033
rect 74763 95977 74849 96033
rect 74905 95977 74991 96033
rect 75047 95977 75133 96033
rect 75189 95977 75275 96033
rect 75331 95977 75416 96033
rect 70000 95941 75416 95977
rect 70000 95885 70047 95941
rect 70103 95885 70171 95941
rect 70227 95885 70295 95941
rect 70351 95885 70419 95941
rect 70475 95891 75416 95941
rect 70475 95885 73855 95891
rect 70000 95835 73855 95885
rect 73911 95835 73997 95891
rect 74053 95835 74139 95891
rect 74195 95835 74281 95891
rect 74337 95835 74423 95891
rect 74479 95835 74565 95891
rect 74621 95835 74707 95891
rect 74763 95835 74849 95891
rect 74905 95835 74991 95891
rect 75047 95835 75133 95891
rect 75189 95835 75275 95891
rect 75331 95835 75416 95891
rect 70000 95817 75416 95835
rect 70000 95761 70047 95817
rect 70103 95761 70171 95817
rect 70227 95761 70295 95817
rect 70351 95761 70419 95817
rect 70475 95761 75416 95817
rect 70000 95749 75416 95761
rect 70000 95693 73855 95749
rect 73911 95693 73997 95749
rect 74053 95693 74139 95749
rect 74195 95693 74281 95749
rect 74337 95693 74423 95749
rect 74479 95693 74565 95749
rect 74621 95693 74707 95749
rect 74763 95693 74849 95749
rect 74905 95693 74991 95749
rect 75047 95693 75133 95749
rect 75189 95693 75275 95749
rect 75331 95693 75416 95749
rect 70000 95637 70047 95693
rect 70103 95637 70171 95693
rect 70227 95637 70295 95693
rect 70351 95637 70419 95693
rect 70475 95637 75416 95693
rect 70000 95607 75416 95637
rect 70000 95569 73855 95607
rect 70000 95513 70047 95569
rect 70103 95513 70171 95569
rect 70227 95513 70295 95569
rect 70351 95513 70419 95569
rect 70475 95551 73855 95569
rect 73911 95551 73997 95607
rect 74053 95551 74139 95607
rect 74195 95551 74281 95607
rect 74337 95551 74423 95607
rect 74479 95551 74565 95607
rect 74621 95551 74707 95607
rect 74763 95551 74849 95607
rect 74905 95551 74991 95607
rect 75047 95551 75133 95607
rect 75189 95551 75275 95607
rect 75331 95551 75416 95607
rect 70475 95513 75416 95551
rect 70000 95465 75416 95513
rect 70000 95445 73855 95465
rect 70000 95389 70047 95445
rect 70103 95389 70171 95445
rect 70227 95389 70295 95445
rect 70351 95389 70419 95445
rect 70475 95409 73855 95445
rect 73911 95409 73997 95465
rect 74053 95409 74139 95465
rect 74195 95409 74281 95465
rect 74337 95409 74423 95465
rect 74479 95409 74565 95465
rect 74621 95409 74707 95465
rect 74763 95409 74849 95465
rect 74905 95409 74991 95465
rect 75047 95409 75133 95465
rect 75189 95409 75275 95465
rect 75331 95409 75416 95465
rect 70475 95389 75416 95409
rect 70000 95323 75416 95389
rect 70000 95321 73855 95323
rect 70000 95265 70047 95321
rect 70103 95265 70171 95321
rect 70227 95265 70295 95321
rect 70351 95265 70419 95321
rect 70475 95267 73855 95321
rect 73911 95267 73997 95323
rect 74053 95267 74139 95323
rect 74195 95267 74281 95323
rect 74337 95267 74423 95323
rect 74479 95267 74565 95323
rect 74621 95267 74707 95323
rect 74763 95267 74849 95323
rect 74905 95267 74991 95323
rect 75047 95267 75133 95323
rect 75189 95267 75275 95323
rect 75331 95267 75416 95323
rect 70475 95265 75416 95267
rect 70000 95198 75416 95265
rect 70000 94811 75416 94878
rect 70000 94755 70047 94811
rect 70103 94755 70171 94811
rect 70227 94755 70295 94811
rect 70351 94755 70419 94811
rect 70475 94799 75416 94811
rect 70475 94755 73855 94799
rect 70000 94743 73855 94755
rect 73911 94743 73997 94799
rect 74053 94743 74139 94799
rect 74195 94743 74281 94799
rect 74337 94743 74423 94799
rect 74479 94743 74565 94799
rect 74621 94743 74707 94799
rect 74763 94743 74849 94799
rect 74905 94743 74991 94799
rect 75047 94743 75133 94799
rect 75189 94743 75275 94799
rect 75331 94743 75416 94799
rect 70000 94687 75416 94743
rect 70000 94631 70047 94687
rect 70103 94631 70171 94687
rect 70227 94631 70295 94687
rect 70351 94631 70419 94687
rect 70475 94657 75416 94687
rect 70475 94631 73855 94657
rect 70000 94601 73855 94631
rect 73911 94601 73997 94657
rect 74053 94601 74139 94657
rect 74195 94601 74281 94657
rect 74337 94601 74423 94657
rect 74479 94601 74565 94657
rect 74621 94601 74707 94657
rect 74763 94601 74849 94657
rect 74905 94601 74991 94657
rect 75047 94601 75133 94657
rect 75189 94601 75275 94657
rect 75331 94601 75416 94657
rect 70000 94563 75416 94601
rect 70000 94507 70047 94563
rect 70103 94507 70171 94563
rect 70227 94507 70295 94563
rect 70351 94507 70419 94563
rect 70475 94515 75416 94563
rect 70475 94507 73855 94515
rect 70000 94459 73855 94507
rect 73911 94459 73997 94515
rect 74053 94459 74139 94515
rect 74195 94459 74281 94515
rect 74337 94459 74423 94515
rect 74479 94459 74565 94515
rect 74621 94459 74707 94515
rect 74763 94459 74849 94515
rect 74905 94459 74991 94515
rect 75047 94459 75133 94515
rect 75189 94459 75275 94515
rect 75331 94459 75416 94515
rect 70000 94439 75416 94459
rect 70000 94383 70047 94439
rect 70103 94383 70171 94439
rect 70227 94383 70295 94439
rect 70351 94383 70419 94439
rect 70475 94383 75416 94439
rect 70000 94373 75416 94383
rect 70000 94317 73855 94373
rect 73911 94317 73997 94373
rect 74053 94317 74139 94373
rect 74195 94317 74281 94373
rect 74337 94317 74423 94373
rect 74479 94317 74565 94373
rect 74621 94317 74707 94373
rect 74763 94317 74849 94373
rect 74905 94317 74991 94373
rect 75047 94317 75133 94373
rect 75189 94317 75275 94373
rect 75331 94317 75416 94373
rect 70000 94315 75416 94317
rect 70000 94259 70047 94315
rect 70103 94259 70171 94315
rect 70227 94259 70295 94315
rect 70351 94259 70419 94315
rect 70475 94259 75416 94315
rect 70000 94231 75416 94259
rect 70000 94191 73855 94231
rect 70000 94135 70047 94191
rect 70103 94135 70171 94191
rect 70227 94135 70295 94191
rect 70351 94135 70419 94191
rect 70475 94175 73855 94191
rect 73911 94175 73997 94231
rect 74053 94175 74139 94231
rect 74195 94175 74281 94231
rect 74337 94175 74423 94231
rect 74479 94175 74565 94231
rect 74621 94175 74707 94231
rect 74763 94175 74849 94231
rect 74905 94175 74991 94231
rect 75047 94175 75133 94231
rect 75189 94175 75275 94231
rect 75331 94175 75416 94231
rect 70475 94135 75416 94175
rect 70000 94089 75416 94135
rect 70000 94067 73855 94089
rect 70000 94011 70047 94067
rect 70103 94011 70171 94067
rect 70227 94011 70295 94067
rect 70351 94011 70419 94067
rect 70475 94033 73855 94067
rect 73911 94033 73997 94089
rect 74053 94033 74139 94089
rect 74195 94033 74281 94089
rect 74337 94033 74423 94089
rect 74479 94033 74565 94089
rect 74621 94033 74707 94089
rect 74763 94033 74849 94089
rect 74905 94033 74991 94089
rect 75047 94033 75133 94089
rect 75189 94033 75275 94089
rect 75331 94033 75416 94089
rect 70475 94011 75416 94033
rect 70000 93947 75416 94011
rect 70000 93943 73855 93947
rect 70000 93887 70047 93943
rect 70103 93887 70171 93943
rect 70227 93887 70295 93943
rect 70351 93887 70419 93943
rect 70475 93891 73855 93943
rect 73911 93891 73997 93947
rect 74053 93891 74139 93947
rect 74195 93891 74281 93947
rect 74337 93891 74423 93947
rect 74479 93891 74565 93947
rect 74621 93891 74707 93947
rect 74763 93891 74849 93947
rect 74905 93891 74991 93947
rect 75047 93891 75133 93947
rect 75189 93891 75275 93947
rect 75331 93891 75416 93947
rect 70475 93887 75416 93891
rect 70000 93819 75416 93887
rect 70000 93763 70047 93819
rect 70103 93763 70171 93819
rect 70227 93763 70295 93819
rect 70351 93763 70419 93819
rect 70475 93805 75416 93819
rect 70475 93763 73855 93805
rect 70000 93749 73855 93763
rect 73911 93749 73997 93805
rect 74053 93749 74139 93805
rect 74195 93749 74281 93805
rect 74337 93749 74423 93805
rect 74479 93749 74565 93805
rect 74621 93749 74707 93805
rect 74763 93749 74849 93805
rect 74905 93749 74991 93805
rect 75047 93749 75133 93805
rect 75189 93749 75275 93805
rect 75331 93749 75416 93805
rect 70000 93695 75416 93749
rect 70000 93639 70047 93695
rect 70103 93639 70171 93695
rect 70227 93639 70295 93695
rect 70351 93639 70419 93695
rect 70475 93663 75416 93695
rect 70475 93639 73855 93663
rect 70000 93607 73855 93639
rect 73911 93607 73997 93663
rect 74053 93607 74139 93663
rect 74195 93607 74281 93663
rect 74337 93607 74423 93663
rect 74479 93607 74565 93663
rect 74621 93607 74707 93663
rect 74763 93607 74849 93663
rect 74905 93607 74991 93663
rect 75047 93607 75133 93663
rect 75189 93607 75275 93663
rect 75331 93607 75416 93663
rect 70000 93571 75416 93607
rect 70000 93515 70047 93571
rect 70103 93515 70171 93571
rect 70227 93515 70295 93571
rect 70351 93515 70419 93571
rect 70475 93521 75416 93571
rect 70475 93515 73855 93521
rect 70000 93465 73855 93515
rect 73911 93465 73997 93521
rect 74053 93465 74139 93521
rect 74195 93465 74281 93521
rect 74337 93465 74423 93521
rect 74479 93465 74565 93521
rect 74621 93465 74707 93521
rect 74763 93465 74849 93521
rect 74905 93465 74991 93521
rect 75047 93465 75133 93521
rect 75189 93465 75275 93521
rect 75331 93465 75416 93521
rect 70000 93447 75416 93465
rect 70000 93391 70047 93447
rect 70103 93391 70171 93447
rect 70227 93391 70295 93447
rect 70351 93391 70419 93447
rect 70475 93391 75416 93447
rect 70000 93379 75416 93391
rect 70000 93323 73855 93379
rect 73911 93323 73997 93379
rect 74053 93323 74139 93379
rect 74195 93323 74281 93379
rect 74337 93323 74423 93379
rect 74479 93323 74565 93379
rect 74621 93323 74707 93379
rect 74763 93323 74849 93379
rect 74905 93323 74991 93379
rect 75047 93323 75133 93379
rect 75189 93323 75275 93379
rect 75331 93323 75416 93379
rect 70000 93267 70047 93323
rect 70103 93267 70171 93323
rect 70227 93267 70295 93323
rect 70351 93267 70419 93323
rect 70475 93267 75416 93323
rect 70000 93237 75416 93267
rect 70000 93199 73855 93237
rect 70000 93143 70047 93199
rect 70103 93143 70171 93199
rect 70227 93143 70295 93199
rect 70351 93143 70419 93199
rect 70475 93181 73855 93199
rect 73911 93181 73997 93237
rect 74053 93181 74139 93237
rect 74195 93181 74281 93237
rect 74337 93181 74423 93237
rect 74479 93181 74565 93237
rect 74621 93181 74707 93237
rect 74763 93181 74849 93237
rect 74905 93181 74991 93237
rect 75047 93181 75133 93237
rect 75189 93181 75275 93237
rect 75331 93181 75416 93237
rect 70475 93143 75416 93181
rect 70000 93095 75416 93143
rect 70000 93075 73855 93095
rect 70000 93019 70047 93075
rect 70103 93019 70171 93075
rect 70227 93019 70295 93075
rect 70351 93019 70419 93075
rect 70475 93039 73855 93075
rect 73911 93039 73997 93095
rect 74053 93039 74139 93095
rect 74195 93039 74281 93095
rect 74337 93039 74423 93095
rect 74479 93039 74565 93095
rect 74621 93039 74707 93095
rect 74763 93039 74849 93095
rect 74905 93039 74991 93095
rect 75047 93039 75133 93095
rect 75189 93039 75275 93095
rect 75331 93039 75416 93095
rect 70475 93019 75416 93039
rect 70000 92953 75416 93019
rect 70000 92951 73855 92953
rect 70000 92895 70047 92951
rect 70103 92895 70171 92951
rect 70227 92895 70295 92951
rect 70351 92895 70419 92951
rect 70475 92897 73855 92951
rect 73911 92897 73997 92953
rect 74053 92897 74139 92953
rect 74195 92897 74281 92953
rect 74337 92897 74423 92953
rect 74479 92897 74565 92953
rect 74621 92897 74707 92953
rect 74763 92897 74849 92953
rect 74905 92897 74991 92953
rect 75047 92897 75133 92953
rect 75189 92897 75275 92953
rect 75331 92897 75416 92953
rect 70475 92895 75416 92897
rect 70000 92828 75416 92895
rect 70000 92105 75416 92172
rect 70000 92049 70047 92105
rect 70103 92049 70171 92105
rect 70227 92049 70295 92105
rect 70351 92049 70419 92105
rect 70475 92093 75416 92105
rect 70475 92049 73855 92093
rect 70000 92037 73855 92049
rect 73911 92037 73997 92093
rect 74053 92037 74139 92093
rect 74195 92037 74281 92093
rect 74337 92037 74423 92093
rect 74479 92037 74565 92093
rect 74621 92037 74707 92093
rect 74763 92037 74849 92093
rect 74905 92037 74991 92093
rect 75047 92037 75133 92093
rect 75189 92037 75275 92093
rect 75331 92037 75416 92093
rect 70000 91981 75416 92037
rect 70000 91925 70047 91981
rect 70103 91925 70171 91981
rect 70227 91925 70295 91981
rect 70351 91925 70419 91981
rect 70475 91951 75416 91981
rect 70475 91925 73855 91951
rect 70000 91895 73855 91925
rect 73911 91895 73997 91951
rect 74053 91895 74139 91951
rect 74195 91895 74281 91951
rect 74337 91895 74423 91951
rect 74479 91895 74565 91951
rect 74621 91895 74707 91951
rect 74763 91895 74849 91951
rect 74905 91895 74991 91951
rect 75047 91895 75133 91951
rect 75189 91895 75275 91951
rect 75331 91895 75416 91951
rect 70000 91857 75416 91895
rect 70000 91801 70047 91857
rect 70103 91801 70171 91857
rect 70227 91801 70295 91857
rect 70351 91801 70419 91857
rect 70475 91809 75416 91857
rect 70475 91801 73855 91809
rect 70000 91753 73855 91801
rect 73911 91753 73997 91809
rect 74053 91753 74139 91809
rect 74195 91753 74281 91809
rect 74337 91753 74423 91809
rect 74479 91753 74565 91809
rect 74621 91753 74707 91809
rect 74763 91753 74849 91809
rect 74905 91753 74991 91809
rect 75047 91753 75133 91809
rect 75189 91753 75275 91809
rect 75331 91753 75416 91809
rect 70000 91733 75416 91753
rect 70000 91677 70047 91733
rect 70103 91677 70171 91733
rect 70227 91677 70295 91733
rect 70351 91677 70419 91733
rect 70475 91677 75416 91733
rect 70000 91667 75416 91677
rect 70000 91611 73855 91667
rect 73911 91611 73997 91667
rect 74053 91611 74139 91667
rect 74195 91611 74281 91667
rect 74337 91611 74423 91667
rect 74479 91611 74565 91667
rect 74621 91611 74707 91667
rect 74763 91611 74849 91667
rect 74905 91611 74991 91667
rect 75047 91611 75133 91667
rect 75189 91611 75275 91667
rect 75331 91611 75416 91667
rect 70000 91609 75416 91611
rect 70000 91553 70047 91609
rect 70103 91553 70171 91609
rect 70227 91553 70295 91609
rect 70351 91553 70419 91609
rect 70475 91553 75416 91609
rect 70000 91525 75416 91553
rect 70000 91485 73855 91525
rect 70000 91429 70047 91485
rect 70103 91429 70171 91485
rect 70227 91429 70295 91485
rect 70351 91429 70419 91485
rect 70475 91469 73855 91485
rect 73911 91469 73997 91525
rect 74053 91469 74139 91525
rect 74195 91469 74281 91525
rect 74337 91469 74423 91525
rect 74479 91469 74565 91525
rect 74621 91469 74707 91525
rect 74763 91469 74849 91525
rect 74905 91469 74991 91525
rect 75047 91469 75133 91525
rect 75189 91469 75275 91525
rect 75331 91469 75416 91525
rect 70475 91429 75416 91469
rect 70000 91383 75416 91429
rect 70000 91361 73855 91383
rect 70000 91305 70047 91361
rect 70103 91305 70171 91361
rect 70227 91305 70295 91361
rect 70351 91305 70419 91361
rect 70475 91327 73855 91361
rect 73911 91327 73997 91383
rect 74053 91327 74139 91383
rect 74195 91327 74281 91383
rect 74337 91327 74423 91383
rect 74479 91327 74565 91383
rect 74621 91327 74707 91383
rect 74763 91327 74849 91383
rect 74905 91327 74991 91383
rect 75047 91327 75133 91383
rect 75189 91327 75275 91383
rect 75331 91327 75416 91383
rect 70475 91305 75416 91327
rect 70000 91241 75416 91305
rect 70000 91237 73855 91241
rect 70000 91181 70047 91237
rect 70103 91181 70171 91237
rect 70227 91181 70295 91237
rect 70351 91181 70419 91237
rect 70475 91185 73855 91237
rect 73911 91185 73997 91241
rect 74053 91185 74139 91241
rect 74195 91185 74281 91241
rect 74337 91185 74423 91241
rect 74479 91185 74565 91241
rect 74621 91185 74707 91241
rect 74763 91185 74849 91241
rect 74905 91185 74991 91241
rect 75047 91185 75133 91241
rect 75189 91185 75275 91241
rect 75331 91185 75416 91241
rect 70475 91181 75416 91185
rect 70000 91113 75416 91181
rect 70000 91057 70047 91113
rect 70103 91057 70171 91113
rect 70227 91057 70295 91113
rect 70351 91057 70419 91113
rect 70475 91099 75416 91113
rect 70475 91057 73855 91099
rect 70000 91043 73855 91057
rect 73911 91043 73997 91099
rect 74053 91043 74139 91099
rect 74195 91043 74281 91099
rect 74337 91043 74423 91099
rect 74479 91043 74565 91099
rect 74621 91043 74707 91099
rect 74763 91043 74849 91099
rect 74905 91043 74991 91099
rect 75047 91043 75133 91099
rect 75189 91043 75275 91099
rect 75331 91043 75416 91099
rect 70000 90989 75416 91043
rect 70000 90933 70047 90989
rect 70103 90933 70171 90989
rect 70227 90933 70295 90989
rect 70351 90933 70419 90989
rect 70475 90957 75416 90989
rect 70475 90933 73855 90957
rect 70000 90901 73855 90933
rect 73911 90901 73997 90957
rect 74053 90901 74139 90957
rect 74195 90901 74281 90957
rect 74337 90901 74423 90957
rect 74479 90901 74565 90957
rect 74621 90901 74707 90957
rect 74763 90901 74849 90957
rect 74905 90901 74991 90957
rect 75047 90901 75133 90957
rect 75189 90901 75275 90957
rect 75331 90901 75416 90957
rect 70000 90865 75416 90901
rect 70000 90809 70047 90865
rect 70103 90809 70171 90865
rect 70227 90809 70295 90865
rect 70351 90809 70419 90865
rect 70475 90815 75416 90865
rect 70475 90809 73855 90815
rect 70000 90759 73855 90809
rect 73911 90759 73997 90815
rect 74053 90759 74139 90815
rect 74195 90759 74281 90815
rect 74337 90759 74423 90815
rect 74479 90759 74565 90815
rect 74621 90759 74707 90815
rect 74763 90759 74849 90815
rect 74905 90759 74991 90815
rect 75047 90759 75133 90815
rect 75189 90759 75275 90815
rect 75331 90759 75416 90815
rect 70000 90741 75416 90759
rect 70000 90685 70047 90741
rect 70103 90685 70171 90741
rect 70227 90685 70295 90741
rect 70351 90685 70419 90741
rect 70475 90685 75416 90741
rect 70000 90673 75416 90685
rect 70000 90617 73855 90673
rect 73911 90617 73997 90673
rect 74053 90617 74139 90673
rect 74195 90617 74281 90673
rect 74337 90617 74423 90673
rect 74479 90617 74565 90673
rect 74621 90617 74707 90673
rect 74763 90617 74849 90673
rect 74905 90617 74991 90673
rect 75047 90617 75133 90673
rect 75189 90617 75275 90673
rect 75331 90617 75416 90673
rect 70000 90561 70047 90617
rect 70103 90561 70171 90617
rect 70227 90561 70295 90617
rect 70351 90561 70419 90617
rect 70475 90561 75416 90617
rect 70000 90531 75416 90561
rect 70000 90493 73855 90531
rect 70000 90437 70047 90493
rect 70103 90437 70171 90493
rect 70227 90437 70295 90493
rect 70351 90437 70419 90493
rect 70475 90475 73855 90493
rect 73911 90475 73997 90531
rect 74053 90475 74139 90531
rect 74195 90475 74281 90531
rect 74337 90475 74423 90531
rect 74479 90475 74565 90531
rect 74621 90475 74707 90531
rect 74763 90475 74849 90531
rect 74905 90475 74991 90531
rect 75047 90475 75133 90531
rect 75189 90475 75275 90531
rect 75331 90475 75416 90531
rect 70475 90437 75416 90475
rect 70000 90389 75416 90437
rect 70000 90369 73855 90389
rect 70000 90313 70047 90369
rect 70103 90313 70171 90369
rect 70227 90313 70295 90369
rect 70351 90313 70419 90369
rect 70475 90333 73855 90369
rect 73911 90333 73997 90389
rect 74053 90333 74139 90389
rect 74195 90333 74281 90389
rect 74337 90333 74423 90389
rect 74479 90333 74565 90389
rect 74621 90333 74707 90389
rect 74763 90333 74849 90389
rect 74905 90333 74991 90389
rect 75047 90333 75133 90389
rect 75189 90333 75275 90389
rect 75331 90333 75416 90389
rect 70475 90313 75416 90333
rect 70000 90247 75416 90313
rect 70000 90245 73855 90247
rect 70000 90189 70047 90245
rect 70103 90189 70171 90245
rect 70227 90189 70295 90245
rect 70351 90189 70419 90245
rect 70475 90191 73855 90245
rect 73911 90191 73997 90247
rect 74053 90191 74139 90247
rect 74195 90191 74281 90247
rect 74337 90191 74423 90247
rect 74479 90191 74565 90247
rect 74621 90191 74707 90247
rect 74763 90191 74849 90247
rect 74905 90191 74991 90247
rect 75047 90191 75133 90247
rect 75189 90191 75275 90247
rect 75331 90191 75416 90247
rect 70475 90189 75416 90191
rect 70000 90122 75416 90189
rect 70000 89735 75416 89802
rect 70000 89679 70047 89735
rect 70103 89679 70171 89735
rect 70227 89679 70295 89735
rect 70351 89679 70419 89735
rect 70475 89723 75416 89735
rect 70475 89679 73855 89723
rect 70000 89667 73855 89679
rect 73911 89667 73997 89723
rect 74053 89667 74139 89723
rect 74195 89667 74281 89723
rect 74337 89667 74423 89723
rect 74479 89667 74565 89723
rect 74621 89667 74707 89723
rect 74763 89667 74849 89723
rect 74905 89667 74991 89723
rect 75047 89667 75133 89723
rect 75189 89667 75275 89723
rect 75331 89667 75416 89723
rect 70000 89611 75416 89667
rect 70000 89555 70047 89611
rect 70103 89555 70171 89611
rect 70227 89555 70295 89611
rect 70351 89555 70419 89611
rect 70475 89581 75416 89611
rect 70475 89555 73855 89581
rect 70000 89525 73855 89555
rect 73911 89525 73997 89581
rect 74053 89525 74139 89581
rect 74195 89525 74281 89581
rect 74337 89525 74423 89581
rect 74479 89525 74565 89581
rect 74621 89525 74707 89581
rect 74763 89525 74849 89581
rect 74905 89525 74991 89581
rect 75047 89525 75133 89581
rect 75189 89525 75275 89581
rect 75331 89525 75416 89581
rect 70000 89487 75416 89525
rect 70000 89431 70047 89487
rect 70103 89431 70171 89487
rect 70227 89431 70295 89487
rect 70351 89431 70419 89487
rect 70475 89439 75416 89487
rect 70475 89431 73855 89439
rect 70000 89383 73855 89431
rect 73911 89383 73997 89439
rect 74053 89383 74139 89439
rect 74195 89383 74281 89439
rect 74337 89383 74423 89439
rect 74479 89383 74565 89439
rect 74621 89383 74707 89439
rect 74763 89383 74849 89439
rect 74905 89383 74991 89439
rect 75047 89383 75133 89439
rect 75189 89383 75275 89439
rect 75331 89383 75416 89439
rect 70000 89363 75416 89383
rect 70000 89307 70047 89363
rect 70103 89307 70171 89363
rect 70227 89307 70295 89363
rect 70351 89307 70419 89363
rect 70475 89307 75416 89363
rect 70000 89297 75416 89307
rect 70000 89241 73855 89297
rect 73911 89241 73997 89297
rect 74053 89241 74139 89297
rect 74195 89241 74281 89297
rect 74337 89241 74423 89297
rect 74479 89241 74565 89297
rect 74621 89241 74707 89297
rect 74763 89241 74849 89297
rect 74905 89241 74991 89297
rect 75047 89241 75133 89297
rect 75189 89241 75275 89297
rect 75331 89241 75416 89297
rect 70000 89239 75416 89241
rect 70000 89183 70047 89239
rect 70103 89183 70171 89239
rect 70227 89183 70295 89239
rect 70351 89183 70419 89239
rect 70475 89183 75416 89239
rect 70000 89155 75416 89183
rect 70000 89115 73855 89155
rect 70000 89059 70047 89115
rect 70103 89059 70171 89115
rect 70227 89059 70295 89115
rect 70351 89059 70419 89115
rect 70475 89099 73855 89115
rect 73911 89099 73997 89155
rect 74053 89099 74139 89155
rect 74195 89099 74281 89155
rect 74337 89099 74423 89155
rect 74479 89099 74565 89155
rect 74621 89099 74707 89155
rect 74763 89099 74849 89155
rect 74905 89099 74991 89155
rect 75047 89099 75133 89155
rect 75189 89099 75275 89155
rect 75331 89099 75416 89155
rect 70475 89059 75416 89099
rect 70000 89013 75416 89059
rect 70000 88991 73855 89013
rect 70000 88935 70047 88991
rect 70103 88935 70171 88991
rect 70227 88935 70295 88991
rect 70351 88935 70419 88991
rect 70475 88957 73855 88991
rect 73911 88957 73997 89013
rect 74053 88957 74139 89013
rect 74195 88957 74281 89013
rect 74337 88957 74423 89013
rect 74479 88957 74565 89013
rect 74621 88957 74707 89013
rect 74763 88957 74849 89013
rect 74905 88957 74991 89013
rect 75047 88957 75133 89013
rect 75189 88957 75275 89013
rect 75331 88957 75416 89013
rect 70475 88935 75416 88957
rect 70000 88871 75416 88935
rect 70000 88867 73855 88871
rect 70000 88811 70047 88867
rect 70103 88811 70171 88867
rect 70227 88811 70295 88867
rect 70351 88811 70419 88867
rect 70475 88815 73855 88867
rect 73911 88815 73997 88871
rect 74053 88815 74139 88871
rect 74195 88815 74281 88871
rect 74337 88815 74423 88871
rect 74479 88815 74565 88871
rect 74621 88815 74707 88871
rect 74763 88815 74849 88871
rect 74905 88815 74991 88871
rect 75047 88815 75133 88871
rect 75189 88815 75275 88871
rect 75331 88815 75416 88871
rect 70475 88811 75416 88815
rect 70000 88743 75416 88811
rect 70000 88687 70047 88743
rect 70103 88687 70171 88743
rect 70227 88687 70295 88743
rect 70351 88687 70419 88743
rect 70475 88729 75416 88743
rect 70475 88687 73855 88729
rect 70000 88673 73855 88687
rect 73911 88673 73997 88729
rect 74053 88673 74139 88729
rect 74195 88673 74281 88729
rect 74337 88673 74423 88729
rect 74479 88673 74565 88729
rect 74621 88673 74707 88729
rect 74763 88673 74849 88729
rect 74905 88673 74991 88729
rect 75047 88673 75133 88729
rect 75189 88673 75275 88729
rect 75331 88673 75416 88729
rect 70000 88619 75416 88673
rect 70000 88563 70047 88619
rect 70103 88563 70171 88619
rect 70227 88563 70295 88619
rect 70351 88563 70419 88619
rect 70475 88587 75416 88619
rect 70475 88563 73855 88587
rect 70000 88531 73855 88563
rect 73911 88531 73997 88587
rect 74053 88531 74139 88587
rect 74195 88531 74281 88587
rect 74337 88531 74423 88587
rect 74479 88531 74565 88587
rect 74621 88531 74707 88587
rect 74763 88531 74849 88587
rect 74905 88531 74991 88587
rect 75047 88531 75133 88587
rect 75189 88531 75275 88587
rect 75331 88531 75416 88587
rect 70000 88495 75416 88531
rect 70000 88439 70047 88495
rect 70103 88439 70171 88495
rect 70227 88439 70295 88495
rect 70351 88439 70419 88495
rect 70475 88445 75416 88495
rect 70475 88439 73855 88445
rect 70000 88389 73855 88439
rect 73911 88389 73997 88445
rect 74053 88389 74139 88445
rect 74195 88389 74281 88445
rect 74337 88389 74423 88445
rect 74479 88389 74565 88445
rect 74621 88389 74707 88445
rect 74763 88389 74849 88445
rect 74905 88389 74991 88445
rect 75047 88389 75133 88445
rect 75189 88389 75275 88445
rect 75331 88389 75416 88445
rect 70000 88371 75416 88389
rect 70000 88315 70047 88371
rect 70103 88315 70171 88371
rect 70227 88315 70295 88371
rect 70351 88315 70419 88371
rect 70475 88315 75416 88371
rect 70000 88303 75416 88315
rect 70000 88247 73855 88303
rect 73911 88247 73997 88303
rect 74053 88247 74139 88303
rect 74195 88247 74281 88303
rect 74337 88247 74423 88303
rect 74479 88247 74565 88303
rect 74621 88247 74707 88303
rect 74763 88247 74849 88303
rect 74905 88247 74991 88303
rect 75047 88247 75133 88303
rect 75189 88247 75275 88303
rect 75331 88247 75416 88303
rect 70000 88191 70047 88247
rect 70103 88191 70171 88247
rect 70227 88191 70295 88247
rect 70351 88191 70419 88247
rect 70475 88191 75416 88247
rect 70000 88161 75416 88191
rect 70000 88123 73855 88161
rect 70000 88067 70047 88123
rect 70103 88067 70171 88123
rect 70227 88067 70295 88123
rect 70351 88067 70419 88123
rect 70475 88105 73855 88123
rect 73911 88105 73997 88161
rect 74053 88105 74139 88161
rect 74195 88105 74281 88161
rect 74337 88105 74423 88161
rect 74479 88105 74565 88161
rect 74621 88105 74707 88161
rect 74763 88105 74849 88161
rect 74905 88105 74991 88161
rect 75047 88105 75133 88161
rect 75189 88105 75275 88161
rect 75331 88105 75416 88161
rect 70475 88067 75416 88105
rect 70000 88019 75416 88067
rect 70000 87999 73855 88019
rect 70000 87943 70047 87999
rect 70103 87943 70171 87999
rect 70227 87943 70295 87999
rect 70351 87943 70419 87999
rect 70475 87963 73855 87999
rect 73911 87963 73997 88019
rect 74053 87963 74139 88019
rect 74195 87963 74281 88019
rect 74337 87963 74423 88019
rect 74479 87963 74565 88019
rect 74621 87963 74707 88019
rect 74763 87963 74849 88019
rect 74905 87963 74991 88019
rect 75047 87963 75133 88019
rect 75189 87963 75275 88019
rect 75331 87963 75416 88019
rect 70475 87943 75416 87963
rect 70000 87877 75416 87943
rect 70000 87875 73855 87877
rect 70000 87819 70047 87875
rect 70103 87819 70171 87875
rect 70227 87819 70295 87875
rect 70351 87819 70419 87875
rect 70475 87821 73855 87875
rect 73911 87821 73997 87877
rect 74053 87821 74139 87877
rect 74195 87821 74281 87877
rect 74337 87821 74423 87877
rect 74479 87821 74565 87877
rect 74621 87821 74707 87877
rect 74763 87821 74849 87877
rect 74905 87821 74991 87877
rect 75047 87821 75133 87877
rect 75189 87821 75275 87877
rect 75331 87821 75416 87877
rect 70475 87819 75416 87821
rect 70000 87752 75416 87819
rect 70000 87105 75416 87172
rect 70000 87049 70047 87105
rect 70103 87049 70171 87105
rect 70227 87049 70295 87105
rect 70351 87049 70419 87105
rect 70475 87094 75416 87105
rect 70475 87049 73866 87094
rect 70000 87038 73866 87049
rect 73922 87038 74008 87094
rect 74064 87038 74150 87094
rect 74206 87038 74292 87094
rect 74348 87038 74434 87094
rect 74490 87038 74576 87094
rect 74632 87038 74718 87094
rect 74774 87038 74860 87094
rect 74916 87038 75002 87094
rect 75058 87038 75144 87094
rect 75200 87038 75286 87094
rect 75342 87038 75416 87094
rect 70000 86981 75416 87038
rect 70000 86925 70047 86981
rect 70103 86925 70171 86981
rect 70227 86925 70295 86981
rect 70351 86925 70419 86981
rect 70475 86952 75416 86981
rect 70475 86925 73866 86952
rect 70000 86896 73866 86925
rect 73922 86896 74008 86952
rect 74064 86896 74150 86952
rect 74206 86896 74292 86952
rect 74348 86896 74434 86952
rect 74490 86896 74576 86952
rect 74632 86896 74718 86952
rect 74774 86896 74860 86952
rect 74916 86896 75002 86952
rect 75058 86896 75144 86952
rect 75200 86896 75286 86952
rect 75342 86896 75416 86952
rect 70000 86857 75416 86896
rect 70000 86801 70047 86857
rect 70103 86801 70171 86857
rect 70227 86801 70295 86857
rect 70351 86801 70419 86857
rect 70475 86810 75416 86857
rect 70475 86801 73866 86810
rect 70000 86754 73866 86801
rect 73922 86754 74008 86810
rect 74064 86754 74150 86810
rect 74206 86754 74292 86810
rect 74348 86754 74434 86810
rect 74490 86754 74576 86810
rect 74632 86754 74718 86810
rect 74774 86754 74860 86810
rect 74916 86754 75002 86810
rect 75058 86754 75144 86810
rect 75200 86754 75286 86810
rect 75342 86754 75416 86810
rect 70000 86733 75416 86754
rect 70000 86677 70047 86733
rect 70103 86677 70171 86733
rect 70227 86677 70295 86733
rect 70351 86677 70419 86733
rect 70475 86677 75416 86733
rect 70000 86668 75416 86677
rect 70000 86612 73866 86668
rect 73922 86612 74008 86668
rect 74064 86612 74150 86668
rect 74206 86612 74292 86668
rect 74348 86612 74434 86668
rect 74490 86612 74576 86668
rect 74632 86612 74718 86668
rect 74774 86612 74860 86668
rect 74916 86612 75002 86668
rect 75058 86612 75144 86668
rect 75200 86612 75286 86668
rect 75342 86612 75416 86668
rect 70000 86609 75416 86612
rect 70000 86553 70047 86609
rect 70103 86553 70171 86609
rect 70227 86553 70295 86609
rect 70351 86553 70419 86609
rect 70475 86553 75416 86609
rect 70000 86526 75416 86553
rect 70000 86485 73866 86526
rect 70000 86429 70047 86485
rect 70103 86429 70171 86485
rect 70227 86429 70295 86485
rect 70351 86429 70419 86485
rect 70475 86470 73866 86485
rect 73922 86470 74008 86526
rect 74064 86470 74150 86526
rect 74206 86470 74292 86526
rect 74348 86470 74434 86526
rect 74490 86470 74576 86526
rect 74632 86470 74718 86526
rect 74774 86470 74860 86526
rect 74916 86470 75002 86526
rect 75058 86470 75144 86526
rect 75200 86470 75286 86526
rect 75342 86470 75416 86526
rect 70475 86429 75416 86470
rect 70000 86384 75416 86429
rect 70000 86361 73866 86384
rect 70000 86305 70047 86361
rect 70103 86305 70171 86361
rect 70227 86305 70295 86361
rect 70351 86305 70419 86361
rect 70475 86328 73866 86361
rect 73922 86328 74008 86384
rect 74064 86328 74150 86384
rect 74206 86328 74292 86384
rect 74348 86328 74434 86384
rect 74490 86328 74576 86384
rect 74632 86328 74718 86384
rect 74774 86328 74860 86384
rect 74916 86328 75002 86384
rect 75058 86328 75144 86384
rect 75200 86328 75286 86384
rect 75342 86328 75416 86384
rect 70475 86305 75416 86328
rect 70000 86242 75416 86305
rect 70000 86237 73866 86242
rect 70000 86181 70047 86237
rect 70103 86181 70171 86237
rect 70227 86181 70295 86237
rect 70351 86181 70419 86237
rect 70475 86186 73866 86237
rect 73922 86186 74008 86242
rect 74064 86186 74150 86242
rect 74206 86186 74292 86242
rect 74348 86186 74434 86242
rect 74490 86186 74576 86242
rect 74632 86186 74718 86242
rect 74774 86186 74860 86242
rect 74916 86186 75002 86242
rect 75058 86186 75144 86242
rect 75200 86186 75286 86242
rect 75342 86186 75416 86242
rect 70475 86181 75416 86186
rect 70000 86113 75416 86181
rect 70000 86057 70047 86113
rect 70103 86057 70171 86113
rect 70227 86057 70295 86113
rect 70351 86057 70419 86113
rect 70475 86100 75416 86113
rect 70475 86057 73866 86100
rect 70000 86044 73866 86057
rect 73922 86044 74008 86100
rect 74064 86044 74150 86100
rect 74206 86044 74292 86100
rect 74348 86044 74434 86100
rect 74490 86044 74576 86100
rect 74632 86044 74718 86100
rect 74774 86044 74860 86100
rect 74916 86044 75002 86100
rect 75058 86044 75144 86100
rect 75200 86044 75286 86100
rect 75342 86044 75416 86100
rect 70000 85989 75416 86044
rect 70000 85933 70047 85989
rect 70103 85933 70171 85989
rect 70227 85933 70295 85989
rect 70351 85933 70419 85989
rect 70475 85958 75416 85989
rect 70475 85933 73866 85958
rect 70000 85902 73866 85933
rect 73922 85902 74008 85958
rect 74064 85902 74150 85958
rect 74206 85902 74292 85958
rect 74348 85902 74434 85958
rect 74490 85902 74576 85958
rect 74632 85902 74718 85958
rect 74774 85902 74860 85958
rect 74916 85902 75002 85958
rect 75058 85902 75144 85958
rect 75200 85902 75286 85958
rect 75342 85902 75416 85958
rect 70000 85865 75416 85902
rect 70000 85809 70047 85865
rect 70103 85809 70171 85865
rect 70227 85809 70295 85865
rect 70351 85809 70419 85865
rect 70475 85816 75416 85865
rect 70475 85809 73866 85816
rect 70000 85760 73866 85809
rect 73922 85760 74008 85816
rect 74064 85760 74150 85816
rect 74206 85760 74292 85816
rect 74348 85760 74434 85816
rect 74490 85760 74576 85816
rect 74632 85760 74718 85816
rect 74774 85760 74860 85816
rect 74916 85760 75002 85816
rect 75058 85760 75144 85816
rect 75200 85760 75286 85816
rect 75342 85760 75416 85816
rect 70000 85741 75416 85760
rect 70000 85685 70047 85741
rect 70103 85685 70171 85741
rect 70227 85685 70295 85741
rect 70351 85685 70419 85741
rect 70475 85685 75416 85741
rect 70000 85674 75416 85685
rect 70000 85618 73866 85674
rect 73922 85618 74008 85674
rect 74064 85618 74150 85674
rect 74206 85618 74292 85674
rect 74348 85618 74434 85674
rect 74490 85618 74576 85674
rect 74632 85618 74718 85674
rect 74774 85618 74860 85674
rect 74916 85618 75002 85674
rect 75058 85618 75144 85674
rect 75200 85618 75286 85674
rect 75342 85618 75416 85674
rect 70000 85617 75416 85618
rect 70000 85561 70047 85617
rect 70103 85561 70171 85617
rect 70227 85561 70295 85617
rect 70351 85561 70419 85617
rect 70475 85561 75416 85617
rect 70000 85532 75416 85561
rect 70000 85493 73866 85532
rect 70000 85437 70047 85493
rect 70103 85437 70171 85493
rect 70227 85437 70295 85493
rect 70351 85437 70419 85493
rect 70475 85476 73866 85493
rect 73922 85476 74008 85532
rect 74064 85476 74150 85532
rect 74206 85476 74292 85532
rect 74348 85476 74434 85532
rect 74490 85476 74576 85532
rect 74632 85476 74718 85532
rect 74774 85476 74860 85532
rect 74916 85476 75002 85532
rect 75058 85476 75144 85532
rect 75200 85476 75286 85532
rect 75342 85476 75416 85532
rect 70475 85437 75416 85476
rect 70000 85390 75416 85437
rect 70000 85369 73866 85390
rect 70000 85313 70047 85369
rect 70103 85313 70171 85369
rect 70227 85313 70295 85369
rect 70351 85313 70419 85369
rect 70475 85334 73866 85369
rect 73922 85334 74008 85390
rect 74064 85334 74150 85390
rect 74206 85334 74292 85390
rect 74348 85334 74434 85390
rect 74490 85334 74576 85390
rect 74632 85334 74718 85390
rect 74774 85334 74860 85390
rect 74916 85334 75002 85390
rect 75058 85334 75144 85390
rect 75200 85334 75286 85390
rect 75342 85334 75416 85390
rect 70475 85313 75416 85334
rect 70000 85272 75416 85313
rect 655272 76035 657172 76088
rect 655272 75979 655343 76035
rect 655399 75979 655485 76035
rect 655541 75979 655627 76035
rect 655683 75979 655769 76035
rect 655825 75979 655911 76035
rect 655967 75979 656053 76035
rect 656109 75979 656195 76035
rect 656251 75979 656337 76035
rect 656393 75979 657172 76035
rect 655272 75945 657172 75979
rect 655272 75889 655326 75945
rect 655382 75893 655450 75945
rect 655506 75893 655574 75945
rect 655630 75893 655698 75945
rect 655399 75889 655450 75893
rect 655541 75889 655574 75893
rect 655683 75889 655698 75893
rect 655754 75893 655822 75945
rect 655878 75893 655946 75945
rect 656002 75893 656070 75945
rect 655754 75889 655769 75893
rect 655878 75889 655911 75893
rect 656002 75889 656053 75893
rect 656126 75889 656194 75945
rect 656250 75893 656318 75945
rect 656374 75893 657172 75945
rect 656251 75889 656318 75893
rect 655272 75837 655343 75889
rect 655399 75837 655485 75889
rect 655541 75837 655627 75889
rect 655683 75837 655769 75889
rect 655825 75837 655911 75889
rect 655967 75837 656053 75889
rect 656109 75837 656195 75889
rect 656251 75837 656337 75889
rect 656393 75837 657172 75893
rect 655272 75821 657172 75837
rect 655272 75765 655326 75821
rect 655382 75765 655450 75821
rect 655506 75765 655574 75821
rect 655630 75765 655698 75821
rect 655754 75765 655822 75821
rect 655878 75765 655946 75821
rect 656002 75765 656070 75821
rect 656126 75765 656194 75821
rect 656250 75765 656318 75821
rect 656374 75765 657172 75821
rect 655272 75751 657172 75765
rect 655272 75697 655343 75751
rect 655399 75697 655485 75751
rect 655541 75697 655627 75751
rect 655683 75697 655769 75751
rect 655825 75697 655911 75751
rect 655967 75697 656053 75751
rect 656109 75697 656195 75751
rect 656251 75697 656337 75751
rect 655272 75641 655326 75697
rect 655399 75695 655450 75697
rect 655541 75695 655574 75697
rect 655683 75695 655698 75697
rect 655382 75641 655450 75695
rect 655506 75641 655574 75695
rect 655630 75641 655698 75695
rect 655754 75695 655769 75697
rect 655878 75695 655911 75697
rect 656002 75695 656053 75697
rect 655754 75641 655822 75695
rect 655878 75641 655946 75695
rect 656002 75641 656070 75695
rect 656126 75641 656194 75697
rect 656251 75695 656318 75697
rect 656393 75695 657172 75751
rect 656250 75641 656318 75695
rect 656374 75641 657172 75695
rect 655272 75609 657172 75641
rect 655272 75573 655343 75609
rect 655399 75573 655485 75609
rect 655541 75573 655627 75609
rect 655683 75573 655769 75609
rect 655825 75573 655911 75609
rect 655967 75573 656053 75609
rect 656109 75573 656195 75609
rect 656251 75573 656337 75609
rect 655272 75517 655326 75573
rect 655399 75553 655450 75573
rect 655541 75553 655574 75573
rect 655683 75553 655698 75573
rect 655382 75517 655450 75553
rect 655506 75517 655574 75553
rect 655630 75517 655698 75553
rect 655754 75553 655769 75573
rect 655878 75553 655911 75573
rect 656002 75553 656053 75573
rect 655754 75517 655822 75553
rect 655878 75517 655946 75553
rect 656002 75517 656070 75553
rect 656126 75517 656194 75573
rect 656251 75553 656318 75573
rect 656393 75553 657172 75609
rect 656250 75517 656318 75553
rect 656374 75517 657172 75553
rect 655272 75467 657172 75517
rect 655272 75449 655343 75467
rect 655399 75449 655485 75467
rect 655541 75449 655627 75467
rect 655683 75449 655769 75467
rect 655825 75449 655911 75467
rect 655967 75449 656053 75467
rect 656109 75449 656195 75467
rect 656251 75449 656337 75467
rect 655272 75393 655326 75449
rect 655399 75411 655450 75449
rect 655541 75411 655574 75449
rect 655683 75411 655698 75449
rect 655382 75393 655450 75411
rect 655506 75393 655574 75411
rect 655630 75393 655698 75411
rect 655754 75411 655769 75449
rect 655878 75411 655911 75449
rect 656002 75411 656053 75449
rect 655754 75393 655822 75411
rect 655878 75393 655946 75411
rect 656002 75393 656070 75411
rect 656126 75393 656194 75449
rect 656251 75411 656318 75449
rect 656393 75411 657172 75467
rect 656250 75393 656318 75411
rect 656374 75393 657172 75411
rect 655272 75325 657172 75393
rect 655272 75269 655326 75325
rect 655399 75269 655450 75325
rect 655541 75269 655574 75325
rect 655683 75269 655698 75325
rect 655754 75269 655769 75325
rect 655878 75269 655911 75325
rect 656002 75269 656053 75325
rect 656126 75269 656194 75325
rect 656251 75269 656318 75325
rect 656393 75269 657172 75325
rect 655272 75201 657172 75269
rect 655272 75145 655326 75201
rect 655382 75183 655450 75201
rect 655506 75183 655574 75201
rect 655630 75183 655698 75201
rect 655399 75145 655450 75183
rect 655541 75145 655574 75183
rect 655683 75145 655698 75183
rect 655754 75183 655822 75201
rect 655878 75183 655946 75201
rect 656002 75183 656070 75201
rect 655754 75145 655769 75183
rect 655878 75145 655911 75183
rect 656002 75145 656053 75183
rect 656126 75145 656194 75201
rect 656250 75183 656318 75201
rect 656374 75183 657172 75201
rect 656251 75145 656318 75183
rect 655272 75127 655343 75145
rect 655399 75127 655485 75145
rect 655541 75127 655627 75145
rect 655683 75127 655769 75145
rect 655825 75127 655911 75145
rect 655967 75127 656053 75145
rect 656109 75127 656195 75145
rect 656251 75127 656337 75145
rect 656393 75127 657172 75183
rect 655272 75077 657172 75127
rect 655272 75021 655326 75077
rect 655382 75041 655450 75077
rect 655506 75041 655574 75077
rect 655630 75041 655698 75077
rect 655399 75021 655450 75041
rect 655541 75021 655574 75041
rect 655683 75021 655698 75041
rect 655754 75041 655822 75077
rect 655878 75041 655946 75077
rect 656002 75041 656070 75077
rect 655754 75021 655769 75041
rect 655878 75021 655911 75041
rect 656002 75021 656053 75041
rect 656126 75021 656194 75077
rect 656250 75041 656318 75077
rect 656374 75041 657172 75077
rect 656251 75021 656318 75041
rect 655272 74985 655343 75021
rect 655399 74985 655485 75021
rect 655541 74985 655627 75021
rect 655683 74985 655769 75021
rect 655825 74985 655911 75021
rect 655967 74985 656053 75021
rect 656109 74985 656195 75021
rect 656251 74985 656337 75021
rect 656393 74985 657172 75041
rect 655272 74953 657172 74985
rect 655272 74897 655326 74953
rect 655382 74899 655450 74953
rect 655506 74899 655574 74953
rect 655630 74899 655698 74953
rect 655399 74897 655450 74899
rect 655541 74897 655574 74899
rect 655683 74897 655698 74899
rect 655754 74899 655822 74953
rect 655878 74899 655946 74953
rect 656002 74899 656070 74953
rect 655754 74897 655769 74899
rect 655878 74897 655911 74899
rect 656002 74897 656053 74899
rect 656126 74897 656194 74953
rect 656250 74899 656318 74953
rect 656374 74899 657172 74953
rect 656251 74897 656318 74899
rect 655272 74843 655343 74897
rect 655399 74843 655485 74897
rect 655541 74843 655627 74897
rect 655683 74843 655769 74897
rect 655825 74843 655911 74897
rect 655967 74843 656053 74897
rect 656109 74843 656195 74897
rect 656251 74843 656337 74897
rect 656393 74843 657172 74899
rect 655272 74829 657172 74843
rect 655272 74773 655326 74829
rect 655382 74773 655450 74829
rect 655506 74773 655574 74829
rect 655630 74773 655698 74829
rect 655754 74773 655822 74829
rect 655878 74773 655946 74829
rect 656002 74773 656070 74829
rect 656126 74773 656194 74829
rect 656250 74773 656318 74829
rect 656374 74773 657172 74829
rect 655272 74757 657172 74773
rect 655272 74705 655343 74757
rect 655399 74705 655485 74757
rect 655541 74705 655627 74757
rect 655683 74705 655769 74757
rect 655825 74705 655911 74757
rect 655967 74705 656053 74757
rect 656109 74705 656195 74757
rect 656251 74705 656337 74757
rect 655272 74649 655326 74705
rect 655399 74701 655450 74705
rect 655541 74701 655574 74705
rect 655683 74701 655698 74705
rect 655382 74649 655450 74701
rect 655506 74649 655574 74701
rect 655630 74649 655698 74701
rect 655754 74701 655769 74705
rect 655878 74701 655911 74705
rect 656002 74701 656053 74705
rect 655754 74649 655822 74701
rect 655878 74649 655946 74701
rect 656002 74649 656070 74701
rect 656126 74649 656194 74705
rect 656251 74701 656318 74705
rect 656393 74701 657172 74757
rect 656250 74649 656318 74701
rect 656374 74649 657172 74701
rect 655272 74615 657172 74649
rect 655272 74581 655343 74615
rect 655399 74581 655485 74615
rect 655541 74581 655627 74615
rect 655683 74581 655769 74615
rect 655825 74581 655911 74615
rect 655967 74581 656053 74615
rect 656109 74581 656195 74615
rect 656251 74581 656337 74615
rect 655272 74525 655326 74581
rect 655399 74559 655450 74581
rect 655541 74559 655574 74581
rect 655683 74559 655698 74581
rect 655382 74525 655450 74559
rect 655506 74525 655574 74559
rect 655630 74525 655698 74559
rect 655754 74559 655769 74581
rect 655878 74559 655911 74581
rect 656002 74559 656053 74581
rect 655754 74525 655822 74559
rect 655878 74525 655946 74559
rect 656002 74525 656070 74559
rect 656126 74525 656194 74581
rect 656251 74559 656318 74581
rect 656393 74559 657172 74615
rect 656250 74525 656318 74559
rect 656374 74525 657172 74559
rect 655272 74488 657172 74525
rect 657752 76035 659802 76088
rect 657752 75979 657823 76035
rect 657879 75979 657965 76035
rect 658021 75979 658107 76035
rect 658163 75979 658249 76035
rect 658305 75979 658391 76035
rect 658447 75979 658533 76035
rect 658589 75979 658675 76035
rect 658731 75979 658817 76035
rect 658873 75979 658959 76035
rect 659015 75979 659101 76035
rect 659157 75979 659243 76035
rect 659299 75979 659385 76035
rect 659441 75979 659527 76035
rect 659583 75979 659669 76035
rect 659725 75979 659802 76035
rect 657752 75945 659802 75979
rect 657752 75889 657806 75945
rect 657862 75893 657930 75945
rect 657986 75893 658054 75945
rect 658110 75893 658178 75945
rect 657879 75889 657930 75893
rect 658021 75889 658054 75893
rect 658163 75889 658178 75893
rect 658234 75893 658302 75945
rect 658358 75893 658426 75945
rect 658482 75893 658550 75945
rect 658234 75889 658249 75893
rect 658358 75889 658391 75893
rect 658482 75889 658533 75893
rect 658606 75889 658674 75945
rect 658730 75893 658798 75945
rect 658854 75893 658922 75945
rect 658978 75893 659046 75945
rect 659102 75893 659170 75945
rect 658731 75889 658798 75893
rect 658873 75889 658922 75893
rect 659015 75889 659046 75893
rect 659157 75889 659170 75893
rect 659226 75893 659294 75945
rect 659350 75893 659418 75945
rect 659474 75893 659542 75945
rect 659226 75889 659243 75893
rect 659350 75889 659385 75893
rect 659474 75889 659527 75893
rect 659598 75889 659666 75945
rect 659722 75893 659802 75945
rect 657752 75837 657823 75889
rect 657879 75837 657965 75889
rect 658021 75837 658107 75889
rect 658163 75837 658249 75889
rect 658305 75837 658391 75889
rect 658447 75837 658533 75889
rect 658589 75837 658675 75889
rect 658731 75837 658817 75889
rect 658873 75837 658959 75889
rect 659015 75837 659101 75889
rect 659157 75837 659243 75889
rect 659299 75837 659385 75889
rect 659441 75837 659527 75889
rect 659583 75837 659669 75889
rect 659725 75837 659802 75893
rect 657752 75821 659802 75837
rect 657752 75765 657806 75821
rect 657862 75765 657930 75821
rect 657986 75765 658054 75821
rect 658110 75765 658178 75821
rect 658234 75765 658302 75821
rect 658358 75765 658426 75821
rect 658482 75765 658550 75821
rect 658606 75765 658674 75821
rect 658730 75765 658798 75821
rect 658854 75765 658922 75821
rect 658978 75765 659046 75821
rect 659102 75765 659170 75821
rect 659226 75765 659294 75821
rect 659350 75765 659418 75821
rect 659474 75765 659542 75821
rect 659598 75765 659666 75821
rect 659722 75765 659802 75821
rect 657752 75751 659802 75765
rect 657752 75697 657823 75751
rect 657879 75697 657965 75751
rect 658021 75697 658107 75751
rect 658163 75697 658249 75751
rect 658305 75697 658391 75751
rect 658447 75697 658533 75751
rect 658589 75697 658675 75751
rect 658731 75697 658817 75751
rect 658873 75697 658959 75751
rect 659015 75697 659101 75751
rect 659157 75697 659243 75751
rect 659299 75697 659385 75751
rect 659441 75697 659527 75751
rect 659583 75697 659669 75751
rect 657752 75641 657806 75697
rect 657879 75695 657930 75697
rect 658021 75695 658054 75697
rect 658163 75695 658178 75697
rect 657862 75641 657930 75695
rect 657986 75641 658054 75695
rect 658110 75641 658178 75695
rect 658234 75695 658249 75697
rect 658358 75695 658391 75697
rect 658482 75695 658533 75697
rect 658234 75641 658302 75695
rect 658358 75641 658426 75695
rect 658482 75641 658550 75695
rect 658606 75641 658674 75697
rect 658731 75695 658798 75697
rect 658873 75695 658922 75697
rect 659015 75695 659046 75697
rect 659157 75695 659170 75697
rect 658730 75641 658798 75695
rect 658854 75641 658922 75695
rect 658978 75641 659046 75695
rect 659102 75641 659170 75695
rect 659226 75695 659243 75697
rect 659350 75695 659385 75697
rect 659474 75695 659527 75697
rect 659226 75641 659294 75695
rect 659350 75641 659418 75695
rect 659474 75641 659542 75695
rect 659598 75641 659666 75697
rect 659725 75695 659802 75751
rect 659722 75641 659802 75695
rect 657752 75609 659802 75641
rect 657752 75573 657823 75609
rect 657879 75573 657965 75609
rect 658021 75573 658107 75609
rect 658163 75573 658249 75609
rect 658305 75573 658391 75609
rect 658447 75573 658533 75609
rect 658589 75573 658675 75609
rect 658731 75573 658817 75609
rect 658873 75573 658959 75609
rect 659015 75573 659101 75609
rect 659157 75573 659243 75609
rect 659299 75573 659385 75609
rect 659441 75573 659527 75609
rect 659583 75573 659669 75609
rect 657752 75517 657806 75573
rect 657879 75553 657930 75573
rect 658021 75553 658054 75573
rect 658163 75553 658178 75573
rect 657862 75517 657930 75553
rect 657986 75517 658054 75553
rect 658110 75517 658178 75553
rect 658234 75553 658249 75573
rect 658358 75553 658391 75573
rect 658482 75553 658533 75573
rect 658234 75517 658302 75553
rect 658358 75517 658426 75553
rect 658482 75517 658550 75553
rect 658606 75517 658674 75573
rect 658731 75553 658798 75573
rect 658873 75553 658922 75573
rect 659015 75553 659046 75573
rect 659157 75553 659170 75573
rect 658730 75517 658798 75553
rect 658854 75517 658922 75553
rect 658978 75517 659046 75553
rect 659102 75517 659170 75553
rect 659226 75553 659243 75573
rect 659350 75553 659385 75573
rect 659474 75553 659527 75573
rect 659226 75517 659294 75553
rect 659350 75517 659418 75553
rect 659474 75517 659542 75553
rect 659598 75517 659666 75573
rect 659725 75553 659802 75609
rect 659722 75517 659802 75553
rect 657752 75467 659802 75517
rect 657752 75449 657823 75467
rect 657879 75449 657965 75467
rect 658021 75449 658107 75467
rect 658163 75449 658249 75467
rect 658305 75449 658391 75467
rect 658447 75449 658533 75467
rect 658589 75449 658675 75467
rect 658731 75449 658817 75467
rect 658873 75449 658959 75467
rect 659015 75449 659101 75467
rect 659157 75449 659243 75467
rect 659299 75449 659385 75467
rect 659441 75449 659527 75467
rect 659583 75449 659669 75467
rect 657752 75393 657806 75449
rect 657879 75411 657930 75449
rect 658021 75411 658054 75449
rect 658163 75411 658178 75449
rect 657862 75393 657930 75411
rect 657986 75393 658054 75411
rect 658110 75393 658178 75411
rect 658234 75411 658249 75449
rect 658358 75411 658391 75449
rect 658482 75411 658533 75449
rect 658234 75393 658302 75411
rect 658358 75393 658426 75411
rect 658482 75393 658550 75411
rect 658606 75393 658674 75449
rect 658731 75411 658798 75449
rect 658873 75411 658922 75449
rect 659015 75411 659046 75449
rect 659157 75411 659170 75449
rect 658730 75393 658798 75411
rect 658854 75393 658922 75411
rect 658978 75393 659046 75411
rect 659102 75393 659170 75411
rect 659226 75411 659243 75449
rect 659350 75411 659385 75449
rect 659474 75411 659527 75449
rect 659226 75393 659294 75411
rect 659350 75393 659418 75411
rect 659474 75393 659542 75411
rect 659598 75393 659666 75449
rect 659725 75411 659802 75467
rect 659722 75393 659802 75411
rect 657752 75325 659802 75393
rect 657752 75269 657806 75325
rect 657879 75269 657930 75325
rect 658021 75269 658054 75325
rect 658163 75269 658178 75325
rect 658234 75269 658249 75325
rect 658358 75269 658391 75325
rect 658482 75269 658533 75325
rect 658606 75269 658674 75325
rect 658731 75269 658798 75325
rect 658873 75269 658922 75325
rect 659015 75269 659046 75325
rect 659157 75269 659170 75325
rect 659226 75269 659243 75325
rect 659350 75269 659385 75325
rect 659474 75269 659527 75325
rect 659598 75269 659666 75325
rect 659725 75269 659802 75325
rect 657752 75201 659802 75269
rect 657752 75145 657806 75201
rect 657862 75183 657930 75201
rect 657986 75183 658054 75201
rect 658110 75183 658178 75201
rect 657879 75145 657930 75183
rect 658021 75145 658054 75183
rect 658163 75145 658178 75183
rect 658234 75183 658302 75201
rect 658358 75183 658426 75201
rect 658482 75183 658550 75201
rect 658234 75145 658249 75183
rect 658358 75145 658391 75183
rect 658482 75145 658533 75183
rect 658606 75145 658674 75201
rect 658730 75183 658798 75201
rect 658854 75183 658922 75201
rect 658978 75183 659046 75201
rect 659102 75183 659170 75201
rect 658731 75145 658798 75183
rect 658873 75145 658922 75183
rect 659015 75145 659046 75183
rect 659157 75145 659170 75183
rect 659226 75183 659294 75201
rect 659350 75183 659418 75201
rect 659474 75183 659542 75201
rect 659226 75145 659243 75183
rect 659350 75145 659385 75183
rect 659474 75145 659527 75183
rect 659598 75145 659666 75201
rect 659722 75183 659802 75201
rect 657752 75127 657823 75145
rect 657879 75127 657965 75145
rect 658021 75127 658107 75145
rect 658163 75127 658249 75145
rect 658305 75127 658391 75145
rect 658447 75127 658533 75145
rect 658589 75127 658675 75145
rect 658731 75127 658817 75145
rect 658873 75127 658959 75145
rect 659015 75127 659101 75145
rect 659157 75127 659243 75145
rect 659299 75127 659385 75145
rect 659441 75127 659527 75145
rect 659583 75127 659669 75145
rect 659725 75127 659802 75183
rect 657752 75077 659802 75127
rect 657752 75021 657806 75077
rect 657862 75041 657930 75077
rect 657986 75041 658054 75077
rect 658110 75041 658178 75077
rect 657879 75021 657930 75041
rect 658021 75021 658054 75041
rect 658163 75021 658178 75041
rect 658234 75041 658302 75077
rect 658358 75041 658426 75077
rect 658482 75041 658550 75077
rect 658234 75021 658249 75041
rect 658358 75021 658391 75041
rect 658482 75021 658533 75041
rect 658606 75021 658674 75077
rect 658730 75041 658798 75077
rect 658854 75041 658922 75077
rect 658978 75041 659046 75077
rect 659102 75041 659170 75077
rect 658731 75021 658798 75041
rect 658873 75021 658922 75041
rect 659015 75021 659046 75041
rect 659157 75021 659170 75041
rect 659226 75041 659294 75077
rect 659350 75041 659418 75077
rect 659474 75041 659542 75077
rect 659226 75021 659243 75041
rect 659350 75021 659385 75041
rect 659474 75021 659527 75041
rect 659598 75021 659666 75077
rect 659722 75041 659802 75077
rect 657752 74985 657823 75021
rect 657879 74985 657965 75021
rect 658021 74985 658107 75021
rect 658163 74985 658249 75021
rect 658305 74985 658391 75021
rect 658447 74985 658533 75021
rect 658589 74985 658675 75021
rect 658731 74985 658817 75021
rect 658873 74985 658959 75021
rect 659015 74985 659101 75021
rect 659157 74985 659243 75021
rect 659299 74985 659385 75021
rect 659441 74985 659527 75021
rect 659583 74985 659669 75021
rect 659725 74985 659802 75041
rect 657752 74953 659802 74985
rect 657752 74897 657806 74953
rect 657862 74899 657930 74953
rect 657986 74899 658054 74953
rect 658110 74899 658178 74953
rect 657879 74897 657930 74899
rect 658021 74897 658054 74899
rect 658163 74897 658178 74899
rect 658234 74899 658302 74953
rect 658358 74899 658426 74953
rect 658482 74899 658550 74953
rect 658234 74897 658249 74899
rect 658358 74897 658391 74899
rect 658482 74897 658533 74899
rect 658606 74897 658674 74953
rect 658730 74899 658798 74953
rect 658854 74899 658922 74953
rect 658978 74899 659046 74953
rect 659102 74899 659170 74953
rect 658731 74897 658798 74899
rect 658873 74897 658922 74899
rect 659015 74897 659046 74899
rect 659157 74897 659170 74899
rect 659226 74899 659294 74953
rect 659350 74899 659418 74953
rect 659474 74899 659542 74953
rect 659226 74897 659243 74899
rect 659350 74897 659385 74899
rect 659474 74897 659527 74899
rect 659598 74897 659666 74953
rect 659722 74899 659802 74953
rect 657752 74843 657823 74897
rect 657879 74843 657965 74897
rect 658021 74843 658107 74897
rect 658163 74843 658249 74897
rect 658305 74843 658391 74897
rect 658447 74843 658533 74897
rect 658589 74843 658675 74897
rect 658731 74843 658817 74897
rect 658873 74843 658959 74897
rect 659015 74843 659101 74897
rect 659157 74843 659243 74897
rect 659299 74843 659385 74897
rect 659441 74843 659527 74897
rect 659583 74843 659669 74897
rect 659725 74843 659802 74899
rect 657752 74829 659802 74843
rect 657752 74773 657806 74829
rect 657862 74773 657930 74829
rect 657986 74773 658054 74829
rect 658110 74773 658178 74829
rect 658234 74773 658302 74829
rect 658358 74773 658426 74829
rect 658482 74773 658550 74829
rect 658606 74773 658674 74829
rect 658730 74773 658798 74829
rect 658854 74773 658922 74829
rect 658978 74773 659046 74829
rect 659102 74773 659170 74829
rect 659226 74773 659294 74829
rect 659350 74773 659418 74829
rect 659474 74773 659542 74829
rect 659598 74773 659666 74829
rect 659722 74773 659802 74829
rect 657752 74757 659802 74773
rect 657752 74705 657823 74757
rect 657879 74705 657965 74757
rect 658021 74705 658107 74757
rect 658163 74705 658249 74757
rect 658305 74705 658391 74757
rect 658447 74705 658533 74757
rect 658589 74705 658675 74757
rect 658731 74705 658817 74757
rect 658873 74705 658959 74757
rect 659015 74705 659101 74757
rect 659157 74705 659243 74757
rect 659299 74705 659385 74757
rect 659441 74705 659527 74757
rect 659583 74705 659669 74757
rect 657752 74649 657806 74705
rect 657879 74701 657930 74705
rect 658021 74701 658054 74705
rect 658163 74701 658178 74705
rect 657862 74649 657930 74701
rect 657986 74649 658054 74701
rect 658110 74649 658178 74701
rect 658234 74701 658249 74705
rect 658358 74701 658391 74705
rect 658482 74701 658533 74705
rect 658234 74649 658302 74701
rect 658358 74649 658426 74701
rect 658482 74649 658550 74701
rect 658606 74649 658674 74705
rect 658731 74701 658798 74705
rect 658873 74701 658922 74705
rect 659015 74701 659046 74705
rect 659157 74701 659170 74705
rect 658730 74649 658798 74701
rect 658854 74649 658922 74701
rect 658978 74649 659046 74701
rect 659102 74649 659170 74701
rect 659226 74701 659243 74705
rect 659350 74701 659385 74705
rect 659474 74701 659527 74705
rect 659226 74649 659294 74701
rect 659350 74649 659418 74701
rect 659474 74649 659542 74701
rect 659598 74649 659666 74705
rect 659725 74701 659802 74757
rect 659722 74649 659802 74701
rect 657752 74615 659802 74649
rect 657752 74581 657823 74615
rect 657879 74581 657965 74615
rect 658021 74581 658107 74615
rect 658163 74581 658249 74615
rect 658305 74581 658391 74615
rect 658447 74581 658533 74615
rect 658589 74581 658675 74615
rect 658731 74581 658817 74615
rect 658873 74581 658959 74615
rect 659015 74581 659101 74615
rect 659157 74581 659243 74615
rect 659299 74581 659385 74615
rect 659441 74581 659527 74615
rect 659583 74581 659669 74615
rect 657752 74525 657806 74581
rect 657879 74559 657930 74581
rect 658021 74559 658054 74581
rect 658163 74559 658178 74581
rect 657862 74525 657930 74559
rect 657986 74525 658054 74559
rect 658110 74525 658178 74559
rect 658234 74559 658249 74581
rect 658358 74559 658391 74581
rect 658482 74559 658533 74581
rect 658234 74525 658302 74559
rect 658358 74525 658426 74559
rect 658482 74525 658550 74559
rect 658606 74525 658674 74581
rect 658731 74559 658798 74581
rect 658873 74559 658922 74581
rect 659015 74559 659046 74581
rect 659157 74559 659170 74581
rect 658730 74525 658798 74559
rect 658854 74525 658922 74559
rect 658978 74525 659046 74559
rect 659102 74525 659170 74559
rect 659226 74559 659243 74581
rect 659350 74559 659385 74581
rect 659474 74559 659527 74581
rect 659226 74525 659294 74559
rect 659350 74525 659418 74559
rect 659474 74525 659542 74559
rect 659598 74525 659666 74581
rect 659725 74559 659802 74615
rect 659722 74525 659802 74559
rect 657752 74488 659802 74525
rect 660122 76035 662172 76088
rect 660122 75979 660193 76035
rect 660249 75979 660335 76035
rect 660391 75979 660477 76035
rect 660533 75979 660619 76035
rect 660675 75979 660761 76035
rect 660817 75979 660903 76035
rect 660959 75979 661045 76035
rect 661101 75979 661187 76035
rect 661243 75979 661329 76035
rect 661385 75979 661471 76035
rect 661527 75979 661613 76035
rect 661669 75979 661755 76035
rect 661811 75979 661897 76035
rect 661953 75979 662039 76035
rect 662095 75979 662172 76035
rect 660122 75945 662172 75979
rect 660122 75889 660176 75945
rect 660232 75893 660300 75945
rect 660356 75893 660424 75945
rect 660480 75893 660548 75945
rect 660249 75889 660300 75893
rect 660391 75889 660424 75893
rect 660533 75889 660548 75893
rect 660604 75893 660672 75945
rect 660728 75893 660796 75945
rect 660852 75893 660920 75945
rect 660604 75889 660619 75893
rect 660728 75889 660761 75893
rect 660852 75889 660903 75893
rect 660976 75889 661044 75945
rect 661100 75893 661168 75945
rect 661224 75893 661292 75945
rect 661348 75893 661416 75945
rect 661472 75893 661540 75945
rect 661101 75889 661168 75893
rect 661243 75889 661292 75893
rect 661385 75889 661416 75893
rect 661527 75889 661540 75893
rect 661596 75893 661664 75945
rect 661720 75893 661788 75945
rect 661844 75893 661912 75945
rect 661596 75889 661613 75893
rect 661720 75889 661755 75893
rect 661844 75889 661897 75893
rect 661968 75889 662036 75945
rect 662092 75893 662172 75945
rect 660122 75837 660193 75889
rect 660249 75837 660335 75889
rect 660391 75837 660477 75889
rect 660533 75837 660619 75889
rect 660675 75837 660761 75889
rect 660817 75837 660903 75889
rect 660959 75837 661045 75889
rect 661101 75837 661187 75889
rect 661243 75837 661329 75889
rect 661385 75837 661471 75889
rect 661527 75837 661613 75889
rect 661669 75837 661755 75889
rect 661811 75837 661897 75889
rect 661953 75837 662039 75889
rect 662095 75837 662172 75893
rect 660122 75821 662172 75837
rect 660122 75765 660176 75821
rect 660232 75765 660300 75821
rect 660356 75765 660424 75821
rect 660480 75765 660548 75821
rect 660604 75765 660672 75821
rect 660728 75765 660796 75821
rect 660852 75765 660920 75821
rect 660976 75765 661044 75821
rect 661100 75765 661168 75821
rect 661224 75765 661292 75821
rect 661348 75765 661416 75821
rect 661472 75765 661540 75821
rect 661596 75765 661664 75821
rect 661720 75765 661788 75821
rect 661844 75765 661912 75821
rect 661968 75765 662036 75821
rect 662092 75765 662172 75821
rect 660122 75751 662172 75765
rect 660122 75697 660193 75751
rect 660249 75697 660335 75751
rect 660391 75697 660477 75751
rect 660533 75697 660619 75751
rect 660675 75697 660761 75751
rect 660817 75697 660903 75751
rect 660959 75697 661045 75751
rect 661101 75697 661187 75751
rect 661243 75697 661329 75751
rect 661385 75697 661471 75751
rect 661527 75697 661613 75751
rect 661669 75697 661755 75751
rect 661811 75697 661897 75751
rect 661953 75697 662039 75751
rect 660122 75641 660176 75697
rect 660249 75695 660300 75697
rect 660391 75695 660424 75697
rect 660533 75695 660548 75697
rect 660232 75641 660300 75695
rect 660356 75641 660424 75695
rect 660480 75641 660548 75695
rect 660604 75695 660619 75697
rect 660728 75695 660761 75697
rect 660852 75695 660903 75697
rect 660604 75641 660672 75695
rect 660728 75641 660796 75695
rect 660852 75641 660920 75695
rect 660976 75641 661044 75697
rect 661101 75695 661168 75697
rect 661243 75695 661292 75697
rect 661385 75695 661416 75697
rect 661527 75695 661540 75697
rect 661100 75641 661168 75695
rect 661224 75641 661292 75695
rect 661348 75641 661416 75695
rect 661472 75641 661540 75695
rect 661596 75695 661613 75697
rect 661720 75695 661755 75697
rect 661844 75695 661897 75697
rect 661596 75641 661664 75695
rect 661720 75641 661788 75695
rect 661844 75641 661912 75695
rect 661968 75641 662036 75697
rect 662095 75695 662172 75751
rect 662092 75641 662172 75695
rect 660122 75609 662172 75641
rect 660122 75573 660193 75609
rect 660249 75573 660335 75609
rect 660391 75573 660477 75609
rect 660533 75573 660619 75609
rect 660675 75573 660761 75609
rect 660817 75573 660903 75609
rect 660959 75573 661045 75609
rect 661101 75573 661187 75609
rect 661243 75573 661329 75609
rect 661385 75573 661471 75609
rect 661527 75573 661613 75609
rect 661669 75573 661755 75609
rect 661811 75573 661897 75609
rect 661953 75573 662039 75609
rect 660122 75517 660176 75573
rect 660249 75553 660300 75573
rect 660391 75553 660424 75573
rect 660533 75553 660548 75573
rect 660232 75517 660300 75553
rect 660356 75517 660424 75553
rect 660480 75517 660548 75553
rect 660604 75553 660619 75573
rect 660728 75553 660761 75573
rect 660852 75553 660903 75573
rect 660604 75517 660672 75553
rect 660728 75517 660796 75553
rect 660852 75517 660920 75553
rect 660976 75517 661044 75573
rect 661101 75553 661168 75573
rect 661243 75553 661292 75573
rect 661385 75553 661416 75573
rect 661527 75553 661540 75573
rect 661100 75517 661168 75553
rect 661224 75517 661292 75553
rect 661348 75517 661416 75553
rect 661472 75517 661540 75553
rect 661596 75553 661613 75573
rect 661720 75553 661755 75573
rect 661844 75553 661897 75573
rect 661596 75517 661664 75553
rect 661720 75517 661788 75553
rect 661844 75517 661912 75553
rect 661968 75517 662036 75573
rect 662095 75553 662172 75609
rect 662092 75517 662172 75553
rect 660122 75467 662172 75517
rect 660122 75449 660193 75467
rect 660249 75449 660335 75467
rect 660391 75449 660477 75467
rect 660533 75449 660619 75467
rect 660675 75449 660761 75467
rect 660817 75449 660903 75467
rect 660959 75449 661045 75467
rect 661101 75449 661187 75467
rect 661243 75449 661329 75467
rect 661385 75449 661471 75467
rect 661527 75449 661613 75467
rect 661669 75449 661755 75467
rect 661811 75449 661897 75467
rect 661953 75449 662039 75467
rect 660122 75393 660176 75449
rect 660249 75411 660300 75449
rect 660391 75411 660424 75449
rect 660533 75411 660548 75449
rect 660232 75393 660300 75411
rect 660356 75393 660424 75411
rect 660480 75393 660548 75411
rect 660604 75411 660619 75449
rect 660728 75411 660761 75449
rect 660852 75411 660903 75449
rect 660604 75393 660672 75411
rect 660728 75393 660796 75411
rect 660852 75393 660920 75411
rect 660976 75393 661044 75449
rect 661101 75411 661168 75449
rect 661243 75411 661292 75449
rect 661385 75411 661416 75449
rect 661527 75411 661540 75449
rect 661100 75393 661168 75411
rect 661224 75393 661292 75411
rect 661348 75393 661416 75411
rect 661472 75393 661540 75411
rect 661596 75411 661613 75449
rect 661720 75411 661755 75449
rect 661844 75411 661897 75449
rect 661596 75393 661664 75411
rect 661720 75393 661788 75411
rect 661844 75393 661912 75411
rect 661968 75393 662036 75449
rect 662095 75411 662172 75467
rect 662092 75393 662172 75411
rect 660122 75325 662172 75393
rect 660122 75269 660176 75325
rect 660249 75269 660300 75325
rect 660391 75269 660424 75325
rect 660533 75269 660548 75325
rect 660604 75269 660619 75325
rect 660728 75269 660761 75325
rect 660852 75269 660903 75325
rect 660976 75269 661044 75325
rect 661101 75269 661168 75325
rect 661243 75269 661292 75325
rect 661385 75269 661416 75325
rect 661527 75269 661540 75325
rect 661596 75269 661613 75325
rect 661720 75269 661755 75325
rect 661844 75269 661897 75325
rect 661968 75269 662036 75325
rect 662095 75269 662172 75325
rect 660122 75201 662172 75269
rect 660122 75145 660176 75201
rect 660232 75183 660300 75201
rect 660356 75183 660424 75201
rect 660480 75183 660548 75201
rect 660249 75145 660300 75183
rect 660391 75145 660424 75183
rect 660533 75145 660548 75183
rect 660604 75183 660672 75201
rect 660728 75183 660796 75201
rect 660852 75183 660920 75201
rect 660604 75145 660619 75183
rect 660728 75145 660761 75183
rect 660852 75145 660903 75183
rect 660976 75145 661044 75201
rect 661100 75183 661168 75201
rect 661224 75183 661292 75201
rect 661348 75183 661416 75201
rect 661472 75183 661540 75201
rect 661101 75145 661168 75183
rect 661243 75145 661292 75183
rect 661385 75145 661416 75183
rect 661527 75145 661540 75183
rect 661596 75183 661664 75201
rect 661720 75183 661788 75201
rect 661844 75183 661912 75201
rect 661596 75145 661613 75183
rect 661720 75145 661755 75183
rect 661844 75145 661897 75183
rect 661968 75145 662036 75201
rect 662092 75183 662172 75201
rect 660122 75127 660193 75145
rect 660249 75127 660335 75145
rect 660391 75127 660477 75145
rect 660533 75127 660619 75145
rect 660675 75127 660761 75145
rect 660817 75127 660903 75145
rect 660959 75127 661045 75145
rect 661101 75127 661187 75145
rect 661243 75127 661329 75145
rect 661385 75127 661471 75145
rect 661527 75127 661613 75145
rect 661669 75127 661755 75145
rect 661811 75127 661897 75145
rect 661953 75127 662039 75145
rect 662095 75127 662172 75183
rect 660122 75077 662172 75127
rect 660122 75021 660176 75077
rect 660232 75041 660300 75077
rect 660356 75041 660424 75077
rect 660480 75041 660548 75077
rect 660249 75021 660300 75041
rect 660391 75021 660424 75041
rect 660533 75021 660548 75041
rect 660604 75041 660672 75077
rect 660728 75041 660796 75077
rect 660852 75041 660920 75077
rect 660604 75021 660619 75041
rect 660728 75021 660761 75041
rect 660852 75021 660903 75041
rect 660976 75021 661044 75077
rect 661100 75041 661168 75077
rect 661224 75041 661292 75077
rect 661348 75041 661416 75077
rect 661472 75041 661540 75077
rect 661101 75021 661168 75041
rect 661243 75021 661292 75041
rect 661385 75021 661416 75041
rect 661527 75021 661540 75041
rect 661596 75041 661664 75077
rect 661720 75041 661788 75077
rect 661844 75041 661912 75077
rect 661596 75021 661613 75041
rect 661720 75021 661755 75041
rect 661844 75021 661897 75041
rect 661968 75021 662036 75077
rect 662092 75041 662172 75077
rect 660122 74985 660193 75021
rect 660249 74985 660335 75021
rect 660391 74985 660477 75021
rect 660533 74985 660619 75021
rect 660675 74985 660761 75021
rect 660817 74985 660903 75021
rect 660959 74985 661045 75021
rect 661101 74985 661187 75021
rect 661243 74985 661329 75021
rect 661385 74985 661471 75021
rect 661527 74985 661613 75021
rect 661669 74985 661755 75021
rect 661811 74985 661897 75021
rect 661953 74985 662039 75021
rect 662095 74985 662172 75041
rect 660122 74953 662172 74985
rect 660122 74897 660176 74953
rect 660232 74899 660300 74953
rect 660356 74899 660424 74953
rect 660480 74899 660548 74953
rect 660249 74897 660300 74899
rect 660391 74897 660424 74899
rect 660533 74897 660548 74899
rect 660604 74899 660672 74953
rect 660728 74899 660796 74953
rect 660852 74899 660920 74953
rect 660604 74897 660619 74899
rect 660728 74897 660761 74899
rect 660852 74897 660903 74899
rect 660976 74897 661044 74953
rect 661100 74899 661168 74953
rect 661224 74899 661292 74953
rect 661348 74899 661416 74953
rect 661472 74899 661540 74953
rect 661101 74897 661168 74899
rect 661243 74897 661292 74899
rect 661385 74897 661416 74899
rect 661527 74897 661540 74899
rect 661596 74899 661664 74953
rect 661720 74899 661788 74953
rect 661844 74899 661912 74953
rect 661596 74897 661613 74899
rect 661720 74897 661755 74899
rect 661844 74897 661897 74899
rect 661968 74897 662036 74953
rect 662092 74899 662172 74953
rect 660122 74843 660193 74897
rect 660249 74843 660335 74897
rect 660391 74843 660477 74897
rect 660533 74843 660619 74897
rect 660675 74843 660761 74897
rect 660817 74843 660903 74897
rect 660959 74843 661045 74897
rect 661101 74843 661187 74897
rect 661243 74843 661329 74897
rect 661385 74843 661471 74897
rect 661527 74843 661613 74897
rect 661669 74843 661755 74897
rect 661811 74843 661897 74897
rect 661953 74843 662039 74897
rect 662095 74843 662172 74899
rect 660122 74829 662172 74843
rect 660122 74773 660176 74829
rect 660232 74773 660300 74829
rect 660356 74773 660424 74829
rect 660480 74773 660548 74829
rect 660604 74773 660672 74829
rect 660728 74773 660796 74829
rect 660852 74773 660920 74829
rect 660976 74773 661044 74829
rect 661100 74773 661168 74829
rect 661224 74773 661292 74829
rect 661348 74773 661416 74829
rect 661472 74773 661540 74829
rect 661596 74773 661664 74829
rect 661720 74773 661788 74829
rect 661844 74773 661912 74829
rect 661968 74773 662036 74829
rect 662092 74773 662172 74829
rect 660122 74757 662172 74773
rect 660122 74705 660193 74757
rect 660249 74705 660335 74757
rect 660391 74705 660477 74757
rect 660533 74705 660619 74757
rect 660675 74705 660761 74757
rect 660817 74705 660903 74757
rect 660959 74705 661045 74757
rect 661101 74705 661187 74757
rect 661243 74705 661329 74757
rect 661385 74705 661471 74757
rect 661527 74705 661613 74757
rect 661669 74705 661755 74757
rect 661811 74705 661897 74757
rect 661953 74705 662039 74757
rect 660122 74649 660176 74705
rect 660249 74701 660300 74705
rect 660391 74701 660424 74705
rect 660533 74701 660548 74705
rect 660232 74649 660300 74701
rect 660356 74649 660424 74701
rect 660480 74649 660548 74701
rect 660604 74701 660619 74705
rect 660728 74701 660761 74705
rect 660852 74701 660903 74705
rect 660604 74649 660672 74701
rect 660728 74649 660796 74701
rect 660852 74649 660920 74701
rect 660976 74649 661044 74705
rect 661101 74701 661168 74705
rect 661243 74701 661292 74705
rect 661385 74701 661416 74705
rect 661527 74701 661540 74705
rect 661100 74649 661168 74701
rect 661224 74649 661292 74701
rect 661348 74649 661416 74701
rect 661472 74649 661540 74701
rect 661596 74701 661613 74705
rect 661720 74701 661755 74705
rect 661844 74701 661897 74705
rect 661596 74649 661664 74701
rect 661720 74649 661788 74701
rect 661844 74649 661912 74701
rect 661968 74649 662036 74705
rect 662095 74701 662172 74757
rect 662092 74649 662172 74701
rect 660122 74615 662172 74649
rect 660122 74581 660193 74615
rect 660249 74581 660335 74615
rect 660391 74581 660477 74615
rect 660533 74581 660619 74615
rect 660675 74581 660761 74615
rect 660817 74581 660903 74615
rect 660959 74581 661045 74615
rect 661101 74581 661187 74615
rect 661243 74581 661329 74615
rect 661385 74581 661471 74615
rect 661527 74581 661613 74615
rect 661669 74581 661755 74615
rect 661811 74581 661897 74615
rect 661953 74581 662039 74615
rect 660122 74525 660176 74581
rect 660249 74559 660300 74581
rect 660391 74559 660424 74581
rect 660533 74559 660548 74581
rect 660232 74525 660300 74559
rect 660356 74525 660424 74559
rect 660480 74525 660548 74559
rect 660604 74559 660619 74581
rect 660728 74559 660761 74581
rect 660852 74559 660903 74581
rect 660604 74525 660672 74559
rect 660728 74525 660796 74559
rect 660852 74525 660920 74559
rect 660976 74525 661044 74581
rect 661101 74559 661168 74581
rect 661243 74559 661292 74581
rect 661385 74559 661416 74581
rect 661527 74559 661540 74581
rect 661100 74525 661168 74559
rect 661224 74525 661292 74559
rect 661348 74525 661416 74559
rect 661472 74525 661540 74559
rect 661596 74559 661613 74581
rect 661720 74559 661755 74581
rect 661844 74559 661897 74581
rect 661596 74525 661664 74559
rect 661720 74525 661788 74559
rect 661844 74525 661912 74559
rect 661968 74525 662036 74581
rect 662095 74559 662172 74615
rect 662092 74525 662172 74559
rect 660122 74488 662172 74525
rect 662828 76035 664878 76088
rect 662828 75979 662899 76035
rect 662955 75979 663041 76035
rect 663097 75979 663183 76035
rect 663239 75979 663325 76035
rect 663381 75979 663467 76035
rect 663523 75979 663609 76035
rect 663665 75979 663751 76035
rect 663807 75979 663893 76035
rect 663949 75979 664035 76035
rect 664091 75979 664177 76035
rect 664233 75979 664319 76035
rect 664375 75979 664461 76035
rect 664517 75979 664603 76035
rect 664659 75979 664745 76035
rect 664801 75979 664878 76035
rect 662828 75945 664878 75979
rect 662828 75889 662882 75945
rect 662938 75893 663006 75945
rect 663062 75893 663130 75945
rect 663186 75893 663254 75945
rect 662955 75889 663006 75893
rect 663097 75889 663130 75893
rect 663239 75889 663254 75893
rect 663310 75893 663378 75945
rect 663434 75893 663502 75945
rect 663558 75893 663626 75945
rect 663310 75889 663325 75893
rect 663434 75889 663467 75893
rect 663558 75889 663609 75893
rect 663682 75889 663750 75945
rect 663806 75893 663874 75945
rect 663930 75893 663998 75945
rect 664054 75893 664122 75945
rect 664178 75893 664246 75945
rect 663807 75889 663874 75893
rect 663949 75889 663998 75893
rect 664091 75889 664122 75893
rect 664233 75889 664246 75893
rect 664302 75893 664370 75945
rect 664426 75893 664494 75945
rect 664550 75893 664618 75945
rect 664302 75889 664319 75893
rect 664426 75889 664461 75893
rect 664550 75889 664603 75893
rect 664674 75889 664742 75945
rect 664798 75893 664878 75945
rect 662828 75837 662899 75889
rect 662955 75837 663041 75889
rect 663097 75837 663183 75889
rect 663239 75837 663325 75889
rect 663381 75837 663467 75889
rect 663523 75837 663609 75889
rect 663665 75837 663751 75889
rect 663807 75837 663893 75889
rect 663949 75837 664035 75889
rect 664091 75837 664177 75889
rect 664233 75837 664319 75889
rect 664375 75837 664461 75889
rect 664517 75837 664603 75889
rect 664659 75837 664745 75889
rect 664801 75837 664878 75893
rect 662828 75821 664878 75837
rect 662828 75765 662882 75821
rect 662938 75765 663006 75821
rect 663062 75765 663130 75821
rect 663186 75765 663254 75821
rect 663310 75765 663378 75821
rect 663434 75765 663502 75821
rect 663558 75765 663626 75821
rect 663682 75765 663750 75821
rect 663806 75765 663874 75821
rect 663930 75765 663998 75821
rect 664054 75765 664122 75821
rect 664178 75765 664246 75821
rect 664302 75765 664370 75821
rect 664426 75765 664494 75821
rect 664550 75765 664618 75821
rect 664674 75765 664742 75821
rect 664798 75765 664878 75821
rect 662828 75751 664878 75765
rect 662828 75697 662899 75751
rect 662955 75697 663041 75751
rect 663097 75697 663183 75751
rect 663239 75697 663325 75751
rect 663381 75697 663467 75751
rect 663523 75697 663609 75751
rect 663665 75697 663751 75751
rect 663807 75697 663893 75751
rect 663949 75697 664035 75751
rect 664091 75697 664177 75751
rect 664233 75697 664319 75751
rect 664375 75697 664461 75751
rect 664517 75697 664603 75751
rect 664659 75697 664745 75751
rect 662828 75641 662882 75697
rect 662955 75695 663006 75697
rect 663097 75695 663130 75697
rect 663239 75695 663254 75697
rect 662938 75641 663006 75695
rect 663062 75641 663130 75695
rect 663186 75641 663254 75695
rect 663310 75695 663325 75697
rect 663434 75695 663467 75697
rect 663558 75695 663609 75697
rect 663310 75641 663378 75695
rect 663434 75641 663502 75695
rect 663558 75641 663626 75695
rect 663682 75641 663750 75697
rect 663807 75695 663874 75697
rect 663949 75695 663998 75697
rect 664091 75695 664122 75697
rect 664233 75695 664246 75697
rect 663806 75641 663874 75695
rect 663930 75641 663998 75695
rect 664054 75641 664122 75695
rect 664178 75641 664246 75695
rect 664302 75695 664319 75697
rect 664426 75695 664461 75697
rect 664550 75695 664603 75697
rect 664302 75641 664370 75695
rect 664426 75641 664494 75695
rect 664550 75641 664618 75695
rect 664674 75641 664742 75697
rect 664801 75695 664878 75751
rect 664798 75641 664878 75695
rect 662828 75609 664878 75641
rect 662828 75573 662899 75609
rect 662955 75573 663041 75609
rect 663097 75573 663183 75609
rect 663239 75573 663325 75609
rect 663381 75573 663467 75609
rect 663523 75573 663609 75609
rect 663665 75573 663751 75609
rect 663807 75573 663893 75609
rect 663949 75573 664035 75609
rect 664091 75573 664177 75609
rect 664233 75573 664319 75609
rect 664375 75573 664461 75609
rect 664517 75573 664603 75609
rect 664659 75573 664745 75609
rect 662828 75517 662882 75573
rect 662955 75553 663006 75573
rect 663097 75553 663130 75573
rect 663239 75553 663254 75573
rect 662938 75517 663006 75553
rect 663062 75517 663130 75553
rect 663186 75517 663254 75553
rect 663310 75553 663325 75573
rect 663434 75553 663467 75573
rect 663558 75553 663609 75573
rect 663310 75517 663378 75553
rect 663434 75517 663502 75553
rect 663558 75517 663626 75553
rect 663682 75517 663750 75573
rect 663807 75553 663874 75573
rect 663949 75553 663998 75573
rect 664091 75553 664122 75573
rect 664233 75553 664246 75573
rect 663806 75517 663874 75553
rect 663930 75517 663998 75553
rect 664054 75517 664122 75553
rect 664178 75517 664246 75553
rect 664302 75553 664319 75573
rect 664426 75553 664461 75573
rect 664550 75553 664603 75573
rect 664302 75517 664370 75553
rect 664426 75517 664494 75553
rect 664550 75517 664618 75553
rect 664674 75517 664742 75573
rect 664801 75553 664878 75609
rect 664798 75517 664878 75553
rect 662828 75467 664878 75517
rect 662828 75449 662899 75467
rect 662955 75449 663041 75467
rect 663097 75449 663183 75467
rect 663239 75449 663325 75467
rect 663381 75449 663467 75467
rect 663523 75449 663609 75467
rect 663665 75449 663751 75467
rect 663807 75449 663893 75467
rect 663949 75449 664035 75467
rect 664091 75449 664177 75467
rect 664233 75449 664319 75467
rect 664375 75449 664461 75467
rect 664517 75449 664603 75467
rect 664659 75449 664745 75467
rect 662828 75393 662882 75449
rect 662955 75411 663006 75449
rect 663097 75411 663130 75449
rect 663239 75411 663254 75449
rect 662938 75393 663006 75411
rect 663062 75393 663130 75411
rect 663186 75393 663254 75411
rect 663310 75411 663325 75449
rect 663434 75411 663467 75449
rect 663558 75411 663609 75449
rect 663310 75393 663378 75411
rect 663434 75393 663502 75411
rect 663558 75393 663626 75411
rect 663682 75393 663750 75449
rect 663807 75411 663874 75449
rect 663949 75411 663998 75449
rect 664091 75411 664122 75449
rect 664233 75411 664246 75449
rect 663806 75393 663874 75411
rect 663930 75393 663998 75411
rect 664054 75393 664122 75411
rect 664178 75393 664246 75411
rect 664302 75411 664319 75449
rect 664426 75411 664461 75449
rect 664550 75411 664603 75449
rect 664302 75393 664370 75411
rect 664426 75393 664494 75411
rect 664550 75393 664618 75411
rect 664674 75393 664742 75449
rect 664801 75411 664878 75467
rect 664798 75393 664878 75411
rect 662828 75325 664878 75393
rect 662828 75269 662882 75325
rect 662955 75269 663006 75325
rect 663097 75269 663130 75325
rect 663239 75269 663254 75325
rect 663310 75269 663325 75325
rect 663434 75269 663467 75325
rect 663558 75269 663609 75325
rect 663682 75269 663750 75325
rect 663807 75269 663874 75325
rect 663949 75269 663998 75325
rect 664091 75269 664122 75325
rect 664233 75269 664246 75325
rect 664302 75269 664319 75325
rect 664426 75269 664461 75325
rect 664550 75269 664603 75325
rect 664674 75269 664742 75325
rect 664801 75269 664878 75325
rect 662828 75201 664878 75269
rect 662828 75145 662882 75201
rect 662938 75183 663006 75201
rect 663062 75183 663130 75201
rect 663186 75183 663254 75201
rect 662955 75145 663006 75183
rect 663097 75145 663130 75183
rect 663239 75145 663254 75183
rect 663310 75183 663378 75201
rect 663434 75183 663502 75201
rect 663558 75183 663626 75201
rect 663310 75145 663325 75183
rect 663434 75145 663467 75183
rect 663558 75145 663609 75183
rect 663682 75145 663750 75201
rect 663806 75183 663874 75201
rect 663930 75183 663998 75201
rect 664054 75183 664122 75201
rect 664178 75183 664246 75201
rect 663807 75145 663874 75183
rect 663949 75145 663998 75183
rect 664091 75145 664122 75183
rect 664233 75145 664246 75183
rect 664302 75183 664370 75201
rect 664426 75183 664494 75201
rect 664550 75183 664618 75201
rect 664302 75145 664319 75183
rect 664426 75145 664461 75183
rect 664550 75145 664603 75183
rect 664674 75145 664742 75201
rect 664798 75183 664878 75201
rect 662828 75127 662899 75145
rect 662955 75127 663041 75145
rect 663097 75127 663183 75145
rect 663239 75127 663325 75145
rect 663381 75127 663467 75145
rect 663523 75127 663609 75145
rect 663665 75127 663751 75145
rect 663807 75127 663893 75145
rect 663949 75127 664035 75145
rect 664091 75127 664177 75145
rect 664233 75127 664319 75145
rect 664375 75127 664461 75145
rect 664517 75127 664603 75145
rect 664659 75127 664745 75145
rect 664801 75127 664878 75183
rect 662828 75077 664878 75127
rect 662828 75021 662882 75077
rect 662938 75041 663006 75077
rect 663062 75041 663130 75077
rect 663186 75041 663254 75077
rect 662955 75021 663006 75041
rect 663097 75021 663130 75041
rect 663239 75021 663254 75041
rect 663310 75041 663378 75077
rect 663434 75041 663502 75077
rect 663558 75041 663626 75077
rect 663310 75021 663325 75041
rect 663434 75021 663467 75041
rect 663558 75021 663609 75041
rect 663682 75021 663750 75077
rect 663806 75041 663874 75077
rect 663930 75041 663998 75077
rect 664054 75041 664122 75077
rect 664178 75041 664246 75077
rect 663807 75021 663874 75041
rect 663949 75021 663998 75041
rect 664091 75021 664122 75041
rect 664233 75021 664246 75041
rect 664302 75041 664370 75077
rect 664426 75041 664494 75077
rect 664550 75041 664618 75077
rect 664302 75021 664319 75041
rect 664426 75021 664461 75041
rect 664550 75021 664603 75041
rect 664674 75021 664742 75077
rect 664798 75041 664878 75077
rect 662828 74985 662899 75021
rect 662955 74985 663041 75021
rect 663097 74985 663183 75021
rect 663239 74985 663325 75021
rect 663381 74985 663467 75021
rect 663523 74985 663609 75021
rect 663665 74985 663751 75021
rect 663807 74985 663893 75021
rect 663949 74985 664035 75021
rect 664091 74985 664177 75021
rect 664233 74985 664319 75021
rect 664375 74985 664461 75021
rect 664517 74985 664603 75021
rect 664659 74985 664745 75021
rect 664801 74985 664878 75041
rect 662828 74953 664878 74985
rect 662828 74897 662882 74953
rect 662938 74899 663006 74953
rect 663062 74899 663130 74953
rect 663186 74899 663254 74953
rect 662955 74897 663006 74899
rect 663097 74897 663130 74899
rect 663239 74897 663254 74899
rect 663310 74899 663378 74953
rect 663434 74899 663502 74953
rect 663558 74899 663626 74953
rect 663310 74897 663325 74899
rect 663434 74897 663467 74899
rect 663558 74897 663609 74899
rect 663682 74897 663750 74953
rect 663806 74899 663874 74953
rect 663930 74899 663998 74953
rect 664054 74899 664122 74953
rect 664178 74899 664246 74953
rect 663807 74897 663874 74899
rect 663949 74897 663998 74899
rect 664091 74897 664122 74899
rect 664233 74897 664246 74899
rect 664302 74899 664370 74953
rect 664426 74899 664494 74953
rect 664550 74899 664618 74953
rect 664302 74897 664319 74899
rect 664426 74897 664461 74899
rect 664550 74897 664603 74899
rect 664674 74897 664742 74953
rect 664798 74899 664878 74953
rect 662828 74843 662899 74897
rect 662955 74843 663041 74897
rect 663097 74843 663183 74897
rect 663239 74843 663325 74897
rect 663381 74843 663467 74897
rect 663523 74843 663609 74897
rect 663665 74843 663751 74897
rect 663807 74843 663893 74897
rect 663949 74843 664035 74897
rect 664091 74843 664177 74897
rect 664233 74843 664319 74897
rect 664375 74843 664461 74897
rect 664517 74843 664603 74897
rect 664659 74843 664745 74897
rect 664801 74843 664878 74899
rect 662828 74829 664878 74843
rect 662828 74773 662882 74829
rect 662938 74773 663006 74829
rect 663062 74773 663130 74829
rect 663186 74773 663254 74829
rect 663310 74773 663378 74829
rect 663434 74773 663502 74829
rect 663558 74773 663626 74829
rect 663682 74773 663750 74829
rect 663806 74773 663874 74829
rect 663930 74773 663998 74829
rect 664054 74773 664122 74829
rect 664178 74773 664246 74829
rect 664302 74773 664370 74829
rect 664426 74773 664494 74829
rect 664550 74773 664618 74829
rect 664674 74773 664742 74829
rect 664798 74773 664878 74829
rect 662828 74757 664878 74773
rect 662828 74705 662899 74757
rect 662955 74705 663041 74757
rect 663097 74705 663183 74757
rect 663239 74705 663325 74757
rect 663381 74705 663467 74757
rect 663523 74705 663609 74757
rect 663665 74705 663751 74757
rect 663807 74705 663893 74757
rect 663949 74705 664035 74757
rect 664091 74705 664177 74757
rect 664233 74705 664319 74757
rect 664375 74705 664461 74757
rect 664517 74705 664603 74757
rect 664659 74705 664745 74757
rect 662828 74649 662882 74705
rect 662955 74701 663006 74705
rect 663097 74701 663130 74705
rect 663239 74701 663254 74705
rect 662938 74649 663006 74701
rect 663062 74649 663130 74701
rect 663186 74649 663254 74701
rect 663310 74701 663325 74705
rect 663434 74701 663467 74705
rect 663558 74701 663609 74705
rect 663310 74649 663378 74701
rect 663434 74649 663502 74701
rect 663558 74649 663626 74701
rect 663682 74649 663750 74705
rect 663807 74701 663874 74705
rect 663949 74701 663998 74705
rect 664091 74701 664122 74705
rect 664233 74701 664246 74705
rect 663806 74649 663874 74701
rect 663930 74649 663998 74701
rect 664054 74649 664122 74701
rect 664178 74649 664246 74701
rect 664302 74701 664319 74705
rect 664426 74701 664461 74705
rect 664550 74701 664603 74705
rect 664302 74649 664370 74701
rect 664426 74649 664494 74701
rect 664550 74649 664618 74701
rect 664674 74649 664742 74705
rect 664801 74701 664878 74757
rect 664798 74649 664878 74701
rect 662828 74615 664878 74649
rect 662828 74581 662899 74615
rect 662955 74581 663041 74615
rect 663097 74581 663183 74615
rect 663239 74581 663325 74615
rect 663381 74581 663467 74615
rect 663523 74581 663609 74615
rect 663665 74581 663751 74615
rect 663807 74581 663893 74615
rect 663949 74581 664035 74615
rect 664091 74581 664177 74615
rect 664233 74581 664319 74615
rect 664375 74581 664461 74615
rect 664517 74581 664603 74615
rect 664659 74581 664745 74615
rect 662828 74525 662882 74581
rect 662955 74559 663006 74581
rect 663097 74559 663130 74581
rect 663239 74559 663254 74581
rect 662938 74525 663006 74559
rect 663062 74525 663130 74559
rect 663186 74525 663254 74559
rect 663310 74559 663325 74581
rect 663434 74559 663467 74581
rect 663558 74559 663609 74581
rect 663310 74525 663378 74559
rect 663434 74525 663502 74559
rect 663558 74525 663626 74559
rect 663682 74525 663750 74581
rect 663807 74559 663874 74581
rect 663949 74559 663998 74581
rect 664091 74559 664122 74581
rect 664233 74559 664246 74581
rect 663806 74525 663874 74559
rect 663930 74525 663998 74559
rect 664054 74525 664122 74559
rect 664178 74525 664246 74559
rect 664302 74559 664319 74581
rect 664426 74559 664461 74581
rect 664550 74559 664603 74581
rect 664302 74525 664370 74559
rect 664426 74525 664494 74559
rect 664550 74525 664618 74559
rect 664674 74525 664742 74581
rect 664801 74559 664878 74615
rect 664798 74525 664878 74559
rect 662828 74488 664878 74525
rect 665198 76035 667248 76088
rect 665198 75979 665269 76035
rect 665325 75979 665411 76035
rect 665467 75979 665553 76035
rect 665609 75979 665695 76035
rect 665751 75979 665837 76035
rect 665893 75979 665979 76035
rect 666035 75979 666121 76035
rect 666177 75979 666263 76035
rect 666319 75979 666405 76035
rect 666461 75979 666547 76035
rect 666603 75979 666689 76035
rect 666745 75979 666831 76035
rect 666887 75979 666973 76035
rect 667029 75979 667115 76035
rect 667171 75979 667248 76035
rect 665198 75945 667248 75979
rect 665198 75889 665252 75945
rect 665308 75893 665376 75945
rect 665432 75893 665500 75945
rect 665556 75893 665624 75945
rect 665325 75889 665376 75893
rect 665467 75889 665500 75893
rect 665609 75889 665624 75893
rect 665680 75893 665748 75945
rect 665804 75893 665872 75945
rect 665928 75893 665996 75945
rect 665680 75889 665695 75893
rect 665804 75889 665837 75893
rect 665928 75889 665979 75893
rect 666052 75889 666120 75945
rect 666176 75893 666244 75945
rect 666300 75893 666368 75945
rect 666424 75893 666492 75945
rect 666548 75893 666616 75945
rect 666177 75889 666244 75893
rect 666319 75889 666368 75893
rect 666461 75889 666492 75893
rect 666603 75889 666616 75893
rect 666672 75893 666740 75945
rect 666796 75893 666864 75945
rect 666920 75893 666988 75945
rect 666672 75889 666689 75893
rect 666796 75889 666831 75893
rect 666920 75889 666973 75893
rect 667044 75889 667112 75945
rect 667168 75893 667248 75945
rect 665198 75837 665269 75889
rect 665325 75837 665411 75889
rect 665467 75837 665553 75889
rect 665609 75837 665695 75889
rect 665751 75837 665837 75889
rect 665893 75837 665979 75889
rect 666035 75837 666121 75889
rect 666177 75837 666263 75889
rect 666319 75837 666405 75889
rect 666461 75837 666547 75889
rect 666603 75837 666689 75889
rect 666745 75837 666831 75889
rect 666887 75837 666973 75889
rect 667029 75837 667115 75889
rect 667171 75837 667248 75893
rect 665198 75821 667248 75837
rect 665198 75765 665252 75821
rect 665308 75765 665376 75821
rect 665432 75765 665500 75821
rect 665556 75765 665624 75821
rect 665680 75765 665748 75821
rect 665804 75765 665872 75821
rect 665928 75765 665996 75821
rect 666052 75765 666120 75821
rect 666176 75765 666244 75821
rect 666300 75765 666368 75821
rect 666424 75765 666492 75821
rect 666548 75765 666616 75821
rect 666672 75765 666740 75821
rect 666796 75765 666864 75821
rect 666920 75765 666988 75821
rect 667044 75765 667112 75821
rect 667168 75765 667248 75821
rect 665198 75751 667248 75765
rect 665198 75697 665269 75751
rect 665325 75697 665411 75751
rect 665467 75697 665553 75751
rect 665609 75697 665695 75751
rect 665751 75697 665837 75751
rect 665893 75697 665979 75751
rect 666035 75697 666121 75751
rect 666177 75697 666263 75751
rect 666319 75697 666405 75751
rect 666461 75697 666547 75751
rect 666603 75697 666689 75751
rect 666745 75697 666831 75751
rect 666887 75697 666973 75751
rect 667029 75697 667115 75751
rect 665198 75641 665252 75697
rect 665325 75695 665376 75697
rect 665467 75695 665500 75697
rect 665609 75695 665624 75697
rect 665308 75641 665376 75695
rect 665432 75641 665500 75695
rect 665556 75641 665624 75695
rect 665680 75695 665695 75697
rect 665804 75695 665837 75697
rect 665928 75695 665979 75697
rect 665680 75641 665748 75695
rect 665804 75641 665872 75695
rect 665928 75641 665996 75695
rect 666052 75641 666120 75697
rect 666177 75695 666244 75697
rect 666319 75695 666368 75697
rect 666461 75695 666492 75697
rect 666603 75695 666616 75697
rect 666176 75641 666244 75695
rect 666300 75641 666368 75695
rect 666424 75641 666492 75695
rect 666548 75641 666616 75695
rect 666672 75695 666689 75697
rect 666796 75695 666831 75697
rect 666920 75695 666973 75697
rect 666672 75641 666740 75695
rect 666796 75641 666864 75695
rect 666920 75641 666988 75695
rect 667044 75641 667112 75697
rect 667171 75695 667248 75751
rect 667168 75641 667248 75695
rect 665198 75609 667248 75641
rect 665198 75573 665269 75609
rect 665325 75573 665411 75609
rect 665467 75573 665553 75609
rect 665609 75573 665695 75609
rect 665751 75573 665837 75609
rect 665893 75573 665979 75609
rect 666035 75573 666121 75609
rect 666177 75573 666263 75609
rect 666319 75573 666405 75609
rect 666461 75573 666547 75609
rect 666603 75573 666689 75609
rect 666745 75573 666831 75609
rect 666887 75573 666973 75609
rect 667029 75573 667115 75609
rect 665198 75517 665252 75573
rect 665325 75553 665376 75573
rect 665467 75553 665500 75573
rect 665609 75553 665624 75573
rect 665308 75517 665376 75553
rect 665432 75517 665500 75553
rect 665556 75517 665624 75553
rect 665680 75553 665695 75573
rect 665804 75553 665837 75573
rect 665928 75553 665979 75573
rect 665680 75517 665748 75553
rect 665804 75517 665872 75553
rect 665928 75517 665996 75553
rect 666052 75517 666120 75573
rect 666177 75553 666244 75573
rect 666319 75553 666368 75573
rect 666461 75553 666492 75573
rect 666603 75553 666616 75573
rect 666176 75517 666244 75553
rect 666300 75517 666368 75553
rect 666424 75517 666492 75553
rect 666548 75517 666616 75553
rect 666672 75553 666689 75573
rect 666796 75553 666831 75573
rect 666920 75553 666973 75573
rect 666672 75517 666740 75553
rect 666796 75517 666864 75553
rect 666920 75517 666988 75553
rect 667044 75517 667112 75573
rect 667171 75553 667248 75609
rect 667168 75517 667248 75553
rect 665198 75467 667248 75517
rect 665198 75449 665269 75467
rect 665325 75449 665411 75467
rect 665467 75449 665553 75467
rect 665609 75449 665695 75467
rect 665751 75449 665837 75467
rect 665893 75449 665979 75467
rect 666035 75449 666121 75467
rect 666177 75449 666263 75467
rect 666319 75449 666405 75467
rect 666461 75449 666547 75467
rect 666603 75449 666689 75467
rect 666745 75449 666831 75467
rect 666887 75449 666973 75467
rect 667029 75449 667115 75467
rect 665198 75393 665252 75449
rect 665325 75411 665376 75449
rect 665467 75411 665500 75449
rect 665609 75411 665624 75449
rect 665308 75393 665376 75411
rect 665432 75393 665500 75411
rect 665556 75393 665624 75411
rect 665680 75411 665695 75449
rect 665804 75411 665837 75449
rect 665928 75411 665979 75449
rect 665680 75393 665748 75411
rect 665804 75393 665872 75411
rect 665928 75393 665996 75411
rect 666052 75393 666120 75449
rect 666177 75411 666244 75449
rect 666319 75411 666368 75449
rect 666461 75411 666492 75449
rect 666603 75411 666616 75449
rect 666176 75393 666244 75411
rect 666300 75393 666368 75411
rect 666424 75393 666492 75411
rect 666548 75393 666616 75411
rect 666672 75411 666689 75449
rect 666796 75411 666831 75449
rect 666920 75411 666973 75449
rect 666672 75393 666740 75411
rect 666796 75393 666864 75411
rect 666920 75393 666988 75411
rect 667044 75393 667112 75449
rect 667171 75411 667248 75467
rect 667168 75393 667248 75411
rect 665198 75325 667248 75393
rect 665198 75269 665252 75325
rect 665325 75269 665376 75325
rect 665467 75269 665500 75325
rect 665609 75269 665624 75325
rect 665680 75269 665695 75325
rect 665804 75269 665837 75325
rect 665928 75269 665979 75325
rect 666052 75269 666120 75325
rect 666177 75269 666244 75325
rect 666319 75269 666368 75325
rect 666461 75269 666492 75325
rect 666603 75269 666616 75325
rect 666672 75269 666689 75325
rect 666796 75269 666831 75325
rect 666920 75269 666973 75325
rect 667044 75269 667112 75325
rect 667171 75269 667248 75325
rect 665198 75201 667248 75269
rect 665198 75145 665252 75201
rect 665308 75183 665376 75201
rect 665432 75183 665500 75201
rect 665556 75183 665624 75201
rect 665325 75145 665376 75183
rect 665467 75145 665500 75183
rect 665609 75145 665624 75183
rect 665680 75183 665748 75201
rect 665804 75183 665872 75201
rect 665928 75183 665996 75201
rect 665680 75145 665695 75183
rect 665804 75145 665837 75183
rect 665928 75145 665979 75183
rect 666052 75145 666120 75201
rect 666176 75183 666244 75201
rect 666300 75183 666368 75201
rect 666424 75183 666492 75201
rect 666548 75183 666616 75201
rect 666177 75145 666244 75183
rect 666319 75145 666368 75183
rect 666461 75145 666492 75183
rect 666603 75145 666616 75183
rect 666672 75183 666740 75201
rect 666796 75183 666864 75201
rect 666920 75183 666988 75201
rect 666672 75145 666689 75183
rect 666796 75145 666831 75183
rect 666920 75145 666973 75183
rect 667044 75145 667112 75201
rect 667168 75183 667248 75201
rect 665198 75127 665269 75145
rect 665325 75127 665411 75145
rect 665467 75127 665553 75145
rect 665609 75127 665695 75145
rect 665751 75127 665837 75145
rect 665893 75127 665979 75145
rect 666035 75127 666121 75145
rect 666177 75127 666263 75145
rect 666319 75127 666405 75145
rect 666461 75127 666547 75145
rect 666603 75127 666689 75145
rect 666745 75127 666831 75145
rect 666887 75127 666973 75145
rect 667029 75127 667115 75145
rect 667171 75127 667248 75183
rect 665198 75077 667248 75127
rect 665198 75021 665252 75077
rect 665308 75041 665376 75077
rect 665432 75041 665500 75077
rect 665556 75041 665624 75077
rect 665325 75021 665376 75041
rect 665467 75021 665500 75041
rect 665609 75021 665624 75041
rect 665680 75041 665748 75077
rect 665804 75041 665872 75077
rect 665928 75041 665996 75077
rect 665680 75021 665695 75041
rect 665804 75021 665837 75041
rect 665928 75021 665979 75041
rect 666052 75021 666120 75077
rect 666176 75041 666244 75077
rect 666300 75041 666368 75077
rect 666424 75041 666492 75077
rect 666548 75041 666616 75077
rect 666177 75021 666244 75041
rect 666319 75021 666368 75041
rect 666461 75021 666492 75041
rect 666603 75021 666616 75041
rect 666672 75041 666740 75077
rect 666796 75041 666864 75077
rect 666920 75041 666988 75077
rect 666672 75021 666689 75041
rect 666796 75021 666831 75041
rect 666920 75021 666973 75041
rect 667044 75021 667112 75077
rect 667168 75041 667248 75077
rect 665198 74985 665269 75021
rect 665325 74985 665411 75021
rect 665467 74985 665553 75021
rect 665609 74985 665695 75021
rect 665751 74985 665837 75021
rect 665893 74985 665979 75021
rect 666035 74985 666121 75021
rect 666177 74985 666263 75021
rect 666319 74985 666405 75021
rect 666461 74985 666547 75021
rect 666603 74985 666689 75021
rect 666745 74985 666831 75021
rect 666887 74985 666973 75021
rect 667029 74985 667115 75021
rect 667171 74985 667248 75041
rect 665198 74953 667248 74985
rect 665198 74897 665252 74953
rect 665308 74899 665376 74953
rect 665432 74899 665500 74953
rect 665556 74899 665624 74953
rect 665325 74897 665376 74899
rect 665467 74897 665500 74899
rect 665609 74897 665624 74899
rect 665680 74899 665748 74953
rect 665804 74899 665872 74953
rect 665928 74899 665996 74953
rect 665680 74897 665695 74899
rect 665804 74897 665837 74899
rect 665928 74897 665979 74899
rect 666052 74897 666120 74953
rect 666176 74899 666244 74953
rect 666300 74899 666368 74953
rect 666424 74899 666492 74953
rect 666548 74899 666616 74953
rect 666177 74897 666244 74899
rect 666319 74897 666368 74899
rect 666461 74897 666492 74899
rect 666603 74897 666616 74899
rect 666672 74899 666740 74953
rect 666796 74899 666864 74953
rect 666920 74899 666988 74953
rect 666672 74897 666689 74899
rect 666796 74897 666831 74899
rect 666920 74897 666973 74899
rect 667044 74897 667112 74953
rect 667168 74899 667248 74953
rect 665198 74843 665269 74897
rect 665325 74843 665411 74897
rect 665467 74843 665553 74897
rect 665609 74843 665695 74897
rect 665751 74843 665837 74897
rect 665893 74843 665979 74897
rect 666035 74843 666121 74897
rect 666177 74843 666263 74897
rect 666319 74843 666405 74897
rect 666461 74843 666547 74897
rect 666603 74843 666689 74897
rect 666745 74843 666831 74897
rect 666887 74843 666973 74897
rect 667029 74843 667115 74897
rect 667171 74843 667248 74899
rect 665198 74829 667248 74843
rect 665198 74773 665252 74829
rect 665308 74773 665376 74829
rect 665432 74773 665500 74829
rect 665556 74773 665624 74829
rect 665680 74773 665748 74829
rect 665804 74773 665872 74829
rect 665928 74773 665996 74829
rect 666052 74773 666120 74829
rect 666176 74773 666244 74829
rect 666300 74773 666368 74829
rect 666424 74773 666492 74829
rect 666548 74773 666616 74829
rect 666672 74773 666740 74829
rect 666796 74773 666864 74829
rect 666920 74773 666988 74829
rect 667044 74773 667112 74829
rect 667168 74773 667248 74829
rect 665198 74757 667248 74773
rect 665198 74705 665269 74757
rect 665325 74705 665411 74757
rect 665467 74705 665553 74757
rect 665609 74705 665695 74757
rect 665751 74705 665837 74757
rect 665893 74705 665979 74757
rect 666035 74705 666121 74757
rect 666177 74705 666263 74757
rect 666319 74705 666405 74757
rect 666461 74705 666547 74757
rect 666603 74705 666689 74757
rect 666745 74705 666831 74757
rect 666887 74705 666973 74757
rect 667029 74705 667115 74757
rect 665198 74649 665252 74705
rect 665325 74701 665376 74705
rect 665467 74701 665500 74705
rect 665609 74701 665624 74705
rect 665308 74649 665376 74701
rect 665432 74649 665500 74701
rect 665556 74649 665624 74701
rect 665680 74701 665695 74705
rect 665804 74701 665837 74705
rect 665928 74701 665979 74705
rect 665680 74649 665748 74701
rect 665804 74649 665872 74701
rect 665928 74649 665996 74701
rect 666052 74649 666120 74705
rect 666177 74701 666244 74705
rect 666319 74701 666368 74705
rect 666461 74701 666492 74705
rect 666603 74701 666616 74705
rect 666176 74649 666244 74701
rect 666300 74649 666368 74701
rect 666424 74649 666492 74701
rect 666548 74649 666616 74701
rect 666672 74701 666689 74705
rect 666796 74701 666831 74705
rect 666920 74701 666973 74705
rect 666672 74649 666740 74701
rect 666796 74649 666864 74701
rect 666920 74649 666988 74701
rect 667044 74649 667112 74705
rect 667171 74701 667248 74757
rect 667168 74649 667248 74701
rect 665198 74615 667248 74649
rect 665198 74581 665269 74615
rect 665325 74581 665411 74615
rect 665467 74581 665553 74615
rect 665609 74581 665695 74615
rect 665751 74581 665837 74615
rect 665893 74581 665979 74615
rect 666035 74581 666121 74615
rect 666177 74581 666263 74615
rect 666319 74581 666405 74615
rect 666461 74581 666547 74615
rect 666603 74581 666689 74615
rect 666745 74581 666831 74615
rect 666887 74581 666973 74615
rect 667029 74581 667115 74615
rect 665198 74525 665252 74581
rect 665325 74559 665376 74581
rect 665467 74559 665500 74581
rect 665609 74559 665624 74581
rect 665308 74525 665376 74559
rect 665432 74525 665500 74559
rect 665556 74525 665624 74559
rect 665680 74559 665695 74581
rect 665804 74559 665837 74581
rect 665928 74559 665979 74581
rect 665680 74525 665748 74559
rect 665804 74525 665872 74559
rect 665928 74525 665996 74559
rect 666052 74525 666120 74581
rect 666177 74559 666244 74581
rect 666319 74559 666368 74581
rect 666461 74559 666492 74581
rect 666603 74559 666616 74581
rect 666176 74525 666244 74559
rect 666300 74525 666368 74559
rect 666424 74525 666492 74559
rect 666548 74525 666616 74559
rect 666672 74559 666689 74581
rect 666796 74559 666831 74581
rect 666920 74559 666973 74581
rect 666672 74525 666740 74559
rect 666796 74525 666864 74559
rect 666920 74525 666988 74559
rect 667044 74525 667112 74581
rect 667171 74559 667248 74615
rect 667168 74525 667248 74559
rect 665198 74488 667248 74525
rect 667828 76035 669728 76088
rect 667828 75979 667899 76035
rect 667955 75979 668041 76035
rect 668097 75979 668183 76035
rect 668239 75979 668325 76035
rect 668381 75979 668467 76035
rect 668523 75979 668609 76035
rect 668665 75979 668751 76035
rect 668807 75979 668893 76035
rect 668949 75979 669035 76035
rect 669091 75979 669177 76035
rect 669233 75979 669319 76035
rect 669375 75979 669461 76035
rect 669517 75979 669603 76035
rect 669659 75979 669728 76035
rect 667828 75945 669728 75979
rect 667828 75889 667882 75945
rect 667938 75893 668006 75945
rect 668062 75893 668130 75945
rect 668186 75893 668254 75945
rect 667955 75889 668006 75893
rect 668097 75889 668130 75893
rect 668239 75889 668254 75893
rect 668310 75893 668378 75945
rect 668434 75893 668502 75945
rect 668558 75893 668626 75945
rect 668310 75889 668325 75893
rect 668434 75889 668467 75893
rect 668558 75889 668609 75893
rect 668682 75889 668750 75945
rect 668806 75893 668874 75945
rect 668930 75893 668998 75945
rect 669054 75893 669122 75945
rect 669178 75893 669246 75945
rect 668807 75889 668874 75893
rect 668949 75889 668998 75893
rect 669091 75889 669122 75893
rect 669233 75889 669246 75893
rect 669302 75893 669370 75945
rect 669426 75893 669494 75945
rect 669550 75893 669618 75945
rect 669302 75889 669319 75893
rect 669426 75889 669461 75893
rect 669550 75889 669603 75893
rect 669674 75889 669728 75945
rect 667828 75837 667899 75889
rect 667955 75837 668041 75889
rect 668097 75837 668183 75889
rect 668239 75837 668325 75889
rect 668381 75837 668467 75889
rect 668523 75837 668609 75889
rect 668665 75837 668751 75889
rect 668807 75837 668893 75889
rect 668949 75837 669035 75889
rect 669091 75837 669177 75889
rect 669233 75837 669319 75889
rect 669375 75837 669461 75889
rect 669517 75837 669603 75889
rect 669659 75837 669728 75889
rect 667828 75821 669728 75837
rect 667828 75765 667882 75821
rect 667938 75765 668006 75821
rect 668062 75765 668130 75821
rect 668186 75765 668254 75821
rect 668310 75765 668378 75821
rect 668434 75765 668502 75821
rect 668558 75765 668626 75821
rect 668682 75765 668750 75821
rect 668806 75765 668874 75821
rect 668930 75765 668998 75821
rect 669054 75765 669122 75821
rect 669178 75765 669246 75821
rect 669302 75765 669370 75821
rect 669426 75765 669494 75821
rect 669550 75765 669618 75821
rect 669674 75765 669728 75821
rect 667828 75751 669728 75765
rect 667828 75697 667899 75751
rect 667955 75697 668041 75751
rect 668097 75697 668183 75751
rect 668239 75697 668325 75751
rect 668381 75697 668467 75751
rect 668523 75697 668609 75751
rect 668665 75697 668751 75751
rect 668807 75697 668893 75751
rect 668949 75697 669035 75751
rect 669091 75697 669177 75751
rect 669233 75697 669319 75751
rect 669375 75697 669461 75751
rect 669517 75697 669603 75751
rect 669659 75697 669728 75751
rect 667828 75641 667882 75697
rect 667955 75695 668006 75697
rect 668097 75695 668130 75697
rect 668239 75695 668254 75697
rect 667938 75641 668006 75695
rect 668062 75641 668130 75695
rect 668186 75641 668254 75695
rect 668310 75695 668325 75697
rect 668434 75695 668467 75697
rect 668558 75695 668609 75697
rect 668310 75641 668378 75695
rect 668434 75641 668502 75695
rect 668558 75641 668626 75695
rect 668682 75641 668750 75697
rect 668807 75695 668874 75697
rect 668949 75695 668998 75697
rect 669091 75695 669122 75697
rect 669233 75695 669246 75697
rect 668806 75641 668874 75695
rect 668930 75641 668998 75695
rect 669054 75641 669122 75695
rect 669178 75641 669246 75695
rect 669302 75695 669319 75697
rect 669426 75695 669461 75697
rect 669550 75695 669603 75697
rect 669302 75641 669370 75695
rect 669426 75641 669494 75695
rect 669550 75641 669618 75695
rect 669674 75641 669728 75697
rect 667828 75609 669728 75641
rect 667828 75573 667899 75609
rect 667955 75573 668041 75609
rect 668097 75573 668183 75609
rect 668239 75573 668325 75609
rect 668381 75573 668467 75609
rect 668523 75573 668609 75609
rect 668665 75573 668751 75609
rect 668807 75573 668893 75609
rect 668949 75573 669035 75609
rect 669091 75573 669177 75609
rect 669233 75573 669319 75609
rect 669375 75573 669461 75609
rect 669517 75573 669603 75609
rect 669659 75573 669728 75609
rect 667828 75517 667882 75573
rect 667955 75553 668006 75573
rect 668097 75553 668130 75573
rect 668239 75553 668254 75573
rect 667938 75517 668006 75553
rect 668062 75517 668130 75553
rect 668186 75517 668254 75553
rect 668310 75553 668325 75573
rect 668434 75553 668467 75573
rect 668558 75553 668609 75573
rect 668310 75517 668378 75553
rect 668434 75517 668502 75553
rect 668558 75517 668626 75553
rect 668682 75517 668750 75573
rect 668807 75553 668874 75573
rect 668949 75553 668998 75573
rect 669091 75553 669122 75573
rect 669233 75553 669246 75573
rect 668806 75517 668874 75553
rect 668930 75517 668998 75553
rect 669054 75517 669122 75553
rect 669178 75517 669246 75553
rect 669302 75553 669319 75573
rect 669426 75553 669461 75573
rect 669550 75553 669603 75573
rect 669302 75517 669370 75553
rect 669426 75517 669494 75553
rect 669550 75517 669618 75553
rect 669674 75517 669728 75573
rect 667828 75467 669728 75517
rect 667828 75449 667899 75467
rect 667955 75449 668041 75467
rect 668097 75449 668183 75467
rect 668239 75449 668325 75467
rect 668381 75449 668467 75467
rect 668523 75449 668609 75467
rect 668665 75449 668751 75467
rect 668807 75449 668893 75467
rect 668949 75449 669035 75467
rect 669091 75449 669177 75467
rect 669233 75449 669319 75467
rect 669375 75449 669461 75467
rect 669517 75449 669603 75467
rect 669659 75449 669728 75467
rect 667828 75393 667882 75449
rect 667955 75411 668006 75449
rect 668097 75411 668130 75449
rect 668239 75411 668254 75449
rect 667938 75393 668006 75411
rect 668062 75393 668130 75411
rect 668186 75393 668254 75411
rect 668310 75411 668325 75449
rect 668434 75411 668467 75449
rect 668558 75411 668609 75449
rect 668310 75393 668378 75411
rect 668434 75393 668502 75411
rect 668558 75393 668626 75411
rect 668682 75393 668750 75449
rect 668807 75411 668874 75449
rect 668949 75411 668998 75449
rect 669091 75411 669122 75449
rect 669233 75411 669246 75449
rect 668806 75393 668874 75411
rect 668930 75393 668998 75411
rect 669054 75393 669122 75411
rect 669178 75393 669246 75411
rect 669302 75411 669319 75449
rect 669426 75411 669461 75449
rect 669550 75411 669603 75449
rect 669302 75393 669370 75411
rect 669426 75393 669494 75411
rect 669550 75393 669618 75411
rect 669674 75393 669728 75449
rect 667828 75325 669728 75393
rect 667828 75269 667882 75325
rect 667955 75269 668006 75325
rect 668097 75269 668130 75325
rect 668239 75269 668254 75325
rect 668310 75269 668325 75325
rect 668434 75269 668467 75325
rect 668558 75269 668609 75325
rect 668682 75269 668750 75325
rect 668807 75269 668874 75325
rect 668949 75269 668998 75325
rect 669091 75269 669122 75325
rect 669233 75269 669246 75325
rect 669302 75269 669319 75325
rect 669426 75269 669461 75325
rect 669550 75269 669603 75325
rect 669674 75269 669728 75325
rect 667828 75201 669728 75269
rect 667828 75145 667882 75201
rect 667938 75183 668006 75201
rect 668062 75183 668130 75201
rect 668186 75183 668254 75201
rect 667955 75145 668006 75183
rect 668097 75145 668130 75183
rect 668239 75145 668254 75183
rect 668310 75183 668378 75201
rect 668434 75183 668502 75201
rect 668558 75183 668626 75201
rect 668310 75145 668325 75183
rect 668434 75145 668467 75183
rect 668558 75145 668609 75183
rect 668682 75145 668750 75201
rect 668806 75183 668874 75201
rect 668930 75183 668998 75201
rect 669054 75183 669122 75201
rect 669178 75183 669246 75201
rect 668807 75145 668874 75183
rect 668949 75145 668998 75183
rect 669091 75145 669122 75183
rect 669233 75145 669246 75183
rect 669302 75183 669370 75201
rect 669426 75183 669494 75201
rect 669550 75183 669618 75201
rect 669302 75145 669319 75183
rect 669426 75145 669461 75183
rect 669550 75145 669603 75183
rect 669674 75145 669728 75201
rect 667828 75127 667899 75145
rect 667955 75127 668041 75145
rect 668097 75127 668183 75145
rect 668239 75127 668325 75145
rect 668381 75127 668467 75145
rect 668523 75127 668609 75145
rect 668665 75127 668751 75145
rect 668807 75127 668893 75145
rect 668949 75127 669035 75145
rect 669091 75127 669177 75145
rect 669233 75127 669319 75145
rect 669375 75127 669461 75145
rect 669517 75127 669603 75145
rect 669659 75127 669728 75145
rect 667828 75077 669728 75127
rect 667828 75021 667882 75077
rect 667938 75041 668006 75077
rect 668062 75041 668130 75077
rect 668186 75041 668254 75077
rect 667955 75021 668006 75041
rect 668097 75021 668130 75041
rect 668239 75021 668254 75041
rect 668310 75041 668378 75077
rect 668434 75041 668502 75077
rect 668558 75041 668626 75077
rect 668310 75021 668325 75041
rect 668434 75021 668467 75041
rect 668558 75021 668609 75041
rect 668682 75021 668750 75077
rect 668806 75041 668874 75077
rect 668930 75041 668998 75077
rect 669054 75041 669122 75077
rect 669178 75041 669246 75077
rect 668807 75021 668874 75041
rect 668949 75021 668998 75041
rect 669091 75021 669122 75041
rect 669233 75021 669246 75041
rect 669302 75041 669370 75077
rect 669426 75041 669494 75077
rect 669550 75041 669618 75077
rect 669302 75021 669319 75041
rect 669426 75021 669461 75041
rect 669550 75021 669603 75041
rect 669674 75021 669728 75077
rect 667828 74985 667899 75021
rect 667955 74985 668041 75021
rect 668097 74985 668183 75021
rect 668239 74985 668325 75021
rect 668381 74985 668467 75021
rect 668523 74985 668609 75021
rect 668665 74985 668751 75021
rect 668807 74985 668893 75021
rect 668949 74985 669035 75021
rect 669091 74985 669177 75021
rect 669233 74985 669319 75021
rect 669375 74985 669461 75021
rect 669517 74985 669603 75021
rect 669659 74985 669728 75021
rect 667828 74953 669728 74985
rect 667828 74897 667882 74953
rect 667938 74899 668006 74953
rect 668062 74899 668130 74953
rect 668186 74899 668254 74953
rect 667955 74897 668006 74899
rect 668097 74897 668130 74899
rect 668239 74897 668254 74899
rect 668310 74899 668378 74953
rect 668434 74899 668502 74953
rect 668558 74899 668626 74953
rect 668310 74897 668325 74899
rect 668434 74897 668467 74899
rect 668558 74897 668609 74899
rect 668682 74897 668750 74953
rect 668806 74899 668874 74953
rect 668930 74899 668998 74953
rect 669054 74899 669122 74953
rect 669178 74899 669246 74953
rect 668807 74897 668874 74899
rect 668949 74897 668998 74899
rect 669091 74897 669122 74899
rect 669233 74897 669246 74899
rect 669302 74899 669370 74953
rect 669426 74899 669494 74953
rect 669550 74899 669618 74953
rect 669302 74897 669319 74899
rect 669426 74897 669461 74899
rect 669550 74897 669603 74899
rect 669674 74897 669728 74953
rect 667828 74843 667899 74897
rect 667955 74843 668041 74897
rect 668097 74843 668183 74897
rect 668239 74843 668325 74897
rect 668381 74843 668467 74897
rect 668523 74843 668609 74897
rect 668665 74843 668751 74897
rect 668807 74843 668893 74897
rect 668949 74843 669035 74897
rect 669091 74843 669177 74897
rect 669233 74843 669319 74897
rect 669375 74843 669461 74897
rect 669517 74843 669603 74897
rect 669659 74843 669728 74897
rect 667828 74829 669728 74843
rect 667828 74773 667882 74829
rect 667938 74773 668006 74829
rect 668062 74773 668130 74829
rect 668186 74773 668254 74829
rect 668310 74773 668378 74829
rect 668434 74773 668502 74829
rect 668558 74773 668626 74829
rect 668682 74773 668750 74829
rect 668806 74773 668874 74829
rect 668930 74773 668998 74829
rect 669054 74773 669122 74829
rect 669178 74773 669246 74829
rect 669302 74773 669370 74829
rect 669426 74773 669494 74829
rect 669550 74773 669618 74829
rect 669674 74773 669728 74829
rect 667828 74757 669728 74773
rect 667828 74705 667899 74757
rect 667955 74705 668041 74757
rect 668097 74705 668183 74757
rect 668239 74705 668325 74757
rect 668381 74705 668467 74757
rect 668523 74705 668609 74757
rect 668665 74705 668751 74757
rect 668807 74705 668893 74757
rect 668949 74705 669035 74757
rect 669091 74705 669177 74757
rect 669233 74705 669319 74757
rect 669375 74705 669461 74757
rect 669517 74705 669603 74757
rect 669659 74705 669728 74757
rect 667828 74649 667882 74705
rect 667955 74701 668006 74705
rect 668097 74701 668130 74705
rect 668239 74701 668254 74705
rect 667938 74649 668006 74701
rect 668062 74649 668130 74701
rect 668186 74649 668254 74701
rect 668310 74701 668325 74705
rect 668434 74701 668467 74705
rect 668558 74701 668609 74705
rect 668310 74649 668378 74701
rect 668434 74649 668502 74701
rect 668558 74649 668626 74701
rect 668682 74649 668750 74705
rect 668807 74701 668874 74705
rect 668949 74701 668998 74705
rect 669091 74701 669122 74705
rect 669233 74701 669246 74705
rect 668806 74649 668874 74701
rect 668930 74649 668998 74701
rect 669054 74649 669122 74701
rect 669178 74649 669246 74701
rect 669302 74701 669319 74705
rect 669426 74701 669461 74705
rect 669550 74701 669603 74705
rect 669302 74649 669370 74701
rect 669426 74649 669494 74701
rect 669550 74649 669618 74701
rect 669674 74649 669728 74705
rect 667828 74615 669728 74649
rect 667828 74581 667899 74615
rect 667955 74581 668041 74615
rect 668097 74581 668183 74615
rect 668239 74581 668325 74615
rect 668381 74581 668467 74615
rect 668523 74581 668609 74615
rect 668665 74581 668751 74615
rect 668807 74581 668893 74615
rect 668949 74581 669035 74615
rect 669091 74581 669177 74615
rect 669233 74581 669319 74615
rect 669375 74581 669461 74615
rect 669517 74581 669603 74615
rect 669659 74581 669728 74615
rect 667828 74525 667882 74581
rect 667955 74559 668006 74581
rect 668097 74559 668130 74581
rect 668239 74559 668254 74581
rect 667938 74525 668006 74559
rect 668062 74525 668130 74559
rect 668186 74525 668254 74559
rect 668310 74559 668325 74581
rect 668434 74559 668467 74581
rect 668558 74559 668609 74581
rect 668310 74525 668378 74559
rect 668434 74525 668502 74559
rect 668558 74525 668626 74559
rect 668682 74525 668750 74581
rect 668807 74559 668874 74581
rect 668949 74559 668998 74581
rect 669091 74559 669122 74581
rect 669233 74559 669246 74581
rect 668806 74525 668874 74559
rect 668930 74525 668998 74559
rect 669054 74525 669122 74559
rect 669178 74525 669246 74559
rect 669302 74559 669319 74581
rect 669426 74559 669461 74581
rect 669550 74559 669603 74581
rect 669302 74525 669370 74559
rect 669426 74525 669494 74559
rect 669550 74525 669618 74559
rect 669674 74525 669728 74581
rect 667828 74488 669728 74525
rect 105272 74035 107172 74088
rect 105272 73979 105343 74035
rect 105399 73979 105485 74035
rect 105541 73979 105627 74035
rect 105683 73979 105769 74035
rect 105825 73979 105911 74035
rect 105967 73979 106053 74035
rect 106109 73979 106195 74035
rect 106251 73979 106337 74035
rect 106393 73979 106479 74035
rect 106535 73979 106621 74035
rect 106677 73979 106763 74035
rect 106819 73979 106905 74035
rect 106961 73979 107047 74035
rect 107103 73979 107172 74035
rect 105272 73945 107172 73979
rect 105272 73889 105326 73945
rect 105382 73893 105450 73945
rect 105506 73893 105574 73945
rect 105630 73893 105698 73945
rect 105399 73889 105450 73893
rect 105541 73889 105574 73893
rect 105683 73889 105698 73893
rect 105754 73893 105822 73945
rect 105878 73893 105946 73945
rect 106002 73893 106070 73945
rect 105754 73889 105769 73893
rect 105878 73889 105911 73893
rect 106002 73889 106053 73893
rect 106126 73889 106194 73945
rect 106250 73893 106318 73945
rect 106374 73893 106442 73945
rect 106498 73893 106566 73945
rect 106622 73893 106690 73945
rect 106251 73889 106318 73893
rect 106393 73889 106442 73893
rect 106535 73889 106566 73893
rect 106677 73889 106690 73893
rect 106746 73893 106814 73945
rect 106870 73893 106938 73945
rect 106994 73893 107062 73945
rect 106746 73889 106763 73893
rect 106870 73889 106905 73893
rect 106994 73889 107047 73893
rect 107118 73889 107172 73945
rect 105272 73837 105343 73889
rect 105399 73837 105485 73889
rect 105541 73837 105627 73889
rect 105683 73837 105769 73889
rect 105825 73837 105911 73889
rect 105967 73837 106053 73889
rect 106109 73837 106195 73889
rect 106251 73837 106337 73889
rect 106393 73837 106479 73889
rect 106535 73837 106621 73889
rect 106677 73837 106763 73889
rect 106819 73837 106905 73889
rect 106961 73837 107047 73889
rect 107103 73837 107172 73889
rect 105272 73821 107172 73837
rect 105272 73765 105326 73821
rect 105382 73765 105450 73821
rect 105506 73765 105574 73821
rect 105630 73765 105698 73821
rect 105754 73765 105822 73821
rect 105878 73765 105946 73821
rect 106002 73765 106070 73821
rect 106126 73765 106194 73821
rect 106250 73765 106318 73821
rect 106374 73765 106442 73821
rect 106498 73765 106566 73821
rect 106622 73765 106690 73821
rect 106746 73765 106814 73821
rect 106870 73765 106938 73821
rect 106994 73765 107062 73821
rect 107118 73765 107172 73821
rect 105272 73751 107172 73765
rect 105272 73697 105343 73751
rect 105399 73697 105485 73751
rect 105541 73697 105627 73751
rect 105683 73697 105769 73751
rect 105825 73697 105911 73751
rect 105967 73697 106053 73751
rect 106109 73697 106195 73751
rect 106251 73697 106337 73751
rect 106393 73697 106479 73751
rect 106535 73697 106621 73751
rect 106677 73697 106763 73751
rect 106819 73697 106905 73751
rect 106961 73697 107047 73751
rect 107103 73697 107172 73751
rect 105272 73641 105326 73697
rect 105399 73695 105450 73697
rect 105541 73695 105574 73697
rect 105683 73695 105698 73697
rect 105382 73641 105450 73695
rect 105506 73641 105574 73695
rect 105630 73641 105698 73695
rect 105754 73695 105769 73697
rect 105878 73695 105911 73697
rect 106002 73695 106053 73697
rect 105754 73641 105822 73695
rect 105878 73641 105946 73695
rect 106002 73641 106070 73695
rect 106126 73641 106194 73697
rect 106251 73695 106318 73697
rect 106393 73695 106442 73697
rect 106535 73695 106566 73697
rect 106677 73695 106690 73697
rect 106250 73641 106318 73695
rect 106374 73641 106442 73695
rect 106498 73641 106566 73695
rect 106622 73641 106690 73695
rect 106746 73695 106763 73697
rect 106870 73695 106905 73697
rect 106994 73695 107047 73697
rect 106746 73641 106814 73695
rect 106870 73641 106938 73695
rect 106994 73641 107062 73695
rect 107118 73641 107172 73697
rect 105272 73609 107172 73641
rect 105272 73573 105343 73609
rect 105399 73573 105485 73609
rect 105541 73573 105627 73609
rect 105683 73573 105769 73609
rect 105825 73573 105911 73609
rect 105967 73573 106053 73609
rect 106109 73573 106195 73609
rect 106251 73573 106337 73609
rect 106393 73573 106479 73609
rect 106535 73573 106621 73609
rect 106677 73573 106763 73609
rect 106819 73573 106905 73609
rect 106961 73573 107047 73609
rect 107103 73573 107172 73609
rect 105272 73517 105326 73573
rect 105399 73553 105450 73573
rect 105541 73553 105574 73573
rect 105683 73553 105698 73573
rect 105382 73517 105450 73553
rect 105506 73517 105574 73553
rect 105630 73517 105698 73553
rect 105754 73553 105769 73573
rect 105878 73553 105911 73573
rect 106002 73553 106053 73573
rect 105754 73517 105822 73553
rect 105878 73517 105946 73553
rect 106002 73517 106070 73553
rect 106126 73517 106194 73573
rect 106251 73553 106318 73573
rect 106393 73553 106442 73573
rect 106535 73553 106566 73573
rect 106677 73553 106690 73573
rect 106250 73517 106318 73553
rect 106374 73517 106442 73553
rect 106498 73517 106566 73553
rect 106622 73517 106690 73553
rect 106746 73553 106763 73573
rect 106870 73553 106905 73573
rect 106994 73553 107047 73573
rect 106746 73517 106814 73553
rect 106870 73517 106938 73553
rect 106994 73517 107062 73553
rect 107118 73517 107172 73573
rect 105272 73467 107172 73517
rect 105272 73449 105343 73467
rect 105399 73449 105485 73467
rect 105541 73449 105627 73467
rect 105683 73449 105769 73467
rect 105825 73449 105911 73467
rect 105967 73449 106053 73467
rect 106109 73449 106195 73467
rect 106251 73449 106337 73467
rect 106393 73449 106479 73467
rect 106535 73449 106621 73467
rect 106677 73449 106763 73467
rect 106819 73449 106905 73467
rect 106961 73449 107047 73467
rect 107103 73449 107172 73467
rect 105272 73393 105326 73449
rect 105399 73411 105450 73449
rect 105541 73411 105574 73449
rect 105683 73411 105698 73449
rect 105382 73393 105450 73411
rect 105506 73393 105574 73411
rect 105630 73393 105698 73411
rect 105754 73411 105769 73449
rect 105878 73411 105911 73449
rect 106002 73411 106053 73449
rect 105754 73393 105822 73411
rect 105878 73393 105946 73411
rect 106002 73393 106070 73411
rect 106126 73393 106194 73449
rect 106251 73411 106318 73449
rect 106393 73411 106442 73449
rect 106535 73411 106566 73449
rect 106677 73411 106690 73449
rect 106250 73393 106318 73411
rect 106374 73393 106442 73411
rect 106498 73393 106566 73411
rect 106622 73393 106690 73411
rect 106746 73411 106763 73449
rect 106870 73411 106905 73449
rect 106994 73411 107047 73449
rect 106746 73393 106814 73411
rect 106870 73393 106938 73411
rect 106994 73393 107062 73411
rect 107118 73393 107172 73449
rect 105272 73325 107172 73393
rect 105272 73269 105326 73325
rect 105399 73269 105450 73325
rect 105541 73269 105574 73325
rect 105683 73269 105698 73325
rect 105754 73269 105769 73325
rect 105878 73269 105911 73325
rect 106002 73269 106053 73325
rect 106126 73269 106194 73325
rect 106251 73269 106318 73325
rect 106393 73269 106442 73325
rect 106535 73269 106566 73325
rect 106677 73269 106690 73325
rect 106746 73269 106763 73325
rect 106870 73269 106905 73325
rect 106994 73269 107047 73325
rect 107118 73269 107172 73325
rect 105272 73201 107172 73269
rect 105272 73145 105326 73201
rect 105382 73183 105450 73201
rect 105506 73183 105574 73201
rect 105630 73183 105698 73201
rect 105399 73145 105450 73183
rect 105541 73145 105574 73183
rect 105683 73145 105698 73183
rect 105754 73183 105822 73201
rect 105878 73183 105946 73201
rect 106002 73183 106070 73201
rect 105754 73145 105769 73183
rect 105878 73145 105911 73183
rect 106002 73145 106053 73183
rect 106126 73145 106194 73201
rect 106250 73183 106318 73201
rect 106374 73183 106442 73201
rect 106498 73183 106566 73201
rect 106622 73183 106690 73201
rect 106251 73145 106318 73183
rect 106393 73145 106442 73183
rect 106535 73145 106566 73183
rect 106677 73145 106690 73183
rect 106746 73183 106814 73201
rect 106870 73183 106938 73201
rect 106994 73183 107062 73201
rect 106746 73145 106763 73183
rect 106870 73145 106905 73183
rect 106994 73145 107047 73183
rect 107118 73145 107172 73201
rect 105272 73127 105343 73145
rect 105399 73127 105485 73145
rect 105541 73127 105627 73145
rect 105683 73127 105769 73145
rect 105825 73127 105911 73145
rect 105967 73127 106053 73145
rect 106109 73127 106195 73145
rect 106251 73127 106337 73145
rect 106393 73127 106479 73145
rect 106535 73127 106621 73145
rect 106677 73127 106763 73145
rect 106819 73127 106905 73145
rect 106961 73127 107047 73145
rect 107103 73127 107172 73145
rect 105272 73077 107172 73127
rect 105272 73021 105326 73077
rect 105382 73041 105450 73077
rect 105506 73041 105574 73077
rect 105630 73041 105698 73077
rect 105399 73021 105450 73041
rect 105541 73021 105574 73041
rect 105683 73021 105698 73041
rect 105754 73041 105822 73077
rect 105878 73041 105946 73077
rect 106002 73041 106070 73077
rect 105754 73021 105769 73041
rect 105878 73021 105911 73041
rect 106002 73021 106053 73041
rect 106126 73021 106194 73077
rect 106250 73041 106318 73077
rect 106374 73041 106442 73077
rect 106498 73041 106566 73077
rect 106622 73041 106690 73077
rect 106251 73021 106318 73041
rect 106393 73021 106442 73041
rect 106535 73021 106566 73041
rect 106677 73021 106690 73041
rect 106746 73041 106814 73077
rect 106870 73041 106938 73077
rect 106994 73041 107062 73077
rect 106746 73021 106763 73041
rect 106870 73021 106905 73041
rect 106994 73021 107047 73041
rect 107118 73021 107172 73077
rect 105272 72985 105343 73021
rect 105399 72985 105485 73021
rect 105541 72985 105627 73021
rect 105683 72985 105769 73021
rect 105825 72985 105911 73021
rect 105967 72985 106053 73021
rect 106109 72985 106195 73021
rect 106251 72985 106337 73021
rect 106393 72985 106479 73021
rect 106535 72985 106621 73021
rect 106677 72985 106763 73021
rect 106819 72985 106905 73021
rect 106961 72985 107047 73021
rect 107103 72985 107172 73021
rect 105272 72953 107172 72985
rect 105272 72897 105326 72953
rect 105382 72899 105450 72953
rect 105506 72899 105574 72953
rect 105630 72899 105698 72953
rect 105399 72897 105450 72899
rect 105541 72897 105574 72899
rect 105683 72897 105698 72899
rect 105754 72899 105822 72953
rect 105878 72899 105946 72953
rect 106002 72899 106070 72953
rect 105754 72897 105769 72899
rect 105878 72897 105911 72899
rect 106002 72897 106053 72899
rect 106126 72897 106194 72953
rect 106250 72899 106318 72953
rect 106374 72899 106442 72953
rect 106498 72899 106566 72953
rect 106622 72899 106690 72953
rect 106251 72897 106318 72899
rect 106393 72897 106442 72899
rect 106535 72897 106566 72899
rect 106677 72897 106690 72899
rect 106746 72899 106814 72953
rect 106870 72899 106938 72953
rect 106994 72899 107062 72953
rect 106746 72897 106763 72899
rect 106870 72897 106905 72899
rect 106994 72897 107047 72899
rect 107118 72897 107172 72953
rect 105272 72843 105343 72897
rect 105399 72843 105485 72897
rect 105541 72843 105627 72897
rect 105683 72843 105769 72897
rect 105825 72843 105911 72897
rect 105967 72843 106053 72897
rect 106109 72843 106195 72897
rect 106251 72843 106337 72897
rect 106393 72843 106479 72897
rect 106535 72843 106621 72897
rect 106677 72843 106763 72897
rect 106819 72843 106905 72897
rect 106961 72843 107047 72897
rect 107103 72843 107172 72897
rect 105272 72829 107172 72843
rect 105272 72773 105326 72829
rect 105382 72773 105450 72829
rect 105506 72773 105574 72829
rect 105630 72773 105698 72829
rect 105754 72773 105822 72829
rect 105878 72773 105946 72829
rect 106002 72773 106070 72829
rect 106126 72773 106194 72829
rect 106250 72773 106318 72829
rect 106374 72773 106442 72829
rect 106498 72773 106566 72829
rect 106622 72773 106690 72829
rect 106746 72773 106814 72829
rect 106870 72773 106938 72829
rect 106994 72773 107062 72829
rect 107118 72773 107172 72829
rect 105272 72757 107172 72773
rect 105272 72705 105343 72757
rect 105399 72705 105485 72757
rect 105541 72705 105627 72757
rect 105683 72705 105769 72757
rect 105825 72705 105911 72757
rect 105967 72705 106053 72757
rect 106109 72705 106195 72757
rect 106251 72705 106337 72757
rect 106393 72705 106479 72757
rect 106535 72705 106621 72757
rect 106677 72705 106763 72757
rect 106819 72705 106905 72757
rect 106961 72705 107047 72757
rect 107103 72705 107172 72757
rect 105272 72649 105326 72705
rect 105399 72701 105450 72705
rect 105541 72701 105574 72705
rect 105683 72701 105698 72705
rect 105382 72649 105450 72701
rect 105506 72649 105574 72701
rect 105630 72649 105698 72701
rect 105754 72701 105769 72705
rect 105878 72701 105911 72705
rect 106002 72701 106053 72705
rect 105754 72649 105822 72701
rect 105878 72649 105946 72701
rect 106002 72649 106070 72701
rect 106126 72649 106194 72705
rect 106251 72701 106318 72705
rect 106393 72701 106442 72705
rect 106535 72701 106566 72705
rect 106677 72701 106690 72705
rect 106250 72649 106318 72701
rect 106374 72649 106442 72701
rect 106498 72649 106566 72701
rect 106622 72649 106690 72701
rect 106746 72701 106763 72705
rect 106870 72701 106905 72705
rect 106994 72701 107047 72705
rect 106746 72649 106814 72701
rect 106870 72649 106938 72701
rect 106994 72649 107062 72701
rect 107118 72649 107172 72705
rect 105272 72615 107172 72649
rect 105272 72581 105343 72615
rect 105399 72581 105485 72615
rect 105541 72581 105627 72615
rect 105683 72581 105769 72615
rect 105825 72581 105911 72615
rect 105967 72581 106053 72615
rect 106109 72581 106195 72615
rect 106251 72581 106337 72615
rect 106393 72581 106479 72615
rect 106535 72581 106621 72615
rect 106677 72581 106763 72615
rect 106819 72581 106905 72615
rect 106961 72581 107047 72615
rect 107103 72581 107172 72615
rect 105272 72525 105326 72581
rect 105399 72559 105450 72581
rect 105541 72559 105574 72581
rect 105683 72559 105698 72581
rect 105382 72525 105450 72559
rect 105506 72525 105574 72559
rect 105630 72525 105698 72559
rect 105754 72559 105769 72581
rect 105878 72559 105911 72581
rect 106002 72559 106053 72581
rect 105754 72525 105822 72559
rect 105878 72525 105946 72559
rect 106002 72525 106070 72559
rect 106126 72525 106194 72581
rect 106251 72559 106318 72581
rect 106393 72559 106442 72581
rect 106535 72559 106566 72581
rect 106677 72559 106690 72581
rect 106250 72525 106318 72559
rect 106374 72525 106442 72559
rect 106498 72525 106566 72559
rect 106622 72525 106690 72559
rect 106746 72559 106763 72581
rect 106870 72559 106905 72581
rect 106994 72559 107047 72581
rect 106746 72525 106814 72559
rect 106870 72525 106938 72559
rect 106994 72525 107062 72559
rect 107118 72525 107172 72581
rect 105272 72473 107172 72525
rect 105272 72457 105343 72473
rect 105399 72457 105485 72473
rect 105541 72457 105627 72473
rect 105683 72457 105769 72473
rect 105825 72457 105911 72473
rect 105967 72457 106053 72473
rect 106109 72457 106195 72473
rect 106251 72457 106337 72473
rect 106393 72457 106479 72473
rect 106535 72457 106621 72473
rect 106677 72457 106763 72473
rect 106819 72457 106905 72473
rect 106961 72457 107047 72473
rect 107103 72457 107172 72473
rect 105272 72401 105326 72457
rect 105399 72417 105450 72457
rect 105541 72417 105574 72457
rect 105683 72417 105698 72457
rect 105382 72401 105450 72417
rect 105506 72401 105574 72417
rect 105630 72401 105698 72417
rect 105754 72417 105769 72457
rect 105878 72417 105911 72457
rect 106002 72417 106053 72457
rect 105754 72401 105822 72417
rect 105878 72401 105946 72417
rect 106002 72401 106070 72417
rect 106126 72401 106194 72457
rect 106251 72417 106318 72457
rect 106393 72417 106442 72457
rect 106535 72417 106566 72457
rect 106677 72417 106690 72457
rect 106250 72401 106318 72417
rect 106374 72401 106442 72417
rect 106498 72401 106566 72417
rect 106622 72401 106690 72417
rect 106746 72417 106763 72457
rect 106870 72417 106905 72457
rect 106994 72417 107047 72457
rect 106746 72401 106814 72417
rect 106870 72401 106938 72417
rect 106994 72401 107062 72417
rect 107118 72401 107172 72457
rect 105272 72333 107172 72401
rect 105272 72277 105326 72333
rect 105382 72331 105450 72333
rect 105506 72331 105574 72333
rect 105630 72331 105698 72333
rect 105399 72277 105450 72331
rect 105541 72277 105574 72331
rect 105683 72277 105698 72331
rect 105754 72331 105822 72333
rect 105878 72331 105946 72333
rect 106002 72331 106070 72333
rect 105754 72277 105769 72331
rect 105878 72277 105911 72331
rect 106002 72277 106053 72331
rect 106126 72277 106194 72333
rect 106250 72331 106318 72333
rect 106374 72331 106442 72333
rect 106498 72331 106566 72333
rect 106622 72331 106690 72333
rect 106251 72277 106318 72331
rect 106393 72277 106442 72331
rect 106535 72277 106566 72331
rect 106677 72277 106690 72331
rect 106746 72331 106814 72333
rect 106870 72331 106938 72333
rect 106994 72331 107062 72333
rect 106746 72277 106763 72331
rect 106870 72277 106905 72331
rect 106994 72277 107047 72331
rect 107118 72277 107172 72333
rect 105272 72275 105343 72277
rect 105399 72275 105485 72277
rect 105541 72275 105627 72277
rect 105683 72275 105769 72277
rect 105825 72275 105911 72277
rect 105967 72275 106053 72277
rect 106109 72275 106195 72277
rect 106251 72275 106337 72277
rect 106393 72275 106479 72277
rect 106535 72275 106621 72277
rect 106677 72275 106763 72277
rect 106819 72275 106905 72277
rect 106961 72275 107047 72277
rect 107103 72275 107172 72277
rect 105272 72209 107172 72275
rect 105272 72153 105326 72209
rect 105382 72189 105450 72209
rect 105506 72189 105574 72209
rect 105630 72189 105698 72209
rect 105399 72153 105450 72189
rect 105541 72153 105574 72189
rect 105683 72153 105698 72189
rect 105754 72189 105822 72209
rect 105878 72189 105946 72209
rect 106002 72189 106070 72209
rect 105754 72153 105769 72189
rect 105878 72153 105911 72189
rect 106002 72153 106053 72189
rect 106126 72153 106194 72209
rect 106250 72189 106318 72209
rect 106374 72189 106442 72209
rect 106498 72189 106566 72209
rect 106622 72189 106690 72209
rect 106251 72153 106318 72189
rect 106393 72153 106442 72189
rect 106535 72153 106566 72189
rect 106677 72153 106690 72189
rect 106746 72189 106814 72209
rect 106870 72189 106938 72209
rect 106994 72189 107062 72209
rect 106746 72153 106763 72189
rect 106870 72153 106905 72189
rect 106994 72153 107047 72189
rect 107118 72153 107172 72209
rect 105272 72133 105343 72153
rect 105399 72133 105485 72153
rect 105541 72133 105627 72153
rect 105683 72133 105769 72153
rect 105825 72133 105911 72153
rect 105967 72133 106053 72153
rect 106109 72133 106195 72153
rect 106251 72133 106337 72153
rect 106393 72133 106479 72153
rect 106535 72133 106621 72153
rect 106677 72133 106763 72153
rect 106819 72133 106905 72153
rect 106961 72133 107047 72153
rect 107103 72133 107172 72153
rect 105272 72088 107172 72133
rect 107752 74035 109802 74088
rect 107752 73979 108995 74035
rect 109051 73979 109137 74035
rect 109193 73979 109279 74035
rect 109335 73979 109421 74035
rect 109477 73979 109563 74035
rect 109619 73979 109705 74035
rect 109761 73979 109802 74035
rect 107752 73945 109802 73979
rect 107752 73893 109046 73945
rect 109102 73893 109170 73945
rect 109226 73893 109294 73945
rect 107752 73837 108995 73893
rect 109102 73889 109137 73893
rect 109226 73889 109279 73893
rect 109350 73889 109418 73945
rect 109474 73893 109542 73945
rect 109598 73893 109666 73945
rect 109722 73893 109802 73945
rect 109477 73889 109542 73893
rect 109619 73889 109666 73893
rect 109051 73837 109137 73889
rect 109193 73837 109279 73889
rect 109335 73837 109421 73889
rect 109477 73837 109563 73889
rect 109619 73837 109705 73889
rect 109761 73837 109802 73893
rect 107752 73821 109802 73837
rect 107752 73765 109046 73821
rect 109102 73765 109170 73821
rect 109226 73765 109294 73821
rect 109350 73765 109418 73821
rect 109474 73765 109542 73821
rect 109598 73765 109666 73821
rect 109722 73765 109802 73821
rect 107752 73751 109802 73765
rect 107752 73695 108995 73751
rect 109051 73697 109137 73751
rect 109193 73697 109279 73751
rect 109335 73697 109421 73751
rect 109477 73697 109563 73751
rect 109619 73697 109705 73751
rect 109102 73695 109137 73697
rect 109226 73695 109279 73697
rect 107752 73641 109046 73695
rect 109102 73641 109170 73695
rect 109226 73641 109294 73695
rect 109350 73641 109418 73697
rect 109477 73695 109542 73697
rect 109619 73695 109666 73697
rect 109761 73695 109802 73751
rect 109474 73641 109542 73695
rect 109598 73641 109666 73695
rect 109722 73641 109802 73695
rect 107752 73609 109802 73641
rect 107752 73553 108995 73609
rect 109051 73573 109137 73609
rect 109193 73573 109279 73609
rect 109335 73573 109421 73609
rect 109477 73573 109563 73609
rect 109619 73573 109705 73609
rect 109102 73553 109137 73573
rect 109226 73553 109279 73573
rect 107752 73517 109046 73553
rect 109102 73517 109170 73553
rect 109226 73517 109294 73553
rect 109350 73517 109418 73573
rect 109477 73553 109542 73573
rect 109619 73553 109666 73573
rect 109761 73553 109802 73609
rect 109474 73517 109542 73553
rect 109598 73517 109666 73553
rect 109722 73517 109802 73553
rect 107752 73467 109802 73517
rect 107752 73411 108995 73467
rect 109051 73449 109137 73467
rect 109193 73449 109279 73467
rect 109335 73449 109421 73467
rect 109477 73449 109563 73467
rect 109619 73449 109705 73467
rect 109102 73411 109137 73449
rect 109226 73411 109279 73449
rect 107752 73393 109046 73411
rect 109102 73393 109170 73411
rect 109226 73393 109294 73411
rect 109350 73393 109418 73449
rect 109477 73411 109542 73449
rect 109619 73411 109666 73449
rect 109761 73411 109802 73467
rect 109474 73393 109542 73411
rect 109598 73393 109666 73411
rect 109722 73393 109802 73411
rect 107752 73325 109802 73393
rect 107752 73269 108995 73325
rect 109102 73269 109137 73325
rect 109226 73269 109279 73325
rect 109350 73269 109418 73325
rect 109477 73269 109542 73325
rect 109619 73269 109666 73325
rect 109761 73269 109802 73325
rect 107752 73201 109802 73269
rect 107752 73183 109046 73201
rect 109102 73183 109170 73201
rect 109226 73183 109294 73201
rect 107752 73127 108995 73183
rect 109102 73145 109137 73183
rect 109226 73145 109279 73183
rect 109350 73145 109418 73201
rect 109474 73183 109542 73201
rect 109598 73183 109666 73201
rect 109722 73183 109802 73201
rect 109477 73145 109542 73183
rect 109619 73145 109666 73183
rect 109051 73127 109137 73145
rect 109193 73127 109279 73145
rect 109335 73127 109421 73145
rect 109477 73127 109563 73145
rect 109619 73127 109705 73145
rect 109761 73127 109802 73183
rect 107752 73077 109802 73127
rect 107752 73041 109046 73077
rect 109102 73041 109170 73077
rect 109226 73041 109294 73077
rect 107752 72985 108995 73041
rect 109102 73021 109137 73041
rect 109226 73021 109279 73041
rect 109350 73021 109418 73077
rect 109474 73041 109542 73077
rect 109598 73041 109666 73077
rect 109722 73041 109802 73077
rect 109477 73021 109542 73041
rect 109619 73021 109666 73041
rect 109051 72985 109137 73021
rect 109193 72985 109279 73021
rect 109335 72985 109421 73021
rect 109477 72985 109563 73021
rect 109619 72985 109705 73021
rect 109761 72985 109802 73041
rect 107752 72953 109802 72985
rect 107752 72899 109046 72953
rect 109102 72899 109170 72953
rect 109226 72899 109294 72953
rect 107752 72843 108995 72899
rect 109102 72897 109137 72899
rect 109226 72897 109279 72899
rect 109350 72897 109418 72953
rect 109474 72899 109542 72953
rect 109598 72899 109666 72953
rect 109722 72899 109802 72953
rect 109477 72897 109542 72899
rect 109619 72897 109666 72899
rect 109051 72843 109137 72897
rect 109193 72843 109279 72897
rect 109335 72843 109421 72897
rect 109477 72843 109563 72897
rect 109619 72843 109705 72897
rect 109761 72843 109802 72899
rect 107752 72829 109802 72843
rect 107752 72773 109046 72829
rect 109102 72773 109170 72829
rect 109226 72773 109294 72829
rect 109350 72773 109418 72829
rect 109474 72773 109542 72829
rect 109598 72773 109666 72829
rect 109722 72773 109802 72829
rect 107752 72757 109802 72773
rect 107752 72701 108995 72757
rect 109051 72705 109137 72757
rect 109193 72705 109279 72757
rect 109335 72705 109421 72757
rect 109477 72705 109563 72757
rect 109619 72705 109705 72757
rect 109102 72701 109137 72705
rect 109226 72701 109279 72705
rect 107752 72649 109046 72701
rect 109102 72649 109170 72701
rect 109226 72649 109294 72701
rect 109350 72649 109418 72705
rect 109477 72701 109542 72705
rect 109619 72701 109666 72705
rect 109761 72701 109802 72757
rect 109474 72649 109542 72701
rect 109598 72649 109666 72701
rect 109722 72649 109802 72701
rect 107752 72615 109802 72649
rect 107752 72559 108995 72615
rect 109051 72581 109137 72615
rect 109193 72581 109279 72615
rect 109335 72581 109421 72615
rect 109477 72581 109563 72615
rect 109619 72581 109705 72615
rect 109102 72559 109137 72581
rect 109226 72559 109279 72581
rect 107752 72525 109046 72559
rect 109102 72525 109170 72559
rect 109226 72525 109294 72559
rect 109350 72525 109418 72581
rect 109477 72559 109542 72581
rect 109619 72559 109666 72581
rect 109761 72559 109802 72615
rect 109474 72525 109542 72559
rect 109598 72525 109666 72559
rect 109722 72525 109802 72559
rect 107752 72473 109802 72525
rect 107752 72417 108995 72473
rect 109051 72457 109137 72473
rect 109193 72457 109279 72473
rect 109335 72457 109421 72473
rect 109477 72457 109563 72473
rect 109619 72457 109705 72473
rect 109102 72417 109137 72457
rect 109226 72417 109279 72457
rect 107752 72401 109046 72417
rect 109102 72401 109170 72417
rect 109226 72401 109294 72417
rect 109350 72401 109418 72457
rect 109477 72417 109542 72457
rect 109619 72417 109666 72457
rect 109761 72417 109802 72473
rect 109474 72401 109542 72417
rect 109598 72401 109666 72417
rect 109722 72401 109802 72417
rect 107752 72333 109802 72401
rect 107752 72331 109046 72333
rect 109102 72331 109170 72333
rect 109226 72331 109294 72333
rect 107752 72275 108995 72331
rect 109102 72277 109137 72331
rect 109226 72277 109279 72331
rect 109350 72277 109418 72333
rect 109474 72331 109542 72333
rect 109598 72331 109666 72333
rect 109722 72331 109802 72333
rect 109477 72277 109542 72331
rect 109619 72277 109666 72331
rect 109051 72275 109137 72277
rect 109193 72275 109279 72277
rect 109335 72275 109421 72277
rect 109477 72275 109563 72277
rect 109619 72275 109705 72277
rect 109761 72275 109802 72331
rect 107752 72209 109802 72275
rect 107752 72189 109046 72209
rect 109102 72189 109170 72209
rect 109226 72189 109294 72209
rect 107752 72133 108995 72189
rect 109102 72153 109137 72189
rect 109226 72153 109279 72189
rect 109350 72153 109418 72209
rect 109474 72189 109542 72209
rect 109598 72189 109666 72209
rect 109722 72189 109802 72209
rect 109477 72153 109542 72189
rect 109619 72153 109666 72189
rect 109051 72133 109137 72153
rect 109193 72133 109279 72153
rect 109335 72133 109421 72153
rect 109477 72133 109563 72153
rect 109619 72133 109705 72153
rect 109761 72133 109802 72189
rect 107752 72088 109802 72133
rect 110122 74035 112172 74088
rect 110122 73979 110193 74035
rect 110249 73979 110335 74035
rect 110391 73979 110477 74035
rect 110533 73979 110619 74035
rect 110675 73979 110761 74035
rect 110817 73979 110903 74035
rect 110959 73979 111045 74035
rect 111101 73979 111187 74035
rect 111243 73979 111329 74035
rect 111385 73979 111471 74035
rect 111527 73979 111613 74035
rect 111669 73979 111755 74035
rect 111811 73979 111897 74035
rect 111953 73979 112039 74035
rect 112095 73979 112172 74035
rect 110122 73945 112172 73979
rect 110122 73889 110176 73945
rect 110232 73893 110300 73945
rect 110356 73893 110424 73945
rect 110480 73893 110548 73945
rect 110249 73889 110300 73893
rect 110391 73889 110424 73893
rect 110533 73889 110548 73893
rect 110604 73893 110672 73945
rect 110728 73893 110796 73945
rect 110852 73893 110920 73945
rect 110604 73889 110619 73893
rect 110728 73889 110761 73893
rect 110852 73889 110903 73893
rect 110976 73889 111044 73945
rect 111100 73893 111168 73945
rect 111224 73893 111292 73945
rect 111348 73893 111416 73945
rect 111472 73893 111540 73945
rect 111101 73889 111168 73893
rect 111243 73889 111292 73893
rect 111385 73889 111416 73893
rect 111527 73889 111540 73893
rect 111596 73893 111664 73945
rect 111720 73893 111788 73945
rect 111844 73893 111912 73945
rect 111596 73889 111613 73893
rect 111720 73889 111755 73893
rect 111844 73889 111897 73893
rect 111968 73889 112036 73945
rect 112092 73893 112172 73945
rect 110122 73837 110193 73889
rect 110249 73837 110335 73889
rect 110391 73837 110477 73889
rect 110533 73837 110619 73889
rect 110675 73837 110761 73889
rect 110817 73837 110903 73889
rect 110959 73837 111045 73889
rect 111101 73837 111187 73889
rect 111243 73837 111329 73889
rect 111385 73837 111471 73889
rect 111527 73837 111613 73889
rect 111669 73837 111755 73889
rect 111811 73837 111897 73889
rect 111953 73837 112039 73889
rect 112095 73837 112172 73893
rect 110122 73821 112172 73837
rect 110122 73765 110176 73821
rect 110232 73765 110300 73821
rect 110356 73765 110424 73821
rect 110480 73765 110548 73821
rect 110604 73765 110672 73821
rect 110728 73765 110796 73821
rect 110852 73765 110920 73821
rect 110976 73765 111044 73821
rect 111100 73765 111168 73821
rect 111224 73765 111292 73821
rect 111348 73765 111416 73821
rect 111472 73765 111540 73821
rect 111596 73765 111664 73821
rect 111720 73765 111788 73821
rect 111844 73765 111912 73821
rect 111968 73765 112036 73821
rect 112092 73765 112172 73821
rect 110122 73751 112172 73765
rect 110122 73697 110193 73751
rect 110249 73697 110335 73751
rect 110391 73697 110477 73751
rect 110533 73697 110619 73751
rect 110675 73697 110761 73751
rect 110817 73697 110903 73751
rect 110959 73697 111045 73751
rect 111101 73697 111187 73751
rect 111243 73697 111329 73751
rect 111385 73697 111471 73751
rect 111527 73697 111613 73751
rect 111669 73697 111755 73751
rect 111811 73697 111897 73751
rect 111953 73697 112039 73751
rect 110122 73641 110176 73697
rect 110249 73695 110300 73697
rect 110391 73695 110424 73697
rect 110533 73695 110548 73697
rect 110232 73641 110300 73695
rect 110356 73641 110424 73695
rect 110480 73641 110548 73695
rect 110604 73695 110619 73697
rect 110728 73695 110761 73697
rect 110852 73695 110903 73697
rect 110604 73641 110672 73695
rect 110728 73641 110796 73695
rect 110852 73641 110920 73695
rect 110976 73641 111044 73697
rect 111101 73695 111168 73697
rect 111243 73695 111292 73697
rect 111385 73695 111416 73697
rect 111527 73695 111540 73697
rect 111100 73641 111168 73695
rect 111224 73641 111292 73695
rect 111348 73641 111416 73695
rect 111472 73641 111540 73695
rect 111596 73695 111613 73697
rect 111720 73695 111755 73697
rect 111844 73695 111897 73697
rect 111596 73641 111664 73695
rect 111720 73641 111788 73695
rect 111844 73641 111912 73695
rect 111968 73641 112036 73697
rect 112095 73695 112172 73751
rect 112092 73641 112172 73695
rect 110122 73609 112172 73641
rect 110122 73573 110193 73609
rect 110249 73573 110335 73609
rect 110391 73573 110477 73609
rect 110533 73573 110619 73609
rect 110675 73573 110761 73609
rect 110817 73573 110903 73609
rect 110959 73573 111045 73609
rect 111101 73573 111187 73609
rect 111243 73573 111329 73609
rect 111385 73573 111471 73609
rect 111527 73573 111613 73609
rect 111669 73573 111755 73609
rect 111811 73573 111897 73609
rect 111953 73573 112039 73609
rect 110122 73517 110176 73573
rect 110249 73553 110300 73573
rect 110391 73553 110424 73573
rect 110533 73553 110548 73573
rect 110232 73517 110300 73553
rect 110356 73517 110424 73553
rect 110480 73517 110548 73553
rect 110604 73553 110619 73573
rect 110728 73553 110761 73573
rect 110852 73553 110903 73573
rect 110604 73517 110672 73553
rect 110728 73517 110796 73553
rect 110852 73517 110920 73553
rect 110976 73517 111044 73573
rect 111101 73553 111168 73573
rect 111243 73553 111292 73573
rect 111385 73553 111416 73573
rect 111527 73553 111540 73573
rect 111100 73517 111168 73553
rect 111224 73517 111292 73553
rect 111348 73517 111416 73553
rect 111472 73517 111540 73553
rect 111596 73553 111613 73573
rect 111720 73553 111755 73573
rect 111844 73553 111897 73573
rect 111596 73517 111664 73553
rect 111720 73517 111788 73553
rect 111844 73517 111912 73553
rect 111968 73517 112036 73573
rect 112095 73553 112172 73609
rect 112092 73517 112172 73553
rect 110122 73467 112172 73517
rect 110122 73449 110193 73467
rect 110249 73449 110335 73467
rect 110391 73449 110477 73467
rect 110533 73449 110619 73467
rect 110675 73449 110761 73467
rect 110817 73449 110903 73467
rect 110959 73449 111045 73467
rect 111101 73449 111187 73467
rect 111243 73449 111329 73467
rect 111385 73449 111471 73467
rect 111527 73449 111613 73467
rect 111669 73449 111755 73467
rect 111811 73449 111897 73467
rect 111953 73449 112039 73467
rect 110122 73393 110176 73449
rect 110249 73411 110300 73449
rect 110391 73411 110424 73449
rect 110533 73411 110548 73449
rect 110232 73393 110300 73411
rect 110356 73393 110424 73411
rect 110480 73393 110548 73411
rect 110604 73411 110619 73449
rect 110728 73411 110761 73449
rect 110852 73411 110903 73449
rect 110604 73393 110672 73411
rect 110728 73393 110796 73411
rect 110852 73393 110920 73411
rect 110976 73393 111044 73449
rect 111101 73411 111168 73449
rect 111243 73411 111292 73449
rect 111385 73411 111416 73449
rect 111527 73411 111540 73449
rect 111100 73393 111168 73411
rect 111224 73393 111292 73411
rect 111348 73393 111416 73411
rect 111472 73393 111540 73411
rect 111596 73411 111613 73449
rect 111720 73411 111755 73449
rect 111844 73411 111897 73449
rect 111596 73393 111664 73411
rect 111720 73393 111788 73411
rect 111844 73393 111912 73411
rect 111968 73393 112036 73449
rect 112095 73411 112172 73467
rect 112092 73393 112172 73411
rect 110122 73325 112172 73393
rect 110122 73269 110176 73325
rect 110249 73269 110300 73325
rect 110391 73269 110424 73325
rect 110533 73269 110548 73325
rect 110604 73269 110619 73325
rect 110728 73269 110761 73325
rect 110852 73269 110903 73325
rect 110976 73269 111044 73325
rect 111101 73269 111168 73325
rect 111243 73269 111292 73325
rect 111385 73269 111416 73325
rect 111527 73269 111540 73325
rect 111596 73269 111613 73325
rect 111720 73269 111755 73325
rect 111844 73269 111897 73325
rect 111968 73269 112036 73325
rect 112095 73269 112172 73325
rect 110122 73201 112172 73269
rect 110122 73145 110176 73201
rect 110232 73183 110300 73201
rect 110356 73183 110424 73201
rect 110480 73183 110548 73201
rect 110249 73145 110300 73183
rect 110391 73145 110424 73183
rect 110533 73145 110548 73183
rect 110604 73183 110672 73201
rect 110728 73183 110796 73201
rect 110852 73183 110920 73201
rect 110604 73145 110619 73183
rect 110728 73145 110761 73183
rect 110852 73145 110903 73183
rect 110976 73145 111044 73201
rect 111100 73183 111168 73201
rect 111224 73183 111292 73201
rect 111348 73183 111416 73201
rect 111472 73183 111540 73201
rect 111101 73145 111168 73183
rect 111243 73145 111292 73183
rect 111385 73145 111416 73183
rect 111527 73145 111540 73183
rect 111596 73183 111664 73201
rect 111720 73183 111788 73201
rect 111844 73183 111912 73201
rect 111596 73145 111613 73183
rect 111720 73145 111755 73183
rect 111844 73145 111897 73183
rect 111968 73145 112036 73201
rect 112092 73183 112172 73201
rect 110122 73127 110193 73145
rect 110249 73127 110335 73145
rect 110391 73127 110477 73145
rect 110533 73127 110619 73145
rect 110675 73127 110761 73145
rect 110817 73127 110903 73145
rect 110959 73127 111045 73145
rect 111101 73127 111187 73145
rect 111243 73127 111329 73145
rect 111385 73127 111471 73145
rect 111527 73127 111613 73145
rect 111669 73127 111755 73145
rect 111811 73127 111897 73145
rect 111953 73127 112039 73145
rect 112095 73127 112172 73183
rect 110122 73077 112172 73127
rect 110122 73021 110176 73077
rect 110232 73041 110300 73077
rect 110356 73041 110424 73077
rect 110480 73041 110548 73077
rect 110249 73021 110300 73041
rect 110391 73021 110424 73041
rect 110533 73021 110548 73041
rect 110604 73041 110672 73077
rect 110728 73041 110796 73077
rect 110852 73041 110920 73077
rect 110604 73021 110619 73041
rect 110728 73021 110761 73041
rect 110852 73021 110903 73041
rect 110976 73021 111044 73077
rect 111100 73041 111168 73077
rect 111224 73041 111292 73077
rect 111348 73041 111416 73077
rect 111472 73041 111540 73077
rect 111101 73021 111168 73041
rect 111243 73021 111292 73041
rect 111385 73021 111416 73041
rect 111527 73021 111540 73041
rect 111596 73041 111664 73077
rect 111720 73041 111788 73077
rect 111844 73041 111912 73077
rect 111596 73021 111613 73041
rect 111720 73021 111755 73041
rect 111844 73021 111897 73041
rect 111968 73021 112036 73077
rect 112092 73041 112172 73077
rect 110122 72985 110193 73021
rect 110249 72985 110335 73021
rect 110391 72985 110477 73021
rect 110533 72985 110619 73021
rect 110675 72985 110761 73021
rect 110817 72985 110903 73021
rect 110959 72985 111045 73021
rect 111101 72985 111187 73021
rect 111243 72985 111329 73021
rect 111385 72985 111471 73021
rect 111527 72985 111613 73021
rect 111669 72985 111755 73021
rect 111811 72985 111897 73021
rect 111953 72985 112039 73021
rect 112095 72985 112172 73041
rect 110122 72953 112172 72985
rect 110122 72897 110176 72953
rect 110232 72899 110300 72953
rect 110356 72899 110424 72953
rect 110480 72899 110548 72953
rect 110249 72897 110300 72899
rect 110391 72897 110424 72899
rect 110533 72897 110548 72899
rect 110604 72899 110672 72953
rect 110728 72899 110796 72953
rect 110852 72899 110920 72953
rect 110604 72897 110619 72899
rect 110728 72897 110761 72899
rect 110852 72897 110903 72899
rect 110976 72897 111044 72953
rect 111100 72899 111168 72953
rect 111224 72899 111292 72953
rect 111348 72899 111416 72953
rect 111472 72899 111540 72953
rect 111101 72897 111168 72899
rect 111243 72897 111292 72899
rect 111385 72897 111416 72899
rect 111527 72897 111540 72899
rect 111596 72899 111664 72953
rect 111720 72899 111788 72953
rect 111844 72899 111912 72953
rect 111596 72897 111613 72899
rect 111720 72897 111755 72899
rect 111844 72897 111897 72899
rect 111968 72897 112036 72953
rect 112092 72899 112172 72953
rect 110122 72843 110193 72897
rect 110249 72843 110335 72897
rect 110391 72843 110477 72897
rect 110533 72843 110619 72897
rect 110675 72843 110761 72897
rect 110817 72843 110903 72897
rect 110959 72843 111045 72897
rect 111101 72843 111187 72897
rect 111243 72843 111329 72897
rect 111385 72843 111471 72897
rect 111527 72843 111613 72897
rect 111669 72843 111755 72897
rect 111811 72843 111897 72897
rect 111953 72843 112039 72897
rect 112095 72843 112172 72899
rect 110122 72829 112172 72843
rect 110122 72773 110176 72829
rect 110232 72773 110300 72829
rect 110356 72773 110424 72829
rect 110480 72773 110548 72829
rect 110604 72773 110672 72829
rect 110728 72773 110796 72829
rect 110852 72773 110920 72829
rect 110976 72773 111044 72829
rect 111100 72773 111168 72829
rect 111224 72773 111292 72829
rect 111348 72773 111416 72829
rect 111472 72773 111540 72829
rect 111596 72773 111664 72829
rect 111720 72773 111788 72829
rect 111844 72773 111912 72829
rect 111968 72773 112036 72829
rect 112092 72773 112172 72829
rect 110122 72757 112172 72773
rect 110122 72705 110193 72757
rect 110249 72705 110335 72757
rect 110391 72705 110477 72757
rect 110533 72705 110619 72757
rect 110675 72705 110761 72757
rect 110817 72705 110903 72757
rect 110959 72705 111045 72757
rect 111101 72705 111187 72757
rect 111243 72705 111329 72757
rect 111385 72705 111471 72757
rect 111527 72705 111613 72757
rect 111669 72705 111755 72757
rect 111811 72705 111897 72757
rect 111953 72705 112039 72757
rect 110122 72649 110176 72705
rect 110249 72701 110300 72705
rect 110391 72701 110424 72705
rect 110533 72701 110548 72705
rect 110232 72649 110300 72701
rect 110356 72649 110424 72701
rect 110480 72649 110548 72701
rect 110604 72701 110619 72705
rect 110728 72701 110761 72705
rect 110852 72701 110903 72705
rect 110604 72649 110672 72701
rect 110728 72649 110796 72701
rect 110852 72649 110920 72701
rect 110976 72649 111044 72705
rect 111101 72701 111168 72705
rect 111243 72701 111292 72705
rect 111385 72701 111416 72705
rect 111527 72701 111540 72705
rect 111100 72649 111168 72701
rect 111224 72649 111292 72701
rect 111348 72649 111416 72701
rect 111472 72649 111540 72701
rect 111596 72701 111613 72705
rect 111720 72701 111755 72705
rect 111844 72701 111897 72705
rect 111596 72649 111664 72701
rect 111720 72649 111788 72701
rect 111844 72649 111912 72701
rect 111968 72649 112036 72705
rect 112095 72701 112172 72757
rect 112092 72649 112172 72701
rect 110122 72615 112172 72649
rect 110122 72581 110193 72615
rect 110249 72581 110335 72615
rect 110391 72581 110477 72615
rect 110533 72581 110619 72615
rect 110675 72581 110761 72615
rect 110817 72581 110903 72615
rect 110959 72581 111045 72615
rect 111101 72581 111187 72615
rect 111243 72581 111329 72615
rect 111385 72581 111471 72615
rect 111527 72581 111613 72615
rect 111669 72581 111755 72615
rect 111811 72581 111897 72615
rect 111953 72581 112039 72615
rect 110122 72525 110176 72581
rect 110249 72559 110300 72581
rect 110391 72559 110424 72581
rect 110533 72559 110548 72581
rect 110232 72525 110300 72559
rect 110356 72525 110424 72559
rect 110480 72525 110548 72559
rect 110604 72559 110619 72581
rect 110728 72559 110761 72581
rect 110852 72559 110903 72581
rect 110604 72525 110672 72559
rect 110728 72525 110796 72559
rect 110852 72525 110920 72559
rect 110976 72525 111044 72581
rect 111101 72559 111168 72581
rect 111243 72559 111292 72581
rect 111385 72559 111416 72581
rect 111527 72559 111540 72581
rect 111100 72525 111168 72559
rect 111224 72525 111292 72559
rect 111348 72525 111416 72559
rect 111472 72525 111540 72559
rect 111596 72559 111613 72581
rect 111720 72559 111755 72581
rect 111844 72559 111897 72581
rect 111596 72525 111664 72559
rect 111720 72525 111788 72559
rect 111844 72525 111912 72559
rect 111968 72525 112036 72581
rect 112095 72559 112172 72615
rect 112092 72525 112172 72559
rect 110122 72473 112172 72525
rect 110122 72457 110193 72473
rect 110249 72457 110335 72473
rect 110391 72457 110477 72473
rect 110533 72457 110619 72473
rect 110675 72457 110761 72473
rect 110817 72457 110903 72473
rect 110959 72457 111045 72473
rect 111101 72457 111187 72473
rect 111243 72457 111329 72473
rect 111385 72457 111471 72473
rect 111527 72457 111613 72473
rect 111669 72457 111755 72473
rect 111811 72457 111897 72473
rect 111953 72457 112039 72473
rect 110122 72401 110176 72457
rect 110249 72417 110300 72457
rect 110391 72417 110424 72457
rect 110533 72417 110548 72457
rect 110232 72401 110300 72417
rect 110356 72401 110424 72417
rect 110480 72401 110548 72417
rect 110604 72417 110619 72457
rect 110728 72417 110761 72457
rect 110852 72417 110903 72457
rect 110604 72401 110672 72417
rect 110728 72401 110796 72417
rect 110852 72401 110920 72417
rect 110976 72401 111044 72457
rect 111101 72417 111168 72457
rect 111243 72417 111292 72457
rect 111385 72417 111416 72457
rect 111527 72417 111540 72457
rect 111100 72401 111168 72417
rect 111224 72401 111292 72417
rect 111348 72401 111416 72417
rect 111472 72401 111540 72417
rect 111596 72417 111613 72457
rect 111720 72417 111755 72457
rect 111844 72417 111897 72457
rect 111596 72401 111664 72417
rect 111720 72401 111788 72417
rect 111844 72401 111912 72417
rect 111968 72401 112036 72457
rect 112095 72417 112172 72473
rect 112092 72401 112172 72417
rect 110122 72333 112172 72401
rect 110122 72277 110176 72333
rect 110232 72331 110300 72333
rect 110356 72331 110424 72333
rect 110480 72331 110548 72333
rect 110249 72277 110300 72331
rect 110391 72277 110424 72331
rect 110533 72277 110548 72331
rect 110604 72331 110672 72333
rect 110728 72331 110796 72333
rect 110852 72331 110920 72333
rect 110604 72277 110619 72331
rect 110728 72277 110761 72331
rect 110852 72277 110903 72331
rect 110976 72277 111044 72333
rect 111100 72331 111168 72333
rect 111224 72331 111292 72333
rect 111348 72331 111416 72333
rect 111472 72331 111540 72333
rect 111101 72277 111168 72331
rect 111243 72277 111292 72331
rect 111385 72277 111416 72331
rect 111527 72277 111540 72331
rect 111596 72331 111664 72333
rect 111720 72331 111788 72333
rect 111844 72331 111912 72333
rect 111596 72277 111613 72331
rect 111720 72277 111755 72331
rect 111844 72277 111897 72331
rect 111968 72277 112036 72333
rect 112092 72331 112172 72333
rect 110122 72275 110193 72277
rect 110249 72275 110335 72277
rect 110391 72275 110477 72277
rect 110533 72275 110619 72277
rect 110675 72275 110761 72277
rect 110817 72275 110903 72277
rect 110959 72275 111045 72277
rect 111101 72275 111187 72277
rect 111243 72275 111329 72277
rect 111385 72275 111471 72277
rect 111527 72275 111613 72277
rect 111669 72275 111755 72277
rect 111811 72275 111897 72277
rect 111953 72275 112039 72277
rect 112095 72275 112172 72331
rect 110122 72209 112172 72275
rect 110122 72153 110176 72209
rect 110232 72189 110300 72209
rect 110356 72189 110424 72209
rect 110480 72189 110548 72209
rect 110249 72153 110300 72189
rect 110391 72153 110424 72189
rect 110533 72153 110548 72189
rect 110604 72189 110672 72209
rect 110728 72189 110796 72209
rect 110852 72189 110920 72209
rect 110604 72153 110619 72189
rect 110728 72153 110761 72189
rect 110852 72153 110903 72189
rect 110976 72153 111044 72209
rect 111100 72189 111168 72209
rect 111224 72189 111292 72209
rect 111348 72189 111416 72209
rect 111472 72189 111540 72209
rect 111101 72153 111168 72189
rect 111243 72153 111292 72189
rect 111385 72153 111416 72189
rect 111527 72153 111540 72189
rect 111596 72189 111664 72209
rect 111720 72189 111788 72209
rect 111844 72189 111912 72209
rect 111596 72153 111613 72189
rect 111720 72153 111755 72189
rect 111844 72153 111897 72189
rect 111968 72153 112036 72209
rect 112092 72189 112172 72209
rect 110122 72133 110193 72153
rect 110249 72133 110335 72153
rect 110391 72133 110477 72153
rect 110533 72133 110619 72153
rect 110675 72133 110761 72153
rect 110817 72133 110903 72153
rect 110959 72133 111045 72153
rect 111101 72133 111187 72153
rect 111243 72133 111329 72153
rect 111385 72133 111471 72153
rect 111527 72133 111613 72153
rect 111669 72133 111755 72153
rect 111811 72133 111897 72153
rect 111953 72133 112039 72153
rect 112095 72133 112172 72189
rect 110122 72088 112172 72133
rect 112828 74035 114878 74088
rect 112828 73979 113325 74035
rect 113381 73979 113467 74035
rect 113523 73979 113609 74035
rect 113665 73979 113751 74035
rect 113807 73979 113893 74035
rect 113949 73979 114035 74035
rect 114091 73979 114177 74035
rect 114233 73979 114319 74035
rect 114375 73979 114461 74035
rect 114517 73979 114603 74035
rect 114659 73979 114745 74035
rect 114801 73979 114878 74035
rect 112828 73945 114878 73979
rect 112828 73889 112882 73945
rect 112938 73889 113006 73945
rect 113062 73889 113130 73945
rect 113186 73889 113254 73945
rect 113310 73893 113378 73945
rect 113434 73893 113502 73945
rect 113558 73893 113626 73945
rect 113310 73889 113325 73893
rect 113434 73889 113467 73893
rect 113558 73889 113609 73893
rect 113682 73889 113750 73945
rect 113806 73893 113874 73945
rect 113930 73893 113998 73945
rect 114054 73893 114122 73945
rect 114178 73893 114246 73945
rect 113807 73889 113874 73893
rect 113949 73889 113998 73893
rect 114091 73889 114122 73893
rect 114233 73889 114246 73893
rect 114302 73893 114370 73945
rect 114426 73893 114494 73945
rect 114550 73893 114618 73945
rect 114302 73889 114319 73893
rect 114426 73889 114461 73893
rect 114550 73889 114603 73893
rect 114674 73889 114742 73945
rect 114798 73893 114878 73945
rect 112828 73837 113325 73889
rect 113381 73837 113467 73889
rect 113523 73837 113609 73889
rect 113665 73837 113751 73889
rect 113807 73837 113893 73889
rect 113949 73837 114035 73889
rect 114091 73837 114177 73889
rect 114233 73837 114319 73889
rect 114375 73837 114461 73889
rect 114517 73837 114603 73889
rect 114659 73837 114745 73889
rect 114801 73837 114878 73893
rect 112828 73821 114878 73837
rect 112828 73765 112882 73821
rect 112938 73765 113006 73821
rect 113062 73765 113130 73821
rect 113186 73765 113254 73821
rect 113310 73765 113378 73821
rect 113434 73765 113502 73821
rect 113558 73765 113626 73821
rect 113682 73765 113750 73821
rect 113806 73765 113874 73821
rect 113930 73765 113998 73821
rect 114054 73765 114122 73821
rect 114178 73765 114246 73821
rect 114302 73765 114370 73821
rect 114426 73765 114494 73821
rect 114550 73765 114618 73821
rect 114674 73765 114742 73821
rect 114798 73765 114878 73821
rect 112828 73751 114878 73765
rect 112828 73697 113325 73751
rect 113381 73697 113467 73751
rect 113523 73697 113609 73751
rect 113665 73697 113751 73751
rect 113807 73697 113893 73751
rect 113949 73697 114035 73751
rect 114091 73697 114177 73751
rect 114233 73697 114319 73751
rect 114375 73697 114461 73751
rect 114517 73697 114603 73751
rect 114659 73697 114745 73751
rect 112828 73641 112882 73697
rect 112938 73641 113006 73697
rect 113062 73641 113130 73697
rect 113186 73641 113254 73697
rect 113310 73695 113325 73697
rect 113434 73695 113467 73697
rect 113558 73695 113609 73697
rect 113310 73641 113378 73695
rect 113434 73641 113502 73695
rect 113558 73641 113626 73695
rect 113682 73641 113750 73697
rect 113807 73695 113874 73697
rect 113949 73695 113998 73697
rect 114091 73695 114122 73697
rect 114233 73695 114246 73697
rect 113806 73641 113874 73695
rect 113930 73641 113998 73695
rect 114054 73641 114122 73695
rect 114178 73641 114246 73695
rect 114302 73695 114319 73697
rect 114426 73695 114461 73697
rect 114550 73695 114603 73697
rect 114302 73641 114370 73695
rect 114426 73641 114494 73695
rect 114550 73641 114618 73695
rect 114674 73641 114742 73697
rect 114801 73695 114878 73751
rect 114798 73641 114878 73695
rect 112828 73609 114878 73641
rect 112828 73573 113325 73609
rect 113381 73573 113467 73609
rect 113523 73573 113609 73609
rect 113665 73573 113751 73609
rect 113807 73573 113893 73609
rect 113949 73573 114035 73609
rect 114091 73573 114177 73609
rect 114233 73573 114319 73609
rect 114375 73573 114461 73609
rect 114517 73573 114603 73609
rect 114659 73573 114745 73609
rect 112828 73517 112882 73573
rect 112938 73517 113006 73573
rect 113062 73517 113130 73573
rect 113186 73517 113254 73573
rect 113310 73553 113325 73573
rect 113434 73553 113467 73573
rect 113558 73553 113609 73573
rect 113310 73517 113378 73553
rect 113434 73517 113502 73553
rect 113558 73517 113626 73553
rect 113682 73517 113750 73573
rect 113807 73553 113874 73573
rect 113949 73553 113998 73573
rect 114091 73553 114122 73573
rect 114233 73553 114246 73573
rect 113806 73517 113874 73553
rect 113930 73517 113998 73553
rect 114054 73517 114122 73553
rect 114178 73517 114246 73553
rect 114302 73553 114319 73573
rect 114426 73553 114461 73573
rect 114550 73553 114603 73573
rect 114302 73517 114370 73553
rect 114426 73517 114494 73553
rect 114550 73517 114618 73553
rect 114674 73517 114742 73573
rect 114801 73553 114878 73609
rect 114798 73517 114878 73553
rect 112828 73467 114878 73517
rect 112828 73449 113325 73467
rect 113381 73449 113467 73467
rect 113523 73449 113609 73467
rect 113665 73449 113751 73467
rect 113807 73449 113893 73467
rect 113949 73449 114035 73467
rect 114091 73449 114177 73467
rect 114233 73449 114319 73467
rect 114375 73449 114461 73467
rect 114517 73449 114603 73467
rect 114659 73449 114745 73467
rect 112828 73393 112882 73449
rect 112938 73393 113006 73449
rect 113062 73393 113130 73449
rect 113186 73393 113254 73449
rect 113310 73411 113325 73449
rect 113434 73411 113467 73449
rect 113558 73411 113609 73449
rect 113310 73393 113378 73411
rect 113434 73393 113502 73411
rect 113558 73393 113626 73411
rect 113682 73393 113750 73449
rect 113807 73411 113874 73449
rect 113949 73411 113998 73449
rect 114091 73411 114122 73449
rect 114233 73411 114246 73449
rect 113806 73393 113874 73411
rect 113930 73393 113998 73411
rect 114054 73393 114122 73411
rect 114178 73393 114246 73411
rect 114302 73411 114319 73449
rect 114426 73411 114461 73449
rect 114550 73411 114603 73449
rect 114302 73393 114370 73411
rect 114426 73393 114494 73411
rect 114550 73393 114618 73411
rect 114674 73393 114742 73449
rect 114801 73411 114878 73467
rect 114798 73393 114878 73411
rect 112828 73325 114878 73393
rect 112828 73269 112882 73325
rect 112938 73269 113006 73325
rect 113062 73269 113130 73325
rect 113186 73269 113254 73325
rect 113310 73269 113325 73325
rect 113434 73269 113467 73325
rect 113558 73269 113609 73325
rect 113682 73269 113750 73325
rect 113807 73269 113874 73325
rect 113949 73269 113998 73325
rect 114091 73269 114122 73325
rect 114233 73269 114246 73325
rect 114302 73269 114319 73325
rect 114426 73269 114461 73325
rect 114550 73269 114603 73325
rect 114674 73269 114742 73325
rect 114801 73269 114878 73325
rect 112828 73201 114878 73269
rect 112828 73145 112882 73201
rect 112938 73145 113006 73201
rect 113062 73145 113130 73201
rect 113186 73145 113254 73201
rect 113310 73183 113378 73201
rect 113434 73183 113502 73201
rect 113558 73183 113626 73201
rect 113310 73145 113325 73183
rect 113434 73145 113467 73183
rect 113558 73145 113609 73183
rect 113682 73145 113750 73201
rect 113806 73183 113874 73201
rect 113930 73183 113998 73201
rect 114054 73183 114122 73201
rect 114178 73183 114246 73201
rect 113807 73145 113874 73183
rect 113949 73145 113998 73183
rect 114091 73145 114122 73183
rect 114233 73145 114246 73183
rect 114302 73183 114370 73201
rect 114426 73183 114494 73201
rect 114550 73183 114618 73201
rect 114302 73145 114319 73183
rect 114426 73145 114461 73183
rect 114550 73145 114603 73183
rect 114674 73145 114742 73201
rect 114798 73183 114878 73201
rect 112828 73127 113325 73145
rect 113381 73127 113467 73145
rect 113523 73127 113609 73145
rect 113665 73127 113751 73145
rect 113807 73127 113893 73145
rect 113949 73127 114035 73145
rect 114091 73127 114177 73145
rect 114233 73127 114319 73145
rect 114375 73127 114461 73145
rect 114517 73127 114603 73145
rect 114659 73127 114745 73145
rect 114801 73127 114878 73183
rect 112828 73077 114878 73127
rect 112828 73021 112882 73077
rect 112938 73021 113006 73077
rect 113062 73021 113130 73077
rect 113186 73021 113254 73077
rect 113310 73041 113378 73077
rect 113434 73041 113502 73077
rect 113558 73041 113626 73077
rect 113310 73021 113325 73041
rect 113434 73021 113467 73041
rect 113558 73021 113609 73041
rect 113682 73021 113750 73077
rect 113806 73041 113874 73077
rect 113930 73041 113998 73077
rect 114054 73041 114122 73077
rect 114178 73041 114246 73077
rect 113807 73021 113874 73041
rect 113949 73021 113998 73041
rect 114091 73021 114122 73041
rect 114233 73021 114246 73041
rect 114302 73041 114370 73077
rect 114426 73041 114494 73077
rect 114550 73041 114618 73077
rect 114302 73021 114319 73041
rect 114426 73021 114461 73041
rect 114550 73021 114603 73041
rect 114674 73021 114742 73077
rect 114798 73041 114878 73077
rect 112828 72985 113325 73021
rect 113381 72985 113467 73021
rect 113523 72985 113609 73021
rect 113665 72985 113751 73021
rect 113807 72985 113893 73021
rect 113949 72985 114035 73021
rect 114091 72985 114177 73021
rect 114233 72985 114319 73021
rect 114375 72985 114461 73021
rect 114517 72985 114603 73021
rect 114659 72985 114745 73021
rect 114801 72985 114878 73041
rect 112828 72953 114878 72985
rect 112828 72897 112882 72953
rect 112938 72897 113006 72953
rect 113062 72897 113130 72953
rect 113186 72897 113254 72953
rect 113310 72899 113378 72953
rect 113434 72899 113502 72953
rect 113558 72899 113626 72953
rect 113310 72897 113325 72899
rect 113434 72897 113467 72899
rect 113558 72897 113609 72899
rect 113682 72897 113750 72953
rect 113806 72899 113874 72953
rect 113930 72899 113998 72953
rect 114054 72899 114122 72953
rect 114178 72899 114246 72953
rect 113807 72897 113874 72899
rect 113949 72897 113998 72899
rect 114091 72897 114122 72899
rect 114233 72897 114246 72899
rect 114302 72899 114370 72953
rect 114426 72899 114494 72953
rect 114550 72899 114618 72953
rect 114302 72897 114319 72899
rect 114426 72897 114461 72899
rect 114550 72897 114603 72899
rect 114674 72897 114742 72953
rect 114798 72899 114878 72953
rect 112828 72843 113325 72897
rect 113381 72843 113467 72897
rect 113523 72843 113609 72897
rect 113665 72843 113751 72897
rect 113807 72843 113893 72897
rect 113949 72843 114035 72897
rect 114091 72843 114177 72897
rect 114233 72843 114319 72897
rect 114375 72843 114461 72897
rect 114517 72843 114603 72897
rect 114659 72843 114745 72897
rect 114801 72843 114878 72899
rect 112828 72829 114878 72843
rect 112828 72773 112882 72829
rect 112938 72773 113006 72829
rect 113062 72773 113130 72829
rect 113186 72773 113254 72829
rect 113310 72773 113378 72829
rect 113434 72773 113502 72829
rect 113558 72773 113626 72829
rect 113682 72773 113750 72829
rect 113806 72773 113874 72829
rect 113930 72773 113998 72829
rect 114054 72773 114122 72829
rect 114178 72773 114246 72829
rect 114302 72773 114370 72829
rect 114426 72773 114494 72829
rect 114550 72773 114618 72829
rect 114674 72773 114742 72829
rect 114798 72773 114878 72829
rect 112828 72757 114878 72773
rect 112828 72705 113325 72757
rect 113381 72705 113467 72757
rect 113523 72705 113609 72757
rect 113665 72705 113751 72757
rect 113807 72705 113893 72757
rect 113949 72705 114035 72757
rect 114091 72705 114177 72757
rect 114233 72705 114319 72757
rect 114375 72705 114461 72757
rect 114517 72705 114603 72757
rect 114659 72705 114745 72757
rect 112828 72649 112882 72705
rect 112938 72649 113006 72705
rect 113062 72649 113130 72705
rect 113186 72649 113254 72705
rect 113310 72701 113325 72705
rect 113434 72701 113467 72705
rect 113558 72701 113609 72705
rect 113310 72649 113378 72701
rect 113434 72649 113502 72701
rect 113558 72649 113626 72701
rect 113682 72649 113750 72705
rect 113807 72701 113874 72705
rect 113949 72701 113998 72705
rect 114091 72701 114122 72705
rect 114233 72701 114246 72705
rect 113806 72649 113874 72701
rect 113930 72649 113998 72701
rect 114054 72649 114122 72701
rect 114178 72649 114246 72701
rect 114302 72701 114319 72705
rect 114426 72701 114461 72705
rect 114550 72701 114603 72705
rect 114302 72649 114370 72701
rect 114426 72649 114494 72701
rect 114550 72649 114618 72701
rect 114674 72649 114742 72705
rect 114801 72701 114878 72757
rect 114798 72649 114878 72701
rect 112828 72615 114878 72649
rect 112828 72581 113325 72615
rect 113381 72581 113467 72615
rect 113523 72581 113609 72615
rect 113665 72581 113751 72615
rect 113807 72581 113893 72615
rect 113949 72581 114035 72615
rect 114091 72581 114177 72615
rect 114233 72581 114319 72615
rect 114375 72581 114461 72615
rect 114517 72581 114603 72615
rect 114659 72581 114745 72615
rect 112828 72525 112882 72581
rect 112938 72525 113006 72581
rect 113062 72525 113130 72581
rect 113186 72525 113254 72581
rect 113310 72559 113325 72581
rect 113434 72559 113467 72581
rect 113558 72559 113609 72581
rect 113310 72525 113378 72559
rect 113434 72525 113502 72559
rect 113558 72525 113626 72559
rect 113682 72525 113750 72581
rect 113807 72559 113874 72581
rect 113949 72559 113998 72581
rect 114091 72559 114122 72581
rect 114233 72559 114246 72581
rect 113806 72525 113874 72559
rect 113930 72525 113998 72559
rect 114054 72525 114122 72559
rect 114178 72525 114246 72559
rect 114302 72559 114319 72581
rect 114426 72559 114461 72581
rect 114550 72559 114603 72581
rect 114302 72525 114370 72559
rect 114426 72525 114494 72559
rect 114550 72525 114618 72559
rect 114674 72525 114742 72581
rect 114801 72559 114878 72615
rect 114798 72525 114878 72559
rect 112828 72473 114878 72525
rect 112828 72457 113325 72473
rect 113381 72457 113467 72473
rect 113523 72457 113609 72473
rect 113665 72457 113751 72473
rect 113807 72457 113893 72473
rect 113949 72457 114035 72473
rect 114091 72457 114177 72473
rect 114233 72457 114319 72473
rect 114375 72457 114461 72473
rect 114517 72457 114603 72473
rect 114659 72457 114745 72473
rect 112828 72401 112882 72457
rect 112938 72401 113006 72457
rect 113062 72401 113130 72457
rect 113186 72401 113254 72457
rect 113310 72417 113325 72457
rect 113434 72417 113467 72457
rect 113558 72417 113609 72457
rect 113310 72401 113378 72417
rect 113434 72401 113502 72417
rect 113558 72401 113626 72417
rect 113682 72401 113750 72457
rect 113807 72417 113874 72457
rect 113949 72417 113998 72457
rect 114091 72417 114122 72457
rect 114233 72417 114246 72457
rect 113806 72401 113874 72417
rect 113930 72401 113998 72417
rect 114054 72401 114122 72417
rect 114178 72401 114246 72417
rect 114302 72417 114319 72457
rect 114426 72417 114461 72457
rect 114550 72417 114603 72457
rect 114302 72401 114370 72417
rect 114426 72401 114494 72417
rect 114550 72401 114618 72417
rect 114674 72401 114742 72457
rect 114801 72417 114878 72473
rect 114798 72401 114878 72417
rect 112828 72333 114878 72401
rect 112828 72277 112882 72333
rect 112938 72277 113006 72333
rect 113062 72277 113130 72333
rect 113186 72277 113254 72333
rect 113310 72331 113378 72333
rect 113434 72331 113502 72333
rect 113558 72331 113626 72333
rect 113310 72277 113325 72331
rect 113434 72277 113467 72331
rect 113558 72277 113609 72331
rect 113682 72277 113750 72333
rect 113806 72331 113874 72333
rect 113930 72331 113998 72333
rect 114054 72331 114122 72333
rect 114178 72331 114246 72333
rect 113807 72277 113874 72331
rect 113949 72277 113998 72331
rect 114091 72277 114122 72331
rect 114233 72277 114246 72331
rect 114302 72331 114370 72333
rect 114426 72331 114494 72333
rect 114550 72331 114618 72333
rect 114302 72277 114319 72331
rect 114426 72277 114461 72331
rect 114550 72277 114603 72331
rect 114674 72277 114742 72333
rect 114798 72331 114878 72333
rect 112828 72275 113325 72277
rect 113381 72275 113467 72277
rect 113523 72275 113609 72277
rect 113665 72275 113751 72277
rect 113807 72275 113893 72277
rect 113949 72275 114035 72277
rect 114091 72275 114177 72277
rect 114233 72275 114319 72277
rect 114375 72275 114461 72277
rect 114517 72275 114603 72277
rect 114659 72275 114745 72277
rect 114801 72275 114878 72331
rect 112828 72209 114878 72275
rect 112828 72153 112882 72209
rect 112938 72153 113006 72209
rect 113062 72153 113130 72209
rect 113186 72153 113254 72209
rect 113310 72189 113378 72209
rect 113434 72189 113502 72209
rect 113558 72189 113626 72209
rect 113310 72153 113325 72189
rect 113434 72153 113467 72189
rect 113558 72153 113609 72189
rect 113682 72153 113750 72209
rect 113806 72189 113874 72209
rect 113930 72189 113998 72209
rect 114054 72189 114122 72209
rect 114178 72189 114246 72209
rect 113807 72153 113874 72189
rect 113949 72153 113998 72189
rect 114091 72153 114122 72189
rect 114233 72153 114246 72189
rect 114302 72189 114370 72209
rect 114426 72189 114494 72209
rect 114550 72189 114618 72209
rect 114302 72153 114319 72189
rect 114426 72153 114461 72189
rect 114550 72153 114603 72189
rect 114674 72153 114742 72209
rect 114798 72189 114878 72209
rect 112828 72133 113325 72153
rect 113381 72133 113467 72153
rect 113523 72133 113609 72153
rect 113665 72133 113751 72153
rect 113807 72133 113893 72153
rect 113949 72133 114035 72153
rect 114091 72133 114177 72153
rect 114233 72133 114319 72153
rect 114375 72133 114461 72153
rect 114517 72133 114603 72153
rect 114659 72133 114745 72153
rect 114801 72133 114878 72189
rect 112828 72088 114878 72133
rect 115198 74035 117248 74088
rect 115198 73979 115269 74035
rect 115325 73979 115411 74035
rect 115467 73979 115553 74035
rect 115609 73979 115695 74035
rect 115751 73979 115837 74035
rect 115893 73979 115979 74035
rect 116035 73979 116121 74035
rect 116177 73979 116263 74035
rect 116319 73979 116405 74035
rect 116461 73979 116547 74035
rect 116603 73979 116689 74035
rect 116745 73979 116831 74035
rect 116887 73979 116973 74035
rect 117029 73979 117115 74035
rect 117171 73979 117248 74035
rect 115198 73945 117248 73979
rect 115198 73889 115252 73945
rect 115308 73893 115376 73945
rect 115432 73893 115500 73945
rect 115556 73893 115624 73945
rect 115325 73889 115376 73893
rect 115467 73889 115500 73893
rect 115609 73889 115624 73893
rect 115680 73893 115748 73945
rect 115804 73893 115872 73945
rect 115928 73893 115996 73945
rect 115680 73889 115695 73893
rect 115804 73889 115837 73893
rect 115928 73889 115979 73893
rect 116052 73889 116120 73945
rect 116176 73893 116244 73945
rect 116300 73893 116368 73945
rect 116424 73893 116492 73945
rect 116548 73893 116616 73945
rect 116177 73889 116244 73893
rect 116319 73889 116368 73893
rect 116461 73889 116492 73893
rect 116603 73889 116616 73893
rect 116672 73893 116740 73945
rect 116796 73893 116864 73945
rect 116920 73893 116988 73945
rect 116672 73889 116689 73893
rect 116796 73889 116831 73893
rect 116920 73889 116973 73893
rect 117044 73889 117112 73945
rect 117168 73893 117248 73945
rect 115198 73837 115269 73889
rect 115325 73837 115411 73889
rect 115467 73837 115553 73889
rect 115609 73837 115695 73889
rect 115751 73837 115837 73889
rect 115893 73837 115979 73889
rect 116035 73837 116121 73889
rect 116177 73837 116263 73889
rect 116319 73837 116405 73889
rect 116461 73837 116547 73889
rect 116603 73837 116689 73889
rect 116745 73837 116831 73889
rect 116887 73837 116973 73889
rect 117029 73837 117115 73889
rect 117171 73837 117248 73893
rect 115198 73821 117248 73837
rect 115198 73765 115252 73821
rect 115308 73765 115376 73821
rect 115432 73765 115500 73821
rect 115556 73765 115624 73821
rect 115680 73765 115748 73821
rect 115804 73765 115872 73821
rect 115928 73765 115996 73821
rect 116052 73765 116120 73821
rect 116176 73765 116244 73821
rect 116300 73765 116368 73821
rect 116424 73765 116492 73821
rect 116548 73765 116616 73821
rect 116672 73765 116740 73821
rect 116796 73765 116864 73821
rect 116920 73765 116988 73821
rect 117044 73765 117112 73821
rect 117168 73765 117248 73821
rect 115198 73751 117248 73765
rect 115198 73697 115269 73751
rect 115325 73697 115411 73751
rect 115467 73697 115553 73751
rect 115609 73697 115695 73751
rect 115751 73697 115837 73751
rect 115893 73697 115979 73751
rect 116035 73697 116121 73751
rect 116177 73697 116263 73751
rect 116319 73697 116405 73751
rect 116461 73697 116547 73751
rect 116603 73697 116689 73751
rect 116745 73697 116831 73751
rect 116887 73697 116973 73751
rect 117029 73697 117115 73751
rect 115198 73641 115252 73697
rect 115325 73695 115376 73697
rect 115467 73695 115500 73697
rect 115609 73695 115624 73697
rect 115308 73641 115376 73695
rect 115432 73641 115500 73695
rect 115556 73641 115624 73695
rect 115680 73695 115695 73697
rect 115804 73695 115837 73697
rect 115928 73695 115979 73697
rect 115680 73641 115748 73695
rect 115804 73641 115872 73695
rect 115928 73641 115996 73695
rect 116052 73641 116120 73697
rect 116177 73695 116244 73697
rect 116319 73695 116368 73697
rect 116461 73695 116492 73697
rect 116603 73695 116616 73697
rect 116176 73641 116244 73695
rect 116300 73641 116368 73695
rect 116424 73641 116492 73695
rect 116548 73641 116616 73695
rect 116672 73695 116689 73697
rect 116796 73695 116831 73697
rect 116920 73695 116973 73697
rect 116672 73641 116740 73695
rect 116796 73641 116864 73695
rect 116920 73641 116988 73695
rect 117044 73641 117112 73697
rect 117171 73695 117248 73751
rect 117168 73641 117248 73695
rect 115198 73609 117248 73641
rect 115198 73573 115269 73609
rect 115325 73573 115411 73609
rect 115467 73573 115553 73609
rect 115609 73573 115695 73609
rect 115751 73573 115837 73609
rect 115893 73573 115979 73609
rect 116035 73573 116121 73609
rect 116177 73573 116263 73609
rect 116319 73573 116405 73609
rect 116461 73573 116547 73609
rect 116603 73573 116689 73609
rect 116745 73573 116831 73609
rect 116887 73573 116973 73609
rect 117029 73573 117115 73609
rect 115198 73517 115252 73573
rect 115325 73553 115376 73573
rect 115467 73553 115500 73573
rect 115609 73553 115624 73573
rect 115308 73517 115376 73553
rect 115432 73517 115500 73553
rect 115556 73517 115624 73553
rect 115680 73553 115695 73573
rect 115804 73553 115837 73573
rect 115928 73553 115979 73573
rect 115680 73517 115748 73553
rect 115804 73517 115872 73553
rect 115928 73517 115996 73553
rect 116052 73517 116120 73573
rect 116177 73553 116244 73573
rect 116319 73553 116368 73573
rect 116461 73553 116492 73573
rect 116603 73553 116616 73573
rect 116176 73517 116244 73553
rect 116300 73517 116368 73553
rect 116424 73517 116492 73553
rect 116548 73517 116616 73553
rect 116672 73553 116689 73573
rect 116796 73553 116831 73573
rect 116920 73553 116973 73573
rect 116672 73517 116740 73553
rect 116796 73517 116864 73553
rect 116920 73517 116988 73553
rect 117044 73517 117112 73573
rect 117171 73553 117248 73609
rect 117168 73517 117248 73553
rect 115198 73467 117248 73517
rect 115198 73449 115269 73467
rect 115325 73449 115411 73467
rect 115467 73449 115553 73467
rect 115609 73449 115695 73467
rect 115751 73449 115837 73467
rect 115893 73449 115979 73467
rect 116035 73449 116121 73467
rect 116177 73449 116263 73467
rect 116319 73449 116405 73467
rect 116461 73449 116547 73467
rect 116603 73449 116689 73467
rect 116745 73449 116831 73467
rect 116887 73449 116973 73467
rect 117029 73449 117115 73467
rect 115198 73393 115252 73449
rect 115325 73411 115376 73449
rect 115467 73411 115500 73449
rect 115609 73411 115624 73449
rect 115308 73393 115376 73411
rect 115432 73393 115500 73411
rect 115556 73393 115624 73411
rect 115680 73411 115695 73449
rect 115804 73411 115837 73449
rect 115928 73411 115979 73449
rect 115680 73393 115748 73411
rect 115804 73393 115872 73411
rect 115928 73393 115996 73411
rect 116052 73393 116120 73449
rect 116177 73411 116244 73449
rect 116319 73411 116368 73449
rect 116461 73411 116492 73449
rect 116603 73411 116616 73449
rect 116176 73393 116244 73411
rect 116300 73393 116368 73411
rect 116424 73393 116492 73411
rect 116548 73393 116616 73411
rect 116672 73411 116689 73449
rect 116796 73411 116831 73449
rect 116920 73411 116973 73449
rect 116672 73393 116740 73411
rect 116796 73393 116864 73411
rect 116920 73393 116988 73411
rect 117044 73393 117112 73449
rect 117171 73411 117248 73467
rect 117168 73393 117248 73411
rect 115198 73325 117248 73393
rect 115198 73269 115252 73325
rect 115325 73269 115376 73325
rect 115467 73269 115500 73325
rect 115609 73269 115624 73325
rect 115680 73269 115695 73325
rect 115804 73269 115837 73325
rect 115928 73269 115979 73325
rect 116052 73269 116120 73325
rect 116177 73269 116244 73325
rect 116319 73269 116368 73325
rect 116461 73269 116492 73325
rect 116603 73269 116616 73325
rect 116672 73269 116689 73325
rect 116796 73269 116831 73325
rect 116920 73269 116973 73325
rect 117044 73269 117112 73325
rect 117171 73269 117248 73325
rect 115198 73201 117248 73269
rect 115198 73145 115252 73201
rect 115308 73183 115376 73201
rect 115432 73183 115500 73201
rect 115556 73183 115624 73201
rect 115325 73145 115376 73183
rect 115467 73145 115500 73183
rect 115609 73145 115624 73183
rect 115680 73183 115748 73201
rect 115804 73183 115872 73201
rect 115928 73183 115996 73201
rect 115680 73145 115695 73183
rect 115804 73145 115837 73183
rect 115928 73145 115979 73183
rect 116052 73145 116120 73201
rect 116176 73183 116244 73201
rect 116300 73183 116368 73201
rect 116424 73183 116492 73201
rect 116548 73183 116616 73201
rect 116177 73145 116244 73183
rect 116319 73145 116368 73183
rect 116461 73145 116492 73183
rect 116603 73145 116616 73183
rect 116672 73183 116740 73201
rect 116796 73183 116864 73201
rect 116920 73183 116988 73201
rect 116672 73145 116689 73183
rect 116796 73145 116831 73183
rect 116920 73145 116973 73183
rect 117044 73145 117112 73201
rect 117168 73183 117248 73201
rect 115198 73127 115269 73145
rect 115325 73127 115411 73145
rect 115467 73127 115553 73145
rect 115609 73127 115695 73145
rect 115751 73127 115837 73145
rect 115893 73127 115979 73145
rect 116035 73127 116121 73145
rect 116177 73127 116263 73145
rect 116319 73127 116405 73145
rect 116461 73127 116547 73145
rect 116603 73127 116689 73145
rect 116745 73127 116831 73145
rect 116887 73127 116973 73145
rect 117029 73127 117115 73145
rect 117171 73127 117248 73183
rect 115198 73077 117248 73127
rect 115198 73021 115252 73077
rect 115308 73041 115376 73077
rect 115432 73041 115500 73077
rect 115556 73041 115624 73077
rect 115325 73021 115376 73041
rect 115467 73021 115500 73041
rect 115609 73021 115624 73041
rect 115680 73041 115748 73077
rect 115804 73041 115872 73077
rect 115928 73041 115996 73077
rect 115680 73021 115695 73041
rect 115804 73021 115837 73041
rect 115928 73021 115979 73041
rect 116052 73021 116120 73077
rect 116176 73041 116244 73077
rect 116300 73041 116368 73077
rect 116424 73041 116492 73077
rect 116548 73041 116616 73077
rect 116177 73021 116244 73041
rect 116319 73021 116368 73041
rect 116461 73021 116492 73041
rect 116603 73021 116616 73041
rect 116672 73041 116740 73077
rect 116796 73041 116864 73077
rect 116920 73041 116988 73077
rect 116672 73021 116689 73041
rect 116796 73021 116831 73041
rect 116920 73021 116973 73041
rect 117044 73021 117112 73077
rect 117168 73041 117248 73077
rect 115198 72985 115269 73021
rect 115325 72985 115411 73021
rect 115467 72985 115553 73021
rect 115609 72985 115695 73021
rect 115751 72985 115837 73021
rect 115893 72985 115979 73021
rect 116035 72985 116121 73021
rect 116177 72985 116263 73021
rect 116319 72985 116405 73021
rect 116461 72985 116547 73021
rect 116603 72985 116689 73021
rect 116745 72985 116831 73021
rect 116887 72985 116973 73021
rect 117029 72985 117115 73021
rect 117171 72985 117248 73041
rect 115198 72953 117248 72985
rect 115198 72897 115252 72953
rect 115308 72899 115376 72953
rect 115432 72899 115500 72953
rect 115556 72899 115624 72953
rect 115325 72897 115376 72899
rect 115467 72897 115500 72899
rect 115609 72897 115624 72899
rect 115680 72899 115748 72953
rect 115804 72899 115872 72953
rect 115928 72899 115996 72953
rect 115680 72897 115695 72899
rect 115804 72897 115837 72899
rect 115928 72897 115979 72899
rect 116052 72897 116120 72953
rect 116176 72899 116244 72953
rect 116300 72899 116368 72953
rect 116424 72899 116492 72953
rect 116548 72899 116616 72953
rect 116177 72897 116244 72899
rect 116319 72897 116368 72899
rect 116461 72897 116492 72899
rect 116603 72897 116616 72899
rect 116672 72899 116740 72953
rect 116796 72899 116864 72953
rect 116920 72899 116988 72953
rect 116672 72897 116689 72899
rect 116796 72897 116831 72899
rect 116920 72897 116973 72899
rect 117044 72897 117112 72953
rect 117168 72899 117248 72953
rect 115198 72843 115269 72897
rect 115325 72843 115411 72897
rect 115467 72843 115553 72897
rect 115609 72843 115695 72897
rect 115751 72843 115837 72897
rect 115893 72843 115979 72897
rect 116035 72843 116121 72897
rect 116177 72843 116263 72897
rect 116319 72843 116405 72897
rect 116461 72843 116547 72897
rect 116603 72843 116689 72897
rect 116745 72843 116831 72897
rect 116887 72843 116973 72897
rect 117029 72843 117115 72897
rect 117171 72843 117248 72899
rect 115198 72829 117248 72843
rect 115198 72773 115252 72829
rect 115308 72773 115376 72829
rect 115432 72773 115500 72829
rect 115556 72773 115624 72829
rect 115680 72773 115748 72829
rect 115804 72773 115872 72829
rect 115928 72773 115996 72829
rect 116052 72773 116120 72829
rect 116176 72773 116244 72829
rect 116300 72773 116368 72829
rect 116424 72773 116492 72829
rect 116548 72773 116616 72829
rect 116672 72773 116740 72829
rect 116796 72773 116864 72829
rect 116920 72773 116988 72829
rect 117044 72773 117112 72829
rect 117168 72773 117248 72829
rect 115198 72757 117248 72773
rect 115198 72705 115269 72757
rect 115325 72705 115411 72757
rect 115467 72705 115553 72757
rect 115609 72705 115695 72757
rect 115751 72705 115837 72757
rect 115893 72705 115979 72757
rect 116035 72705 116121 72757
rect 116177 72705 116263 72757
rect 116319 72705 116405 72757
rect 116461 72705 116547 72757
rect 116603 72705 116689 72757
rect 116745 72705 116831 72757
rect 116887 72705 116973 72757
rect 117029 72705 117115 72757
rect 115198 72649 115252 72705
rect 115325 72701 115376 72705
rect 115467 72701 115500 72705
rect 115609 72701 115624 72705
rect 115308 72649 115376 72701
rect 115432 72649 115500 72701
rect 115556 72649 115624 72701
rect 115680 72701 115695 72705
rect 115804 72701 115837 72705
rect 115928 72701 115979 72705
rect 115680 72649 115748 72701
rect 115804 72649 115872 72701
rect 115928 72649 115996 72701
rect 116052 72649 116120 72705
rect 116177 72701 116244 72705
rect 116319 72701 116368 72705
rect 116461 72701 116492 72705
rect 116603 72701 116616 72705
rect 116176 72649 116244 72701
rect 116300 72649 116368 72701
rect 116424 72649 116492 72701
rect 116548 72649 116616 72701
rect 116672 72701 116689 72705
rect 116796 72701 116831 72705
rect 116920 72701 116973 72705
rect 116672 72649 116740 72701
rect 116796 72649 116864 72701
rect 116920 72649 116988 72701
rect 117044 72649 117112 72705
rect 117171 72701 117248 72757
rect 117168 72649 117248 72701
rect 115198 72615 117248 72649
rect 115198 72581 115269 72615
rect 115325 72581 115411 72615
rect 115467 72581 115553 72615
rect 115609 72581 115695 72615
rect 115751 72581 115837 72615
rect 115893 72581 115979 72615
rect 116035 72581 116121 72615
rect 116177 72581 116263 72615
rect 116319 72581 116405 72615
rect 116461 72581 116547 72615
rect 116603 72581 116689 72615
rect 116745 72581 116831 72615
rect 116887 72581 116973 72615
rect 117029 72581 117115 72615
rect 115198 72525 115252 72581
rect 115325 72559 115376 72581
rect 115467 72559 115500 72581
rect 115609 72559 115624 72581
rect 115308 72525 115376 72559
rect 115432 72525 115500 72559
rect 115556 72525 115624 72559
rect 115680 72559 115695 72581
rect 115804 72559 115837 72581
rect 115928 72559 115979 72581
rect 115680 72525 115748 72559
rect 115804 72525 115872 72559
rect 115928 72525 115996 72559
rect 116052 72525 116120 72581
rect 116177 72559 116244 72581
rect 116319 72559 116368 72581
rect 116461 72559 116492 72581
rect 116603 72559 116616 72581
rect 116176 72525 116244 72559
rect 116300 72525 116368 72559
rect 116424 72525 116492 72559
rect 116548 72525 116616 72559
rect 116672 72559 116689 72581
rect 116796 72559 116831 72581
rect 116920 72559 116973 72581
rect 116672 72525 116740 72559
rect 116796 72525 116864 72559
rect 116920 72525 116988 72559
rect 117044 72525 117112 72581
rect 117171 72559 117248 72615
rect 117168 72525 117248 72559
rect 115198 72473 117248 72525
rect 115198 72457 115269 72473
rect 115325 72457 115411 72473
rect 115467 72457 115553 72473
rect 115609 72457 115695 72473
rect 115751 72457 115837 72473
rect 115893 72457 115979 72473
rect 116035 72457 116121 72473
rect 116177 72457 116263 72473
rect 116319 72457 116405 72473
rect 116461 72457 116547 72473
rect 116603 72457 116689 72473
rect 116745 72457 116831 72473
rect 116887 72457 116973 72473
rect 117029 72457 117115 72473
rect 115198 72401 115252 72457
rect 115325 72417 115376 72457
rect 115467 72417 115500 72457
rect 115609 72417 115624 72457
rect 115308 72401 115376 72417
rect 115432 72401 115500 72417
rect 115556 72401 115624 72417
rect 115680 72417 115695 72457
rect 115804 72417 115837 72457
rect 115928 72417 115979 72457
rect 115680 72401 115748 72417
rect 115804 72401 115872 72417
rect 115928 72401 115996 72417
rect 116052 72401 116120 72457
rect 116177 72417 116244 72457
rect 116319 72417 116368 72457
rect 116461 72417 116492 72457
rect 116603 72417 116616 72457
rect 116176 72401 116244 72417
rect 116300 72401 116368 72417
rect 116424 72401 116492 72417
rect 116548 72401 116616 72417
rect 116672 72417 116689 72457
rect 116796 72417 116831 72457
rect 116920 72417 116973 72457
rect 116672 72401 116740 72417
rect 116796 72401 116864 72417
rect 116920 72401 116988 72417
rect 117044 72401 117112 72457
rect 117171 72417 117248 72473
rect 117168 72401 117248 72417
rect 115198 72333 117248 72401
rect 115198 72277 115252 72333
rect 115308 72331 115376 72333
rect 115432 72331 115500 72333
rect 115556 72331 115624 72333
rect 115325 72277 115376 72331
rect 115467 72277 115500 72331
rect 115609 72277 115624 72331
rect 115680 72331 115748 72333
rect 115804 72331 115872 72333
rect 115928 72331 115996 72333
rect 115680 72277 115695 72331
rect 115804 72277 115837 72331
rect 115928 72277 115979 72331
rect 116052 72277 116120 72333
rect 116176 72331 116244 72333
rect 116300 72331 116368 72333
rect 116424 72331 116492 72333
rect 116548 72331 116616 72333
rect 116177 72277 116244 72331
rect 116319 72277 116368 72331
rect 116461 72277 116492 72331
rect 116603 72277 116616 72331
rect 116672 72331 116740 72333
rect 116796 72331 116864 72333
rect 116920 72331 116988 72333
rect 116672 72277 116689 72331
rect 116796 72277 116831 72331
rect 116920 72277 116973 72331
rect 117044 72277 117112 72333
rect 117168 72331 117248 72333
rect 115198 72275 115269 72277
rect 115325 72275 115411 72277
rect 115467 72275 115553 72277
rect 115609 72275 115695 72277
rect 115751 72275 115837 72277
rect 115893 72275 115979 72277
rect 116035 72275 116121 72277
rect 116177 72275 116263 72277
rect 116319 72275 116405 72277
rect 116461 72275 116547 72277
rect 116603 72275 116689 72277
rect 116745 72275 116831 72277
rect 116887 72275 116973 72277
rect 117029 72275 117115 72277
rect 117171 72275 117248 72331
rect 115198 72209 117248 72275
rect 115198 72153 115252 72209
rect 115308 72189 115376 72209
rect 115432 72189 115500 72209
rect 115556 72189 115624 72209
rect 115325 72153 115376 72189
rect 115467 72153 115500 72189
rect 115609 72153 115624 72189
rect 115680 72189 115748 72209
rect 115804 72189 115872 72209
rect 115928 72189 115996 72209
rect 115680 72153 115695 72189
rect 115804 72153 115837 72189
rect 115928 72153 115979 72189
rect 116052 72153 116120 72209
rect 116176 72189 116244 72209
rect 116300 72189 116368 72209
rect 116424 72189 116492 72209
rect 116548 72189 116616 72209
rect 116177 72153 116244 72189
rect 116319 72153 116368 72189
rect 116461 72153 116492 72189
rect 116603 72153 116616 72189
rect 116672 72189 116740 72209
rect 116796 72189 116864 72209
rect 116920 72189 116988 72209
rect 116672 72153 116689 72189
rect 116796 72153 116831 72189
rect 116920 72153 116973 72189
rect 117044 72153 117112 72209
rect 117168 72189 117248 72209
rect 115198 72133 115269 72153
rect 115325 72133 115411 72153
rect 115467 72133 115553 72153
rect 115609 72133 115695 72153
rect 115751 72133 115837 72153
rect 115893 72133 115979 72153
rect 116035 72133 116121 72153
rect 116177 72133 116263 72153
rect 116319 72133 116405 72153
rect 116461 72133 116547 72153
rect 116603 72133 116689 72153
rect 116745 72133 116831 72153
rect 116887 72133 116973 72153
rect 117029 72133 117115 72153
rect 117171 72133 117248 72189
rect 115198 72088 117248 72133
rect 117828 74035 119728 74088
rect 117828 73979 117899 74035
rect 117955 73979 118041 74035
rect 118097 73979 118183 74035
rect 118239 73979 118325 74035
rect 118381 73979 118467 74035
rect 118523 73979 118609 74035
rect 118665 73979 118751 74035
rect 118807 73979 118893 74035
rect 118949 73979 119035 74035
rect 119091 73979 119177 74035
rect 119233 73979 119319 74035
rect 119375 73979 119461 74035
rect 119517 73979 119603 74035
rect 119659 73979 119728 74035
rect 117828 73945 119728 73979
rect 117828 73889 117882 73945
rect 117938 73893 118006 73945
rect 118062 73893 118130 73945
rect 118186 73893 118254 73945
rect 117955 73889 118006 73893
rect 118097 73889 118130 73893
rect 118239 73889 118254 73893
rect 118310 73893 118378 73945
rect 118434 73893 118502 73945
rect 118558 73893 118626 73945
rect 118310 73889 118325 73893
rect 118434 73889 118467 73893
rect 118558 73889 118609 73893
rect 118682 73889 118750 73945
rect 118806 73893 118874 73945
rect 118930 73893 118998 73945
rect 119054 73893 119122 73945
rect 119178 73893 119246 73945
rect 118807 73889 118874 73893
rect 118949 73889 118998 73893
rect 119091 73889 119122 73893
rect 119233 73889 119246 73893
rect 119302 73893 119370 73945
rect 119426 73893 119494 73945
rect 119550 73893 119618 73945
rect 119302 73889 119319 73893
rect 119426 73889 119461 73893
rect 119550 73889 119603 73893
rect 119674 73889 119728 73945
rect 117828 73837 117899 73889
rect 117955 73837 118041 73889
rect 118097 73837 118183 73889
rect 118239 73837 118325 73889
rect 118381 73837 118467 73889
rect 118523 73837 118609 73889
rect 118665 73837 118751 73889
rect 118807 73837 118893 73889
rect 118949 73837 119035 73889
rect 119091 73837 119177 73889
rect 119233 73837 119319 73889
rect 119375 73837 119461 73889
rect 119517 73837 119603 73889
rect 119659 73837 119728 73889
rect 117828 73821 119728 73837
rect 117828 73765 117882 73821
rect 117938 73765 118006 73821
rect 118062 73765 118130 73821
rect 118186 73765 118254 73821
rect 118310 73765 118378 73821
rect 118434 73765 118502 73821
rect 118558 73765 118626 73821
rect 118682 73765 118750 73821
rect 118806 73765 118874 73821
rect 118930 73765 118998 73821
rect 119054 73765 119122 73821
rect 119178 73765 119246 73821
rect 119302 73765 119370 73821
rect 119426 73765 119494 73821
rect 119550 73765 119618 73821
rect 119674 73765 119728 73821
rect 117828 73751 119728 73765
rect 117828 73697 117899 73751
rect 117955 73697 118041 73751
rect 118097 73697 118183 73751
rect 118239 73697 118325 73751
rect 118381 73697 118467 73751
rect 118523 73697 118609 73751
rect 118665 73697 118751 73751
rect 118807 73697 118893 73751
rect 118949 73697 119035 73751
rect 119091 73697 119177 73751
rect 119233 73697 119319 73751
rect 119375 73697 119461 73751
rect 119517 73697 119603 73751
rect 119659 73697 119728 73751
rect 117828 73641 117882 73697
rect 117955 73695 118006 73697
rect 118097 73695 118130 73697
rect 118239 73695 118254 73697
rect 117938 73641 118006 73695
rect 118062 73641 118130 73695
rect 118186 73641 118254 73695
rect 118310 73695 118325 73697
rect 118434 73695 118467 73697
rect 118558 73695 118609 73697
rect 118310 73641 118378 73695
rect 118434 73641 118502 73695
rect 118558 73641 118626 73695
rect 118682 73641 118750 73697
rect 118807 73695 118874 73697
rect 118949 73695 118998 73697
rect 119091 73695 119122 73697
rect 119233 73695 119246 73697
rect 118806 73641 118874 73695
rect 118930 73641 118998 73695
rect 119054 73641 119122 73695
rect 119178 73641 119246 73695
rect 119302 73695 119319 73697
rect 119426 73695 119461 73697
rect 119550 73695 119603 73697
rect 119302 73641 119370 73695
rect 119426 73641 119494 73695
rect 119550 73641 119618 73695
rect 119674 73641 119728 73697
rect 117828 73609 119728 73641
rect 117828 73573 117899 73609
rect 117955 73573 118041 73609
rect 118097 73573 118183 73609
rect 118239 73573 118325 73609
rect 118381 73573 118467 73609
rect 118523 73573 118609 73609
rect 118665 73573 118751 73609
rect 118807 73573 118893 73609
rect 118949 73573 119035 73609
rect 119091 73573 119177 73609
rect 119233 73573 119319 73609
rect 119375 73573 119461 73609
rect 119517 73573 119603 73609
rect 119659 73573 119728 73609
rect 117828 73517 117882 73573
rect 117955 73553 118006 73573
rect 118097 73553 118130 73573
rect 118239 73553 118254 73573
rect 117938 73517 118006 73553
rect 118062 73517 118130 73553
rect 118186 73517 118254 73553
rect 118310 73553 118325 73573
rect 118434 73553 118467 73573
rect 118558 73553 118609 73573
rect 118310 73517 118378 73553
rect 118434 73517 118502 73553
rect 118558 73517 118626 73553
rect 118682 73517 118750 73573
rect 118807 73553 118874 73573
rect 118949 73553 118998 73573
rect 119091 73553 119122 73573
rect 119233 73553 119246 73573
rect 118806 73517 118874 73553
rect 118930 73517 118998 73553
rect 119054 73517 119122 73553
rect 119178 73517 119246 73553
rect 119302 73553 119319 73573
rect 119426 73553 119461 73573
rect 119550 73553 119603 73573
rect 119302 73517 119370 73553
rect 119426 73517 119494 73553
rect 119550 73517 119618 73553
rect 119674 73517 119728 73573
rect 117828 73467 119728 73517
rect 117828 73449 117899 73467
rect 117955 73449 118041 73467
rect 118097 73449 118183 73467
rect 118239 73449 118325 73467
rect 118381 73449 118467 73467
rect 118523 73449 118609 73467
rect 118665 73449 118751 73467
rect 118807 73449 118893 73467
rect 118949 73449 119035 73467
rect 119091 73449 119177 73467
rect 119233 73449 119319 73467
rect 119375 73449 119461 73467
rect 119517 73449 119603 73467
rect 119659 73449 119728 73467
rect 117828 73393 117882 73449
rect 117955 73411 118006 73449
rect 118097 73411 118130 73449
rect 118239 73411 118254 73449
rect 117938 73393 118006 73411
rect 118062 73393 118130 73411
rect 118186 73393 118254 73411
rect 118310 73411 118325 73449
rect 118434 73411 118467 73449
rect 118558 73411 118609 73449
rect 118310 73393 118378 73411
rect 118434 73393 118502 73411
rect 118558 73393 118626 73411
rect 118682 73393 118750 73449
rect 118807 73411 118874 73449
rect 118949 73411 118998 73449
rect 119091 73411 119122 73449
rect 119233 73411 119246 73449
rect 118806 73393 118874 73411
rect 118930 73393 118998 73411
rect 119054 73393 119122 73411
rect 119178 73393 119246 73411
rect 119302 73411 119319 73449
rect 119426 73411 119461 73449
rect 119550 73411 119603 73449
rect 119302 73393 119370 73411
rect 119426 73393 119494 73411
rect 119550 73393 119618 73411
rect 119674 73393 119728 73449
rect 117828 73325 119728 73393
rect 117828 73269 117882 73325
rect 117955 73269 118006 73325
rect 118097 73269 118130 73325
rect 118239 73269 118254 73325
rect 118310 73269 118325 73325
rect 118434 73269 118467 73325
rect 118558 73269 118609 73325
rect 118682 73269 118750 73325
rect 118807 73269 118874 73325
rect 118949 73269 118998 73325
rect 119091 73269 119122 73325
rect 119233 73269 119246 73325
rect 119302 73269 119319 73325
rect 119426 73269 119461 73325
rect 119550 73269 119603 73325
rect 119674 73269 119728 73325
rect 117828 73201 119728 73269
rect 117828 73145 117882 73201
rect 117938 73183 118006 73201
rect 118062 73183 118130 73201
rect 118186 73183 118254 73201
rect 117955 73145 118006 73183
rect 118097 73145 118130 73183
rect 118239 73145 118254 73183
rect 118310 73183 118378 73201
rect 118434 73183 118502 73201
rect 118558 73183 118626 73201
rect 118310 73145 118325 73183
rect 118434 73145 118467 73183
rect 118558 73145 118609 73183
rect 118682 73145 118750 73201
rect 118806 73183 118874 73201
rect 118930 73183 118998 73201
rect 119054 73183 119122 73201
rect 119178 73183 119246 73201
rect 118807 73145 118874 73183
rect 118949 73145 118998 73183
rect 119091 73145 119122 73183
rect 119233 73145 119246 73183
rect 119302 73183 119370 73201
rect 119426 73183 119494 73201
rect 119550 73183 119618 73201
rect 119302 73145 119319 73183
rect 119426 73145 119461 73183
rect 119550 73145 119603 73183
rect 119674 73145 119728 73201
rect 117828 73127 117899 73145
rect 117955 73127 118041 73145
rect 118097 73127 118183 73145
rect 118239 73127 118325 73145
rect 118381 73127 118467 73145
rect 118523 73127 118609 73145
rect 118665 73127 118751 73145
rect 118807 73127 118893 73145
rect 118949 73127 119035 73145
rect 119091 73127 119177 73145
rect 119233 73127 119319 73145
rect 119375 73127 119461 73145
rect 119517 73127 119603 73145
rect 119659 73127 119728 73145
rect 117828 73077 119728 73127
rect 117828 73021 117882 73077
rect 117938 73041 118006 73077
rect 118062 73041 118130 73077
rect 118186 73041 118254 73077
rect 117955 73021 118006 73041
rect 118097 73021 118130 73041
rect 118239 73021 118254 73041
rect 118310 73041 118378 73077
rect 118434 73041 118502 73077
rect 118558 73041 118626 73077
rect 118310 73021 118325 73041
rect 118434 73021 118467 73041
rect 118558 73021 118609 73041
rect 118682 73021 118750 73077
rect 118806 73041 118874 73077
rect 118930 73041 118998 73077
rect 119054 73041 119122 73077
rect 119178 73041 119246 73077
rect 118807 73021 118874 73041
rect 118949 73021 118998 73041
rect 119091 73021 119122 73041
rect 119233 73021 119246 73041
rect 119302 73041 119370 73077
rect 119426 73041 119494 73077
rect 119550 73041 119618 73077
rect 119302 73021 119319 73041
rect 119426 73021 119461 73041
rect 119550 73021 119603 73041
rect 119674 73021 119728 73077
rect 117828 72985 117899 73021
rect 117955 72985 118041 73021
rect 118097 72985 118183 73021
rect 118239 72985 118325 73021
rect 118381 72985 118467 73021
rect 118523 72985 118609 73021
rect 118665 72985 118751 73021
rect 118807 72985 118893 73021
rect 118949 72985 119035 73021
rect 119091 72985 119177 73021
rect 119233 72985 119319 73021
rect 119375 72985 119461 73021
rect 119517 72985 119603 73021
rect 119659 72985 119728 73021
rect 117828 72953 119728 72985
rect 117828 72897 117882 72953
rect 117938 72899 118006 72953
rect 118062 72899 118130 72953
rect 118186 72899 118254 72953
rect 117955 72897 118006 72899
rect 118097 72897 118130 72899
rect 118239 72897 118254 72899
rect 118310 72899 118378 72953
rect 118434 72899 118502 72953
rect 118558 72899 118626 72953
rect 118310 72897 118325 72899
rect 118434 72897 118467 72899
rect 118558 72897 118609 72899
rect 118682 72897 118750 72953
rect 118806 72899 118874 72953
rect 118930 72899 118998 72953
rect 119054 72899 119122 72953
rect 119178 72899 119246 72953
rect 118807 72897 118874 72899
rect 118949 72897 118998 72899
rect 119091 72897 119122 72899
rect 119233 72897 119246 72899
rect 119302 72899 119370 72953
rect 119426 72899 119494 72953
rect 119550 72899 119618 72953
rect 119302 72897 119319 72899
rect 119426 72897 119461 72899
rect 119550 72897 119603 72899
rect 119674 72897 119728 72953
rect 117828 72843 117899 72897
rect 117955 72843 118041 72897
rect 118097 72843 118183 72897
rect 118239 72843 118325 72897
rect 118381 72843 118467 72897
rect 118523 72843 118609 72897
rect 118665 72843 118751 72897
rect 118807 72843 118893 72897
rect 118949 72843 119035 72897
rect 119091 72843 119177 72897
rect 119233 72843 119319 72897
rect 119375 72843 119461 72897
rect 119517 72843 119603 72897
rect 119659 72843 119728 72897
rect 117828 72829 119728 72843
rect 117828 72773 117882 72829
rect 117938 72773 118006 72829
rect 118062 72773 118130 72829
rect 118186 72773 118254 72829
rect 118310 72773 118378 72829
rect 118434 72773 118502 72829
rect 118558 72773 118626 72829
rect 118682 72773 118750 72829
rect 118806 72773 118874 72829
rect 118930 72773 118998 72829
rect 119054 72773 119122 72829
rect 119178 72773 119246 72829
rect 119302 72773 119370 72829
rect 119426 72773 119494 72829
rect 119550 72773 119618 72829
rect 119674 72773 119728 72829
rect 117828 72757 119728 72773
rect 117828 72705 117899 72757
rect 117955 72705 118041 72757
rect 118097 72705 118183 72757
rect 118239 72705 118325 72757
rect 118381 72705 118467 72757
rect 118523 72705 118609 72757
rect 118665 72705 118751 72757
rect 118807 72705 118893 72757
rect 118949 72705 119035 72757
rect 119091 72705 119177 72757
rect 119233 72705 119319 72757
rect 119375 72705 119461 72757
rect 119517 72705 119603 72757
rect 119659 72705 119728 72757
rect 117828 72649 117882 72705
rect 117955 72701 118006 72705
rect 118097 72701 118130 72705
rect 118239 72701 118254 72705
rect 117938 72649 118006 72701
rect 118062 72649 118130 72701
rect 118186 72649 118254 72701
rect 118310 72701 118325 72705
rect 118434 72701 118467 72705
rect 118558 72701 118609 72705
rect 118310 72649 118378 72701
rect 118434 72649 118502 72701
rect 118558 72649 118626 72701
rect 118682 72649 118750 72705
rect 118807 72701 118874 72705
rect 118949 72701 118998 72705
rect 119091 72701 119122 72705
rect 119233 72701 119246 72705
rect 118806 72649 118874 72701
rect 118930 72649 118998 72701
rect 119054 72649 119122 72701
rect 119178 72649 119246 72701
rect 119302 72701 119319 72705
rect 119426 72701 119461 72705
rect 119550 72701 119603 72705
rect 119302 72649 119370 72701
rect 119426 72649 119494 72701
rect 119550 72649 119618 72701
rect 119674 72649 119728 72705
rect 117828 72615 119728 72649
rect 117828 72581 117899 72615
rect 117955 72581 118041 72615
rect 118097 72581 118183 72615
rect 118239 72581 118325 72615
rect 118381 72581 118467 72615
rect 118523 72581 118609 72615
rect 118665 72581 118751 72615
rect 118807 72581 118893 72615
rect 118949 72581 119035 72615
rect 119091 72581 119177 72615
rect 119233 72581 119319 72615
rect 119375 72581 119461 72615
rect 119517 72581 119603 72615
rect 119659 72581 119728 72615
rect 117828 72525 117882 72581
rect 117955 72559 118006 72581
rect 118097 72559 118130 72581
rect 118239 72559 118254 72581
rect 117938 72525 118006 72559
rect 118062 72525 118130 72559
rect 118186 72525 118254 72559
rect 118310 72559 118325 72581
rect 118434 72559 118467 72581
rect 118558 72559 118609 72581
rect 118310 72525 118378 72559
rect 118434 72525 118502 72559
rect 118558 72525 118626 72559
rect 118682 72525 118750 72581
rect 118807 72559 118874 72581
rect 118949 72559 118998 72581
rect 119091 72559 119122 72581
rect 119233 72559 119246 72581
rect 118806 72525 118874 72559
rect 118930 72525 118998 72559
rect 119054 72525 119122 72559
rect 119178 72525 119246 72559
rect 119302 72559 119319 72581
rect 119426 72559 119461 72581
rect 119550 72559 119603 72581
rect 119302 72525 119370 72559
rect 119426 72525 119494 72559
rect 119550 72525 119618 72559
rect 119674 72525 119728 72581
rect 117828 72473 119728 72525
rect 117828 72457 117899 72473
rect 117955 72457 118041 72473
rect 118097 72457 118183 72473
rect 118239 72457 118325 72473
rect 118381 72457 118467 72473
rect 118523 72457 118609 72473
rect 118665 72457 118751 72473
rect 118807 72457 118893 72473
rect 118949 72457 119035 72473
rect 119091 72457 119177 72473
rect 119233 72457 119319 72473
rect 119375 72457 119461 72473
rect 119517 72457 119603 72473
rect 119659 72457 119728 72473
rect 117828 72401 117882 72457
rect 117955 72417 118006 72457
rect 118097 72417 118130 72457
rect 118239 72417 118254 72457
rect 117938 72401 118006 72417
rect 118062 72401 118130 72417
rect 118186 72401 118254 72417
rect 118310 72417 118325 72457
rect 118434 72417 118467 72457
rect 118558 72417 118609 72457
rect 118310 72401 118378 72417
rect 118434 72401 118502 72417
rect 118558 72401 118626 72417
rect 118682 72401 118750 72457
rect 118807 72417 118874 72457
rect 118949 72417 118998 72457
rect 119091 72417 119122 72457
rect 119233 72417 119246 72457
rect 118806 72401 118874 72417
rect 118930 72401 118998 72417
rect 119054 72401 119122 72417
rect 119178 72401 119246 72417
rect 119302 72417 119319 72457
rect 119426 72417 119461 72457
rect 119550 72417 119603 72457
rect 119302 72401 119370 72417
rect 119426 72401 119494 72417
rect 119550 72401 119618 72417
rect 119674 72401 119728 72457
rect 117828 72333 119728 72401
rect 117828 72277 117882 72333
rect 117938 72331 118006 72333
rect 118062 72331 118130 72333
rect 118186 72331 118254 72333
rect 117955 72277 118006 72331
rect 118097 72277 118130 72331
rect 118239 72277 118254 72331
rect 118310 72331 118378 72333
rect 118434 72331 118502 72333
rect 118558 72331 118626 72333
rect 118310 72277 118325 72331
rect 118434 72277 118467 72331
rect 118558 72277 118609 72331
rect 118682 72277 118750 72333
rect 118806 72331 118874 72333
rect 118930 72331 118998 72333
rect 119054 72331 119122 72333
rect 119178 72331 119246 72333
rect 118807 72277 118874 72331
rect 118949 72277 118998 72331
rect 119091 72277 119122 72331
rect 119233 72277 119246 72331
rect 119302 72331 119370 72333
rect 119426 72331 119494 72333
rect 119550 72331 119618 72333
rect 119302 72277 119319 72331
rect 119426 72277 119461 72331
rect 119550 72277 119603 72331
rect 119674 72277 119728 72333
rect 117828 72275 117899 72277
rect 117955 72275 118041 72277
rect 118097 72275 118183 72277
rect 118239 72275 118325 72277
rect 118381 72275 118467 72277
rect 118523 72275 118609 72277
rect 118665 72275 118751 72277
rect 118807 72275 118893 72277
rect 118949 72275 119035 72277
rect 119091 72275 119177 72277
rect 119233 72275 119319 72277
rect 119375 72275 119461 72277
rect 119517 72275 119603 72277
rect 119659 72275 119728 72277
rect 117828 72209 119728 72275
rect 117828 72153 117882 72209
rect 117938 72189 118006 72209
rect 118062 72189 118130 72209
rect 118186 72189 118254 72209
rect 117955 72153 118006 72189
rect 118097 72153 118130 72189
rect 118239 72153 118254 72189
rect 118310 72189 118378 72209
rect 118434 72189 118502 72209
rect 118558 72189 118626 72209
rect 118310 72153 118325 72189
rect 118434 72153 118467 72189
rect 118558 72153 118609 72189
rect 118682 72153 118750 72209
rect 118806 72189 118874 72209
rect 118930 72189 118998 72209
rect 119054 72189 119122 72209
rect 119178 72189 119246 72209
rect 118807 72153 118874 72189
rect 118949 72153 118998 72189
rect 119091 72153 119122 72189
rect 119233 72153 119246 72189
rect 119302 72189 119370 72209
rect 119426 72189 119494 72209
rect 119550 72189 119618 72209
rect 119302 72153 119319 72189
rect 119426 72153 119461 72189
rect 119550 72153 119603 72189
rect 119674 72153 119728 72209
rect 117828 72133 117899 72153
rect 117955 72133 118041 72153
rect 118097 72133 118183 72153
rect 118239 72133 118325 72153
rect 118381 72133 118467 72153
rect 118523 72133 118609 72153
rect 118665 72133 118751 72153
rect 118807 72133 118893 72153
rect 118949 72133 119035 72153
rect 119091 72133 119177 72153
rect 119233 72133 119319 72153
rect 119375 72133 119461 72153
rect 119517 72133 119603 72153
rect 119659 72133 119728 72153
rect 117828 72088 119728 72133
rect 270272 74035 272172 74088
rect 270272 73979 270343 74035
rect 270399 73979 270485 74035
rect 270541 73979 270627 74035
rect 270683 73979 270769 74035
rect 270825 73979 270911 74035
rect 270967 73979 271053 74035
rect 271109 73979 271195 74035
rect 271251 73979 271337 74035
rect 271393 73979 271479 74035
rect 271535 73979 271621 74035
rect 271677 73979 271763 74035
rect 271819 73979 271905 74035
rect 271961 73979 272047 74035
rect 272103 73979 272172 74035
rect 270272 73945 272172 73979
rect 270272 73889 270326 73945
rect 270382 73893 270450 73945
rect 270506 73893 270574 73945
rect 270630 73893 270698 73945
rect 270399 73889 270450 73893
rect 270541 73889 270574 73893
rect 270683 73889 270698 73893
rect 270754 73893 270822 73945
rect 270878 73893 270946 73945
rect 271002 73893 271070 73945
rect 270754 73889 270769 73893
rect 270878 73889 270911 73893
rect 271002 73889 271053 73893
rect 271126 73889 271194 73945
rect 271250 73893 271318 73945
rect 271374 73893 271442 73945
rect 271498 73893 271566 73945
rect 271622 73893 271690 73945
rect 271251 73889 271318 73893
rect 271393 73889 271442 73893
rect 271535 73889 271566 73893
rect 271677 73889 271690 73893
rect 271746 73893 271814 73945
rect 271870 73893 271938 73945
rect 271994 73893 272062 73945
rect 271746 73889 271763 73893
rect 271870 73889 271905 73893
rect 271994 73889 272047 73893
rect 272118 73889 272172 73945
rect 270272 73837 270343 73889
rect 270399 73837 270485 73889
rect 270541 73837 270627 73889
rect 270683 73837 270769 73889
rect 270825 73837 270911 73889
rect 270967 73837 271053 73889
rect 271109 73837 271195 73889
rect 271251 73837 271337 73889
rect 271393 73837 271479 73889
rect 271535 73837 271621 73889
rect 271677 73837 271763 73889
rect 271819 73837 271905 73889
rect 271961 73837 272047 73889
rect 272103 73837 272172 73889
rect 270272 73821 272172 73837
rect 270272 73765 270326 73821
rect 270382 73765 270450 73821
rect 270506 73765 270574 73821
rect 270630 73765 270698 73821
rect 270754 73765 270822 73821
rect 270878 73765 270946 73821
rect 271002 73765 271070 73821
rect 271126 73765 271194 73821
rect 271250 73765 271318 73821
rect 271374 73765 271442 73821
rect 271498 73765 271566 73821
rect 271622 73765 271690 73821
rect 271746 73765 271814 73821
rect 271870 73765 271938 73821
rect 271994 73765 272062 73821
rect 272118 73765 272172 73821
rect 270272 73751 272172 73765
rect 270272 73697 270343 73751
rect 270399 73697 270485 73751
rect 270541 73697 270627 73751
rect 270683 73697 270769 73751
rect 270825 73697 270911 73751
rect 270967 73697 271053 73751
rect 271109 73697 271195 73751
rect 271251 73697 271337 73751
rect 271393 73697 271479 73751
rect 271535 73697 271621 73751
rect 271677 73697 271763 73751
rect 271819 73697 271905 73751
rect 271961 73697 272047 73751
rect 272103 73697 272172 73751
rect 270272 73641 270326 73697
rect 270399 73695 270450 73697
rect 270541 73695 270574 73697
rect 270683 73695 270698 73697
rect 270382 73641 270450 73695
rect 270506 73641 270574 73695
rect 270630 73641 270698 73695
rect 270754 73695 270769 73697
rect 270878 73695 270911 73697
rect 271002 73695 271053 73697
rect 270754 73641 270822 73695
rect 270878 73641 270946 73695
rect 271002 73641 271070 73695
rect 271126 73641 271194 73697
rect 271251 73695 271318 73697
rect 271393 73695 271442 73697
rect 271535 73695 271566 73697
rect 271677 73695 271690 73697
rect 271250 73641 271318 73695
rect 271374 73641 271442 73695
rect 271498 73641 271566 73695
rect 271622 73641 271690 73695
rect 271746 73695 271763 73697
rect 271870 73695 271905 73697
rect 271994 73695 272047 73697
rect 271746 73641 271814 73695
rect 271870 73641 271938 73695
rect 271994 73641 272062 73695
rect 272118 73641 272172 73697
rect 270272 73609 272172 73641
rect 270272 73573 270343 73609
rect 270399 73573 270485 73609
rect 270541 73573 270627 73609
rect 270683 73573 270769 73609
rect 270825 73573 270911 73609
rect 270967 73573 271053 73609
rect 271109 73573 271195 73609
rect 271251 73573 271337 73609
rect 271393 73573 271479 73609
rect 271535 73573 271621 73609
rect 271677 73573 271763 73609
rect 271819 73573 271905 73609
rect 271961 73573 272047 73609
rect 272103 73573 272172 73609
rect 270272 73517 270326 73573
rect 270399 73553 270450 73573
rect 270541 73553 270574 73573
rect 270683 73553 270698 73573
rect 270382 73517 270450 73553
rect 270506 73517 270574 73553
rect 270630 73517 270698 73553
rect 270754 73553 270769 73573
rect 270878 73553 270911 73573
rect 271002 73553 271053 73573
rect 270754 73517 270822 73553
rect 270878 73517 270946 73553
rect 271002 73517 271070 73553
rect 271126 73517 271194 73573
rect 271251 73553 271318 73573
rect 271393 73553 271442 73573
rect 271535 73553 271566 73573
rect 271677 73553 271690 73573
rect 271250 73517 271318 73553
rect 271374 73517 271442 73553
rect 271498 73517 271566 73553
rect 271622 73517 271690 73553
rect 271746 73553 271763 73573
rect 271870 73553 271905 73573
rect 271994 73553 272047 73573
rect 271746 73517 271814 73553
rect 271870 73517 271938 73553
rect 271994 73517 272062 73553
rect 272118 73517 272172 73573
rect 270272 73467 272172 73517
rect 270272 73449 270343 73467
rect 270399 73449 270485 73467
rect 270541 73449 270627 73467
rect 270683 73449 270769 73467
rect 270825 73449 270911 73467
rect 270967 73449 271053 73467
rect 271109 73449 271195 73467
rect 271251 73449 271337 73467
rect 271393 73449 271479 73467
rect 271535 73449 271621 73467
rect 271677 73449 271763 73467
rect 271819 73449 271905 73467
rect 271961 73449 272047 73467
rect 272103 73449 272172 73467
rect 270272 73393 270326 73449
rect 270399 73411 270450 73449
rect 270541 73411 270574 73449
rect 270683 73411 270698 73449
rect 270382 73393 270450 73411
rect 270506 73393 270574 73411
rect 270630 73393 270698 73411
rect 270754 73411 270769 73449
rect 270878 73411 270911 73449
rect 271002 73411 271053 73449
rect 270754 73393 270822 73411
rect 270878 73393 270946 73411
rect 271002 73393 271070 73411
rect 271126 73393 271194 73449
rect 271251 73411 271318 73449
rect 271393 73411 271442 73449
rect 271535 73411 271566 73449
rect 271677 73411 271690 73449
rect 271250 73393 271318 73411
rect 271374 73393 271442 73411
rect 271498 73393 271566 73411
rect 271622 73393 271690 73411
rect 271746 73411 271763 73449
rect 271870 73411 271905 73449
rect 271994 73411 272047 73449
rect 271746 73393 271814 73411
rect 271870 73393 271938 73411
rect 271994 73393 272062 73411
rect 272118 73393 272172 73449
rect 270272 73325 272172 73393
rect 270272 73269 270326 73325
rect 270399 73269 270450 73325
rect 270541 73269 270574 73325
rect 270683 73269 270698 73325
rect 270754 73269 270769 73325
rect 270878 73269 270911 73325
rect 271002 73269 271053 73325
rect 271126 73269 271194 73325
rect 271251 73269 271318 73325
rect 271393 73269 271442 73325
rect 271535 73269 271566 73325
rect 271677 73269 271690 73325
rect 271746 73269 271763 73325
rect 271870 73269 271905 73325
rect 271994 73269 272047 73325
rect 272118 73269 272172 73325
rect 270272 73201 272172 73269
rect 270272 73145 270326 73201
rect 270382 73183 270450 73201
rect 270506 73183 270574 73201
rect 270630 73183 270698 73201
rect 270399 73145 270450 73183
rect 270541 73145 270574 73183
rect 270683 73145 270698 73183
rect 270754 73183 270822 73201
rect 270878 73183 270946 73201
rect 271002 73183 271070 73201
rect 270754 73145 270769 73183
rect 270878 73145 270911 73183
rect 271002 73145 271053 73183
rect 271126 73145 271194 73201
rect 271250 73183 271318 73201
rect 271374 73183 271442 73201
rect 271498 73183 271566 73201
rect 271622 73183 271690 73201
rect 271251 73145 271318 73183
rect 271393 73145 271442 73183
rect 271535 73145 271566 73183
rect 271677 73145 271690 73183
rect 271746 73183 271814 73201
rect 271870 73183 271938 73201
rect 271994 73183 272062 73201
rect 271746 73145 271763 73183
rect 271870 73145 271905 73183
rect 271994 73145 272047 73183
rect 272118 73145 272172 73201
rect 270272 73127 270343 73145
rect 270399 73127 270485 73145
rect 270541 73127 270627 73145
rect 270683 73127 270769 73145
rect 270825 73127 270911 73145
rect 270967 73127 271053 73145
rect 271109 73127 271195 73145
rect 271251 73127 271337 73145
rect 271393 73127 271479 73145
rect 271535 73127 271621 73145
rect 271677 73127 271763 73145
rect 271819 73127 271905 73145
rect 271961 73127 272047 73145
rect 272103 73127 272172 73145
rect 270272 73077 272172 73127
rect 270272 73021 270326 73077
rect 270382 73041 270450 73077
rect 270506 73041 270574 73077
rect 270630 73041 270698 73077
rect 270399 73021 270450 73041
rect 270541 73021 270574 73041
rect 270683 73021 270698 73041
rect 270754 73041 270822 73077
rect 270878 73041 270946 73077
rect 271002 73041 271070 73077
rect 270754 73021 270769 73041
rect 270878 73021 270911 73041
rect 271002 73021 271053 73041
rect 271126 73021 271194 73077
rect 271250 73041 271318 73077
rect 271374 73041 271442 73077
rect 271498 73041 271566 73077
rect 271622 73041 271690 73077
rect 271251 73021 271318 73041
rect 271393 73021 271442 73041
rect 271535 73021 271566 73041
rect 271677 73021 271690 73041
rect 271746 73041 271814 73077
rect 271870 73041 271938 73077
rect 271994 73041 272062 73077
rect 271746 73021 271763 73041
rect 271870 73021 271905 73041
rect 271994 73021 272047 73041
rect 272118 73021 272172 73077
rect 270272 72985 270343 73021
rect 270399 72985 270485 73021
rect 270541 72985 270627 73021
rect 270683 72985 270769 73021
rect 270825 72985 270911 73021
rect 270967 72985 271053 73021
rect 271109 72985 271195 73021
rect 271251 72985 271337 73021
rect 271393 72985 271479 73021
rect 271535 72985 271621 73021
rect 271677 72985 271763 73021
rect 271819 72985 271905 73021
rect 271961 72985 272047 73021
rect 272103 72985 272172 73021
rect 270272 72953 272172 72985
rect 270272 72897 270326 72953
rect 270382 72899 270450 72953
rect 270506 72899 270574 72953
rect 270630 72899 270698 72953
rect 270399 72897 270450 72899
rect 270541 72897 270574 72899
rect 270683 72897 270698 72899
rect 270754 72899 270822 72953
rect 270878 72899 270946 72953
rect 271002 72899 271070 72953
rect 270754 72897 270769 72899
rect 270878 72897 270911 72899
rect 271002 72897 271053 72899
rect 271126 72897 271194 72953
rect 271250 72899 271318 72953
rect 271374 72899 271442 72953
rect 271498 72899 271566 72953
rect 271622 72899 271690 72953
rect 271251 72897 271318 72899
rect 271393 72897 271442 72899
rect 271535 72897 271566 72899
rect 271677 72897 271690 72899
rect 271746 72899 271814 72953
rect 271870 72899 271938 72953
rect 271994 72899 272062 72953
rect 271746 72897 271763 72899
rect 271870 72897 271905 72899
rect 271994 72897 272047 72899
rect 272118 72897 272172 72953
rect 270272 72843 270343 72897
rect 270399 72843 270485 72897
rect 270541 72843 270627 72897
rect 270683 72843 270769 72897
rect 270825 72843 270911 72897
rect 270967 72843 271053 72897
rect 271109 72843 271195 72897
rect 271251 72843 271337 72897
rect 271393 72843 271479 72897
rect 271535 72843 271621 72897
rect 271677 72843 271763 72897
rect 271819 72843 271905 72897
rect 271961 72843 272047 72897
rect 272103 72843 272172 72897
rect 270272 72829 272172 72843
rect 270272 72773 270326 72829
rect 270382 72773 270450 72829
rect 270506 72773 270574 72829
rect 270630 72773 270698 72829
rect 270754 72773 270822 72829
rect 270878 72773 270946 72829
rect 271002 72773 271070 72829
rect 271126 72773 271194 72829
rect 271250 72773 271318 72829
rect 271374 72773 271442 72829
rect 271498 72773 271566 72829
rect 271622 72773 271690 72829
rect 271746 72773 271814 72829
rect 271870 72773 271938 72829
rect 271994 72773 272062 72829
rect 272118 72773 272172 72829
rect 270272 72757 272172 72773
rect 270272 72705 270343 72757
rect 270399 72705 270485 72757
rect 270541 72705 270627 72757
rect 270683 72705 270769 72757
rect 270825 72705 270911 72757
rect 270967 72705 271053 72757
rect 271109 72705 271195 72757
rect 271251 72705 271337 72757
rect 271393 72705 271479 72757
rect 271535 72705 271621 72757
rect 271677 72705 271763 72757
rect 271819 72705 271905 72757
rect 271961 72705 272047 72757
rect 272103 72705 272172 72757
rect 270272 72649 270326 72705
rect 270399 72701 270450 72705
rect 270541 72701 270574 72705
rect 270683 72701 270698 72705
rect 270382 72649 270450 72701
rect 270506 72649 270574 72701
rect 270630 72649 270698 72701
rect 270754 72701 270769 72705
rect 270878 72701 270911 72705
rect 271002 72701 271053 72705
rect 270754 72649 270822 72701
rect 270878 72649 270946 72701
rect 271002 72649 271070 72701
rect 271126 72649 271194 72705
rect 271251 72701 271318 72705
rect 271393 72701 271442 72705
rect 271535 72701 271566 72705
rect 271677 72701 271690 72705
rect 271250 72649 271318 72701
rect 271374 72649 271442 72701
rect 271498 72649 271566 72701
rect 271622 72649 271690 72701
rect 271746 72701 271763 72705
rect 271870 72701 271905 72705
rect 271994 72701 272047 72705
rect 271746 72649 271814 72701
rect 271870 72649 271938 72701
rect 271994 72649 272062 72701
rect 272118 72649 272172 72705
rect 270272 72615 272172 72649
rect 270272 72581 270343 72615
rect 270399 72581 270485 72615
rect 270541 72581 270627 72615
rect 270683 72581 270769 72615
rect 270825 72581 270911 72615
rect 270967 72581 271053 72615
rect 271109 72581 271195 72615
rect 271251 72581 271337 72615
rect 271393 72581 271479 72615
rect 271535 72581 271621 72615
rect 271677 72581 271763 72615
rect 271819 72581 271905 72615
rect 271961 72581 272047 72615
rect 272103 72581 272172 72615
rect 270272 72525 270326 72581
rect 270399 72559 270450 72581
rect 270541 72559 270574 72581
rect 270683 72559 270698 72581
rect 270382 72525 270450 72559
rect 270506 72525 270574 72559
rect 270630 72525 270698 72559
rect 270754 72559 270769 72581
rect 270878 72559 270911 72581
rect 271002 72559 271053 72581
rect 270754 72525 270822 72559
rect 270878 72525 270946 72559
rect 271002 72525 271070 72559
rect 271126 72525 271194 72581
rect 271251 72559 271318 72581
rect 271393 72559 271442 72581
rect 271535 72559 271566 72581
rect 271677 72559 271690 72581
rect 271250 72525 271318 72559
rect 271374 72525 271442 72559
rect 271498 72525 271566 72559
rect 271622 72525 271690 72559
rect 271746 72559 271763 72581
rect 271870 72559 271905 72581
rect 271994 72559 272047 72581
rect 271746 72525 271814 72559
rect 271870 72525 271938 72559
rect 271994 72525 272062 72559
rect 272118 72525 272172 72581
rect 270272 72473 272172 72525
rect 270272 72457 270343 72473
rect 270399 72457 270485 72473
rect 270541 72457 270627 72473
rect 270683 72457 270769 72473
rect 270825 72457 270911 72473
rect 270967 72457 271053 72473
rect 271109 72457 271195 72473
rect 271251 72457 271337 72473
rect 271393 72457 271479 72473
rect 271535 72457 271621 72473
rect 271677 72457 271763 72473
rect 271819 72457 271905 72473
rect 271961 72457 272047 72473
rect 272103 72457 272172 72473
rect 270272 72401 270326 72457
rect 270399 72417 270450 72457
rect 270541 72417 270574 72457
rect 270683 72417 270698 72457
rect 270382 72401 270450 72417
rect 270506 72401 270574 72417
rect 270630 72401 270698 72417
rect 270754 72417 270769 72457
rect 270878 72417 270911 72457
rect 271002 72417 271053 72457
rect 270754 72401 270822 72417
rect 270878 72401 270946 72417
rect 271002 72401 271070 72417
rect 271126 72401 271194 72457
rect 271251 72417 271318 72457
rect 271393 72417 271442 72457
rect 271535 72417 271566 72457
rect 271677 72417 271690 72457
rect 271250 72401 271318 72417
rect 271374 72401 271442 72417
rect 271498 72401 271566 72417
rect 271622 72401 271690 72417
rect 271746 72417 271763 72457
rect 271870 72417 271905 72457
rect 271994 72417 272047 72457
rect 271746 72401 271814 72417
rect 271870 72401 271938 72417
rect 271994 72401 272062 72417
rect 272118 72401 272172 72457
rect 270272 72333 272172 72401
rect 270272 72277 270326 72333
rect 270382 72331 270450 72333
rect 270506 72331 270574 72333
rect 270630 72331 270698 72333
rect 270399 72277 270450 72331
rect 270541 72277 270574 72331
rect 270683 72277 270698 72331
rect 270754 72331 270822 72333
rect 270878 72331 270946 72333
rect 271002 72331 271070 72333
rect 270754 72277 270769 72331
rect 270878 72277 270911 72331
rect 271002 72277 271053 72331
rect 271126 72277 271194 72333
rect 271250 72331 271318 72333
rect 271374 72331 271442 72333
rect 271498 72331 271566 72333
rect 271622 72331 271690 72333
rect 271251 72277 271318 72331
rect 271393 72277 271442 72331
rect 271535 72277 271566 72331
rect 271677 72277 271690 72331
rect 271746 72331 271814 72333
rect 271870 72331 271938 72333
rect 271994 72331 272062 72333
rect 271746 72277 271763 72331
rect 271870 72277 271905 72331
rect 271994 72277 272047 72331
rect 272118 72277 272172 72333
rect 270272 72275 270343 72277
rect 270399 72275 270485 72277
rect 270541 72275 270627 72277
rect 270683 72275 270769 72277
rect 270825 72275 270911 72277
rect 270967 72275 271053 72277
rect 271109 72275 271195 72277
rect 271251 72275 271337 72277
rect 271393 72275 271479 72277
rect 271535 72275 271621 72277
rect 271677 72275 271763 72277
rect 271819 72275 271905 72277
rect 271961 72275 272047 72277
rect 272103 72275 272172 72277
rect 270272 72209 272172 72275
rect 270272 72153 270326 72209
rect 270382 72189 270450 72209
rect 270506 72189 270574 72209
rect 270630 72189 270698 72209
rect 270399 72153 270450 72189
rect 270541 72153 270574 72189
rect 270683 72153 270698 72189
rect 270754 72189 270822 72209
rect 270878 72189 270946 72209
rect 271002 72189 271070 72209
rect 270754 72153 270769 72189
rect 270878 72153 270911 72189
rect 271002 72153 271053 72189
rect 271126 72153 271194 72209
rect 271250 72189 271318 72209
rect 271374 72189 271442 72209
rect 271498 72189 271566 72209
rect 271622 72189 271690 72209
rect 271251 72153 271318 72189
rect 271393 72153 271442 72189
rect 271535 72153 271566 72189
rect 271677 72153 271690 72189
rect 271746 72189 271814 72209
rect 271870 72189 271938 72209
rect 271994 72189 272062 72209
rect 271746 72153 271763 72189
rect 271870 72153 271905 72189
rect 271994 72153 272047 72189
rect 272118 72153 272172 72209
rect 270272 72133 270343 72153
rect 270399 72133 270485 72153
rect 270541 72133 270627 72153
rect 270683 72133 270769 72153
rect 270825 72133 270911 72153
rect 270967 72133 271053 72153
rect 271109 72133 271195 72153
rect 271251 72133 271337 72153
rect 271393 72133 271479 72153
rect 271535 72133 271621 72153
rect 271677 72133 271763 72153
rect 271819 72133 271905 72153
rect 271961 72133 272047 72153
rect 272103 72133 272172 72153
rect 270272 72088 272172 72133
rect 272752 74035 274802 74088
rect 272752 73979 272823 74035
rect 272879 73979 272965 74035
rect 273021 73979 273107 74035
rect 273163 73979 273249 74035
rect 273305 73979 273391 74035
rect 273447 73979 273533 74035
rect 273589 73979 273675 74035
rect 273731 73979 273817 74035
rect 273873 73979 273959 74035
rect 274015 73979 274101 74035
rect 274157 73979 274243 74035
rect 274299 73979 274385 74035
rect 274441 73979 274527 74035
rect 274583 73979 274669 74035
rect 274725 73979 274802 74035
rect 272752 73945 274802 73979
rect 272752 73889 272806 73945
rect 272862 73893 272930 73945
rect 272986 73893 273054 73945
rect 273110 73893 273178 73945
rect 272879 73889 272930 73893
rect 273021 73889 273054 73893
rect 273163 73889 273178 73893
rect 273234 73893 273302 73945
rect 273358 73893 273426 73945
rect 273482 73893 273550 73945
rect 273234 73889 273249 73893
rect 273358 73889 273391 73893
rect 273482 73889 273533 73893
rect 273606 73889 273674 73945
rect 273730 73893 273798 73945
rect 273854 73893 273922 73945
rect 273978 73893 274046 73945
rect 274102 73893 274170 73945
rect 273731 73889 273798 73893
rect 273873 73889 273922 73893
rect 274015 73889 274046 73893
rect 274157 73889 274170 73893
rect 274226 73893 274294 73945
rect 274350 73893 274418 73945
rect 274474 73893 274542 73945
rect 274226 73889 274243 73893
rect 274350 73889 274385 73893
rect 274474 73889 274527 73893
rect 274598 73889 274666 73945
rect 274722 73893 274802 73945
rect 272752 73837 272823 73889
rect 272879 73837 272965 73889
rect 273021 73837 273107 73889
rect 273163 73837 273249 73889
rect 273305 73837 273391 73889
rect 273447 73837 273533 73889
rect 273589 73837 273675 73889
rect 273731 73837 273817 73889
rect 273873 73837 273959 73889
rect 274015 73837 274101 73889
rect 274157 73837 274243 73889
rect 274299 73837 274385 73889
rect 274441 73837 274527 73889
rect 274583 73837 274669 73889
rect 274725 73837 274802 73893
rect 272752 73821 274802 73837
rect 272752 73765 272806 73821
rect 272862 73765 272930 73821
rect 272986 73765 273054 73821
rect 273110 73765 273178 73821
rect 273234 73765 273302 73821
rect 273358 73765 273426 73821
rect 273482 73765 273550 73821
rect 273606 73765 273674 73821
rect 273730 73765 273798 73821
rect 273854 73765 273922 73821
rect 273978 73765 274046 73821
rect 274102 73765 274170 73821
rect 274226 73765 274294 73821
rect 274350 73765 274418 73821
rect 274474 73765 274542 73821
rect 274598 73765 274666 73821
rect 274722 73765 274802 73821
rect 272752 73751 274802 73765
rect 272752 73697 272823 73751
rect 272879 73697 272965 73751
rect 273021 73697 273107 73751
rect 273163 73697 273249 73751
rect 273305 73697 273391 73751
rect 273447 73697 273533 73751
rect 273589 73697 273675 73751
rect 273731 73697 273817 73751
rect 273873 73697 273959 73751
rect 274015 73697 274101 73751
rect 274157 73697 274243 73751
rect 274299 73697 274385 73751
rect 274441 73697 274527 73751
rect 274583 73697 274669 73751
rect 272752 73641 272806 73697
rect 272879 73695 272930 73697
rect 273021 73695 273054 73697
rect 273163 73695 273178 73697
rect 272862 73641 272930 73695
rect 272986 73641 273054 73695
rect 273110 73641 273178 73695
rect 273234 73695 273249 73697
rect 273358 73695 273391 73697
rect 273482 73695 273533 73697
rect 273234 73641 273302 73695
rect 273358 73641 273426 73695
rect 273482 73641 273550 73695
rect 273606 73641 273674 73697
rect 273731 73695 273798 73697
rect 273873 73695 273922 73697
rect 274015 73695 274046 73697
rect 274157 73695 274170 73697
rect 273730 73641 273798 73695
rect 273854 73641 273922 73695
rect 273978 73641 274046 73695
rect 274102 73641 274170 73695
rect 274226 73695 274243 73697
rect 274350 73695 274385 73697
rect 274474 73695 274527 73697
rect 274226 73641 274294 73695
rect 274350 73641 274418 73695
rect 274474 73641 274542 73695
rect 274598 73641 274666 73697
rect 274725 73695 274802 73751
rect 274722 73641 274802 73695
rect 272752 73609 274802 73641
rect 272752 73573 272823 73609
rect 272879 73573 272965 73609
rect 273021 73573 273107 73609
rect 273163 73573 273249 73609
rect 273305 73573 273391 73609
rect 273447 73573 273533 73609
rect 273589 73573 273675 73609
rect 273731 73573 273817 73609
rect 273873 73573 273959 73609
rect 274015 73573 274101 73609
rect 274157 73573 274243 73609
rect 274299 73573 274385 73609
rect 274441 73573 274527 73609
rect 274583 73573 274669 73609
rect 272752 73517 272806 73573
rect 272879 73553 272930 73573
rect 273021 73553 273054 73573
rect 273163 73553 273178 73573
rect 272862 73517 272930 73553
rect 272986 73517 273054 73553
rect 273110 73517 273178 73553
rect 273234 73553 273249 73573
rect 273358 73553 273391 73573
rect 273482 73553 273533 73573
rect 273234 73517 273302 73553
rect 273358 73517 273426 73553
rect 273482 73517 273550 73553
rect 273606 73517 273674 73573
rect 273731 73553 273798 73573
rect 273873 73553 273922 73573
rect 274015 73553 274046 73573
rect 274157 73553 274170 73573
rect 273730 73517 273798 73553
rect 273854 73517 273922 73553
rect 273978 73517 274046 73553
rect 274102 73517 274170 73553
rect 274226 73553 274243 73573
rect 274350 73553 274385 73573
rect 274474 73553 274527 73573
rect 274226 73517 274294 73553
rect 274350 73517 274418 73553
rect 274474 73517 274542 73553
rect 274598 73517 274666 73573
rect 274725 73553 274802 73609
rect 274722 73517 274802 73553
rect 272752 73467 274802 73517
rect 272752 73449 272823 73467
rect 272879 73449 272965 73467
rect 273021 73449 273107 73467
rect 273163 73449 273249 73467
rect 273305 73449 273391 73467
rect 273447 73449 273533 73467
rect 273589 73449 273675 73467
rect 273731 73449 273817 73467
rect 273873 73449 273959 73467
rect 274015 73449 274101 73467
rect 274157 73449 274243 73467
rect 274299 73449 274385 73467
rect 274441 73449 274527 73467
rect 274583 73449 274669 73467
rect 272752 73393 272806 73449
rect 272879 73411 272930 73449
rect 273021 73411 273054 73449
rect 273163 73411 273178 73449
rect 272862 73393 272930 73411
rect 272986 73393 273054 73411
rect 273110 73393 273178 73411
rect 273234 73411 273249 73449
rect 273358 73411 273391 73449
rect 273482 73411 273533 73449
rect 273234 73393 273302 73411
rect 273358 73393 273426 73411
rect 273482 73393 273550 73411
rect 273606 73393 273674 73449
rect 273731 73411 273798 73449
rect 273873 73411 273922 73449
rect 274015 73411 274046 73449
rect 274157 73411 274170 73449
rect 273730 73393 273798 73411
rect 273854 73393 273922 73411
rect 273978 73393 274046 73411
rect 274102 73393 274170 73411
rect 274226 73411 274243 73449
rect 274350 73411 274385 73449
rect 274474 73411 274527 73449
rect 274226 73393 274294 73411
rect 274350 73393 274418 73411
rect 274474 73393 274542 73411
rect 274598 73393 274666 73449
rect 274725 73411 274802 73467
rect 274722 73393 274802 73411
rect 272752 73325 274802 73393
rect 272752 73269 272806 73325
rect 272879 73269 272930 73325
rect 273021 73269 273054 73325
rect 273163 73269 273178 73325
rect 273234 73269 273249 73325
rect 273358 73269 273391 73325
rect 273482 73269 273533 73325
rect 273606 73269 273674 73325
rect 273731 73269 273798 73325
rect 273873 73269 273922 73325
rect 274015 73269 274046 73325
rect 274157 73269 274170 73325
rect 274226 73269 274243 73325
rect 274350 73269 274385 73325
rect 274474 73269 274527 73325
rect 274598 73269 274666 73325
rect 274725 73269 274802 73325
rect 272752 73201 274802 73269
rect 272752 73145 272806 73201
rect 272862 73183 272930 73201
rect 272986 73183 273054 73201
rect 273110 73183 273178 73201
rect 272879 73145 272930 73183
rect 273021 73145 273054 73183
rect 273163 73145 273178 73183
rect 273234 73183 273302 73201
rect 273358 73183 273426 73201
rect 273482 73183 273550 73201
rect 273234 73145 273249 73183
rect 273358 73145 273391 73183
rect 273482 73145 273533 73183
rect 273606 73145 273674 73201
rect 273730 73183 273798 73201
rect 273854 73183 273922 73201
rect 273978 73183 274046 73201
rect 274102 73183 274170 73201
rect 273731 73145 273798 73183
rect 273873 73145 273922 73183
rect 274015 73145 274046 73183
rect 274157 73145 274170 73183
rect 274226 73183 274294 73201
rect 274350 73183 274418 73201
rect 274474 73183 274542 73201
rect 274226 73145 274243 73183
rect 274350 73145 274385 73183
rect 274474 73145 274527 73183
rect 274598 73145 274666 73201
rect 274722 73183 274802 73201
rect 272752 73127 272823 73145
rect 272879 73127 272965 73145
rect 273021 73127 273107 73145
rect 273163 73127 273249 73145
rect 273305 73127 273391 73145
rect 273447 73127 273533 73145
rect 273589 73127 273675 73145
rect 273731 73127 273817 73145
rect 273873 73127 273959 73145
rect 274015 73127 274101 73145
rect 274157 73127 274243 73145
rect 274299 73127 274385 73145
rect 274441 73127 274527 73145
rect 274583 73127 274669 73145
rect 274725 73127 274802 73183
rect 272752 73077 274802 73127
rect 272752 73021 272806 73077
rect 272862 73041 272930 73077
rect 272986 73041 273054 73077
rect 273110 73041 273178 73077
rect 272879 73021 272930 73041
rect 273021 73021 273054 73041
rect 273163 73021 273178 73041
rect 273234 73041 273302 73077
rect 273358 73041 273426 73077
rect 273482 73041 273550 73077
rect 273234 73021 273249 73041
rect 273358 73021 273391 73041
rect 273482 73021 273533 73041
rect 273606 73021 273674 73077
rect 273730 73041 273798 73077
rect 273854 73041 273922 73077
rect 273978 73041 274046 73077
rect 274102 73041 274170 73077
rect 273731 73021 273798 73041
rect 273873 73021 273922 73041
rect 274015 73021 274046 73041
rect 274157 73021 274170 73041
rect 274226 73041 274294 73077
rect 274350 73041 274418 73077
rect 274474 73041 274542 73077
rect 274226 73021 274243 73041
rect 274350 73021 274385 73041
rect 274474 73021 274527 73041
rect 274598 73021 274666 73077
rect 274722 73041 274802 73077
rect 272752 72985 272823 73021
rect 272879 72985 272965 73021
rect 273021 72985 273107 73021
rect 273163 72985 273249 73021
rect 273305 72985 273391 73021
rect 273447 72985 273533 73021
rect 273589 72985 273675 73021
rect 273731 72985 273817 73021
rect 273873 72985 273959 73021
rect 274015 72985 274101 73021
rect 274157 72985 274243 73021
rect 274299 72985 274385 73021
rect 274441 72985 274527 73021
rect 274583 72985 274669 73021
rect 274725 72985 274802 73041
rect 272752 72953 274802 72985
rect 272752 72897 272806 72953
rect 272862 72899 272930 72953
rect 272986 72899 273054 72953
rect 273110 72899 273178 72953
rect 272879 72897 272930 72899
rect 273021 72897 273054 72899
rect 273163 72897 273178 72899
rect 273234 72899 273302 72953
rect 273358 72899 273426 72953
rect 273482 72899 273550 72953
rect 273234 72897 273249 72899
rect 273358 72897 273391 72899
rect 273482 72897 273533 72899
rect 273606 72897 273674 72953
rect 273730 72899 273798 72953
rect 273854 72899 273922 72953
rect 273978 72899 274046 72953
rect 274102 72899 274170 72953
rect 273731 72897 273798 72899
rect 273873 72897 273922 72899
rect 274015 72897 274046 72899
rect 274157 72897 274170 72899
rect 274226 72899 274294 72953
rect 274350 72899 274418 72953
rect 274474 72899 274542 72953
rect 274226 72897 274243 72899
rect 274350 72897 274385 72899
rect 274474 72897 274527 72899
rect 274598 72897 274666 72953
rect 274722 72899 274802 72953
rect 272752 72843 272823 72897
rect 272879 72843 272965 72897
rect 273021 72843 273107 72897
rect 273163 72843 273249 72897
rect 273305 72843 273391 72897
rect 273447 72843 273533 72897
rect 273589 72843 273675 72897
rect 273731 72843 273817 72897
rect 273873 72843 273959 72897
rect 274015 72843 274101 72897
rect 274157 72843 274243 72897
rect 274299 72843 274385 72897
rect 274441 72843 274527 72897
rect 274583 72843 274669 72897
rect 274725 72843 274802 72899
rect 272752 72829 274802 72843
rect 272752 72773 272806 72829
rect 272862 72773 272930 72829
rect 272986 72773 273054 72829
rect 273110 72773 273178 72829
rect 273234 72773 273302 72829
rect 273358 72773 273426 72829
rect 273482 72773 273550 72829
rect 273606 72773 273674 72829
rect 273730 72773 273798 72829
rect 273854 72773 273922 72829
rect 273978 72773 274046 72829
rect 274102 72773 274170 72829
rect 274226 72773 274294 72829
rect 274350 72773 274418 72829
rect 274474 72773 274542 72829
rect 274598 72773 274666 72829
rect 274722 72773 274802 72829
rect 272752 72757 274802 72773
rect 272752 72705 272823 72757
rect 272879 72705 272965 72757
rect 273021 72705 273107 72757
rect 273163 72705 273249 72757
rect 273305 72705 273391 72757
rect 273447 72705 273533 72757
rect 273589 72705 273675 72757
rect 273731 72705 273817 72757
rect 273873 72705 273959 72757
rect 274015 72705 274101 72757
rect 274157 72705 274243 72757
rect 274299 72705 274385 72757
rect 274441 72705 274527 72757
rect 274583 72705 274669 72757
rect 272752 72649 272806 72705
rect 272879 72701 272930 72705
rect 273021 72701 273054 72705
rect 273163 72701 273178 72705
rect 272862 72649 272930 72701
rect 272986 72649 273054 72701
rect 273110 72649 273178 72701
rect 273234 72701 273249 72705
rect 273358 72701 273391 72705
rect 273482 72701 273533 72705
rect 273234 72649 273302 72701
rect 273358 72649 273426 72701
rect 273482 72649 273550 72701
rect 273606 72649 273674 72705
rect 273731 72701 273798 72705
rect 273873 72701 273922 72705
rect 274015 72701 274046 72705
rect 274157 72701 274170 72705
rect 273730 72649 273798 72701
rect 273854 72649 273922 72701
rect 273978 72649 274046 72701
rect 274102 72649 274170 72701
rect 274226 72701 274243 72705
rect 274350 72701 274385 72705
rect 274474 72701 274527 72705
rect 274226 72649 274294 72701
rect 274350 72649 274418 72701
rect 274474 72649 274542 72701
rect 274598 72649 274666 72705
rect 274725 72701 274802 72757
rect 274722 72649 274802 72701
rect 272752 72615 274802 72649
rect 272752 72581 272823 72615
rect 272879 72581 272965 72615
rect 273021 72581 273107 72615
rect 273163 72581 273249 72615
rect 273305 72581 273391 72615
rect 273447 72581 273533 72615
rect 273589 72581 273675 72615
rect 273731 72581 273817 72615
rect 273873 72581 273959 72615
rect 274015 72581 274101 72615
rect 274157 72581 274243 72615
rect 274299 72581 274385 72615
rect 274441 72581 274527 72615
rect 274583 72581 274669 72615
rect 272752 72525 272806 72581
rect 272879 72559 272930 72581
rect 273021 72559 273054 72581
rect 273163 72559 273178 72581
rect 272862 72525 272930 72559
rect 272986 72525 273054 72559
rect 273110 72525 273178 72559
rect 273234 72559 273249 72581
rect 273358 72559 273391 72581
rect 273482 72559 273533 72581
rect 273234 72525 273302 72559
rect 273358 72525 273426 72559
rect 273482 72525 273550 72559
rect 273606 72525 273674 72581
rect 273731 72559 273798 72581
rect 273873 72559 273922 72581
rect 274015 72559 274046 72581
rect 274157 72559 274170 72581
rect 273730 72525 273798 72559
rect 273854 72525 273922 72559
rect 273978 72525 274046 72559
rect 274102 72525 274170 72559
rect 274226 72559 274243 72581
rect 274350 72559 274385 72581
rect 274474 72559 274527 72581
rect 274226 72525 274294 72559
rect 274350 72525 274418 72559
rect 274474 72525 274542 72559
rect 274598 72525 274666 72581
rect 274725 72559 274802 72615
rect 274722 72525 274802 72559
rect 272752 72473 274802 72525
rect 272752 72457 272823 72473
rect 272879 72457 272965 72473
rect 273021 72457 273107 72473
rect 273163 72457 273249 72473
rect 273305 72457 273391 72473
rect 273447 72457 273533 72473
rect 273589 72457 273675 72473
rect 273731 72457 273817 72473
rect 273873 72457 273959 72473
rect 274015 72457 274101 72473
rect 274157 72457 274243 72473
rect 274299 72457 274385 72473
rect 274441 72457 274527 72473
rect 274583 72457 274669 72473
rect 272752 72401 272806 72457
rect 272879 72417 272930 72457
rect 273021 72417 273054 72457
rect 273163 72417 273178 72457
rect 272862 72401 272930 72417
rect 272986 72401 273054 72417
rect 273110 72401 273178 72417
rect 273234 72417 273249 72457
rect 273358 72417 273391 72457
rect 273482 72417 273533 72457
rect 273234 72401 273302 72417
rect 273358 72401 273426 72417
rect 273482 72401 273550 72417
rect 273606 72401 273674 72457
rect 273731 72417 273798 72457
rect 273873 72417 273922 72457
rect 274015 72417 274046 72457
rect 274157 72417 274170 72457
rect 273730 72401 273798 72417
rect 273854 72401 273922 72417
rect 273978 72401 274046 72417
rect 274102 72401 274170 72417
rect 274226 72417 274243 72457
rect 274350 72417 274385 72457
rect 274474 72417 274527 72457
rect 274226 72401 274294 72417
rect 274350 72401 274418 72417
rect 274474 72401 274542 72417
rect 274598 72401 274666 72457
rect 274725 72417 274802 72473
rect 274722 72401 274802 72417
rect 272752 72333 274802 72401
rect 272752 72277 272806 72333
rect 272862 72331 272930 72333
rect 272986 72331 273054 72333
rect 273110 72331 273178 72333
rect 272879 72277 272930 72331
rect 273021 72277 273054 72331
rect 273163 72277 273178 72331
rect 273234 72331 273302 72333
rect 273358 72331 273426 72333
rect 273482 72331 273550 72333
rect 273234 72277 273249 72331
rect 273358 72277 273391 72331
rect 273482 72277 273533 72331
rect 273606 72277 273674 72333
rect 273730 72331 273798 72333
rect 273854 72331 273922 72333
rect 273978 72331 274046 72333
rect 274102 72331 274170 72333
rect 273731 72277 273798 72331
rect 273873 72277 273922 72331
rect 274015 72277 274046 72331
rect 274157 72277 274170 72331
rect 274226 72331 274294 72333
rect 274350 72331 274418 72333
rect 274474 72331 274542 72333
rect 274226 72277 274243 72331
rect 274350 72277 274385 72331
rect 274474 72277 274527 72331
rect 274598 72277 274666 72333
rect 274722 72331 274802 72333
rect 272752 72275 272823 72277
rect 272879 72275 272965 72277
rect 273021 72275 273107 72277
rect 273163 72275 273249 72277
rect 273305 72275 273391 72277
rect 273447 72275 273533 72277
rect 273589 72275 273675 72277
rect 273731 72275 273817 72277
rect 273873 72275 273959 72277
rect 274015 72275 274101 72277
rect 274157 72275 274243 72277
rect 274299 72275 274385 72277
rect 274441 72275 274527 72277
rect 274583 72275 274669 72277
rect 274725 72275 274802 72331
rect 272752 72209 274802 72275
rect 272752 72153 272806 72209
rect 272862 72189 272930 72209
rect 272986 72189 273054 72209
rect 273110 72189 273178 72209
rect 272879 72153 272930 72189
rect 273021 72153 273054 72189
rect 273163 72153 273178 72189
rect 273234 72189 273302 72209
rect 273358 72189 273426 72209
rect 273482 72189 273550 72209
rect 273234 72153 273249 72189
rect 273358 72153 273391 72189
rect 273482 72153 273533 72189
rect 273606 72153 273674 72209
rect 273730 72189 273798 72209
rect 273854 72189 273922 72209
rect 273978 72189 274046 72209
rect 274102 72189 274170 72209
rect 273731 72153 273798 72189
rect 273873 72153 273922 72189
rect 274015 72153 274046 72189
rect 274157 72153 274170 72189
rect 274226 72189 274294 72209
rect 274350 72189 274418 72209
rect 274474 72189 274542 72209
rect 274226 72153 274243 72189
rect 274350 72153 274385 72189
rect 274474 72153 274527 72189
rect 274598 72153 274666 72209
rect 274722 72189 274802 72209
rect 272752 72133 272823 72153
rect 272879 72133 272965 72153
rect 273021 72133 273107 72153
rect 273163 72133 273249 72153
rect 273305 72133 273391 72153
rect 273447 72133 273533 72153
rect 273589 72133 273675 72153
rect 273731 72133 273817 72153
rect 273873 72133 273959 72153
rect 274015 72133 274101 72153
rect 274157 72133 274243 72153
rect 274299 72133 274385 72153
rect 274441 72133 274527 72153
rect 274583 72133 274669 72153
rect 274725 72133 274802 72189
rect 272752 72088 274802 72133
rect 275122 74035 277172 74088
rect 275122 73979 275193 74035
rect 275249 73979 275335 74035
rect 275391 73979 275477 74035
rect 275533 73979 275619 74035
rect 275675 73979 275761 74035
rect 275817 73979 275903 74035
rect 275959 73979 276045 74035
rect 276101 73979 276187 74035
rect 276243 73979 276329 74035
rect 276385 73979 276471 74035
rect 276527 73979 276613 74035
rect 276669 73979 276755 74035
rect 276811 73979 276897 74035
rect 276953 73979 277039 74035
rect 277095 73979 277172 74035
rect 275122 73945 277172 73979
rect 275122 73889 275176 73945
rect 275232 73893 275300 73945
rect 275356 73893 275424 73945
rect 275480 73893 275548 73945
rect 275249 73889 275300 73893
rect 275391 73889 275424 73893
rect 275533 73889 275548 73893
rect 275604 73893 275672 73945
rect 275728 73893 275796 73945
rect 275852 73893 275920 73945
rect 275604 73889 275619 73893
rect 275728 73889 275761 73893
rect 275852 73889 275903 73893
rect 275976 73889 276044 73945
rect 276100 73893 276168 73945
rect 276224 73893 276292 73945
rect 276348 73893 276416 73945
rect 276472 73893 276540 73945
rect 276101 73889 276168 73893
rect 276243 73889 276292 73893
rect 276385 73889 276416 73893
rect 276527 73889 276540 73893
rect 276596 73893 276664 73945
rect 276720 73893 276788 73945
rect 276844 73893 276912 73945
rect 276596 73889 276613 73893
rect 276720 73889 276755 73893
rect 276844 73889 276897 73893
rect 276968 73889 277036 73945
rect 277092 73893 277172 73945
rect 275122 73837 275193 73889
rect 275249 73837 275335 73889
rect 275391 73837 275477 73889
rect 275533 73837 275619 73889
rect 275675 73837 275761 73889
rect 275817 73837 275903 73889
rect 275959 73837 276045 73889
rect 276101 73837 276187 73889
rect 276243 73837 276329 73889
rect 276385 73837 276471 73889
rect 276527 73837 276613 73889
rect 276669 73837 276755 73889
rect 276811 73837 276897 73889
rect 276953 73837 277039 73889
rect 277095 73837 277172 73893
rect 275122 73821 277172 73837
rect 275122 73765 275176 73821
rect 275232 73765 275300 73821
rect 275356 73765 275424 73821
rect 275480 73765 275548 73821
rect 275604 73765 275672 73821
rect 275728 73765 275796 73821
rect 275852 73765 275920 73821
rect 275976 73765 276044 73821
rect 276100 73765 276168 73821
rect 276224 73765 276292 73821
rect 276348 73765 276416 73821
rect 276472 73765 276540 73821
rect 276596 73765 276664 73821
rect 276720 73765 276788 73821
rect 276844 73765 276912 73821
rect 276968 73765 277036 73821
rect 277092 73765 277172 73821
rect 275122 73751 277172 73765
rect 275122 73697 275193 73751
rect 275249 73697 275335 73751
rect 275391 73697 275477 73751
rect 275533 73697 275619 73751
rect 275675 73697 275761 73751
rect 275817 73697 275903 73751
rect 275959 73697 276045 73751
rect 276101 73697 276187 73751
rect 276243 73697 276329 73751
rect 276385 73697 276471 73751
rect 276527 73697 276613 73751
rect 276669 73697 276755 73751
rect 276811 73697 276897 73751
rect 276953 73697 277039 73751
rect 275122 73641 275176 73697
rect 275249 73695 275300 73697
rect 275391 73695 275424 73697
rect 275533 73695 275548 73697
rect 275232 73641 275300 73695
rect 275356 73641 275424 73695
rect 275480 73641 275548 73695
rect 275604 73695 275619 73697
rect 275728 73695 275761 73697
rect 275852 73695 275903 73697
rect 275604 73641 275672 73695
rect 275728 73641 275796 73695
rect 275852 73641 275920 73695
rect 275976 73641 276044 73697
rect 276101 73695 276168 73697
rect 276243 73695 276292 73697
rect 276385 73695 276416 73697
rect 276527 73695 276540 73697
rect 276100 73641 276168 73695
rect 276224 73641 276292 73695
rect 276348 73641 276416 73695
rect 276472 73641 276540 73695
rect 276596 73695 276613 73697
rect 276720 73695 276755 73697
rect 276844 73695 276897 73697
rect 276596 73641 276664 73695
rect 276720 73641 276788 73695
rect 276844 73641 276912 73695
rect 276968 73641 277036 73697
rect 277095 73695 277172 73751
rect 277092 73641 277172 73695
rect 275122 73609 277172 73641
rect 275122 73573 275193 73609
rect 275249 73573 275335 73609
rect 275391 73573 275477 73609
rect 275533 73573 275619 73609
rect 275675 73573 275761 73609
rect 275817 73573 275903 73609
rect 275959 73573 276045 73609
rect 276101 73573 276187 73609
rect 276243 73573 276329 73609
rect 276385 73573 276471 73609
rect 276527 73573 276613 73609
rect 276669 73573 276755 73609
rect 276811 73573 276897 73609
rect 276953 73573 277039 73609
rect 275122 73517 275176 73573
rect 275249 73553 275300 73573
rect 275391 73553 275424 73573
rect 275533 73553 275548 73573
rect 275232 73517 275300 73553
rect 275356 73517 275424 73553
rect 275480 73517 275548 73553
rect 275604 73553 275619 73573
rect 275728 73553 275761 73573
rect 275852 73553 275903 73573
rect 275604 73517 275672 73553
rect 275728 73517 275796 73553
rect 275852 73517 275920 73553
rect 275976 73517 276044 73573
rect 276101 73553 276168 73573
rect 276243 73553 276292 73573
rect 276385 73553 276416 73573
rect 276527 73553 276540 73573
rect 276100 73517 276168 73553
rect 276224 73517 276292 73553
rect 276348 73517 276416 73553
rect 276472 73517 276540 73553
rect 276596 73553 276613 73573
rect 276720 73553 276755 73573
rect 276844 73553 276897 73573
rect 276596 73517 276664 73553
rect 276720 73517 276788 73553
rect 276844 73517 276912 73553
rect 276968 73517 277036 73573
rect 277095 73553 277172 73609
rect 277092 73517 277172 73553
rect 275122 73467 277172 73517
rect 275122 73449 275193 73467
rect 275249 73449 275335 73467
rect 275391 73449 275477 73467
rect 275533 73449 275619 73467
rect 275675 73449 275761 73467
rect 275817 73449 275903 73467
rect 275959 73449 276045 73467
rect 276101 73449 276187 73467
rect 276243 73449 276329 73467
rect 276385 73449 276471 73467
rect 276527 73449 276613 73467
rect 276669 73449 276755 73467
rect 276811 73449 276897 73467
rect 276953 73449 277039 73467
rect 275122 73393 275176 73449
rect 275249 73411 275300 73449
rect 275391 73411 275424 73449
rect 275533 73411 275548 73449
rect 275232 73393 275300 73411
rect 275356 73393 275424 73411
rect 275480 73393 275548 73411
rect 275604 73411 275619 73449
rect 275728 73411 275761 73449
rect 275852 73411 275903 73449
rect 275604 73393 275672 73411
rect 275728 73393 275796 73411
rect 275852 73393 275920 73411
rect 275976 73393 276044 73449
rect 276101 73411 276168 73449
rect 276243 73411 276292 73449
rect 276385 73411 276416 73449
rect 276527 73411 276540 73449
rect 276100 73393 276168 73411
rect 276224 73393 276292 73411
rect 276348 73393 276416 73411
rect 276472 73393 276540 73411
rect 276596 73411 276613 73449
rect 276720 73411 276755 73449
rect 276844 73411 276897 73449
rect 276596 73393 276664 73411
rect 276720 73393 276788 73411
rect 276844 73393 276912 73411
rect 276968 73393 277036 73449
rect 277095 73411 277172 73467
rect 277092 73393 277172 73411
rect 275122 73325 277172 73393
rect 275122 73269 275176 73325
rect 275249 73269 275300 73325
rect 275391 73269 275424 73325
rect 275533 73269 275548 73325
rect 275604 73269 275619 73325
rect 275728 73269 275761 73325
rect 275852 73269 275903 73325
rect 275976 73269 276044 73325
rect 276101 73269 276168 73325
rect 276243 73269 276292 73325
rect 276385 73269 276416 73325
rect 276527 73269 276540 73325
rect 276596 73269 276613 73325
rect 276720 73269 276755 73325
rect 276844 73269 276897 73325
rect 276968 73269 277036 73325
rect 277095 73269 277172 73325
rect 275122 73201 277172 73269
rect 275122 73145 275176 73201
rect 275232 73183 275300 73201
rect 275356 73183 275424 73201
rect 275480 73183 275548 73201
rect 275249 73145 275300 73183
rect 275391 73145 275424 73183
rect 275533 73145 275548 73183
rect 275604 73183 275672 73201
rect 275728 73183 275796 73201
rect 275852 73183 275920 73201
rect 275604 73145 275619 73183
rect 275728 73145 275761 73183
rect 275852 73145 275903 73183
rect 275976 73145 276044 73201
rect 276100 73183 276168 73201
rect 276224 73183 276292 73201
rect 276348 73183 276416 73201
rect 276472 73183 276540 73201
rect 276101 73145 276168 73183
rect 276243 73145 276292 73183
rect 276385 73145 276416 73183
rect 276527 73145 276540 73183
rect 276596 73183 276664 73201
rect 276720 73183 276788 73201
rect 276844 73183 276912 73201
rect 276596 73145 276613 73183
rect 276720 73145 276755 73183
rect 276844 73145 276897 73183
rect 276968 73145 277036 73201
rect 277092 73183 277172 73201
rect 275122 73127 275193 73145
rect 275249 73127 275335 73145
rect 275391 73127 275477 73145
rect 275533 73127 275619 73145
rect 275675 73127 275761 73145
rect 275817 73127 275903 73145
rect 275959 73127 276045 73145
rect 276101 73127 276187 73145
rect 276243 73127 276329 73145
rect 276385 73127 276471 73145
rect 276527 73127 276613 73145
rect 276669 73127 276755 73145
rect 276811 73127 276897 73145
rect 276953 73127 277039 73145
rect 277095 73127 277172 73183
rect 275122 73077 277172 73127
rect 275122 73021 275176 73077
rect 275232 73041 275300 73077
rect 275356 73041 275424 73077
rect 275480 73041 275548 73077
rect 275249 73021 275300 73041
rect 275391 73021 275424 73041
rect 275533 73021 275548 73041
rect 275604 73041 275672 73077
rect 275728 73041 275796 73077
rect 275852 73041 275920 73077
rect 275604 73021 275619 73041
rect 275728 73021 275761 73041
rect 275852 73021 275903 73041
rect 275976 73021 276044 73077
rect 276100 73041 276168 73077
rect 276224 73041 276292 73077
rect 276348 73041 276416 73077
rect 276472 73041 276540 73077
rect 276101 73021 276168 73041
rect 276243 73021 276292 73041
rect 276385 73021 276416 73041
rect 276527 73021 276540 73041
rect 276596 73041 276664 73077
rect 276720 73041 276788 73077
rect 276844 73041 276912 73077
rect 276596 73021 276613 73041
rect 276720 73021 276755 73041
rect 276844 73021 276897 73041
rect 276968 73021 277036 73077
rect 277092 73041 277172 73077
rect 275122 72985 275193 73021
rect 275249 72985 275335 73021
rect 275391 72985 275477 73021
rect 275533 72985 275619 73021
rect 275675 72985 275761 73021
rect 275817 72985 275903 73021
rect 275959 72985 276045 73021
rect 276101 72985 276187 73021
rect 276243 72985 276329 73021
rect 276385 72985 276471 73021
rect 276527 72985 276613 73021
rect 276669 72985 276755 73021
rect 276811 72985 276897 73021
rect 276953 72985 277039 73021
rect 277095 72985 277172 73041
rect 275122 72953 277172 72985
rect 275122 72897 275176 72953
rect 275232 72899 275300 72953
rect 275356 72899 275424 72953
rect 275480 72899 275548 72953
rect 275249 72897 275300 72899
rect 275391 72897 275424 72899
rect 275533 72897 275548 72899
rect 275604 72899 275672 72953
rect 275728 72899 275796 72953
rect 275852 72899 275920 72953
rect 275604 72897 275619 72899
rect 275728 72897 275761 72899
rect 275852 72897 275903 72899
rect 275976 72897 276044 72953
rect 276100 72899 276168 72953
rect 276224 72899 276292 72953
rect 276348 72899 276416 72953
rect 276472 72899 276540 72953
rect 276101 72897 276168 72899
rect 276243 72897 276292 72899
rect 276385 72897 276416 72899
rect 276527 72897 276540 72899
rect 276596 72899 276664 72953
rect 276720 72899 276788 72953
rect 276844 72899 276912 72953
rect 276596 72897 276613 72899
rect 276720 72897 276755 72899
rect 276844 72897 276897 72899
rect 276968 72897 277036 72953
rect 277092 72899 277172 72953
rect 275122 72843 275193 72897
rect 275249 72843 275335 72897
rect 275391 72843 275477 72897
rect 275533 72843 275619 72897
rect 275675 72843 275761 72897
rect 275817 72843 275903 72897
rect 275959 72843 276045 72897
rect 276101 72843 276187 72897
rect 276243 72843 276329 72897
rect 276385 72843 276471 72897
rect 276527 72843 276613 72897
rect 276669 72843 276755 72897
rect 276811 72843 276897 72897
rect 276953 72843 277039 72897
rect 277095 72843 277172 72899
rect 275122 72829 277172 72843
rect 275122 72773 275176 72829
rect 275232 72773 275300 72829
rect 275356 72773 275424 72829
rect 275480 72773 275548 72829
rect 275604 72773 275672 72829
rect 275728 72773 275796 72829
rect 275852 72773 275920 72829
rect 275976 72773 276044 72829
rect 276100 72773 276168 72829
rect 276224 72773 276292 72829
rect 276348 72773 276416 72829
rect 276472 72773 276540 72829
rect 276596 72773 276664 72829
rect 276720 72773 276788 72829
rect 276844 72773 276912 72829
rect 276968 72773 277036 72829
rect 277092 72773 277172 72829
rect 275122 72757 277172 72773
rect 275122 72705 275193 72757
rect 275249 72705 275335 72757
rect 275391 72705 275477 72757
rect 275533 72705 275619 72757
rect 275675 72705 275761 72757
rect 275817 72705 275903 72757
rect 275959 72705 276045 72757
rect 276101 72705 276187 72757
rect 276243 72705 276329 72757
rect 276385 72705 276471 72757
rect 276527 72705 276613 72757
rect 276669 72705 276755 72757
rect 276811 72705 276897 72757
rect 276953 72705 277039 72757
rect 275122 72649 275176 72705
rect 275249 72701 275300 72705
rect 275391 72701 275424 72705
rect 275533 72701 275548 72705
rect 275232 72649 275300 72701
rect 275356 72649 275424 72701
rect 275480 72649 275548 72701
rect 275604 72701 275619 72705
rect 275728 72701 275761 72705
rect 275852 72701 275903 72705
rect 275604 72649 275672 72701
rect 275728 72649 275796 72701
rect 275852 72649 275920 72701
rect 275976 72649 276044 72705
rect 276101 72701 276168 72705
rect 276243 72701 276292 72705
rect 276385 72701 276416 72705
rect 276527 72701 276540 72705
rect 276100 72649 276168 72701
rect 276224 72649 276292 72701
rect 276348 72649 276416 72701
rect 276472 72649 276540 72701
rect 276596 72701 276613 72705
rect 276720 72701 276755 72705
rect 276844 72701 276897 72705
rect 276596 72649 276664 72701
rect 276720 72649 276788 72701
rect 276844 72649 276912 72701
rect 276968 72649 277036 72705
rect 277095 72701 277172 72757
rect 277092 72649 277172 72701
rect 275122 72615 277172 72649
rect 275122 72581 275193 72615
rect 275249 72581 275335 72615
rect 275391 72581 275477 72615
rect 275533 72581 275619 72615
rect 275675 72581 275761 72615
rect 275817 72581 275903 72615
rect 275959 72581 276045 72615
rect 276101 72581 276187 72615
rect 276243 72581 276329 72615
rect 276385 72581 276471 72615
rect 276527 72581 276613 72615
rect 276669 72581 276755 72615
rect 276811 72581 276897 72615
rect 276953 72581 277039 72615
rect 275122 72525 275176 72581
rect 275249 72559 275300 72581
rect 275391 72559 275424 72581
rect 275533 72559 275548 72581
rect 275232 72525 275300 72559
rect 275356 72525 275424 72559
rect 275480 72525 275548 72559
rect 275604 72559 275619 72581
rect 275728 72559 275761 72581
rect 275852 72559 275903 72581
rect 275604 72525 275672 72559
rect 275728 72525 275796 72559
rect 275852 72525 275920 72559
rect 275976 72525 276044 72581
rect 276101 72559 276168 72581
rect 276243 72559 276292 72581
rect 276385 72559 276416 72581
rect 276527 72559 276540 72581
rect 276100 72525 276168 72559
rect 276224 72525 276292 72559
rect 276348 72525 276416 72559
rect 276472 72525 276540 72559
rect 276596 72559 276613 72581
rect 276720 72559 276755 72581
rect 276844 72559 276897 72581
rect 276596 72525 276664 72559
rect 276720 72525 276788 72559
rect 276844 72525 276912 72559
rect 276968 72525 277036 72581
rect 277095 72559 277172 72615
rect 277092 72525 277172 72559
rect 275122 72473 277172 72525
rect 275122 72457 275193 72473
rect 275249 72457 275335 72473
rect 275391 72457 275477 72473
rect 275533 72457 275619 72473
rect 275675 72457 275761 72473
rect 275817 72457 275903 72473
rect 275959 72457 276045 72473
rect 276101 72457 276187 72473
rect 276243 72457 276329 72473
rect 276385 72457 276471 72473
rect 276527 72457 276613 72473
rect 276669 72457 276755 72473
rect 276811 72457 276897 72473
rect 276953 72457 277039 72473
rect 275122 72401 275176 72457
rect 275249 72417 275300 72457
rect 275391 72417 275424 72457
rect 275533 72417 275548 72457
rect 275232 72401 275300 72417
rect 275356 72401 275424 72417
rect 275480 72401 275548 72417
rect 275604 72417 275619 72457
rect 275728 72417 275761 72457
rect 275852 72417 275903 72457
rect 275604 72401 275672 72417
rect 275728 72401 275796 72417
rect 275852 72401 275920 72417
rect 275976 72401 276044 72457
rect 276101 72417 276168 72457
rect 276243 72417 276292 72457
rect 276385 72417 276416 72457
rect 276527 72417 276540 72457
rect 276100 72401 276168 72417
rect 276224 72401 276292 72417
rect 276348 72401 276416 72417
rect 276472 72401 276540 72417
rect 276596 72417 276613 72457
rect 276720 72417 276755 72457
rect 276844 72417 276897 72457
rect 276596 72401 276664 72417
rect 276720 72401 276788 72417
rect 276844 72401 276912 72417
rect 276968 72401 277036 72457
rect 277095 72417 277172 72473
rect 277092 72401 277172 72417
rect 275122 72333 277172 72401
rect 275122 72277 275176 72333
rect 275232 72331 275300 72333
rect 275356 72331 275424 72333
rect 275480 72331 275548 72333
rect 275249 72277 275300 72331
rect 275391 72277 275424 72331
rect 275533 72277 275548 72331
rect 275604 72331 275672 72333
rect 275728 72331 275796 72333
rect 275852 72331 275920 72333
rect 275604 72277 275619 72331
rect 275728 72277 275761 72331
rect 275852 72277 275903 72331
rect 275976 72277 276044 72333
rect 276100 72331 276168 72333
rect 276224 72331 276292 72333
rect 276348 72331 276416 72333
rect 276472 72331 276540 72333
rect 276101 72277 276168 72331
rect 276243 72277 276292 72331
rect 276385 72277 276416 72331
rect 276527 72277 276540 72331
rect 276596 72331 276664 72333
rect 276720 72331 276788 72333
rect 276844 72331 276912 72333
rect 276596 72277 276613 72331
rect 276720 72277 276755 72331
rect 276844 72277 276897 72331
rect 276968 72277 277036 72333
rect 277092 72331 277172 72333
rect 275122 72275 275193 72277
rect 275249 72275 275335 72277
rect 275391 72275 275477 72277
rect 275533 72275 275619 72277
rect 275675 72275 275761 72277
rect 275817 72275 275903 72277
rect 275959 72275 276045 72277
rect 276101 72275 276187 72277
rect 276243 72275 276329 72277
rect 276385 72275 276471 72277
rect 276527 72275 276613 72277
rect 276669 72275 276755 72277
rect 276811 72275 276897 72277
rect 276953 72275 277039 72277
rect 277095 72275 277172 72331
rect 275122 72209 277172 72275
rect 275122 72153 275176 72209
rect 275232 72189 275300 72209
rect 275356 72189 275424 72209
rect 275480 72189 275548 72209
rect 275249 72153 275300 72189
rect 275391 72153 275424 72189
rect 275533 72153 275548 72189
rect 275604 72189 275672 72209
rect 275728 72189 275796 72209
rect 275852 72189 275920 72209
rect 275604 72153 275619 72189
rect 275728 72153 275761 72189
rect 275852 72153 275903 72189
rect 275976 72153 276044 72209
rect 276100 72189 276168 72209
rect 276224 72189 276292 72209
rect 276348 72189 276416 72209
rect 276472 72189 276540 72209
rect 276101 72153 276168 72189
rect 276243 72153 276292 72189
rect 276385 72153 276416 72189
rect 276527 72153 276540 72189
rect 276596 72189 276664 72209
rect 276720 72189 276788 72209
rect 276844 72189 276912 72209
rect 276596 72153 276613 72189
rect 276720 72153 276755 72189
rect 276844 72153 276897 72189
rect 276968 72153 277036 72209
rect 277092 72189 277172 72209
rect 275122 72133 275193 72153
rect 275249 72133 275335 72153
rect 275391 72133 275477 72153
rect 275533 72133 275619 72153
rect 275675 72133 275761 72153
rect 275817 72133 275903 72153
rect 275959 72133 276045 72153
rect 276101 72133 276187 72153
rect 276243 72133 276329 72153
rect 276385 72133 276471 72153
rect 276527 72133 276613 72153
rect 276669 72133 276755 72153
rect 276811 72133 276897 72153
rect 276953 72133 277039 72153
rect 277095 72133 277172 72189
rect 275122 72088 277172 72133
rect 277828 74035 279878 74088
rect 277828 73979 277899 74035
rect 277955 73979 278041 74035
rect 278097 73979 278183 74035
rect 278239 73979 278325 74035
rect 278381 73979 278467 74035
rect 278523 73979 278609 74035
rect 278665 73979 278751 74035
rect 278807 73979 278893 74035
rect 278949 73979 279035 74035
rect 279091 73979 279177 74035
rect 279233 73979 279319 74035
rect 279375 73979 279461 74035
rect 279517 73979 279603 74035
rect 279659 73979 279745 74035
rect 279801 73979 279878 74035
rect 277828 73945 279878 73979
rect 277828 73889 277882 73945
rect 277938 73893 278006 73945
rect 278062 73893 278130 73945
rect 278186 73893 278254 73945
rect 277955 73889 278006 73893
rect 278097 73889 278130 73893
rect 278239 73889 278254 73893
rect 278310 73893 278378 73945
rect 278434 73893 278502 73945
rect 278558 73893 278626 73945
rect 278310 73889 278325 73893
rect 278434 73889 278467 73893
rect 278558 73889 278609 73893
rect 278682 73889 278750 73945
rect 278806 73893 278874 73945
rect 278930 73893 278998 73945
rect 279054 73893 279122 73945
rect 279178 73893 279246 73945
rect 278807 73889 278874 73893
rect 278949 73889 278998 73893
rect 279091 73889 279122 73893
rect 279233 73889 279246 73893
rect 279302 73893 279370 73945
rect 279426 73893 279494 73945
rect 279550 73893 279618 73945
rect 279302 73889 279319 73893
rect 279426 73889 279461 73893
rect 279550 73889 279603 73893
rect 279674 73889 279742 73945
rect 279798 73893 279878 73945
rect 277828 73837 277899 73889
rect 277955 73837 278041 73889
rect 278097 73837 278183 73889
rect 278239 73837 278325 73889
rect 278381 73837 278467 73889
rect 278523 73837 278609 73889
rect 278665 73837 278751 73889
rect 278807 73837 278893 73889
rect 278949 73837 279035 73889
rect 279091 73837 279177 73889
rect 279233 73837 279319 73889
rect 279375 73837 279461 73889
rect 279517 73837 279603 73889
rect 279659 73837 279745 73889
rect 279801 73837 279878 73893
rect 277828 73821 279878 73837
rect 277828 73765 277882 73821
rect 277938 73765 278006 73821
rect 278062 73765 278130 73821
rect 278186 73765 278254 73821
rect 278310 73765 278378 73821
rect 278434 73765 278502 73821
rect 278558 73765 278626 73821
rect 278682 73765 278750 73821
rect 278806 73765 278874 73821
rect 278930 73765 278998 73821
rect 279054 73765 279122 73821
rect 279178 73765 279246 73821
rect 279302 73765 279370 73821
rect 279426 73765 279494 73821
rect 279550 73765 279618 73821
rect 279674 73765 279742 73821
rect 279798 73765 279878 73821
rect 277828 73751 279878 73765
rect 277828 73697 277899 73751
rect 277955 73697 278041 73751
rect 278097 73697 278183 73751
rect 278239 73697 278325 73751
rect 278381 73697 278467 73751
rect 278523 73697 278609 73751
rect 278665 73697 278751 73751
rect 278807 73697 278893 73751
rect 278949 73697 279035 73751
rect 279091 73697 279177 73751
rect 279233 73697 279319 73751
rect 279375 73697 279461 73751
rect 279517 73697 279603 73751
rect 279659 73697 279745 73751
rect 277828 73641 277882 73697
rect 277955 73695 278006 73697
rect 278097 73695 278130 73697
rect 278239 73695 278254 73697
rect 277938 73641 278006 73695
rect 278062 73641 278130 73695
rect 278186 73641 278254 73695
rect 278310 73695 278325 73697
rect 278434 73695 278467 73697
rect 278558 73695 278609 73697
rect 278310 73641 278378 73695
rect 278434 73641 278502 73695
rect 278558 73641 278626 73695
rect 278682 73641 278750 73697
rect 278807 73695 278874 73697
rect 278949 73695 278998 73697
rect 279091 73695 279122 73697
rect 279233 73695 279246 73697
rect 278806 73641 278874 73695
rect 278930 73641 278998 73695
rect 279054 73641 279122 73695
rect 279178 73641 279246 73695
rect 279302 73695 279319 73697
rect 279426 73695 279461 73697
rect 279550 73695 279603 73697
rect 279302 73641 279370 73695
rect 279426 73641 279494 73695
rect 279550 73641 279618 73695
rect 279674 73641 279742 73697
rect 279801 73695 279878 73751
rect 279798 73641 279878 73695
rect 277828 73609 279878 73641
rect 277828 73573 277899 73609
rect 277955 73573 278041 73609
rect 278097 73573 278183 73609
rect 278239 73573 278325 73609
rect 278381 73573 278467 73609
rect 278523 73573 278609 73609
rect 278665 73573 278751 73609
rect 278807 73573 278893 73609
rect 278949 73573 279035 73609
rect 279091 73573 279177 73609
rect 279233 73573 279319 73609
rect 279375 73573 279461 73609
rect 279517 73573 279603 73609
rect 279659 73573 279745 73609
rect 277828 73517 277882 73573
rect 277955 73553 278006 73573
rect 278097 73553 278130 73573
rect 278239 73553 278254 73573
rect 277938 73517 278006 73553
rect 278062 73517 278130 73553
rect 278186 73517 278254 73553
rect 278310 73553 278325 73573
rect 278434 73553 278467 73573
rect 278558 73553 278609 73573
rect 278310 73517 278378 73553
rect 278434 73517 278502 73553
rect 278558 73517 278626 73553
rect 278682 73517 278750 73573
rect 278807 73553 278874 73573
rect 278949 73553 278998 73573
rect 279091 73553 279122 73573
rect 279233 73553 279246 73573
rect 278806 73517 278874 73553
rect 278930 73517 278998 73553
rect 279054 73517 279122 73553
rect 279178 73517 279246 73553
rect 279302 73553 279319 73573
rect 279426 73553 279461 73573
rect 279550 73553 279603 73573
rect 279302 73517 279370 73553
rect 279426 73517 279494 73553
rect 279550 73517 279618 73553
rect 279674 73517 279742 73573
rect 279801 73553 279878 73609
rect 279798 73517 279878 73553
rect 277828 73467 279878 73517
rect 277828 73449 277899 73467
rect 277955 73449 278041 73467
rect 278097 73449 278183 73467
rect 278239 73449 278325 73467
rect 278381 73449 278467 73467
rect 278523 73449 278609 73467
rect 278665 73449 278751 73467
rect 278807 73449 278893 73467
rect 278949 73449 279035 73467
rect 279091 73449 279177 73467
rect 279233 73449 279319 73467
rect 279375 73449 279461 73467
rect 279517 73449 279603 73467
rect 279659 73449 279745 73467
rect 277828 73393 277882 73449
rect 277955 73411 278006 73449
rect 278097 73411 278130 73449
rect 278239 73411 278254 73449
rect 277938 73393 278006 73411
rect 278062 73393 278130 73411
rect 278186 73393 278254 73411
rect 278310 73411 278325 73449
rect 278434 73411 278467 73449
rect 278558 73411 278609 73449
rect 278310 73393 278378 73411
rect 278434 73393 278502 73411
rect 278558 73393 278626 73411
rect 278682 73393 278750 73449
rect 278807 73411 278874 73449
rect 278949 73411 278998 73449
rect 279091 73411 279122 73449
rect 279233 73411 279246 73449
rect 278806 73393 278874 73411
rect 278930 73393 278998 73411
rect 279054 73393 279122 73411
rect 279178 73393 279246 73411
rect 279302 73411 279319 73449
rect 279426 73411 279461 73449
rect 279550 73411 279603 73449
rect 279302 73393 279370 73411
rect 279426 73393 279494 73411
rect 279550 73393 279618 73411
rect 279674 73393 279742 73449
rect 279801 73411 279878 73467
rect 279798 73393 279878 73411
rect 277828 73325 279878 73393
rect 277828 73269 277882 73325
rect 277955 73269 278006 73325
rect 278097 73269 278130 73325
rect 278239 73269 278254 73325
rect 278310 73269 278325 73325
rect 278434 73269 278467 73325
rect 278558 73269 278609 73325
rect 278682 73269 278750 73325
rect 278807 73269 278874 73325
rect 278949 73269 278998 73325
rect 279091 73269 279122 73325
rect 279233 73269 279246 73325
rect 279302 73269 279319 73325
rect 279426 73269 279461 73325
rect 279550 73269 279603 73325
rect 279674 73269 279742 73325
rect 279801 73269 279878 73325
rect 277828 73201 279878 73269
rect 277828 73145 277882 73201
rect 277938 73183 278006 73201
rect 278062 73183 278130 73201
rect 278186 73183 278254 73201
rect 277955 73145 278006 73183
rect 278097 73145 278130 73183
rect 278239 73145 278254 73183
rect 278310 73183 278378 73201
rect 278434 73183 278502 73201
rect 278558 73183 278626 73201
rect 278310 73145 278325 73183
rect 278434 73145 278467 73183
rect 278558 73145 278609 73183
rect 278682 73145 278750 73201
rect 278806 73183 278874 73201
rect 278930 73183 278998 73201
rect 279054 73183 279122 73201
rect 279178 73183 279246 73201
rect 278807 73145 278874 73183
rect 278949 73145 278998 73183
rect 279091 73145 279122 73183
rect 279233 73145 279246 73183
rect 279302 73183 279370 73201
rect 279426 73183 279494 73201
rect 279550 73183 279618 73201
rect 279302 73145 279319 73183
rect 279426 73145 279461 73183
rect 279550 73145 279603 73183
rect 279674 73145 279742 73201
rect 279798 73183 279878 73201
rect 277828 73127 277899 73145
rect 277955 73127 278041 73145
rect 278097 73127 278183 73145
rect 278239 73127 278325 73145
rect 278381 73127 278467 73145
rect 278523 73127 278609 73145
rect 278665 73127 278751 73145
rect 278807 73127 278893 73145
rect 278949 73127 279035 73145
rect 279091 73127 279177 73145
rect 279233 73127 279319 73145
rect 279375 73127 279461 73145
rect 279517 73127 279603 73145
rect 279659 73127 279745 73145
rect 279801 73127 279878 73183
rect 277828 73077 279878 73127
rect 277828 73021 277882 73077
rect 277938 73041 278006 73077
rect 278062 73041 278130 73077
rect 278186 73041 278254 73077
rect 277955 73021 278006 73041
rect 278097 73021 278130 73041
rect 278239 73021 278254 73041
rect 278310 73041 278378 73077
rect 278434 73041 278502 73077
rect 278558 73041 278626 73077
rect 278310 73021 278325 73041
rect 278434 73021 278467 73041
rect 278558 73021 278609 73041
rect 278682 73021 278750 73077
rect 278806 73041 278874 73077
rect 278930 73041 278998 73077
rect 279054 73041 279122 73077
rect 279178 73041 279246 73077
rect 278807 73021 278874 73041
rect 278949 73021 278998 73041
rect 279091 73021 279122 73041
rect 279233 73021 279246 73041
rect 279302 73041 279370 73077
rect 279426 73041 279494 73077
rect 279550 73041 279618 73077
rect 279302 73021 279319 73041
rect 279426 73021 279461 73041
rect 279550 73021 279603 73041
rect 279674 73021 279742 73077
rect 279798 73041 279878 73077
rect 277828 72985 277899 73021
rect 277955 72985 278041 73021
rect 278097 72985 278183 73021
rect 278239 72985 278325 73021
rect 278381 72985 278467 73021
rect 278523 72985 278609 73021
rect 278665 72985 278751 73021
rect 278807 72985 278893 73021
rect 278949 72985 279035 73021
rect 279091 72985 279177 73021
rect 279233 72985 279319 73021
rect 279375 72985 279461 73021
rect 279517 72985 279603 73021
rect 279659 72985 279745 73021
rect 279801 72985 279878 73041
rect 277828 72953 279878 72985
rect 277828 72897 277882 72953
rect 277938 72899 278006 72953
rect 278062 72899 278130 72953
rect 278186 72899 278254 72953
rect 277955 72897 278006 72899
rect 278097 72897 278130 72899
rect 278239 72897 278254 72899
rect 278310 72899 278378 72953
rect 278434 72899 278502 72953
rect 278558 72899 278626 72953
rect 278310 72897 278325 72899
rect 278434 72897 278467 72899
rect 278558 72897 278609 72899
rect 278682 72897 278750 72953
rect 278806 72899 278874 72953
rect 278930 72899 278998 72953
rect 279054 72899 279122 72953
rect 279178 72899 279246 72953
rect 278807 72897 278874 72899
rect 278949 72897 278998 72899
rect 279091 72897 279122 72899
rect 279233 72897 279246 72899
rect 279302 72899 279370 72953
rect 279426 72899 279494 72953
rect 279550 72899 279618 72953
rect 279302 72897 279319 72899
rect 279426 72897 279461 72899
rect 279550 72897 279603 72899
rect 279674 72897 279742 72953
rect 279798 72899 279878 72953
rect 277828 72843 277899 72897
rect 277955 72843 278041 72897
rect 278097 72843 278183 72897
rect 278239 72843 278325 72897
rect 278381 72843 278467 72897
rect 278523 72843 278609 72897
rect 278665 72843 278751 72897
rect 278807 72843 278893 72897
rect 278949 72843 279035 72897
rect 279091 72843 279177 72897
rect 279233 72843 279319 72897
rect 279375 72843 279461 72897
rect 279517 72843 279603 72897
rect 279659 72843 279745 72897
rect 279801 72843 279878 72899
rect 277828 72829 279878 72843
rect 277828 72773 277882 72829
rect 277938 72773 278006 72829
rect 278062 72773 278130 72829
rect 278186 72773 278254 72829
rect 278310 72773 278378 72829
rect 278434 72773 278502 72829
rect 278558 72773 278626 72829
rect 278682 72773 278750 72829
rect 278806 72773 278874 72829
rect 278930 72773 278998 72829
rect 279054 72773 279122 72829
rect 279178 72773 279246 72829
rect 279302 72773 279370 72829
rect 279426 72773 279494 72829
rect 279550 72773 279618 72829
rect 279674 72773 279742 72829
rect 279798 72773 279878 72829
rect 277828 72757 279878 72773
rect 277828 72705 277899 72757
rect 277955 72705 278041 72757
rect 278097 72705 278183 72757
rect 278239 72705 278325 72757
rect 278381 72705 278467 72757
rect 278523 72705 278609 72757
rect 278665 72705 278751 72757
rect 278807 72705 278893 72757
rect 278949 72705 279035 72757
rect 279091 72705 279177 72757
rect 279233 72705 279319 72757
rect 279375 72705 279461 72757
rect 279517 72705 279603 72757
rect 279659 72705 279745 72757
rect 277828 72649 277882 72705
rect 277955 72701 278006 72705
rect 278097 72701 278130 72705
rect 278239 72701 278254 72705
rect 277938 72649 278006 72701
rect 278062 72649 278130 72701
rect 278186 72649 278254 72701
rect 278310 72701 278325 72705
rect 278434 72701 278467 72705
rect 278558 72701 278609 72705
rect 278310 72649 278378 72701
rect 278434 72649 278502 72701
rect 278558 72649 278626 72701
rect 278682 72649 278750 72705
rect 278807 72701 278874 72705
rect 278949 72701 278998 72705
rect 279091 72701 279122 72705
rect 279233 72701 279246 72705
rect 278806 72649 278874 72701
rect 278930 72649 278998 72701
rect 279054 72649 279122 72701
rect 279178 72649 279246 72701
rect 279302 72701 279319 72705
rect 279426 72701 279461 72705
rect 279550 72701 279603 72705
rect 279302 72649 279370 72701
rect 279426 72649 279494 72701
rect 279550 72649 279618 72701
rect 279674 72649 279742 72705
rect 279801 72701 279878 72757
rect 279798 72649 279878 72701
rect 277828 72615 279878 72649
rect 277828 72581 277899 72615
rect 277955 72581 278041 72615
rect 278097 72581 278183 72615
rect 278239 72581 278325 72615
rect 278381 72581 278467 72615
rect 278523 72581 278609 72615
rect 278665 72581 278751 72615
rect 278807 72581 278893 72615
rect 278949 72581 279035 72615
rect 279091 72581 279177 72615
rect 279233 72581 279319 72615
rect 279375 72581 279461 72615
rect 279517 72581 279603 72615
rect 279659 72581 279745 72615
rect 277828 72525 277882 72581
rect 277955 72559 278006 72581
rect 278097 72559 278130 72581
rect 278239 72559 278254 72581
rect 277938 72525 278006 72559
rect 278062 72525 278130 72559
rect 278186 72525 278254 72559
rect 278310 72559 278325 72581
rect 278434 72559 278467 72581
rect 278558 72559 278609 72581
rect 278310 72525 278378 72559
rect 278434 72525 278502 72559
rect 278558 72525 278626 72559
rect 278682 72525 278750 72581
rect 278807 72559 278874 72581
rect 278949 72559 278998 72581
rect 279091 72559 279122 72581
rect 279233 72559 279246 72581
rect 278806 72525 278874 72559
rect 278930 72525 278998 72559
rect 279054 72525 279122 72559
rect 279178 72525 279246 72559
rect 279302 72559 279319 72581
rect 279426 72559 279461 72581
rect 279550 72559 279603 72581
rect 279302 72525 279370 72559
rect 279426 72525 279494 72559
rect 279550 72525 279618 72559
rect 279674 72525 279742 72581
rect 279801 72559 279878 72615
rect 279798 72525 279878 72559
rect 277828 72473 279878 72525
rect 277828 72457 277899 72473
rect 277955 72457 278041 72473
rect 278097 72457 278183 72473
rect 278239 72457 278325 72473
rect 278381 72457 278467 72473
rect 278523 72457 278609 72473
rect 278665 72457 278751 72473
rect 278807 72457 278893 72473
rect 278949 72457 279035 72473
rect 279091 72457 279177 72473
rect 279233 72457 279319 72473
rect 279375 72457 279461 72473
rect 279517 72457 279603 72473
rect 279659 72457 279745 72473
rect 277828 72401 277882 72457
rect 277955 72417 278006 72457
rect 278097 72417 278130 72457
rect 278239 72417 278254 72457
rect 277938 72401 278006 72417
rect 278062 72401 278130 72417
rect 278186 72401 278254 72417
rect 278310 72417 278325 72457
rect 278434 72417 278467 72457
rect 278558 72417 278609 72457
rect 278310 72401 278378 72417
rect 278434 72401 278502 72417
rect 278558 72401 278626 72417
rect 278682 72401 278750 72457
rect 278807 72417 278874 72457
rect 278949 72417 278998 72457
rect 279091 72417 279122 72457
rect 279233 72417 279246 72457
rect 278806 72401 278874 72417
rect 278930 72401 278998 72417
rect 279054 72401 279122 72417
rect 279178 72401 279246 72417
rect 279302 72417 279319 72457
rect 279426 72417 279461 72457
rect 279550 72417 279603 72457
rect 279302 72401 279370 72417
rect 279426 72401 279494 72417
rect 279550 72401 279618 72417
rect 279674 72401 279742 72457
rect 279801 72417 279878 72473
rect 279798 72401 279878 72417
rect 277828 72333 279878 72401
rect 277828 72277 277882 72333
rect 277938 72331 278006 72333
rect 278062 72331 278130 72333
rect 278186 72331 278254 72333
rect 277955 72277 278006 72331
rect 278097 72277 278130 72331
rect 278239 72277 278254 72331
rect 278310 72331 278378 72333
rect 278434 72331 278502 72333
rect 278558 72331 278626 72333
rect 278310 72277 278325 72331
rect 278434 72277 278467 72331
rect 278558 72277 278609 72331
rect 278682 72277 278750 72333
rect 278806 72331 278874 72333
rect 278930 72331 278998 72333
rect 279054 72331 279122 72333
rect 279178 72331 279246 72333
rect 278807 72277 278874 72331
rect 278949 72277 278998 72331
rect 279091 72277 279122 72331
rect 279233 72277 279246 72331
rect 279302 72331 279370 72333
rect 279426 72331 279494 72333
rect 279550 72331 279618 72333
rect 279302 72277 279319 72331
rect 279426 72277 279461 72331
rect 279550 72277 279603 72331
rect 279674 72277 279742 72333
rect 279798 72331 279878 72333
rect 277828 72275 277899 72277
rect 277955 72275 278041 72277
rect 278097 72275 278183 72277
rect 278239 72275 278325 72277
rect 278381 72275 278467 72277
rect 278523 72275 278609 72277
rect 278665 72275 278751 72277
rect 278807 72275 278893 72277
rect 278949 72275 279035 72277
rect 279091 72275 279177 72277
rect 279233 72275 279319 72277
rect 279375 72275 279461 72277
rect 279517 72275 279603 72277
rect 279659 72275 279745 72277
rect 279801 72275 279878 72331
rect 277828 72209 279878 72275
rect 277828 72153 277882 72209
rect 277938 72189 278006 72209
rect 278062 72189 278130 72209
rect 278186 72189 278254 72209
rect 277955 72153 278006 72189
rect 278097 72153 278130 72189
rect 278239 72153 278254 72189
rect 278310 72189 278378 72209
rect 278434 72189 278502 72209
rect 278558 72189 278626 72209
rect 278310 72153 278325 72189
rect 278434 72153 278467 72189
rect 278558 72153 278609 72189
rect 278682 72153 278750 72209
rect 278806 72189 278874 72209
rect 278930 72189 278998 72209
rect 279054 72189 279122 72209
rect 279178 72189 279246 72209
rect 278807 72153 278874 72189
rect 278949 72153 278998 72189
rect 279091 72153 279122 72189
rect 279233 72153 279246 72189
rect 279302 72189 279370 72209
rect 279426 72189 279494 72209
rect 279550 72189 279618 72209
rect 279302 72153 279319 72189
rect 279426 72153 279461 72189
rect 279550 72153 279603 72189
rect 279674 72153 279742 72209
rect 279798 72189 279878 72209
rect 277828 72133 277899 72153
rect 277955 72133 278041 72153
rect 278097 72133 278183 72153
rect 278239 72133 278325 72153
rect 278381 72133 278467 72153
rect 278523 72133 278609 72153
rect 278665 72133 278751 72153
rect 278807 72133 278893 72153
rect 278949 72133 279035 72153
rect 279091 72133 279177 72153
rect 279233 72133 279319 72153
rect 279375 72133 279461 72153
rect 279517 72133 279603 72153
rect 279659 72133 279745 72153
rect 279801 72133 279878 72189
rect 277828 72088 279878 72133
rect 280198 74035 282248 74088
rect 280198 73979 280269 74035
rect 280325 73979 280411 74035
rect 280467 73979 280553 74035
rect 280609 73979 280695 74035
rect 280751 73979 280837 74035
rect 280893 73979 280979 74035
rect 281035 73979 281121 74035
rect 281177 73979 281263 74035
rect 281319 73979 281405 74035
rect 281461 73979 281547 74035
rect 281603 73979 281689 74035
rect 281745 73979 281831 74035
rect 281887 73979 281973 74035
rect 282029 73979 282115 74035
rect 282171 73979 282248 74035
rect 280198 73945 282248 73979
rect 280198 73889 280252 73945
rect 280308 73893 280376 73945
rect 280432 73893 280500 73945
rect 280556 73893 280624 73945
rect 280325 73889 280376 73893
rect 280467 73889 280500 73893
rect 280609 73889 280624 73893
rect 280680 73893 280748 73945
rect 280804 73893 280872 73945
rect 280928 73893 280996 73945
rect 280680 73889 280695 73893
rect 280804 73889 280837 73893
rect 280928 73889 280979 73893
rect 281052 73889 281120 73945
rect 281176 73893 281244 73945
rect 281300 73893 281368 73945
rect 281424 73893 281492 73945
rect 281548 73893 281616 73945
rect 281177 73889 281244 73893
rect 281319 73889 281368 73893
rect 281461 73889 281492 73893
rect 281603 73889 281616 73893
rect 281672 73893 281740 73945
rect 281796 73893 281864 73945
rect 281920 73893 281988 73945
rect 281672 73889 281689 73893
rect 281796 73889 281831 73893
rect 281920 73889 281973 73893
rect 282044 73889 282112 73945
rect 282168 73893 282248 73945
rect 280198 73837 280269 73889
rect 280325 73837 280411 73889
rect 280467 73837 280553 73889
rect 280609 73837 280695 73889
rect 280751 73837 280837 73889
rect 280893 73837 280979 73889
rect 281035 73837 281121 73889
rect 281177 73837 281263 73889
rect 281319 73837 281405 73889
rect 281461 73837 281547 73889
rect 281603 73837 281689 73889
rect 281745 73837 281831 73889
rect 281887 73837 281973 73889
rect 282029 73837 282115 73889
rect 282171 73837 282248 73893
rect 280198 73821 282248 73837
rect 280198 73765 280252 73821
rect 280308 73765 280376 73821
rect 280432 73765 280500 73821
rect 280556 73765 280624 73821
rect 280680 73765 280748 73821
rect 280804 73765 280872 73821
rect 280928 73765 280996 73821
rect 281052 73765 281120 73821
rect 281176 73765 281244 73821
rect 281300 73765 281368 73821
rect 281424 73765 281492 73821
rect 281548 73765 281616 73821
rect 281672 73765 281740 73821
rect 281796 73765 281864 73821
rect 281920 73765 281988 73821
rect 282044 73765 282112 73821
rect 282168 73765 282248 73821
rect 280198 73751 282248 73765
rect 280198 73697 280269 73751
rect 280325 73697 280411 73751
rect 280467 73697 280553 73751
rect 280609 73697 280695 73751
rect 280751 73697 280837 73751
rect 280893 73697 280979 73751
rect 281035 73697 281121 73751
rect 281177 73697 281263 73751
rect 281319 73697 281405 73751
rect 281461 73697 281547 73751
rect 281603 73697 281689 73751
rect 281745 73697 281831 73751
rect 281887 73697 281973 73751
rect 282029 73697 282115 73751
rect 280198 73641 280252 73697
rect 280325 73695 280376 73697
rect 280467 73695 280500 73697
rect 280609 73695 280624 73697
rect 280308 73641 280376 73695
rect 280432 73641 280500 73695
rect 280556 73641 280624 73695
rect 280680 73695 280695 73697
rect 280804 73695 280837 73697
rect 280928 73695 280979 73697
rect 280680 73641 280748 73695
rect 280804 73641 280872 73695
rect 280928 73641 280996 73695
rect 281052 73641 281120 73697
rect 281177 73695 281244 73697
rect 281319 73695 281368 73697
rect 281461 73695 281492 73697
rect 281603 73695 281616 73697
rect 281176 73641 281244 73695
rect 281300 73641 281368 73695
rect 281424 73641 281492 73695
rect 281548 73641 281616 73695
rect 281672 73695 281689 73697
rect 281796 73695 281831 73697
rect 281920 73695 281973 73697
rect 281672 73641 281740 73695
rect 281796 73641 281864 73695
rect 281920 73641 281988 73695
rect 282044 73641 282112 73697
rect 282171 73695 282248 73751
rect 282168 73641 282248 73695
rect 280198 73609 282248 73641
rect 280198 73573 280269 73609
rect 280325 73573 280411 73609
rect 280467 73573 280553 73609
rect 280609 73573 280695 73609
rect 280751 73573 280837 73609
rect 280893 73573 280979 73609
rect 281035 73573 281121 73609
rect 281177 73573 281263 73609
rect 281319 73573 281405 73609
rect 281461 73573 281547 73609
rect 281603 73573 281689 73609
rect 281745 73573 281831 73609
rect 281887 73573 281973 73609
rect 282029 73573 282115 73609
rect 280198 73517 280252 73573
rect 280325 73553 280376 73573
rect 280467 73553 280500 73573
rect 280609 73553 280624 73573
rect 280308 73517 280376 73553
rect 280432 73517 280500 73553
rect 280556 73517 280624 73553
rect 280680 73553 280695 73573
rect 280804 73553 280837 73573
rect 280928 73553 280979 73573
rect 280680 73517 280748 73553
rect 280804 73517 280872 73553
rect 280928 73517 280996 73553
rect 281052 73517 281120 73573
rect 281177 73553 281244 73573
rect 281319 73553 281368 73573
rect 281461 73553 281492 73573
rect 281603 73553 281616 73573
rect 281176 73517 281244 73553
rect 281300 73517 281368 73553
rect 281424 73517 281492 73553
rect 281548 73517 281616 73553
rect 281672 73553 281689 73573
rect 281796 73553 281831 73573
rect 281920 73553 281973 73573
rect 281672 73517 281740 73553
rect 281796 73517 281864 73553
rect 281920 73517 281988 73553
rect 282044 73517 282112 73573
rect 282171 73553 282248 73609
rect 282168 73517 282248 73553
rect 280198 73467 282248 73517
rect 280198 73449 280269 73467
rect 280325 73449 280411 73467
rect 280467 73449 280553 73467
rect 280609 73449 280695 73467
rect 280751 73449 280837 73467
rect 280893 73449 280979 73467
rect 281035 73449 281121 73467
rect 281177 73449 281263 73467
rect 281319 73449 281405 73467
rect 281461 73449 281547 73467
rect 281603 73449 281689 73467
rect 281745 73449 281831 73467
rect 281887 73449 281973 73467
rect 282029 73449 282115 73467
rect 280198 73393 280252 73449
rect 280325 73411 280376 73449
rect 280467 73411 280500 73449
rect 280609 73411 280624 73449
rect 280308 73393 280376 73411
rect 280432 73393 280500 73411
rect 280556 73393 280624 73411
rect 280680 73411 280695 73449
rect 280804 73411 280837 73449
rect 280928 73411 280979 73449
rect 280680 73393 280748 73411
rect 280804 73393 280872 73411
rect 280928 73393 280996 73411
rect 281052 73393 281120 73449
rect 281177 73411 281244 73449
rect 281319 73411 281368 73449
rect 281461 73411 281492 73449
rect 281603 73411 281616 73449
rect 281176 73393 281244 73411
rect 281300 73393 281368 73411
rect 281424 73393 281492 73411
rect 281548 73393 281616 73411
rect 281672 73411 281689 73449
rect 281796 73411 281831 73449
rect 281920 73411 281973 73449
rect 281672 73393 281740 73411
rect 281796 73393 281864 73411
rect 281920 73393 281988 73411
rect 282044 73393 282112 73449
rect 282171 73411 282248 73467
rect 282168 73393 282248 73411
rect 280198 73325 282248 73393
rect 280198 73269 280252 73325
rect 280325 73269 280376 73325
rect 280467 73269 280500 73325
rect 280609 73269 280624 73325
rect 280680 73269 280695 73325
rect 280804 73269 280837 73325
rect 280928 73269 280979 73325
rect 281052 73269 281120 73325
rect 281177 73269 281244 73325
rect 281319 73269 281368 73325
rect 281461 73269 281492 73325
rect 281603 73269 281616 73325
rect 281672 73269 281689 73325
rect 281796 73269 281831 73325
rect 281920 73269 281973 73325
rect 282044 73269 282112 73325
rect 282171 73269 282248 73325
rect 280198 73201 282248 73269
rect 280198 73145 280252 73201
rect 280308 73183 280376 73201
rect 280432 73183 280500 73201
rect 280556 73183 280624 73201
rect 280325 73145 280376 73183
rect 280467 73145 280500 73183
rect 280609 73145 280624 73183
rect 280680 73183 280748 73201
rect 280804 73183 280872 73201
rect 280928 73183 280996 73201
rect 280680 73145 280695 73183
rect 280804 73145 280837 73183
rect 280928 73145 280979 73183
rect 281052 73145 281120 73201
rect 281176 73183 281244 73201
rect 281300 73183 281368 73201
rect 281424 73183 281492 73201
rect 281548 73183 281616 73201
rect 281177 73145 281244 73183
rect 281319 73145 281368 73183
rect 281461 73145 281492 73183
rect 281603 73145 281616 73183
rect 281672 73183 281740 73201
rect 281796 73183 281864 73201
rect 281920 73183 281988 73201
rect 281672 73145 281689 73183
rect 281796 73145 281831 73183
rect 281920 73145 281973 73183
rect 282044 73145 282112 73201
rect 282168 73183 282248 73201
rect 280198 73127 280269 73145
rect 280325 73127 280411 73145
rect 280467 73127 280553 73145
rect 280609 73127 280695 73145
rect 280751 73127 280837 73145
rect 280893 73127 280979 73145
rect 281035 73127 281121 73145
rect 281177 73127 281263 73145
rect 281319 73127 281405 73145
rect 281461 73127 281547 73145
rect 281603 73127 281689 73145
rect 281745 73127 281831 73145
rect 281887 73127 281973 73145
rect 282029 73127 282115 73145
rect 282171 73127 282248 73183
rect 280198 73077 282248 73127
rect 280198 73021 280252 73077
rect 280308 73041 280376 73077
rect 280432 73041 280500 73077
rect 280556 73041 280624 73077
rect 280325 73021 280376 73041
rect 280467 73021 280500 73041
rect 280609 73021 280624 73041
rect 280680 73041 280748 73077
rect 280804 73041 280872 73077
rect 280928 73041 280996 73077
rect 280680 73021 280695 73041
rect 280804 73021 280837 73041
rect 280928 73021 280979 73041
rect 281052 73021 281120 73077
rect 281176 73041 281244 73077
rect 281300 73041 281368 73077
rect 281424 73041 281492 73077
rect 281548 73041 281616 73077
rect 281177 73021 281244 73041
rect 281319 73021 281368 73041
rect 281461 73021 281492 73041
rect 281603 73021 281616 73041
rect 281672 73041 281740 73077
rect 281796 73041 281864 73077
rect 281920 73041 281988 73077
rect 281672 73021 281689 73041
rect 281796 73021 281831 73041
rect 281920 73021 281973 73041
rect 282044 73021 282112 73077
rect 282168 73041 282248 73077
rect 280198 72985 280269 73021
rect 280325 72985 280411 73021
rect 280467 72985 280553 73021
rect 280609 72985 280695 73021
rect 280751 72985 280837 73021
rect 280893 72985 280979 73021
rect 281035 72985 281121 73021
rect 281177 72985 281263 73021
rect 281319 72985 281405 73021
rect 281461 72985 281547 73021
rect 281603 72985 281689 73021
rect 281745 72985 281831 73021
rect 281887 72985 281973 73021
rect 282029 72985 282115 73021
rect 282171 72985 282248 73041
rect 280198 72953 282248 72985
rect 280198 72897 280252 72953
rect 280308 72899 280376 72953
rect 280432 72899 280500 72953
rect 280556 72899 280624 72953
rect 280325 72897 280376 72899
rect 280467 72897 280500 72899
rect 280609 72897 280624 72899
rect 280680 72899 280748 72953
rect 280804 72899 280872 72953
rect 280928 72899 280996 72953
rect 280680 72897 280695 72899
rect 280804 72897 280837 72899
rect 280928 72897 280979 72899
rect 281052 72897 281120 72953
rect 281176 72899 281244 72953
rect 281300 72899 281368 72953
rect 281424 72899 281492 72953
rect 281548 72899 281616 72953
rect 281177 72897 281244 72899
rect 281319 72897 281368 72899
rect 281461 72897 281492 72899
rect 281603 72897 281616 72899
rect 281672 72899 281740 72953
rect 281796 72899 281864 72953
rect 281920 72899 281988 72953
rect 281672 72897 281689 72899
rect 281796 72897 281831 72899
rect 281920 72897 281973 72899
rect 282044 72897 282112 72953
rect 282168 72899 282248 72953
rect 280198 72843 280269 72897
rect 280325 72843 280411 72897
rect 280467 72843 280553 72897
rect 280609 72843 280695 72897
rect 280751 72843 280837 72897
rect 280893 72843 280979 72897
rect 281035 72843 281121 72897
rect 281177 72843 281263 72897
rect 281319 72843 281405 72897
rect 281461 72843 281547 72897
rect 281603 72843 281689 72897
rect 281745 72843 281831 72897
rect 281887 72843 281973 72897
rect 282029 72843 282115 72897
rect 282171 72843 282248 72899
rect 280198 72829 282248 72843
rect 280198 72773 280252 72829
rect 280308 72773 280376 72829
rect 280432 72773 280500 72829
rect 280556 72773 280624 72829
rect 280680 72773 280748 72829
rect 280804 72773 280872 72829
rect 280928 72773 280996 72829
rect 281052 72773 281120 72829
rect 281176 72773 281244 72829
rect 281300 72773 281368 72829
rect 281424 72773 281492 72829
rect 281548 72773 281616 72829
rect 281672 72773 281740 72829
rect 281796 72773 281864 72829
rect 281920 72773 281988 72829
rect 282044 72773 282112 72829
rect 282168 72773 282248 72829
rect 280198 72757 282248 72773
rect 280198 72705 280269 72757
rect 280325 72705 280411 72757
rect 280467 72705 280553 72757
rect 280609 72705 280695 72757
rect 280751 72705 280837 72757
rect 280893 72705 280979 72757
rect 281035 72705 281121 72757
rect 281177 72705 281263 72757
rect 281319 72705 281405 72757
rect 281461 72705 281547 72757
rect 281603 72705 281689 72757
rect 281745 72705 281831 72757
rect 281887 72705 281973 72757
rect 282029 72705 282115 72757
rect 280198 72649 280252 72705
rect 280325 72701 280376 72705
rect 280467 72701 280500 72705
rect 280609 72701 280624 72705
rect 280308 72649 280376 72701
rect 280432 72649 280500 72701
rect 280556 72649 280624 72701
rect 280680 72701 280695 72705
rect 280804 72701 280837 72705
rect 280928 72701 280979 72705
rect 280680 72649 280748 72701
rect 280804 72649 280872 72701
rect 280928 72649 280996 72701
rect 281052 72649 281120 72705
rect 281177 72701 281244 72705
rect 281319 72701 281368 72705
rect 281461 72701 281492 72705
rect 281603 72701 281616 72705
rect 281176 72649 281244 72701
rect 281300 72649 281368 72701
rect 281424 72649 281492 72701
rect 281548 72649 281616 72701
rect 281672 72701 281689 72705
rect 281796 72701 281831 72705
rect 281920 72701 281973 72705
rect 281672 72649 281740 72701
rect 281796 72649 281864 72701
rect 281920 72649 281988 72701
rect 282044 72649 282112 72705
rect 282171 72701 282248 72757
rect 282168 72649 282248 72701
rect 280198 72615 282248 72649
rect 280198 72581 280269 72615
rect 280325 72581 280411 72615
rect 280467 72581 280553 72615
rect 280609 72581 280695 72615
rect 280751 72581 280837 72615
rect 280893 72581 280979 72615
rect 281035 72581 281121 72615
rect 281177 72581 281263 72615
rect 281319 72581 281405 72615
rect 281461 72581 281547 72615
rect 281603 72581 281689 72615
rect 281745 72581 281831 72615
rect 281887 72581 281973 72615
rect 282029 72581 282115 72615
rect 280198 72525 280252 72581
rect 280325 72559 280376 72581
rect 280467 72559 280500 72581
rect 280609 72559 280624 72581
rect 280308 72525 280376 72559
rect 280432 72525 280500 72559
rect 280556 72525 280624 72559
rect 280680 72559 280695 72581
rect 280804 72559 280837 72581
rect 280928 72559 280979 72581
rect 280680 72525 280748 72559
rect 280804 72525 280872 72559
rect 280928 72525 280996 72559
rect 281052 72525 281120 72581
rect 281177 72559 281244 72581
rect 281319 72559 281368 72581
rect 281461 72559 281492 72581
rect 281603 72559 281616 72581
rect 281176 72525 281244 72559
rect 281300 72525 281368 72559
rect 281424 72525 281492 72559
rect 281548 72525 281616 72559
rect 281672 72559 281689 72581
rect 281796 72559 281831 72581
rect 281920 72559 281973 72581
rect 281672 72525 281740 72559
rect 281796 72525 281864 72559
rect 281920 72525 281988 72559
rect 282044 72525 282112 72581
rect 282171 72559 282248 72615
rect 282168 72525 282248 72559
rect 280198 72473 282248 72525
rect 280198 72457 280269 72473
rect 280325 72457 280411 72473
rect 280467 72457 280553 72473
rect 280609 72457 280695 72473
rect 280751 72457 280837 72473
rect 280893 72457 280979 72473
rect 281035 72457 281121 72473
rect 281177 72457 281263 72473
rect 281319 72457 281405 72473
rect 281461 72457 281547 72473
rect 281603 72457 281689 72473
rect 281745 72457 281831 72473
rect 281887 72457 281973 72473
rect 282029 72457 282115 72473
rect 280198 72401 280252 72457
rect 280325 72417 280376 72457
rect 280467 72417 280500 72457
rect 280609 72417 280624 72457
rect 280308 72401 280376 72417
rect 280432 72401 280500 72417
rect 280556 72401 280624 72417
rect 280680 72417 280695 72457
rect 280804 72417 280837 72457
rect 280928 72417 280979 72457
rect 280680 72401 280748 72417
rect 280804 72401 280872 72417
rect 280928 72401 280996 72417
rect 281052 72401 281120 72457
rect 281177 72417 281244 72457
rect 281319 72417 281368 72457
rect 281461 72417 281492 72457
rect 281603 72417 281616 72457
rect 281176 72401 281244 72417
rect 281300 72401 281368 72417
rect 281424 72401 281492 72417
rect 281548 72401 281616 72417
rect 281672 72417 281689 72457
rect 281796 72417 281831 72457
rect 281920 72417 281973 72457
rect 281672 72401 281740 72417
rect 281796 72401 281864 72417
rect 281920 72401 281988 72417
rect 282044 72401 282112 72457
rect 282171 72417 282248 72473
rect 282168 72401 282248 72417
rect 280198 72333 282248 72401
rect 280198 72277 280252 72333
rect 280308 72331 280376 72333
rect 280432 72331 280500 72333
rect 280556 72331 280624 72333
rect 280325 72277 280376 72331
rect 280467 72277 280500 72331
rect 280609 72277 280624 72331
rect 280680 72331 280748 72333
rect 280804 72331 280872 72333
rect 280928 72331 280996 72333
rect 280680 72277 280695 72331
rect 280804 72277 280837 72331
rect 280928 72277 280979 72331
rect 281052 72277 281120 72333
rect 281176 72331 281244 72333
rect 281300 72331 281368 72333
rect 281424 72331 281492 72333
rect 281548 72331 281616 72333
rect 281177 72277 281244 72331
rect 281319 72277 281368 72331
rect 281461 72277 281492 72331
rect 281603 72277 281616 72331
rect 281672 72331 281740 72333
rect 281796 72331 281864 72333
rect 281920 72331 281988 72333
rect 281672 72277 281689 72331
rect 281796 72277 281831 72331
rect 281920 72277 281973 72331
rect 282044 72277 282112 72333
rect 282168 72331 282248 72333
rect 280198 72275 280269 72277
rect 280325 72275 280411 72277
rect 280467 72275 280553 72277
rect 280609 72275 280695 72277
rect 280751 72275 280837 72277
rect 280893 72275 280979 72277
rect 281035 72275 281121 72277
rect 281177 72275 281263 72277
rect 281319 72275 281405 72277
rect 281461 72275 281547 72277
rect 281603 72275 281689 72277
rect 281745 72275 281831 72277
rect 281887 72275 281973 72277
rect 282029 72275 282115 72277
rect 282171 72275 282248 72331
rect 280198 72209 282248 72275
rect 280198 72153 280252 72209
rect 280308 72189 280376 72209
rect 280432 72189 280500 72209
rect 280556 72189 280624 72209
rect 280325 72153 280376 72189
rect 280467 72153 280500 72189
rect 280609 72153 280624 72189
rect 280680 72189 280748 72209
rect 280804 72189 280872 72209
rect 280928 72189 280996 72209
rect 280680 72153 280695 72189
rect 280804 72153 280837 72189
rect 280928 72153 280979 72189
rect 281052 72153 281120 72209
rect 281176 72189 281244 72209
rect 281300 72189 281368 72209
rect 281424 72189 281492 72209
rect 281548 72189 281616 72209
rect 281177 72153 281244 72189
rect 281319 72153 281368 72189
rect 281461 72153 281492 72189
rect 281603 72153 281616 72189
rect 281672 72189 281740 72209
rect 281796 72189 281864 72209
rect 281920 72189 281988 72209
rect 281672 72153 281689 72189
rect 281796 72153 281831 72189
rect 281920 72153 281973 72189
rect 282044 72153 282112 72209
rect 282168 72189 282248 72209
rect 280198 72133 280269 72153
rect 280325 72133 280411 72153
rect 280467 72133 280553 72153
rect 280609 72133 280695 72153
rect 280751 72133 280837 72153
rect 280893 72133 280979 72153
rect 281035 72133 281121 72153
rect 281177 72133 281263 72153
rect 281319 72133 281405 72153
rect 281461 72133 281547 72153
rect 281603 72133 281689 72153
rect 281745 72133 281831 72153
rect 281887 72133 281973 72153
rect 282029 72133 282115 72153
rect 282171 72133 282248 72189
rect 280198 72088 282248 72133
rect 282828 74035 284728 74088
rect 282828 73979 282899 74035
rect 282955 73979 283041 74035
rect 283097 73979 283183 74035
rect 283239 73979 283325 74035
rect 283381 73979 283467 74035
rect 283523 73979 283609 74035
rect 283665 73979 283751 74035
rect 283807 73979 283893 74035
rect 283949 73979 284728 74035
rect 282828 73945 284728 73979
rect 282828 73889 282882 73945
rect 282938 73893 283006 73945
rect 283062 73893 283130 73945
rect 283186 73893 283254 73945
rect 282955 73889 283006 73893
rect 283097 73889 283130 73893
rect 283239 73889 283254 73893
rect 283310 73893 283378 73945
rect 283434 73893 283502 73945
rect 283558 73893 283626 73945
rect 283310 73889 283325 73893
rect 283434 73889 283467 73893
rect 283558 73889 283609 73893
rect 283682 73889 283750 73945
rect 283806 73893 283874 73945
rect 283930 73893 284728 73945
rect 283807 73889 283874 73893
rect 282828 73837 282899 73889
rect 282955 73837 283041 73889
rect 283097 73837 283183 73889
rect 283239 73837 283325 73889
rect 283381 73837 283467 73889
rect 283523 73837 283609 73889
rect 283665 73837 283751 73889
rect 283807 73837 283893 73889
rect 283949 73837 284728 73893
rect 282828 73821 284728 73837
rect 282828 73765 282882 73821
rect 282938 73765 283006 73821
rect 283062 73765 283130 73821
rect 283186 73765 283254 73821
rect 283310 73765 283378 73821
rect 283434 73765 283502 73821
rect 283558 73765 283626 73821
rect 283682 73765 283750 73821
rect 283806 73765 283874 73821
rect 283930 73765 284728 73821
rect 282828 73751 284728 73765
rect 282828 73697 282899 73751
rect 282955 73697 283041 73751
rect 283097 73697 283183 73751
rect 283239 73697 283325 73751
rect 283381 73697 283467 73751
rect 283523 73697 283609 73751
rect 283665 73697 283751 73751
rect 283807 73697 283893 73751
rect 282828 73641 282882 73697
rect 282955 73695 283006 73697
rect 283097 73695 283130 73697
rect 283239 73695 283254 73697
rect 282938 73641 283006 73695
rect 283062 73641 283130 73695
rect 283186 73641 283254 73695
rect 283310 73695 283325 73697
rect 283434 73695 283467 73697
rect 283558 73695 283609 73697
rect 283310 73641 283378 73695
rect 283434 73641 283502 73695
rect 283558 73641 283626 73695
rect 283682 73641 283750 73697
rect 283807 73695 283874 73697
rect 283949 73695 284728 73751
rect 283806 73641 283874 73695
rect 283930 73641 284728 73695
rect 282828 73609 284728 73641
rect 282828 73573 282899 73609
rect 282955 73573 283041 73609
rect 283097 73573 283183 73609
rect 283239 73573 283325 73609
rect 283381 73573 283467 73609
rect 283523 73573 283609 73609
rect 283665 73573 283751 73609
rect 283807 73573 283893 73609
rect 282828 73517 282882 73573
rect 282955 73553 283006 73573
rect 283097 73553 283130 73573
rect 283239 73553 283254 73573
rect 282938 73517 283006 73553
rect 283062 73517 283130 73553
rect 283186 73517 283254 73553
rect 283310 73553 283325 73573
rect 283434 73553 283467 73573
rect 283558 73553 283609 73573
rect 283310 73517 283378 73553
rect 283434 73517 283502 73553
rect 283558 73517 283626 73553
rect 283682 73517 283750 73573
rect 283807 73553 283874 73573
rect 283949 73553 284728 73609
rect 283806 73517 283874 73553
rect 283930 73517 284728 73553
rect 282828 73467 284728 73517
rect 282828 73449 282899 73467
rect 282955 73449 283041 73467
rect 283097 73449 283183 73467
rect 283239 73449 283325 73467
rect 283381 73449 283467 73467
rect 283523 73449 283609 73467
rect 283665 73449 283751 73467
rect 283807 73449 283893 73467
rect 282828 73393 282882 73449
rect 282955 73411 283006 73449
rect 283097 73411 283130 73449
rect 283239 73411 283254 73449
rect 282938 73393 283006 73411
rect 283062 73393 283130 73411
rect 283186 73393 283254 73411
rect 283310 73411 283325 73449
rect 283434 73411 283467 73449
rect 283558 73411 283609 73449
rect 283310 73393 283378 73411
rect 283434 73393 283502 73411
rect 283558 73393 283626 73411
rect 283682 73393 283750 73449
rect 283807 73411 283874 73449
rect 283949 73411 284728 73467
rect 283806 73393 283874 73411
rect 283930 73393 284728 73411
rect 282828 73325 284728 73393
rect 282828 73269 282882 73325
rect 282955 73269 283006 73325
rect 283097 73269 283130 73325
rect 283239 73269 283254 73325
rect 283310 73269 283325 73325
rect 283434 73269 283467 73325
rect 283558 73269 283609 73325
rect 283682 73269 283750 73325
rect 283807 73269 283874 73325
rect 283949 73269 284728 73325
rect 282828 73201 284728 73269
rect 282828 73145 282882 73201
rect 282938 73183 283006 73201
rect 283062 73183 283130 73201
rect 283186 73183 283254 73201
rect 282955 73145 283006 73183
rect 283097 73145 283130 73183
rect 283239 73145 283254 73183
rect 283310 73183 283378 73201
rect 283434 73183 283502 73201
rect 283558 73183 283626 73201
rect 283310 73145 283325 73183
rect 283434 73145 283467 73183
rect 283558 73145 283609 73183
rect 283682 73145 283750 73201
rect 283806 73183 283874 73201
rect 283930 73183 284728 73201
rect 283807 73145 283874 73183
rect 282828 73127 282899 73145
rect 282955 73127 283041 73145
rect 283097 73127 283183 73145
rect 283239 73127 283325 73145
rect 283381 73127 283467 73145
rect 283523 73127 283609 73145
rect 283665 73127 283751 73145
rect 283807 73127 283893 73145
rect 283949 73127 284728 73183
rect 282828 73077 284728 73127
rect 282828 73021 282882 73077
rect 282938 73041 283006 73077
rect 283062 73041 283130 73077
rect 283186 73041 283254 73077
rect 282955 73021 283006 73041
rect 283097 73021 283130 73041
rect 283239 73021 283254 73041
rect 283310 73041 283378 73077
rect 283434 73041 283502 73077
rect 283558 73041 283626 73077
rect 283310 73021 283325 73041
rect 283434 73021 283467 73041
rect 283558 73021 283609 73041
rect 283682 73021 283750 73077
rect 283806 73041 283874 73077
rect 283930 73041 284728 73077
rect 283807 73021 283874 73041
rect 282828 72985 282899 73021
rect 282955 72985 283041 73021
rect 283097 72985 283183 73021
rect 283239 72985 283325 73021
rect 283381 72985 283467 73021
rect 283523 72985 283609 73021
rect 283665 72985 283751 73021
rect 283807 72985 283893 73021
rect 283949 72985 284728 73041
rect 282828 72953 284728 72985
rect 282828 72897 282882 72953
rect 282938 72899 283006 72953
rect 283062 72899 283130 72953
rect 283186 72899 283254 72953
rect 282955 72897 283006 72899
rect 283097 72897 283130 72899
rect 283239 72897 283254 72899
rect 283310 72899 283378 72953
rect 283434 72899 283502 72953
rect 283558 72899 283626 72953
rect 283310 72897 283325 72899
rect 283434 72897 283467 72899
rect 283558 72897 283609 72899
rect 283682 72897 283750 72953
rect 283806 72899 283874 72953
rect 283930 72899 284728 72953
rect 283807 72897 283874 72899
rect 282828 72843 282899 72897
rect 282955 72843 283041 72897
rect 283097 72843 283183 72897
rect 283239 72843 283325 72897
rect 283381 72843 283467 72897
rect 283523 72843 283609 72897
rect 283665 72843 283751 72897
rect 283807 72843 283893 72897
rect 283949 72843 284728 72899
rect 282828 72829 284728 72843
rect 282828 72773 282882 72829
rect 282938 72773 283006 72829
rect 283062 72773 283130 72829
rect 283186 72773 283254 72829
rect 283310 72773 283378 72829
rect 283434 72773 283502 72829
rect 283558 72773 283626 72829
rect 283682 72773 283750 72829
rect 283806 72773 283874 72829
rect 283930 72773 284728 72829
rect 282828 72757 284728 72773
rect 282828 72705 282899 72757
rect 282955 72705 283041 72757
rect 283097 72705 283183 72757
rect 283239 72705 283325 72757
rect 283381 72705 283467 72757
rect 283523 72705 283609 72757
rect 283665 72705 283751 72757
rect 283807 72705 283893 72757
rect 282828 72649 282882 72705
rect 282955 72701 283006 72705
rect 283097 72701 283130 72705
rect 283239 72701 283254 72705
rect 282938 72649 283006 72701
rect 283062 72649 283130 72701
rect 283186 72649 283254 72701
rect 283310 72701 283325 72705
rect 283434 72701 283467 72705
rect 283558 72701 283609 72705
rect 283310 72649 283378 72701
rect 283434 72649 283502 72701
rect 283558 72649 283626 72701
rect 283682 72649 283750 72705
rect 283807 72701 283874 72705
rect 283949 72701 284728 72757
rect 283806 72649 283874 72701
rect 283930 72649 284728 72701
rect 282828 72615 284728 72649
rect 282828 72581 282899 72615
rect 282955 72581 283041 72615
rect 283097 72581 283183 72615
rect 283239 72581 283325 72615
rect 283381 72581 283467 72615
rect 283523 72581 283609 72615
rect 283665 72581 283751 72615
rect 283807 72581 283893 72615
rect 282828 72525 282882 72581
rect 282955 72559 283006 72581
rect 283097 72559 283130 72581
rect 283239 72559 283254 72581
rect 282938 72525 283006 72559
rect 283062 72525 283130 72559
rect 283186 72525 283254 72559
rect 283310 72559 283325 72581
rect 283434 72559 283467 72581
rect 283558 72559 283609 72581
rect 283310 72525 283378 72559
rect 283434 72525 283502 72559
rect 283558 72525 283626 72559
rect 283682 72525 283750 72581
rect 283807 72559 283874 72581
rect 283949 72559 284728 72615
rect 283806 72525 283874 72559
rect 283930 72525 284728 72559
rect 282828 72473 284728 72525
rect 282828 72457 282899 72473
rect 282955 72457 283041 72473
rect 283097 72457 283183 72473
rect 283239 72457 283325 72473
rect 283381 72457 283467 72473
rect 283523 72457 283609 72473
rect 283665 72457 283751 72473
rect 283807 72457 283893 72473
rect 282828 72401 282882 72457
rect 282955 72417 283006 72457
rect 283097 72417 283130 72457
rect 283239 72417 283254 72457
rect 282938 72401 283006 72417
rect 283062 72401 283130 72417
rect 283186 72401 283254 72417
rect 283310 72417 283325 72457
rect 283434 72417 283467 72457
rect 283558 72417 283609 72457
rect 283310 72401 283378 72417
rect 283434 72401 283502 72417
rect 283558 72401 283626 72417
rect 283682 72401 283750 72457
rect 283807 72417 283874 72457
rect 283949 72417 284728 72473
rect 283806 72401 283874 72417
rect 283930 72401 284728 72417
rect 282828 72333 284728 72401
rect 282828 72277 282882 72333
rect 282938 72331 283006 72333
rect 283062 72331 283130 72333
rect 283186 72331 283254 72333
rect 282955 72277 283006 72331
rect 283097 72277 283130 72331
rect 283239 72277 283254 72331
rect 283310 72331 283378 72333
rect 283434 72331 283502 72333
rect 283558 72331 283626 72333
rect 283310 72277 283325 72331
rect 283434 72277 283467 72331
rect 283558 72277 283609 72331
rect 283682 72277 283750 72333
rect 283806 72331 283874 72333
rect 283930 72331 284728 72333
rect 283807 72277 283874 72331
rect 282828 72275 282899 72277
rect 282955 72275 283041 72277
rect 283097 72275 283183 72277
rect 283239 72275 283325 72277
rect 283381 72275 283467 72277
rect 283523 72275 283609 72277
rect 283665 72275 283751 72277
rect 283807 72275 283893 72277
rect 283949 72275 284728 72331
rect 282828 72209 284728 72275
rect 282828 72153 282882 72209
rect 282938 72189 283006 72209
rect 283062 72189 283130 72209
rect 283186 72189 283254 72209
rect 282955 72153 283006 72189
rect 283097 72153 283130 72189
rect 283239 72153 283254 72189
rect 283310 72189 283378 72209
rect 283434 72189 283502 72209
rect 283558 72189 283626 72209
rect 283310 72153 283325 72189
rect 283434 72153 283467 72189
rect 283558 72153 283609 72189
rect 283682 72153 283750 72209
rect 283806 72189 283874 72209
rect 283930 72189 284728 72209
rect 283807 72153 283874 72189
rect 282828 72133 282899 72153
rect 282955 72133 283041 72153
rect 283097 72133 283183 72153
rect 283239 72133 283325 72153
rect 283381 72133 283467 72153
rect 283523 72133 283609 72153
rect 283665 72133 283751 72153
rect 283807 72133 283893 72153
rect 283949 72133 284728 72189
rect 282828 72088 284728 72133
rect 600272 74035 602172 74088
rect 600272 73979 600343 74035
rect 600399 73979 600485 74035
rect 600541 73979 600627 74035
rect 600683 73979 600769 74035
rect 600825 73979 600911 74035
rect 600967 73979 601053 74035
rect 601109 73979 601195 74035
rect 601251 73979 601337 74035
rect 601393 73979 601479 74035
rect 601535 73979 601621 74035
rect 601677 73979 601763 74035
rect 601819 73979 601905 74035
rect 601961 73979 602047 74035
rect 602103 73979 602172 74035
rect 600272 73945 602172 73979
rect 600272 73889 600326 73945
rect 600382 73893 600450 73945
rect 600506 73893 600574 73945
rect 600630 73893 600698 73945
rect 600399 73889 600450 73893
rect 600541 73889 600574 73893
rect 600683 73889 600698 73893
rect 600754 73893 600822 73945
rect 600878 73893 600946 73945
rect 601002 73893 601070 73945
rect 600754 73889 600769 73893
rect 600878 73889 600911 73893
rect 601002 73889 601053 73893
rect 601126 73889 601194 73945
rect 601250 73893 601318 73945
rect 601374 73893 601442 73945
rect 601498 73893 601566 73945
rect 601622 73893 601690 73945
rect 601251 73889 601318 73893
rect 601393 73889 601442 73893
rect 601535 73889 601566 73893
rect 601677 73889 601690 73893
rect 601746 73893 601814 73945
rect 601870 73893 601938 73945
rect 601994 73893 602062 73945
rect 601746 73889 601763 73893
rect 601870 73889 601905 73893
rect 601994 73889 602047 73893
rect 602118 73889 602172 73945
rect 600272 73837 600343 73889
rect 600399 73837 600485 73889
rect 600541 73837 600627 73889
rect 600683 73837 600769 73889
rect 600825 73837 600911 73889
rect 600967 73837 601053 73889
rect 601109 73837 601195 73889
rect 601251 73837 601337 73889
rect 601393 73837 601479 73889
rect 601535 73837 601621 73889
rect 601677 73837 601763 73889
rect 601819 73837 601905 73889
rect 601961 73837 602047 73889
rect 602103 73837 602172 73889
rect 600272 73821 602172 73837
rect 600272 73765 600326 73821
rect 600382 73765 600450 73821
rect 600506 73765 600574 73821
rect 600630 73765 600698 73821
rect 600754 73765 600822 73821
rect 600878 73765 600946 73821
rect 601002 73765 601070 73821
rect 601126 73765 601194 73821
rect 601250 73765 601318 73821
rect 601374 73765 601442 73821
rect 601498 73765 601566 73821
rect 601622 73765 601690 73821
rect 601746 73765 601814 73821
rect 601870 73765 601938 73821
rect 601994 73765 602062 73821
rect 602118 73765 602172 73821
rect 600272 73751 602172 73765
rect 600272 73697 600343 73751
rect 600399 73697 600485 73751
rect 600541 73697 600627 73751
rect 600683 73697 600769 73751
rect 600825 73697 600911 73751
rect 600967 73697 601053 73751
rect 601109 73697 601195 73751
rect 601251 73697 601337 73751
rect 601393 73697 601479 73751
rect 601535 73697 601621 73751
rect 601677 73697 601763 73751
rect 601819 73697 601905 73751
rect 601961 73697 602047 73751
rect 602103 73697 602172 73751
rect 600272 73641 600326 73697
rect 600399 73695 600450 73697
rect 600541 73695 600574 73697
rect 600683 73695 600698 73697
rect 600382 73641 600450 73695
rect 600506 73641 600574 73695
rect 600630 73641 600698 73695
rect 600754 73695 600769 73697
rect 600878 73695 600911 73697
rect 601002 73695 601053 73697
rect 600754 73641 600822 73695
rect 600878 73641 600946 73695
rect 601002 73641 601070 73695
rect 601126 73641 601194 73697
rect 601251 73695 601318 73697
rect 601393 73695 601442 73697
rect 601535 73695 601566 73697
rect 601677 73695 601690 73697
rect 601250 73641 601318 73695
rect 601374 73641 601442 73695
rect 601498 73641 601566 73695
rect 601622 73641 601690 73695
rect 601746 73695 601763 73697
rect 601870 73695 601905 73697
rect 601994 73695 602047 73697
rect 601746 73641 601814 73695
rect 601870 73641 601938 73695
rect 601994 73641 602062 73695
rect 602118 73641 602172 73697
rect 600272 73609 602172 73641
rect 600272 73573 600343 73609
rect 600399 73573 600485 73609
rect 600541 73573 600627 73609
rect 600683 73573 600769 73609
rect 600825 73573 600911 73609
rect 600967 73573 601053 73609
rect 601109 73573 601195 73609
rect 601251 73573 601337 73609
rect 601393 73573 601479 73609
rect 601535 73573 601621 73609
rect 601677 73573 601763 73609
rect 601819 73573 601905 73609
rect 601961 73573 602047 73609
rect 602103 73573 602172 73609
rect 600272 73517 600326 73573
rect 600399 73553 600450 73573
rect 600541 73553 600574 73573
rect 600683 73553 600698 73573
rect 600382 73517 600450 73553
rect 600506 73517 600574 73553
rect 600630 73517 600698 73553
rect 600754 73553 600769 73573
rect 600878 73553 600911 73573
rect 601002 73553 601053 73573
rect 600754 73517 600822 73553
rect 600878 73517 600946 73553
rect 601002 73517 601070 73553
rect 601126 73517 601194 73573
rect 601251 73553 601318 73573
rect 601393 73553 601442 73573
rect 601535 73553 601566 73573
rect 601677 73553 601690 73573
rect 601250 73517 601318 73553
rect 601374 73517 601442 73553
rect 601498 73517 601566 73553
rect 601622 73517 601690 73553
rect 601746 73553 601763 73573
rect 601870 73553 601905 73573
rect 601994 73553 602047 73573
rect 601746 73517 601814 73553
rect 601870 73517 601938 73553
rect 601994 73517 602062 73553
rect 602118 73517 602172 73573
rect 600272 73467 602172 73517
rect 600272 73449 600343 73467
rect 600399 73449 600485 73467
rect 600541 73449 600627 73467
rect 600683 73449 600769 73467
rect 600825 73449 600911 73467
rect 600967 73449 601053 73467
rect 601109 73449 601195 73467
rect 601251 73449 601337 73467
rect 601393 73449 601479 73467
rect 601535 73449 601621 73467
rect 601677 73449 601763 73467
rect 601819 73449 601905 73467
rect 601961 73449 602047 73467
rect 602103 73449 602172 73467
rect 600272 73393 600326 73449
rect 600399 73411 600450 73449
rect 600541 73411 600574 73449
rect 600683 73411 600698 73449
rect 600382 73393 600450 73411
rect 600506 73393 600574 73411
rect 600630 73393 600698 73411
rect 600754 73411 600769 73449
rect 600878 73411 600911 73449
rect 601002 73411 601053 73449
rect 600754 73393 600822 73411
rect 600878 73393 600946 73411
rect 601002 73393 601070 73411
rect 601126 73393 601194 73449
rect 601251 73411 601318 73449
rect 601393 73411 601442 73449
rect 601535 73411 601566 73449
rect 601677 73411 601690 73449
rect 601250 73393 601318 73411
rect 601374 73393 601442 73411
rect 601498 73393 601566 73411
rect 601622 73393 601690 73411
rect 601746 73411 601763 73449
rect 601870 73411 601905 73449
rect 601994 73411 602047 73449
rect 601746 73393 601814 73411
rect 601870 73393 601938 73411
rect 601994 73393 602062 73411
rect 602118 73393 602172 73449
rect 600272 73325 602172 73393
rect 600272 73269 600326 73325
rect 600399 73269 600450 73325
rect 600541 73269 600574 73325
rect 600683 73269 600698 73325
rect 600754 73269 600769 73325
rect 600878 73269 600911 73325
rect 601002 73269 601053 73325
rect 601126 73269 601194 73325
rect 601251 73269 601318 73325
rect 601393 73269 601442 73325
rect 601535 73269 601566 73325
rect 601677 73269 601690 73325
rect 601746 73269 601763 73325
rect 601870 73269 601905 73325
rect 601994 73269 602047 73325
rect 602118 73269 602172 73325
rect 600272 73201 602172 73269
rect 600272 73145 600326 73201
rect 600382 73183 600450 73201
rect 600506 73183 600574 73201
rect 600630 73183 600698 73201
rect 600399 73145 600450 73183
rect 600541 73145 600574 73183
rect 600683 73145 600698 73183
rect 600754 73183 600822 73201
rect 600878 73183 600946 73201
rect 601002 73183 601070 73201
rect 600754 73145 600769 73183
rect 600878 73145 600911 73183
rect 601002 73145 601053 73183
rect 601126 73145 601194 73201
rect 601250 73183 601318 73201
rect 601374 73183 601442 73201
rect 601498 73183 601566 73201
rect 601622 73183 601690 73201
rect 601251 73145 601318 73183
rect 601393 73145 601442 73183
rect 601535 73145 601566 73183
rect 601677 73145 601690 73183
rect 601746 73183 601814 73201
rect 601870 73183 601938 73201
rect 601994 73183 602062 73201
rect 601746 73145 601763 73183
rect 601870 73145 601905 73183
rect 601994 73145 602047 73183
rect 602118 73145 602172 73201
rect 600272 73127 600343 73145
rect 600399 73127 600485 73145
rect 600541 73127 600627 73145
rect 600683 73127 600769 73145
rect 600825 73127 600911 73145
rect 600967 73127 601053 73145
rect 601109 73127 601195 73145
rect 601251 73127 601337 73145
rect 601393 73127 601479 73145
rect 601535 73127 601621 73145
rect 601677 73127 601763 73145
rect 601819 73127 601905 73145
rect 601961 73127 602047 73145
rect 602103 73127 602172 73145
rect 600272 73077 602172 73127
rect 600272 73021 600326 73077
rect 600382 73041 600450 73077
rect 600506 73041 600574 73077
rect 600630 73041 600698 73077
rect 600399 73021 600450 73041
rect 600541 73021 600574 73041
rect 600683 73021 600698 73041
rect 600754 73041 600822 73077
rect 600878 73041 600946 73077
rect 601002 73041 601070 73077
rect 600754 73021 600769 73041
rect 600878 73021 600911 73041
rect 601002 73021 601053 73041
rect 601126 73021 601194 73077
rect 601250 73041 601318 73077
rect 601374 73041 601442 73077
rect 601498 73041 601566 73077
rect 601622 73041 601690 73077
rect 601251 73021 601318 73041
rect 601393 73021 601442 73041
rect 601535 73021 601566 73041
rect 601677 73021 601690 73041
rect 601746 73041 601814 73077
rect 601870 73041 601938 73077
rect 601994 73041 602062 73077
rect 601746 73021 601763 73041
rect 601870 73021 601905 73041
rect 601994 73021 602047 73041
rect 602118 73021 602172 73077
rect 600272 72985 600343 73021
rect 600399 72985 600485 73021
rect 600541 72985 600627 73021
rect 600683 72985 600769 73021
rect 600825 72985 600911 73021
rect 600967 72985 601053 73021
rect 601109 72985 601195 73021
rect 601251 72985 601337 73021
rect 601393 72985 601479 73021
rect 601535 72985 601621 73021
rect 601677 72985 601763 73021
rect 601819 72985 601905 73021
rect 601961 72985 602047 73021
rect 602103 72985 602172 73021
rect 600272 72953 602172 72985
rect 600272 72897 600326 72953
rect 600382 72899 600450 72953
rect 600506 72899 600574 72953
rect 600630 72899 600698 72953
rect 600399 72897 600450 72899
rect 600541 72897 600574 72899
rect 600683 72897 600698 72899
rect 600754 72899 600822 72953
rect 600878 72899 600946 72953
rect 601002 72899 601070 72953
rect 600754 72897 600769 72899
rect 600878 72897 600911 72899
rect 601002 72897 601053 72899
rect 601126 72897 601194 72953
rect 601250 72899 601318 72953
rect 601374 72899 601442 72953
rect 601498 72899 601566 72953
rect 601622 72899 601690 72953
rect 601251 72897 601318 72899
rect 601393 72897 601442 72899
rect 601535 72897 601566 72899
rect 601677 72897 601690 72899
rect 601746 72899 601814 72953
rect 601870 72899 601938 72953
rect 601994 72899 602062 72953
rect 601746 72897 601763 72899
rect 601870 72897 601905 72899
rect 601994 72897 602047 72899
rect 602118 72897 602172 72953
rect 600272 72843 600343 72897
rect 600399 72843 600485 72897
rect 600541 72843 600627 72897
rect 600683 72843 600769 72897
rect 600825 72843 600911 72897
rect 600967 72843 601053 72897
rect 601109 72843 601195 72897
rect 601251 72843 601337 72897
rect 601393 72843 601479 72897
rect 601535 72843 601621 72897
rect 601677 72843 601763 72897
rect 601819 72843 601905 72897
rect 601961 72843 602047 72897
rect 602103 72843 602172 72897
rect 600272 72829 602172 72843
rect 600272 72773 600326 72829
rect 600382 72773 600450 72829
rect 600506 72773 600574 72829
rect 600630 72773 600698 72829
rect 600754 72773 600822 72829
rect 600878 72773 600946 72829
rect 601002 72773 601070 72829
rect 601126 72773 601194 72829
rect 601250 72773 601318 72829
rect 601374 72773 601442 72829
rect 601498 72773 601566 72829
rect 601622 72773 601690 72829
rect 601746 72773 601814 72829
rect 601870 72773 601938 72829
rect 601994 72773 602062 72829
rect 602118 72773 602172 72829
rect 600272 72757 602172 72773
rect 600272 72705 600343 72757
rect 600399 72705 600485 72757
rect 600541 72705 600627 72757
rect 600683 72705 600769 72757
rect 600825 72705 600911 72757
rect 600967 72705 601053 72757
rect 601109 72705 601195 72757
rect 601251 72705 601337 72757
rect 601393 72705 601479 72757
rect 601535 72705 601621 72757
rect 601677 72705 601763 72757
rect 601819 72705 601905 72757
rect 601961 72705 602047 72757
rect 602103 72705 602172 72757
rect 600272 72649 600326 72705
rect 600399 72701 600450 72705
rect 600541 72701 600574 72705
rect 600683 72701 600698 72705
rect 600382 72649 600450 72701
rect 600506 72649 600574 72701
rect 600630 72649 600698 72701
rect 600754 72701 600769 72705
rect 600878 72701 600911 72705
rect 601002 72701 601053 72705
rect 600754 72649 600822 72701
rect 600878 72649 600946 72701
rect 601002 72649 601070 72701
rect 601126 72649 601194 72705
rect 601251 72701 601318 72705
rect 601393 72701 601442 72705
rect 601535 72701 601566 72705
rect 601677 72701 601690 72705
rect 601250 72649 601318 72701
rect 601374 72649 601442 72701
rect 601498 72649 601566 72701
rect 601622 72649 601690 72701
rect 601746 72701 601763 72705
rect 601870 72701 601905 72705
rect 601994 72701 602047 72705
rect 601746 72649 601814 72701
rect 601870 72649 601938 72701
rect 601994 72649 602062 72701
rect 602118 72649 602172 72705
rect 600272 72615 602172 72649
rect 600272 72581 600343 72615
rect 600399 72581 600485 72615
rect 600541 72581 600627 72615
rect 600683 72581 600769 72615
rect 600825 72581 600911 72615
rect 600967 72581 601053 72615
rect 601109 72581 601195 72615
rect 601251 72581 601337 72615
rect 601393 72581 601479 72615
rect 601535 72581 601621 72615
rect 601677 72581 601763 72615
rect 601819 72581 601905 72615
rect 601961 72581 602047 72615
rect 602103 72581 602172 72615
rect 600272 72525 600326 72581
rect 600399 72559 600450 72581
rect 600541 72559 600574 72581
rect 600683 72559 600698 72581
rect 600382 72525 600450 72559
rect 600506 72525 600574 72559
rect 600630 72525 600698 72559
rect 600754 72559 600769 72581
rect 600878 72559 600911 72581
rect 601002 72559 601053 72581
rect 600754 72525 600822 72559
rect 600878 72525 600946 72559
rect 601002 72525 601070 72559
rect 601126 72525 601194 72581
rect 601251 72559 601318 72581
rect 601393 72559 601442 72581
rect 601535 72559 601566 72581
rect 601677 72559 601690 72581
rect 601250 72525 601318 72559
rect 601374 72525 601442 72559
rect 601498 72525 601566 72559
rect 601622 72525 601690 72559
rect 601746 72559 601763 72581
rect 601870 72559 601905 72581
rect 601994 72559 602047 72581
rect 601746 72525 601814 72559
rect 601870 72525 601938 72559
rect 601994 72525 602062 72559
rect 602118 72525 602172 72581
rect 600272 72473 602172 72525
rect 600272 72457 600343 72473
rect 600399 72457 600485 72473
rect 600541 72457 600627 72473
rect 600683 72457 600769 72473
rect 600825 72457 600911 72473
rect 600967 72457 601053 72473
rect 601109 72457 601195 72473
rect 601251 72457 601337 72473
rect 601393 72457 601479 72473
rect 601535 72457 601621 72473
rect 601677 72457 601763 72473
rect 601819 72457 601905 72473
rect 601961 72457 602047 72473
rect 602103 72457 602172 72473
rect 600272 72401 600326 72457
rect 600399 72417 600450 72457
rect 600541 72417 600574 72457
rect 600683 72417 600698 72457
rect 600382 72401 600450 72417
rect 600506 72401 600574 72417
rect 600630 72401 600698 72417
rect 600754 72417 600769 72457
rect 600878 72417 600911 72457
rect 601002 72417 601053 72457
rect 600754 72401 600822 72417
rect 600878 72401 600946 72417
rect 601002 72401 601070 72417
rect 601126 72401 601194 72457
rect 601251 72417 601318 72457
rect 601393 72417 601442 72457
rect 601535 72417 601566 72457
rect 601677 72417 601690 72457
rect 601250 72401 601318 72417
rect 601374 72401 601442 72417
rect 601498 72401 601566 72417
rect 601622 72401 601690 72417
rect 601746 72417 601763 72457
rect 601870 72417 601905 72457
rect 601994 72417 602047 72457
rect 601746 72401 601814 72417
rect 601870 72401 601938 72417
rect 601994 72401 602062 72417
rect 602118 72401 602172 72457
rect 600272 72333 602172 72401
rect 600272 72277 600326 72333
rect 600382 72331 600450 72333
rect 600506 72331 600574 72333
rect 600630 72331 600698 72333
rect 600399 72277 600450 72331
rect 600541 72277 600574 72331
rect 600683 72277 600698 72331
rect 600754 72331 600822 72333
rect 600878 72331 600946 72333
rect 601002 72331 601070 72333
rect 600754 72277 600769 72331
rect 600878 72277 600911 72331
rect 601002 72277 601053 72331
rect 601126 72277 601194 72333
rect 601250 72331 601318 72333
rect 601374 72331 601442 72333
rect 601498 72331 601566 72333
rect 601622 72331 601690 72333
rect 601251 72277 601318 72331
rect 601393 72277 601442 72331
rect 601535 72277 601566 72331
rect 601677 72277 601690 72331
rect 601746 72331 601814 72333
rect 601870 72331 601938 72333
rect 601994 72331 602062 72333
rect 601746 72277 601763 72331
rect 601870 72277 601905 72331
rect 601994 72277 602047 72331
rect 602118 72277 602172 72333
rect 600272 72275 600343 72277
rect 600399 72275 600485 72277
rect 600541 72275 600627 72277
rect 600683 72275 600769 72277
rect 600825 72275 600911 72277
rect 600967 72275 601053 72277
rect 601109 72275 601195 72277
rect 601251 72275 601337 72277
rect 601393 72275 601479 72277
rect 601535 72275 601621 72277
rect 601677 72275 601763 72277
rect 601819 72275 601905 72277
rect 601961 72275 602047 72277
rect 602103 72275 602172 72277
rect 600272 72209 602172 72275
rect 600272 72153 600326 72209
rect 600382 72189 600450 72209
rect 600506 72189 600574 72209
rect 600630 72189 600698 72209
rect 600399 72153 600450 72189
rect 600541 72153 600574 72189
rect 600683 72153 600698 72189
rect 600754 72189 600822 72209
rect 600878 72189 600946 72209
rect 601002 72189 601070 72209
rect 600754 72153 600769 72189
rect 600878 72153 600911 72189
rect 601002 72153 601053 72189
rect 601126 72153 601194 72209
rect 601250 72189 601318 72209
rect 601374 72189 601442 72209
rect 601498 72189 601566 72209
rect 601622 72189 601690 72209
rect 601251 72153 601318 72189
rect 601393 72153 601442 72189
rect 601535 72153 601566 72189
rect 601677 72153 601690 72189
rect 601746 72189 601814 72209
rect 601870 72189 601938 72209
rect 601994 72189 602062 72209
rect 601746 72153 601763 72189
rect 601870 72153 601905 72189
rect 601994 72153 602047 72189
rect 602118 72153 602172 72209
rect 600272 72133 600343 72153
rect 600399 72133 600485 72153
rect 600541 72133 600627 72153
rect 600683 72133 600769 72153
rect 600825 72133 600911 72153
rect 600967 72133 601053 72153
rect 601109 72133 601195 72153
rect 601251 72133 601337 72153
rect 601393 72133 601479 72153
rect 601535 72133 601621 72153
rect 601677 72133 601763 72153
rect 601819 72133 601905 72153
rect 601961 72133 602047 72153
rect 602103 72133 602172 72153
rect 600272 72088 602172 72133
rect 602752 74035 604802 74088
rect 602752 73979 602823 74035
rect 602879 73979 602965 74035
rect 603021 73979 603107 74035
rect 603163 73979 603249 74035
rect 603305 73979 603391 74035
rect 603447 73979 603533 74035
rect 603589 73979 603675 74035
rect 603731 73979 603817 74035
rect 603873 73979 603959 74035
rect 604015 73979 604802 74035
rect 602752 73945 604802 73979
rect 602752 73889 602806 73945
rect 602862 73893 602930 73945
rect 602986 73893 603054 73945
rect 603110 73893 603178 73945
rect 602879 73889 602930 73893
rect 603021 73889 603054 73893
rect 603163 73889 603178 73893
rect 603234 73893 603302 73945
rect 603358 73893 603426 73945
rect 603482 73893 603550 73945
rect 603234 73889 603249 73893
rect 603358 73889 603391 73893
rect 603482 73889 603533 73893
rect 603606 73889 603674 73945
rect 603730 73893 603798 73945
rect 603854 73893 603922 73945
rect 603978 73893 604802 73945
rect 603731 73889 603798 73893
rect 603873 73889 603922 73893
rect 602752 73837 602823 73889
rect 602879 73837 602965 73889
rect 603021 73837 603107 73889
rect 603163 73837 603249 73889
rect 603305 73837 603391 73889
rect 603447 73837 603533 73889
rect 603589 73837 603675 73889
rect 603731 73837 603817 73889
rect 603873 73837 603959 73889
rect 604015 73837 604802 73893
rect 602752 73821 604802 73837
rect 602752 73765 602806 73821
rect 602862 73765 602930 73821
rect 602986 73765 603054 73821
rect 603110 73765 603178 73821
rect 603234 73765 603302 73821
rect 603358 73765 603426 73821
rect 603482 73765 603550 73821
rect 603606 73765 603674 73821
rect 603730 73765 603798 73821
rect 603854 73765 603922 73821
rect 603978 73765 604802 73821
rect 602752 73751 604802 73765
rect 602752 73697 602823 73751
rect 602879 73697 602965 73751
rect 603021 73697 603107 73751
rect 603163 73697 603249 73751
rect 603305 73697 603391 73751
rect 603447 73697 603533 73751
rect 603589 73697 603675 73751
rect 603731 73697 603817 73751
rect 603873 73697 603959 73751
rect 602752 73641 602806 73697
rect 602879 73695 602930 73697
rect 603021 73695 603054 73697
rect 603163 73695 603178 73697
rect 602862 73641 602930 73695
rect 602986 73641 603054 73695
rect 603110 73641 603178 73695
rect 603234 73695 603249 73697
rect 603358 73695 603391 73697
rect 603482 73695 603533 73697
rect 603234 73641 603302 73695
rect 603358 73641 603426 73695
rect 603482 73641 603550 73695
rect 603606 73641 603674 73697
rect 603731 73695 603798 73697
rect 603873 73695 603922 73697
rect 604015 73695 604802 73751
rect 603730 73641 603798 73695
rect 603854 73641 603922 73695
rect 603978 73641 604802 73695
rect 602752 73609 604802 73641
rect 602752 73573 602823 73609
rect 602879 73573 602965 73609
rect 603021 73573 603107 73609
rect 603163 73573 603249 73609
rect 603305 73573 603391 73609
rect 603447 73573 603533 73609
rect 603589 73573 603675 73609
rect 603731 73573 603817 73609
rect 603873 73573 603959 73609
rect 602752 73517 602806 73573
rect 602879 73553 602930 73573
rect 603021 73553 603054 73573
rect 603163 73553 603178 73573
rect 602862 73517 602930 73553
rect 602986 73517 603054 73553
rect 603110 73517 603178 73553
rect 603234 73553 603249 73573
rect 603358 73553 603391 73573
rect 603482 73553 603533 73573
rect 603234 73517 603302 73553
rect 603358 73517 603426 73553
rect 603482 73517 603550 73553
rect 603606 73517 603674 73573
rect 603731 73553 603798 73573
rect 603873 73553 603922 73573
rect 604015 73553 604802 73609
rect 603730 73517 603798 73553
rect 603854 73517 603922 73553
rect 603978 73517 604802 73553
rect 602752 73467 604802 73517
rect 602752 73449 602823 73467
rect 602879 73449 602965 73467
rect 603021 73449 603107 73467
rect 603163 73449 603249 73467
rect 603305 73449 603391 73467
rect 603447 73449 603533 73467
rect 603589 73449 603675 73467
rect 603731 73449 603817 73467
rect 603873 73449 603959 73467
rect 602752 73393 602806 73449
rect 602879 73411 602930 73449
rect 603021 73411 603054 73449
rect 603163 73411 603178 73449
rect 602862 73393 602930 73411
rect 602986 73393 603054 73411
rect 603110 73393 603178 73411
rect 603234 73411 603249 73449
rect 603358 73411 603391 73449
rect 603482 73411 603533 73449
rect 603234 73393 603302 73411
rect 603358 73393 603426 73411
rect 603482 73393 603550 73411
rect 603606 73393 603674 73449
rect 603731 73411 603798 73449
rect 603873 73411 603922 73449
rect 604015 73411 604802 73467
rect 603730 73393 603798 73411
rect 603854 73393 603922 73411
rect 603978 73393 604802 73411
rect 602752 73325 604802 73393
rect 602752 73269 602806 73325
rect 602879 73269 602930 73325
rect 603021 73269 603054 73325
rect 603163 73269 603178 73325
rect 603234 73269 603249 73325
rect 603358 73269 603391 73325
rect 603482 73269 603533 73325
rect 603606 73269 603674 73325
rect 603731 73269 603798 73325
rect 603873 73269 603922 73325
rect 604015 73269 604802 73325
rect 602752 73201 604802 73269
rect 602752 73145 602806 73201
rect 602862 73183 602930 73201
rect 602986 73183 603054 73201
rect 603110 73183 603178 73201
rect 602879 73145 602930 73183
rect 603021 73145 603054 73183
rect 603163 73145 603178 73183
rect 603234 73183 603302 73201
rect 603358 73183 603426 73201
rect 603482 73183 603550 73201
rect 603234 73145 603249 73183
rect 603358 73145 603391 73183
rect 603482 73145 603533 73183
rect 603606 73145 603674 73201
rect 603730 73183 603798 73201
rect 603854 73183 603922 73201
rect 603978 73183 604802 73201
rect 603731 73145 603798 73183
rect 603873 73145 603922 73183
rect 602752 73127 602823 73145
rect 602879 73127 602965 73145
rect 603021 73127 603107 73145
rect 603163 73127 603249 73145
rect 603305 73127 603391 73145
rect 603447 73127 603533 73145
rect 603589 73127 603675 73145
rect 603731 73127 603817 73145
rect 603873 73127 603959 73145
rect 604015 73127 604802 73183
rect 602752 73077 604802 73127
rect 602752 73021 602806 73077
rect 602862 73041 602930 73077
rect 602986 73041 603054 73077
rect 603110 73041 603178 73077
rect 602879 73021 602930 73041
rect 603021 73021 603054 73041
rect 603163 73021 603178 73041
rect 603234 73041 603302 73077
rect 603358 73041 603426 73077
rect 603482 73041 603550 73077
rect 603234 73021 603249 73041
rect 603358 73021 603391 73041
rect 603482 73021 603533 73041
rect 603606 73021 603674 73077
rect 603730 73041 603798 73077
rect 603854 73041 603922 73077
rect 603978 73041 604802 73077
rect 603731 73021 603798 73041
rect 603873 73021 603922 73041
rect 602752 72985 602823 73021
rect 602879 72985 602965 73021
rect 603021 72985 603107 73021
rect 603163 72985 603249 73021
rect 603305 72985 603391 73021
rect 603447 72985 603533 73021
rect 603589 72985 603675 73021
rect 603731 72985 603817 73021
rect 603873 72985 603959 73021
rect 604015 72985 604802 73041
rect 602752 72953 604802 72985
rect 602752 72897 602806 72953
rect 602862 72899 602930 72953
rect 602986 72899 603054 72953
rect 603110 72899 603178 72953
rect 602879 72897 602930 72899
rect 603021 72897 603054 72899
rect 603163 72897 603178 72899
rect 603234 72899 603302 72953
rect 603358 72899 603426 72953
rect 603482 72899 603550 72953
rect 603234 72897 603249 72899
rect 603358 72897 603391 72899
rect 603482 72897 603533 72899
rect 603606 72897 603674 72953
rect 603730 72899 603798 72953
rect 603854 72899 603922 72953
rect 603978 72899 604802 72953
rect 603731 72897 603798 72899
rect 603873 72897 603922 72899
rect 602752 72843 602823 72897
rect 602879 72843 602965 72897
rect 603021 72843 603107 72897
rect 603163 72843 603249 72897
rect 603305 72843 603391 72897
rect 603447 72843 603533 72897
rect 603589 72843 603675 72897
rect 603731 72843 603817 72897
rect 603873 72843 603959 72897
rect 604015 72843 604802 72899
rect 602752 72829 604802 72843
rect 602752 72773 602806 72829
rect 602862 72773 602930 72829
rect 602986 72773 603054 72829
rect 603110 72773 603178 72829
rect 603234 72773 603302 72829
rect 603358 72773 603426 72829
rect 603482 72773 603550 72829
rect 603606 72773 603674 72829
rect 603730 72773 603798 72829
rect 603854 72773 603922 72829
rect 603978 72773 604802 72829
rect 602752 72757 604802 72773
rect 602752 72705 602823 72757
rect 602879 72705 602965 72757
rect 603021 72705 603107 72757
rect 603163 72705 603249 72757
rect 603305 72705 603391 72757
rect 603447 72705 603533 72757
rect 603589 72705 603675 72757
rect 603731 72705 603817 72757
rect 603873 72705 603959 72757
rect 602752 72649 602806 72705
rect 602879 72701 602930 72705
rect 603021 72701 603054 72705
rect 603163 72701 603178 72705
rect 602862 72649 602930 72701
rect 602986 72649 603054 72701
rect 603110 72649 603178 72701
rect 603234 72701 603249 72705
rect 603358 72701 603391 72705
rect 603482 72701 603533 72705
rect 603234 72649 603302 72701
rect 603358 72649 603426 72701
rect 603482 72649 603550 72701
rect 603606 72649 603674 72705
rect 603731 72701 603798 72705
rect 603873 72701 603922 72705
rect 604015 72701 604802 72757
rect 603730 72649 603798 72701
rect 603854 72649 603922 72701
rect 603978 72649 604802 72701
rect 602752 72615 604802 72649
rect 602752 72581 602823 72615
rect 602879 72581 602965 72615
rect 603021 72581 603107 72615
rect 603163 72581 603249 72615
rect 603305 72581 603391 72615
rect 603447 72581 603533 72615
rect 603589 72581 603675 72615
rect 603731 72581 603817 72615
rect 603873 72581 603959 72615
rect 602752 72525 602806 72581
rect 602879 72559 602930 72581
rect 603021 72559 603054 72581
rect 603163 72559 603178 72581
rect 602862 72525 602930 72559
rect 602986 72525 603054 72559
rect 603110 72525 603178 72559
rect 603234 72559 603249 72581
rect 603358 72559 603391 72581
rect 603482 72559 603533 72581
rect 603234 72525 603302 72559
rect 603358 72525 603426 72559
rect 603482 72525 603550 72559
rect 603606 72525 603674 72581
rect 603731 72559 603798 72581
rect 603873 72559 603922 72581
rect 604015 72559 604802 72615
rect 603730 72525 603798 72559
rect 603854 72525 603922 72559
rect 603978 72525 604802 72559
rect 602752 72473 604802 72525
rect 602752 72457 602823 72473
rect 602879 72457 602965 72473
rect 603021 72457 603107 72473
rect 603163 72457 603249 72473
rect 603305 72457 603391 72473
rect 603447 72457 603533 72473
rect 603589 72457 603675 72473
rect 603731 72457 603817 72473
rect 603873 72457 603959 72473
rect 602752 72401 602806 72457
rect 602879 72417 602930 72457
rect 603021 72417 603054 72457
rect 603163 72417 603178 72457
rect 602862 72401 602930 72417
rect 602986 72401 603054 72417
rect 603110 72401 603178 72417
rect 603234 72417 603249 72457
rect 603358 72417 603391 72457
rect 603482 72417 603533 72457
rect 603234 72401 603302 72417
rect 603358 72401 603426 72417
rect 603482 72401 603550 72417
rect 603606 72401 603674 72457
rect 603731 72417 603798 72457
rect 603873 72417 603922 72457
rect 604015 72417 604802 72473
rect 603730 72401 603798 72417
rect 603854 72401 603922 72417
rect 603978 72401 604802 72417
rect 602752 72333 604802 72401
rect 602752 72277 602806 72333
rect 602862 72331 602930 72333
rect 602986 72331 603054 72333
rect 603110 72331 603178 72333
rect 602879 72277 602930 72331
rect 603021 72277 603054 72331
rect 603163 72277 603178 72331
rect 603234 72331 603302 72333
rect 603358 72331 603426 72333
rect 603482 72331 603550 72333
rect 603234 72277 603249 72331
rect 603358 72277 603391 72331
rect 603482 72277 603533 72331
rect 603606 72277 603674 72333
rect 603730 72331 603798 72333
rect 603854 72331 603922 72333
rect 603978 72331 604802 72333
rect 603731 72277 603798 72331
rect 603873 72277 603922 72331
rect 602752 72275 602823 72277
rect 602879 72275 602965 72277
rect 603021 72275 603107 72277
rect 603163 72275 603249 72277
rect 603305 72275 603391 72277
rect 603447 72275 603533 72277
rect 603589 72275 603675 72277
rect 603731 72275 603817 72277
rect 603873 72275 603959 72277
rect 604015 72275 604802 72331
rect 602752 72209 604802 72275
rect 602752 72153 602806 72209
rect 602862 72189 602930 72209
rect 602986 72189 603054 72209
rect 603110 72189 603178 72209
rect 602879 72153 602930 72189
rect 603021 72153 603054 72189
rect 603163 72153 603178 72189
rect 603234 72189 603302 72209
rect 603358 72189 603426 72209
rect 603482 72189 603550 72209
rect 603234 72153 603249 72189
rect 603358 72153 603391 72189
rect 603482 72153 603533 72189
rect 603606 72153 603674 72209
rect 603730 72189 603798 72209
rect 603854 72189 603922 72209
rect 603978 72189 604802 72209
rect 603731 72153 603798 72189
rect 603873 72153 603922 72189
rect 602752 72133 602823 72153
rect 602879 72133 602965 72153
rect 603021 72133 603107 72153
rect 603163 72133 603249 72153
rect 603305 72133 603391 72153
rect 603447 72133 603533 72153
rect 603589 72133 603675 72153
rect 603731 72133 603817 72153
rect 603873 72133 603959 72153
rect 604015 72133 604802 72189
rect 602752 72088 604802 72133
rect 605122 74035 607172 74088
rect 605122 73979 605193 74035
rect 605249 73979 605335 74035
rect 605391 73979 605477 74035
rect 605533 73979 605619 74035
rect 605675 73979 605761 74035
rect 605817 73979 605903 74035
rect 605959 73979 606045 74035
rect 606101 73979 606187 74035
rect 606243 73979 606329 74035
rect 606385 73979 606471 74035
rect 606527 73979 606613 74035
rect 606669 73979 606755 74035
rect 606811 73979 606897 74035
rect 606953 73979 607039 74035
rect 607095 73979 607172 74035
rect 605122 73945 607172 73979
rect 605122 73889 605176 73945
rect 605232 73893 605300 73945
rect 605356 73893 605424 73945
rect 605480 73893 605548 73945
rect 605249 73889 605300 73893
rect 605391 73889 605424 73893
rect 605533 73889 605548 73893
rect 605604 73893 605672 73945
rect 605728 73893 605796 73945
rect 605852 73893 605920 73945
rect 605604 73889 605619 73893
rect 605728 73889 605761 73893
rect 605852 73889 605903 73893
rect 605976 73889 606044 73945
rect 606100 73893 606168 73945
rect 606224 73893 606292 73945
rect 606348 73893 606416 73945
rect 606472 73893 606540 73945
rect 606101 73889 606168 73893
rect 606243 73889 606292 73893
rect 606385 73889 606416 73893
rect 606527 73889 606540 73893
rect 606596 73893 606664 73945
rect 606720 73893 606788 73945
rect 606844 73893 606912 73945
rect 606596 73889 606613 73893
rect 606720 73889 606755 73893
rect 606844 73889 606897 73893
rect 606968 73889 607036 73945
rect 607092 73893 607172 73945
rect 605122 73837 605193 73889
rect 605249 73837 605335 73889
rect 605391 73837 605477 73889
rect 605533 73837 605619 73889
rect 605675 73837 605761 73889
rect 605817 73837 605903 73889
rect 605959 73837 606045 73889
rect 606101 73837 606187 73889
rect 606243 73837 606329 73889
rect 606385 73837 606471 73889
rect 606527 73837 606613 73889
rect 606669 73837 606755 73889
rect 606811 73837 606897 73889
rect 606953 73837 607039 73889
rect 607095 73837 607172 73893
rect 605122 73821 607172 73837
rect 605122 73765 605176 73821
rect 605232 73765 605300 73821
rect 605356 73765 605424 73821
rect 605480 73765 605548 73821
rect 605604 73765 605672 73821
rect 605728 73765 605796 73821
rect 605852 73765 605920 73821
rect 605976 73765 606044 73821
rect 606100 73765 606168 73821
rect 606224 73765 606292 73821
rect 606348 73765 606416 73821
rect 606472 73765 606540 73821
rect 606596 73765 606664 73821
rect 606720 73765 606788 73821
rect 606844 73765 606912 73821
rect 606968 73765 607036 73821
rect 607092 73765 607172 73821
rect 605122 73751 607172 73765
rect 605122 73697 605193 73751
rect 605249 73697 605335 73751
rect 605391 73697 605477 73751
rect 605533 73697 605619 73751
rect 605675 73697 605761 73751
rect 605817 73697 605903 73751
rect 605959 73697 606045 73751
rect 606101 73697 606187 73751
rect 606243 73697 606329 73751
rect 606385 73697 606471 73751
rect 606527 73697 606613 73751
rect 606669 73697 606755 73751
rect 606811 73697 606897 73751
rect 606953 73697 607039 73751
rect 605122 73641 605176 73697
rect 605249 73695 605300 73697
rect 605391 73695 605424 73697
rect 605533 73695 605548 73697
rect 605232 73641 605300 73695
rect 605356 73641 605424 73695
rect 605480 73641 605548 73695
rect 605604 73695 605619 73697
rect 605728 73695 605761 73697
rect 605852 73695 605903 73697
rect 605604 73641 605672 73695
rect 605728 73641 605796 73695
rect 605852 73641 605920 73695
rect 605976 73641 606044 73697
rect 606101 73695 606168 73697
rect 606243 73695 606292 73697
rect 606385 73695 606416 73697
rect 606527 73695 606540 73697
rect 606100 73641 606168 73695
rect 606224 73641 606292 73695
rect 606348 73641 606416 73695
rect 606472 73641 606540 73695
rect 606596 73695 606613 73697
rect 606720 73695 606755 73697
rect 606844 73695 606897 73697
rect 606596 73641 606664 73695
rect 606720 73641 606788 73695
rect 606844 73641 606912 73695
rect 606968 73641 607036 73697
rect 607095 73695 607172 73751
rect 607092 73641 607172 73695
rect 605122 73609 607172 73641
rect 605122 73573 605193 73609
rect 605249 73573 605335 73609
rect 605391 73573 605477 73609
rect 605533 73573 605619 73609
rect 605675 73573 605761 73609
rect 605817 73573 605903 73609
rect 605959 73573 606045 73609
rect 606101 73573 606187 73609
rect 606243 73573 606329 73609
rect 606385 73573 606471 73609
rect 606527 73573 606613 73609
rect 606669 73573 606755 73609
rect 606811 73573 606897 73609
rect 606953 73573 607039 73609
rect 605122 73517 605176 73573
rect 605249 73553 605300 73573
rect 605391 73553 605424 73573
rect 605533 73553 605548 73573
rect 605232 73517 605300 73553
rect 605356 73517 605424 73553
rect 605480 73517 605548 73553
rect 605604 73553 605619 73573
rect 605728 73553 605761 73573
rect 605852 73553 605903 73573
rect 605604 73517 605672 73553
rect 605728 73517 605796 73553
rect 605852 73517 605920 73553
rect 605976 73517 606044 73573
rect 606101 73553 606168 73573
rect 606243 73553 606292 73573
rect 606385 73553 606416 73573
rect 606527 73553 606540 73573
rect 606100 73517 606168 73553
rect 606224 73517 606292 73553
rect 606348 73517 606416 73553
rect 606472 73517 606540 73553
rect 606596 73553 606613 73573
rect 606720 73553 606755 73573
rect 606844 73553 606897 73573
rect 606596 73517 606664 73553
rect 606720 73517 606788 73553
rect 606844 73517 606912 73553
rect 606968 73517 607036 73573
rect 607095 73553 607172 73609
rect 607092 73517 607172 73553
rect 605122 73467 607172 73517
rect 605122 73449 605193 73467
rect 605249 73449 605335 73467
rect 605391 73449 605477 73467
rect 605533 73449 605619 73467
rect 605675 73449 605761 73467
rect 605817 73449 605903 73467
rect 605959 73449 606045 73467
rect 606101 73449 606187 73467
rect 606243 73449 606329 73467
rect 606385 73449 606471 73467
rect 606527 73449 606613 73467
rect 606669 73449 606755 73467
rect 606811 73449 606897 73467
rect 606953 73449 607039 73467
rect 605122 73393 605176 73449
rect 605249 73411 605300 73449
rect 605391 73411 605424 73449
rect 605533 73411 605548 73449
rect 605232 73393 605300 73411
rect 605356 73393 605424 73411
rect 605480 73393 605548 73411
rect 605604 73411 605619 73449
rect 605728 73411 605761 73449
rect 605852 73411 605903 73449
rect 605604 73393 605672 73411
rect 605728 73393 605796 73411
rect 605852 73393 605920 73411
rect 605976 73393 606044 73449
rect 606101 73411 606168 73449
rect 606243 73411 606292 73449
rect 606385 73411 606416 73449
rect 606527 73411 606540 73449
rect 606100 73393 606168 73411
rect 606224 73393 606292 73411
rect 606348 73393 606416 73411
rect 606472 73393 606540 73411
rect 606596 73411 606613 73449
rect 606720 73411 606755 73449
rect 606844 73411 606897 73449
rect 606596 73393 606664 73411
rect 606720 73393 606788 73411
rect 606844 73393 606912 73411
rect 606968 73393 607036 73449
rect 607095 73411 607172 73467
rect 607092 73393 607172 73411
rect 605122 73325 607172 73393
rect 605122 73269 605176 73325
rect 605249 73269 605300 73325
rect 605391 73269 605424 73325
rect 605533 73269 605548 73325
rect 605604 73269 605619 73325
rect 605728 73269 605761 73325
rect 605852 73269 605903 73325
rect 605976 73269 606044 73325
rect 606101 73269 606168 73325
rect 606243 73269 606292 73325
rect 606385 73269 606416 73325
rect 606527 73269 606540 73325
rect 606596 73269 606613 73325
rect 606720 73269 606755 73325
rect 606844 73269 606897 73325
rect 606968 73269 607036 73325
rect 607095 73269 607172 73325
rect 605122 73201 607172 73269
rect 605122 73145 605176 73201
rect 605232 73183 605300 73201
rect 605356 73183 605424 73201
rect 605480 73183 605548 73201
rect 605249 73145 605300 73183
rect 605391 73145 605424 73183
rect 605533 73145 605548 73183
rect 605604 73183 605672 73201
rect 605728 73183 605796 73201
rect 605852 73183 605920 73201
rect 605604 73145 605619 73183
rect 605728 73145 605761 73183
rect 605852 73145 605903 73183
rect 605976 73145 606044 73201
rect 606100 73183 606168 73201
rect 606224 73183 606292 73201
rect 606348 73183 606416 73201
rect 606472 73183 606540 73201
rect 606101 73145 606168 73183
rect 606243 73145 606292 73183
rect 606385 73145 606416 73183
rect 606527 73145 606540 73183
rect 606596 73183 606664 73201
rect 606720 73183 606788 73201
rect 606844 73183 606912 73201
rect 606596 73145 606613 73183
rect 606720 73145 606755 73183
rect 606844 73145 606897 73183
rect 606968 73145 607036 73201
rect 607092 73183 607172 73201
rect 605122 73127 605193 73145
rect 605249 73127 605335 73145
rect 605391 73127 605477 73145
rect 605533 73127 605619 73145
rect 605675 73127 605761 73145
rect 605817 73127 605903 73145
rect 605959 73127 606045 73145
rect 606101 73127 606187 73145
rect 606243 73127 606329 73145
rect 606385 73127 606471 73145
rect 606527 73127 606613 73145
rect 606669 73127 606755 73145
rect 606811 73127 606897 73145
rect 606953 73127 607039 73145
rect 607095 73127 607172 73183
rect 605122 73077 607172 73127
rect 605122 73021 605176 73077
rect 605232 73041 605300 73077
rect 605356 73041 605424 73077
rect 605480 73041 605548 73077
rect 605249 73021 605300 73041
rect 605391 73021 605424 73041
rect 605533 73021 605548 73041
rect 605604 73041 605672 73077
rect 605728 73041 605796 73077
rect 605852 73041 605920 73077
rect 605604 73021 605619 73041
rect 605728 73021 605761 73041
rect 605852 73021 605903 73041
rect 605976 73021 606044 73077
rect 606100 73041 606168 73077
rect 606224 73041 606292 73077
rect 606348 73041 606416 73077
rect 606472 73041 606540 73077
rect 606101 73021 606168 73041
rect 606243 73021 606292 73041
rect 606385 73021 606416 73041
rect 606527 73021 606540 73041
rect 606596 73041 606664 73077
rect 606720 73041 606788 73077
rect 606844 73041 606912 73077
rect 606596 73021 606613 73041
rect 606720 73021 606755 73041
rect 606844 73021 606897 73041
rect 606968 73021 607036 73077
rect 607092 73041 607172 73077
rect 605122 72985 605193 73021
rect 605249 72985 605335 73021
rect 605391 72985 605477 73021
rect 605533 72985 605619 73021
rect 605675 72985 605761 73021
rect 605817 72985 605903 73021
rect 605959 72985 606045 73021
rect 606101 72985 606187 73021
rect 606243 72985 606329 73021
rect 606385 72985 606471 73021
rect 606527 72985 606613 73021
rect 606669 72985 606755 73021
rect 606811 72985 606897 73021
rect 606953 72985 607039 73021
rect 607095 72985 607172 73041
rect 605122 72953 607172 72985
rect 605122 72897 605176 72953
rect 605232 72899 605300 72953
rect 605356 72899 605424 72953
rect 605480 72899 605548 72953
rect 605249 72897 605300 72899
rect 605391 72897 605424 72899
rect 605533 72897 605548 72899
rect 605604 72899 605672 72953
rect 605728 72899 605796 72953
rect 605852 72899 605920 72953
rect 605604 72897 605619 72899
rect 605728 72897 605761 72899
rect 605852 72897 605903 72899
rect 605976 72897 606044 72953
rect 606100 72899 606168 72953
rect 606224 72899 606292 72953
rect 606348 72899 606416 72953
rect 606472 72899 606540 72953
rect 606101 72897 606168 72899
rect 606243 72897 606292 72899
rect 606385 72897 606416 72899
rect 606527 72897 606540 72899
rect 606596 72899 606664 72953
rect 606720 72899 606788 72953
rect 606844 72899 606912 72953
rect 606596 72897 606613 72899
rect 606720 72897 606755 72899
rect 606844 72897 606897 72899
rect 606968 72897 607036 72953
rect 607092 72899 607172 72953
rect 605122 72843 605193 72897
rect 605249 72843 605335 72897
rect 605391 72843 605477 72897
rect 605533 72843 605619 72897
rect 605675 72843 605761 72897
rect 605817 72843 605903 72897
rect 605959 72843 606045 72897
rect 606101 72843 606187 72897
rect 606243 72843 606329 72897
rect 606385 72843 606471 72897
rect 606527 72843 606613 72897
rect 606669 72843 606755 72897
rect 606811 72843 606897 72897
rect 606953 72843 607039 72897
rect 607095 72843 607172 72899
rect 605122 72829 607172 72843
rect 605122 72773 605176 72829
rect 605232 72773 605300 72829
rect 605356 72773 605424 72829
rect 605480 72773 605548 72829
rect 605604 72773 605672 72829
rect 605728 72773 605796 72829
rect 605852 72773 605920 72829
rect 605976 72773 606044 72829
rect 606100 72773 606168 72829
rect 606224 72773 606292 72829
rect 606348 72773 606416 72829
rect 606472 72773 606540 72829
rect 606596 72773 606664 72829
rect 606720 72773 606788 72829
rect 606844 72773 606912 72829
rect 606968 72773 607036 72829
rect 607092 72773 607172 72829
rect 605122 72757 607172 72773
rect 605122 72705 605193 72757
rect 605249 72705 605335 72757
rect 605391 72705 605477 72757
rect 605533 72705 605619 72757
rect 605675 72705 605761 72757
rect 605817 72705 605903 72757
rect 605959 72705 606045 72757
rect 606101 72705 606187 72757
rect 606243 72705 606329 72757
rect 606385 72705 606471 72757
rect 606527 72705 606613 72757
rect 606669 72705 606755 72757
rect 606811 72705 606897 72757
rect 606953 72705 607039 72757
rect 605122 72649 605176 72705
rect 605249 72701 605300 72705
rect 605391 72701 605424 72705
rect 605533 72701 605548 72705
rect 605232 72649 605300 72701
rect 605356 72649 605424 72701
rect 605480 72649 605548 72701
rect 605604 72701 605619 72705
rect 605728 72701 605761 72705
rect 605852 72701 605903 72705
rect 605604 72649 605672 72701
rect 605728 72649 605796 72701
rect 605852 72649 605920 72701
rect 605976 72649 606044 72705
rect 606101 72701 606168 72705
rect 606243 72701 606292 72705
rect 606385 72701 606416 72705
rect 606527 72701 606540 72705
rect 606100 72649 606168 72701
rect 606224 72649 606292 72701
rect 606348 72649 606416 72701
rect 606472 72649 606540 72701
rect 606596 72701 606613 72705
rect 606720 72701 606755 72705
rect 606844 72701 606897 72705
rect 606596 72649 606664 72701
rect 606720 72649 606788 72701
rect 606844 72649 606912 72701
rect 606968 72649 607036 72705
rect 607095 72701 607172 72757
rect 607092 72649 607172 72701
rect 605122 72615 607172 72649
rect 605122 72581 605193 72615
rect 605249 72581 605335 72615
rect 605391 72581 605477 72615
rect 605533 72581 605619 72615
rect 605675 72581 605761 72615
rect 605817 72581 605903 72615
rect 605959 72581 606045 72615
rect 606101 72581 606187 72615
rect 606243 72581 606329 72615
rect 606385 72581 606471 72615
rect 606527 72581 606613 72615
rect 606669 72581 606755 72615
rect 606811 72581 606897 72615
rect 606953 72581 607039 72615
rect 605122 72525 605176 72581
rect 605249 72559 605300 72581
rect 605391 72559 605424 72581
rect 605533 72559 605548 72581
rect 605232 72525 605300 72559
rect 605356 72525 605424 72559
rect 605480 72525 605548 72559
rect 605604 72559 605619 72581
rect 605728 72559 605761 72581
rect 605852 72559 605903 72581
rect 605604 72525 605672 72559
rect 605728 72525 605796 72559
rect 605852 72525 605920 72559
rect 605976 72525 606044 72581
rect 606101 72559 606168 72581
rect 606243 72559 606292 72581
rect 606385 72559 606416 72581
rect 606527 72559 606540 72581
rect 606100 72525 606168 72559
rect 606224 72525 606292 72559
rect 606348 72525 606416 72559
rect 606472 72525 606540 72559
rect 606596 72559 606613 72581
rect 606720 72559 606755 72581
rect 606844 72559 606897 72581
rect 606596 72525 606664 72559
rect 606720 72525 606788 72559
rect 606844 72525 606912 72559
rect 606968 72525 607036 72581
rect 607095 72559 607172 72615
rect 607092 72525 607172 72559
rect 605122 72473 607172 72525
rect 605122 72457 605193 72473
rect 605249 72457 605335 72473
rect 605391 72457 605477 72473
rect 605533 72457 605619 72473
rect 605675 72457 605761 72473
rect 605817 72457 605903 72473
rect 605959 72457 606045 72473
rect 606101 72457 606187 72473
rect 606243 72457 606329 72473
rect 606385 72457 606471 72473
rect 606527 72457 606613 72473
rect 606669 72457 606755 72473
rect 606811 72457 606897 72473
rect 606953 72457 607039 72473
rect 605122 72401 605176 72457
rect 605249 72417 605300 72457
rect 605391 72417 605424 72457
rect 605533 72417 605548 72457
rect 605232 72401 605300 72417
rect 605356 72401 605424 72417
rect 605480 72401 605548 72417
rect 605604 72417 605619 72457
rect 605728 72417 605761 72457
rect 605852 72417 605903 72457
rect 605604 72401 605672 72417
rect 605728 72401 605796 72417
rect 605852 72401 605920 72417
rect 605976 72401 606044 72457
rect 606101 72417 606168 72457
rect 606243 72417 606292 72457
rect 606385 72417 606416 72457
rect 606527 72417 606540 72457
rect 606100 72401 606168 72417
rect 606224 72401 606292 72417
rect 606348 72401 606416 72417
rect 606472 72401 606540 72417
rect 606596 72417 606613 72457
rect 606720 72417 606755 72457
rect 606844 72417 606897 72457
rect 606596 72401 606664 72417
rect 606720 72401 606788 72417
rect 606844 72401 606912 72417
rect 606968 72401 607036 72457
rect 607095 72417 607172 72473
rect 607092 72401 607172 72417
rect 605122 72333 607172 72401
rect 605122 72277 605176 72333
rect 605232 72331 605300 72333
rect 605356 72331 605424 72333
rect 605480 72331 605548 72333
rect 605249 72277 605300 72331
rect 605391 72277 605424 72331
rect 605533 72277 605548 72331
rect 605604 72331 605672 72333
rect 605728 72331 605796 72333
rect 605852 72331 605920 72333
rect 605604 72277 605619 72331
rect 605728 72277 605761 72331
rect 605852 72277 605903 72331
rect 605976 72277 606044 72333
rect 606100 72331 606168 72333
rect 606224 72331 606292 72333
rect 606348 72331 606416 72333
rect 606472 72331 606540 72333
rect 606101 72277 606168 72331
rect 606243 72277 606292 72331
rect 606385 72277 606416 72331
rect 606527 72277 606540 72331
rect 606596 72331 606664 72333
rect 606720 72331 606788 72333
rect 606844 72331 606912 72333
rect 606596 72277 606613 72331
rect 606720 72277 606755 72331
rect 606844 72277 606897 72331
rect 606968 72277 607036 72333
rect 607092 72331 607172 72333
rect 605122 72275 605193 72277
rect 605249 72275 605335 72277
rect 605391 72275 605477 72277
rect 605533 72275 605619 72277
rect 605675 72275 605761 72277
rect 605817 72275 605903 72277
rect 605959 72275 606045 72277
rect 606101 72275 606187 72277
rect 606243 72275 606329 72277
rect 606385 72275 606471 72277
rect 606527 72275 606613 72277
rect 606669 72275 606755 72277
rect 606811 72275 606897 72277
rect 606953 72275 607039 72277
rect 607095 72275 607172 72331
rect 605122 72209 607172 72275
rect 605122 72153 605176 72209
rect 605232 72189 605300 72209
rect 605356 72189 605424 72209
rect 605480 72189 605548 72209
rect 605249 72153 605300 72189
rect 605391 72153 605424 72189
rect 605533 72153 605548 72189
rect 605604 72189 605672 72209
rect 605728 72189 605796 72209
rect 605852 72189 605920 72209
rect 605604 72153 605619 72189
rect 605728 72153 605761 72189
rect 605852 72153 605903 72189
rect 605976 72153 606044 72209
rect 606100 72189 606168 72209
rect 606224 72189 606292 72209
rect 606348 72189 606416 72209
rect 606472 72189 606540 72209
rect 606101 72153 606168 72189
rect 606243 72153 606292 72189
rect 606385 72153 606416 72189
rect 606527 72153 606540 72189
rect 606596 72189 606664 72209
rect 606720 72189 606788 72209
rect 606844 72189 606912 72209
rect 606596 72153 606613 72189
rect 606720 72153 606755 72189
rect 606844 72153 606897 72189
rect 606968 72153 607036 72209
rect 607092 72189 607172 72209
rect 605122 72133 605193 72153
rect 605249 72133 605335 72153
rect 605391 72133 605477 72153
rect 605533 72133 605619 72153
rect 605675 72133 605761 72153
rect 605817 72133 605903 72153
rect 605959 72133 606045 72153
rect 606101 72133 606187 72153
rect 606243 72133 606329 72153
rect 606385 72133 606471 72153
rect 606527 72133 606613 72153
rect 606669 72133 606755 72153
rect 606811 72133 606897 72153
rect 606953 72133 607039 72153
rect 607095 72133 607172 72189
rect 605122 72088 607172 72133
rect 607828 74035 609878 74088
rect 607828 73979 607899 74035
rect 607955 73979 608041 74035
rect 608097 73979 608183 74035
rect 608239 73979 608325 74035
rect 608381 73979 608467 74035
rect 608523 73979 608609 74035
rect 608665 73979 608751 74035
rect 608807 73979 608893 74035
rect 608949 73979 609035 74035
rect 609091 73979 609177 74035
rect 609233 73979 609319 74035
rect 609375 73979 609461 74035
rect 609517 73979 609603 74035
rect 609659 73979 609745 74035
rect 609801 73979 609878 74035
rect 607828 73945 609878 73979
rect 607828 73889 607882 73945
rect 607938 73893 608006 73945
rect 608062 73893 608130 73945
rect 608186 73893 608254 73945
rect 607955 73889 608006 73893
rect 608097 73889 608130 73893
rect 608239 73889 608254 73893
rect 608310 73893 608378 73945
rect 608434 73893 608502 73945
rect 608558 73893 608626 73945
rect 608310 73889 608325 73893
rect 608434 73889 608467 73893
rect 608558 73889 608609 73893
rect 608682 73889 608750 73945
rect 608806 73893 608874 73945
rect 608930 73893 608998 73945
rect 609054 73893 609122 73945
rect 609178 73893 609246 73945
rect 608807 73889 608874 73893
rect 608949 73889 608998 73893
rect 609091 73889 609122 73893
rect 609233 73889 609246 73893
rect 609302 73893 609370 73945
rect 609426 73893 609494 73945
rect 609550 73893 609618 73945
rect 609302 73889 609319 73893
rect 609426 73889 609461 73893
rect 609550 73889 609603 73893
rect 609674 73889 609742 73945
rect 609798 73893 609878 73945
rect 607828 73837 607899 73889
rect 607955 73837 608041 73889
rect 608097 73837 608183 73889
rect 608239 73837 608325 73889
rect 608381 73837 608467 73889
rect 608523 73837 608609 73889
rect 608665 73837 608751 73889
rect 608807 73837 608893 73889
rect 608949 73837 609035 73889
rect 609091 73837 609177 73889
rect 609233 73837 609319 73889
rect 609375 73837 609461 73889
rect 609517 73837 609603 73889
rect 609659 73837 609745 73889
rect 609801 73837 609878 73893
rect 607828 73821 609878 73837
rect 607828 73765 607882 73821
rect 607938 73765 608006 73821
rect 608062 73765 608130 73821
rect 608186 73765 608254 73821
rect 608310 73765 608378 73821
rect 608434 73765 608502 73821
rect 608558 73765 608626 73821
rect 608682 73765 608750 73821
rect 608806 73765 608874 73821
rect 608930 73765 608998 73821
rect 609054 73765 609122 73821
rect 609178 73765 609246 73821
rect 609302 73765 609370 73821
rect 609426 73765 609494 73821
rect 609550 73765 609618 73821
rect 609674 73765 609742 73821
rect 609798 73765 609878 73821
rect 607828 73751 609878 73765
rect 607828 73697 607899 73751
rect 607955 73697 608041 73751
rect 608097 73697 608183 73751
rect 608239 73697 608325 73751
rect 608381 73697 608467 73751
rect 608523 73697 608609 73751
rect 608665 73697 608751 73751
rect 608807 73697 608893 73751
rect 608949 73697 609035 73751
rect 609091 73697 609177 73751
rect 609233 73697 609319 73751
rect 609375 73697 609461 73751
rect 609517 73697 609603 73751
rect 609659 73697 609745 73751
rect 607828 73641 607882 73697
rect 607955 73695 608006 73697
rect 608097 73695 608130 73697
rect 608239 73695 608254 73697
rect 607938 73641 608006 73695
rect 608062 73641 608130 73695
rect 608186 73641 608254 73695
rect 608310 73695 608325 73697
rect 608434 73695 608467 73697
rect 608558 73695 608609 73697
rect 608310 73641 608378 73695
rect 608434 73641 608502 73695
rect 608558 73641 608626 73695
rect 608682 73641 608750 73697
rect 608807 73695 608874 73697
rect 608949 73695 608998 73697
rect 609091 73695 609122 73697
rect 609233 73695 609246 73697
rect 608806 73641 608874 73695
rect 608930 73641 608998 73695
rect 609054 73641 609122 73695
rect 609178 73641 609246 73695
rect 609302 73695 609319 73697
rect 609426 73695 609461 73697
rect 609550 73695 609603 73697
rect 609302 73641 609370 73695
rect 609426 73641 609494 73695
rect 609550 73641 609618 73695
rect 609674 73641 609742 73697
rect 609801 73695 609878 73751
rect 609798 73641 609878 73695
rect 607828 73609 609878 73641
rect 607828 73573 607899 73609
rect 607955 73573 608041 73609
rect 608097 73573 608183 73609
rect 608239 73573 608325 73609
rect 608381 73573 608467 73609
rect 608523 73573 608609 73609
rect 608665 73573 608751 73609
rect 608807 73573 608893 73609
rect 608949 73573 609035 73609
rect 609091 73573 609177 73609
rect 609233 73573 609319 73609
rect 609375 73573 609461 73609
rect 609517 73573 609603 73609
rect 609659 73573 609745 73609
rect 607828 73517 607882 73573
rect 607955 73553 608006 73573
rect 608097 73553 608130 73573
rect 608239 73553 608254 73573
rect 607938 73517 608006 73553
rect 608062 73517 608130 73553
rect 608186 73517 608254 73553
rect 608310 73553 608325 73573
rect 608434 73553 608467 73573
rect 608558 73553 608609 73573
rect 608310 73517 608378 73553
rect 608434 73517 608502 73553
rect 608558 73517 608626 73553
rect 608682 73517 608750 73573
rect 608807 73553 608874 73573
rect 608949 73553 608998 73573
rect 609091 73553 609122 73573
rect 609233 73553 609246 73573
rect 608806 73517 608874 73553
rect 608930 73517 608998 73553
rect 609054 73517 609122 73553
rect 609178 73517 609246 73553
rect 609302 73553 609319 73573
rect 609426 73553 609461 73573
rect 609550 73553 609603 73573
rect 609302 73517 609370 73553
rect 609426 73517 609494 73553
rect 609550 73517 609618 73553
rect 609674 73517 609742 73573
rect 609801 73553 609878 73609
rect 609798 73517 609878 73553
rect 607828 73467 609878 73517
rect 607828 73449 607899 73467
rect 607955 73449 608041 73467
rect 608097 73449 608183 73467
rect 608239 73449 608325 73467
rect 608381 73449 608467 73467
rect 608523 73449 608609 73467
rect 608665 73449 608751 73467
rect 608807 73449 608893 73467
rect 608949 73449 609035 73467
rect 609091 73449 609177 73467
rect 609233 73449 609319 73467
rect 609375 73449 609461 73467
rect 609517 73449 609603 73467
rect 609659 73449 609745 73467
rect 607828 73393 607882 73449
rect 607955 73411 608006 73449
rect 608097 73411 608130 73449
rect 608239 73411 608254 73449
rect 607938 73393 608006 73411
rect 608062 73393 608130 73411
rect 608186 73393 608254 73411
rect 608310 73411 608325 73449
rect 608434 73411 608467 73449
rect 608558 73411 608609 73449
rect 608310 73393 608378 73411
rect 608434 73393 608502 73411
rect 608558 73393 608626 73411
rect 608682 73393 608750 73449
rect 608807 73411 608874 73449
rect 608949 73411 608998 73449
rect 609091 73411 609122 73449
rect 609233 73411 609246 73449
rect 608806 73393 608874 73411
rect 608930 73393 608998 73411
rect 609054 73393 609122 73411
rect 609178 73393 609246 73411
rect 609302 73411 609319 73449
rect 609426 73411 609461 73449
rect 609550 73411 609603 73449
rect 609302 73393 609370 73411
rect 609426 73393 609494 73411
rect 609550 73393 609618 73411
rect 609674 73393 609742 73449
rect 609801 73411 609878 73467
rect 609798 73393 609878 73411
rect 607828 73325 609878 73393
rect 607828 73269 607882 73325
rect 607955 73269 608006 73325
rect 608097 73269 608130 73325
rect 608239 73269 608254 73325
rect 608310 73269 608325 73325
rect 608434 73269 608467 73325
rect 608558 73269 608609 73325
rect 608682 73269 608750 73325
rect 608807 73269 608874 73325
rect 608949 73269 608998 73325
rect 609091 73269 609122 73325
rect 609233 73269 609246 73325
rect 609302 73269 609319 73325
rect 609426 73269 609461 73325
rect 609550 73269 609603 73325
rect 609674 73269 609742 73325
rect 609801 73269 609878 73325
rect 607828 73201 609878 73269
rect 607828 73145 607882 73201
rect 607938 73183 608006 73201
rect 608062 73183 608130 73201
rect 608186 73183 608254 73201
rect 607955 73145 608006 73183
rect 608097 73145 608130 73183
rect 608239 73145 608254 73183
rect 608310 73183 608378 73201
rect 608434 73183 608502 73201
rect 608558 73183 608626 73201
rect 608310 73145 608325 73183
rect 608434 73145 608467 73183
rect 608558 73145 608609 73183
rect 608682 73145 608750 73201
rect 608806 73183 608874 73201
rect 608930 73183 608998 73201
rect 609054 73183 609122 73201
rect 609178 73183 609246 73201
rect 608807 73145 608874 73183
rect 608949 73145 608998 73183
rect 609091 73145 609122 73183
rect 609233 73145 609246 73183
rect 609302 73183 609370 73201
rect 609426 73183 609494 73201
rect 609550 73183 609618 73201
rect 609302 73145 609319 73183
rect 609426 73145 609461 73183
rect 609550 73145 609603 73183
rect 609674 73145 609742 73201
rect 609798 73183 609878 73201
rect 607828 73127 607899 73145
rect 607955 73127 608041 73145
rect 608097 73127 608183 73145
rect 608239 73127 608325 73145
rect 608381 73127 608467 73145
rect 608523 73127 608609 73145
rect 608665 73127 608751 73145
rect 608807 73127 608893 73145
rect 608949 73127 609035 73145
rect 609091 73127 609177 73145
rect 609233 73127 609319 73145
rect 609375 73127 609461 73145
rect 609517 73127 609603 73145
rect 609659 73127 609745 73145
rect 609801 73127 609878 73183
rect 607828 73077 609878 73127
rect 607828 73021 607882 73077
rect 607938 73041 608006 73077
rect 608062 73041 608130 73077
rect 608186 73041 608254 73077
rect 607955 73021 608006 73041
rect 608097 73021 608130 73041
rect 608239 73021 608254 73041
rect 608310 73041 608378 73077
rect 608434 73041 608502 73077
rect 608558 73041 608626 73077
rect 608310 73021 608325 73041
rect 608434 73021 608467 73041
rect 608558 73021 608609 73041
rect 608682 73021 608750 73077
rect 608806 73041 608874 73077
rect 608930 73041 608998 73077
rect 609054 73041 609122 73077
rect 609178 73041 609246 73077
rect 608807 73021 608874 73041
rect 608949 73021 608998 73041
rect 609091 73021 609122 73041
rect 609233 73021 609246 73041
rect 609302 73041 609370 73077
rect 609426 73041 609494 73077
rect 609550 73041 609618 73077
rect 609302 73021 609319 73041
rect 609426 73021 609461 73041
rect 609550 73021 609603 73041
rect 609674 73021 609742 73077
rect 609798 73041 609878 73077
rect 607828 72985 607899 73021
rect 607955 72985 608041 73021
rect 608097 72985 608183 73021
rect 608239 72985 608325 73021
rect 608381 72985 608467 73021
rect 608523 72985 608609 73021
rect 608665 72985 608751 73021
rect 608807 72985 608893 73021
rect 608949 72985 609035 73021
rect 609091 72985 609177 73021
rect 609233 72985 609319 73021
rect 609375 72985 609461 73021
rect 609517 72985 609603 73021
rect 609659 72985 609745 73021
rect 609801 72985 609878 73041
rect 607828 72953 609878 72985
rect 607828 72897 607882 72953
rect 607938 72899 608006 72953
rect 608062 72899 608130 72953
rect 608186 72899 608254 72953
rect 607955 72897 608006 72899
rect 608097 72897 608130 72899
rect 608239 72897 608254 72899
rect 608310 72899 608378 72953
rect 608434 72899 608502 72953
rect 608558 72899 608626 72953
rect 608310 72897 608325 72899
rect 608434 72897 608467 72899
rect 608558 72897 608609 72899
rect 608682 72897 608750 72953
rect 608806 72899 608874 72953
rect 608930 72899 608998 72953
rect 609054 72899 609122 72953
rect 609178 72899 609246 72953
rect 608807 72897 608874 72899
rect 608949 72897 608998 72899
rect 609091 72897 609122 72899
rect 609233 72897 609246 72899
rect 609302 72899 609370 72953
rect 609426 72899 609494 72953
rect 609550 72899 609618 72953
rect 609302 72897 609319 72899
rect 609426 72897 609461 72899
rect 609550 72897 609603 72899
rect 609674 72897 609742 72953
rect 609798 72899 609878 72953
rect 607828 72843 607899 72897
rect 607955 72843 608041 72897
rect 608097 72843 608183 72897
rect 608239 72843 608325 72897
rect 608381 72843 608467 72897
rect 608523 72843 608609 72897
rect 608665 72843 608751 72897
rect 608807 72843 608893 72897
rect 608949 72843 609035 72897
rect 609091 72843 609177 72897
rect 609233 72843 609319 72897
rect 609375 72843 609461 72897
rect 609517 72843 609603 72897
rect 609659 72843 609745 72897
rect 609801 72843 609878 72899
rect 607828 72829 609878 72843
rect 607828 72773 607882 72829
rect 607938 72773 608006 72829
rect 608062 72773 608130 72829
rect 608186 72773 608254 72829
rect 608310 72773 608378 72829
rect 608434 72773 608502 72829
rect 608558 72773 608626 72829
rect 608682 72773 608750 72829
rect 608806 72773 608874 72829
rect 608930 72773 608998 72829
rect 609054 72773 609122 72829
rect 609178 72773 609246 72829
rect 609302 72773 609370 72829
rect 609426 72773 609494 72829
rect 609550 72773 609618 72829
rect 609674 72773 609742 72829
rect 609798 72773 609878 72829
rect 607828 72757 609878 72773
rect 607828 72705 607899 72757
rect 607955 72705 608041 72757
rect 608097 72705 608183 72757
rect 608239 72705 608325 72757
rect 608381 72705 608467 72757
rect 608523 72705 608609 72757
rect 608665 72705 608751 72757
rect 608807 72705 608893 72757
rect 608949 72705 609035 72757
rect 609091 72705 609177 72757
rect 609233 72705 609319 72757
rect 609375 72705 609461 72757
rect 609517 72705 609603 72757
rect 609659 72705 609745 72757
rect 607828 72649 607882 72705
rect 607955 72701 608006 72705
rect 608097 72701 608130 72705
rect 608239 72701 608254 72705
rect 607938 72649 608006 72701
rect 608062 72649 608130 72701
rect 608186 72649 608254 72701
rect 608310 72701 608325 72705
rect 608434 72701 608467 72705
rect 608558 72701 608609 72705
rect 608310 72649 608378 72701
rect 608434 72649 608502 72701
rect 608558 72649 608626 72701
rect 608682 72649 608750 72705
rect 608807 72701 608874 72705
rect 608949 72701 608998 72705
rect 609091 72701 609122 72705
rect 609233 72701 609246 72705
rect 608806 72649 608874 72701
rect 608930 72649 608998 72701
rect 609054 72649 609122 72701
rect 609178 72649 609246 72701
rect 609302 72701 609319 72705
rect 609426 72701 609461 72705
rect 609550 72701 609603 72705
rect 609302 72649 609370 72701
rect 609426 72649 609494 72701
rect 609550 72649 609618 72701
rect 609674 72649 609742 72705
rect 609801 72701 609878 72757
rect 609798 72649 609878 72701
rect 607828 72615 609878 72649
rect 607828 72581 607899 72615
rect 607955 72581 608041 72615
rect 608097 72581 608183 72615
rect 608239 72581 608325 72615
rect 608381 72581 608467 72615
rect 608523 72581 608609 72615
rect 608665 72581 608751 72615
rect 608807 72581 608893 72615
rect 608949 72581 609035 72615
rect 609091 72581 609177 72615
rect 609233 72581 609319 72615
rect 609375 72581 609461 72615
rect 609517 72581 609603 72615
rect 609659 72581 609745 72615
rect 607828 72525 607882 72581
rect 607955 72559 608006 72581
rect 608097 72559 608130 72581
rect 608239 72559 608254 72581
rect 607938 72525 608006 72559
rect 608062 72525 608130 72559
rect 608186 72525 608254 72559
rect 608310 72559 608325 72581
rect 608434 72559 608467 72581
rect 608558 72559 608609 72581
rect 608310 72525 608378 72559
rect 608434 72525 608502 72559
rect 608558 72525 608626 72559
rect 608682 72525 608750 72581
rect 608807 72559 608874 72581
rect 608949 72559 608998 72581
rect 609091 72559 609122 72581
rect 609233 72559 609246 72581
rect 608806 72525 608874 72559
rect 608930 72525 608998 72559
rect 609054 72525 609122 72559
rect 609178 72525 609246 72559
rect 609302 72559 609319 72581
rect 609426 72559 609461 72581
rect 609550 72559 609603 72581
rect 609302 72525 609370 72559
rect 609426 72525 609494 72559
rect 609550 72525 609618 72559
rect 609674 72525 609742 72581
rect 609801 72559 609878 72615
rect 609798 72525 609878 72559
rect 607828 72473 609878 72525
rect 607828 72457 607899 72473
rect 607955 72457 608041 72473
rect 608097 72457 608183 72473
rect 608239 72457 608325 72473
rect 608381 72457 608467 72473
rect 608523 72457 608609 72473
rect 608665 72457 608751 72473
rect 608807 72457 608893 72473
rect 608949 72457 609035 72473
rect 609091 72457 609177 72473
rect 609233 72457 609319 72473
rect 609375 72457 609461 72473
rect 609517 72457 609603 72473
rect 609659 72457 609745 72473
rect 607828 72401 607882 72457
rect 607955 72417 608006 72457
rect 608097 72417 608130 72457
rect 608239 72417 608254 72457
rect 607938 72401 608006 72417
rect 608062 72401 608130 72417
rect 608186 72401 608254 72417
rect 608310 72417 608325 72457
rect 608434 72417 608467 72457
rect 608558 72417 608609 72457
rect 608310 72401 608378 72417
rect 608434 72401 608502 72417
rect 608558 72401 608626 72417
rect 608682 72401 608750 72457
rect 608807 72417 608874 72457
rect 608949 72417 608998 72457
rect 609091 72417 609122 72457
rect 609233 72417 609246 72457
rect 608806 72401 608874 72417
rect 608930 72401 608998 72417
rect 609054 72401 609122 72417
rect 609178 72401 609246 72417
rect 609302 72417 609319 72457
rect 609426 72417 609461 72457
rect 609550 72417 609603 72457
rect 609302 72401 609370 72417
rect 609426 72401 609494 72417
rect 609550 72401 609618 72417
rect 609674 72401 609742 72457
rect 609801 72417 609878 72473
rect 609798 72401 609878 72417
rect 607828 72333 609878 72401
rect 607828 72277 607882 72333
rect 607938 72331 608006 72333
rect 608062 72331 608130 72333
rect 608186 72331 608254 72333
rect 607955 72277 608006 72331
rect 608097 72277 608130 72331
rect 608239 72277 608254 72331
rect 608310 72331 608378 72333
rect 608434 72331 608502 72333
rect 608558 72331 608626 72333
rect 608310 72277 608325 72331
rect 608434 72277 608467 72331
rect 608558 72277 608609 72331
rect 608682 72277 608750 72333
rect 608806 72331 608874 72333
rect 608930 72331 608998 72333
rect 609054 72331 609122 72333
rect 609178 72331 609246 72333
rect 608807 72277 608874 72331
rect 608949 72277 608998 72331
rect 609091 72277 609122 72331
rect 609233 72277 609246 72331
rect 609302 72331 609370 72333
rect 609426 72331 609494 72333
rect 609550 72331 609618 72333
rect 609302 72277 609319 72331
rect 609426 72277 609461 72331
rect 609550 72277 609603 72331
rect 609674 72277 609742 72333
rect 609798 72331 609878 72333
rect 607828 72275 607899 72277
rect 607955 72275 608041 72277
rect 608097 72275 608183 72277
rect 608239 72275 608325 72277
rect 608381 72275 608467 72277
rect 608523 72275 608609 72277
rect 608665 72275 608751 72277
rect 608807 72275 608893 72277
rect 608949 72275 609035 72277
rect 609091 72275 609177 72277
rect 609233 72275 609319 72277
rect 609375 72275 609461 72277
rect 609517 72275 609603 72277
rect 609659 72275 609745 72277
rect 609801 72275 609878 72331
rect 607828 72209 609878 72275
rect 607828 72153 607882 72209
rect 607938 72189 608006 72209
rect 608062 72189 608130 72209
rect 608186 72189 608254 72209
rect 607955 72153 608006 72189
rect 608097 72153 608130 72189
rect 608239 72153 608254 72189
rect 608310 72189 608378 72209
rect 608434 72189 608502 72209
rect 608558 72189 608626 72209
rect 608310 72153 608325 72189
rect 608434 72153 608467 72189
rect 608558 72153 608609 72189
rect 608682 72153 608750 72209
rect 608806 72189 608874 72209
rect 608930 72189 608998 72209
rect 609054 72189 609122 72209
rect 609178 72189 609246 72209
rect 608807 72153 608874 72189
rect 608949 72153 608998 72189
rect 609091 72153 609122 72189
rect 609233 72153 609246 72189
rect 609302 72189 609370 72209
rect 609426 72189 609494 72209
rect 609550 72189 609618 72209
rect 609302 72153 609319 72189
rect 609426 72153 609461 72189
rect 609550 72153 609603 72189
rect 609674 72153 609742 72209
rect 609798 72189 609878 72209
rect 607828 72133 607899 72153
rect 607955 72133 608041 72153
rect 608097 72133 608183 72153
rect 608239 72133 608325 72153
rect 608381 72133 608467 72153
rect 608523 72133 608609 72153
rect 608665 72133 608751 72153
rect 608807 72133 608893 72153
rect 608949 72133 609035 72153
rect 609091 72133 609177 72153
rect 609233 72133 609319 72153
rect 609375 72133 609461 72153
rect 609517 72133 609603 72153
rect 609659 72133 609745 72153
rect 609801 72133 609878 72189
rect 607828 72088 609878 72133
rect 610198 74035 612248 74088
rect 610198 73979 610269 74035
rect 610325 73979 610411 74035
rect 610467 73979 610553 74035
rect 610609 73979 610695 74035
rect 610751 73979 610837 74035
rect 610893 73979 610979 74035
rect 611035 73979 611121 74035
rect 611177 73979 611263 74035
rect 611319 73979 611405 74035
rect 611461 73979 611547 74035
rect 611603 73979 611689 74035
rect 611745 73979 611831 74035
rect 611887 73979 611973 74035
rect 612029 73979 612115 74035
rect 612171 73979 612248 74035
rect 610198 73945 612248 73979
rect 610198 73889 610252 73945
rect 610308 73893 610376 73945
rect 610432 73893 610500 73945
rect 610556 73893 610624 73945
rect 610325 73889 610376 73893
rect 610467 73889 610500 73893
rect 610609 73889 610624 73893
rect 610680 73893 610748 73945
rect 610804 73893 610872 73945
rect 610928 73893 610996 73945
rect 610680 73889 610695 73893
rect 610804 73889 610837 73893
rect 610928 73889 610979 73893
rect 611052 73889 611120 73945
rect 611176 73893 611244 73945
rect 611300 73893 611368 73945
rect 611424 73893 611492 73945
rect 611548 73893 611616 73945
rect 611177 73889 611244 73893
rect 611319 73889 611368 73893
rect 611461 73889 611492 73893
rect 611603 73889 611616 73893
rect 611672 73893 611740 73945
rect 611796 73893 611864 73945
rect 611920 73893 611988 73945
rect 611672 73889 611689 73893
rect 611796 73889 611831 73893
rect 611920 73889 611973 73893
rect 612044 73889 612112 73945
rect 612168 73893 612248 73945
rect 610198 73837 610269 73889
rect 610325 73837 610411 73889
rect 610467 73837 610553 73889
rect 610609 73837 610695 73889
rect 610751 73837 610837 73889
rect 610893 73837 610979 73889
rect 611035 73837 611121 73889
rect 611177 73837 611263 73889
rect 611319 73837 611405 73889
rect 611461 73837 611547 73889
rect 611603 73837 611689 73889
rect 611745 73837 611831 73889
rect 611887 73837 611973 73889
rect 612029 73837 612115 73889
rect 612171 73837 612248 73893
rect 610198 73821 612248 73837
rect 610198 73765 610252 73821
rect 610308 73765 610376 73821
rect 610432 73765 610500 73821
rect 610556 73765 610624 73821
rect 610680 73765 610748 73821
rect 610804 73765 610872 73821
rect 610928 73765 610996 73821
rect 611052 73765 611120 73821
rect 611176 73765 611244 73821
rect 611300 73765 611368 73821
rect 611424 73765 611492 73821
rect 611548 73765 611616 73821
rect 611672 73765 611740 73821
rect 611796 73765 611864 73821
rect 611920 73765 611988 73821
rect 612044 73765 612112 73821
rect 612168 73765 612248 73821
rect 610198 73751 612248 73765
rect 610198 73697 610269 73751
rect 610325 73697 610411 73751
rect 610467 73697 610553 73751
rect 610609 73697 610695 73751
rect 610751 73697 610837 73751
rect 610893 73697 610979 73751
rect 611035 73697 611121 73751
rect 611177 73697 611263 73751
rect 611319 73697 611405 73751
rect 611461 73697 611547 73751
rect 611603 73697 611689 73751
rect 611745 73697 611831 73751
rect 611887 73697 611973 73751
rect 612029 73697 612115 73751
rect 610198 73641 610252 73697
rect 610325 73695 610376 73697
rect 610467 73695 610500 73697
rect 610609 73695 610624 73697
rect 610308 73641 610376 73695
rect 610432 73641 610500 73695
rect 610556 73641 610624 73695
rect 610680 73695 610695 73697
rect 610804 73695 610837 73697
rect 610928 73695 610979 73697
rect 610680 73641 610748 73695
rect 610804 73641 610872 73695
rect 610928 73641 610996 73695
rect 611052 73641 611120 73697
rect 611177 73695 611244 73697
rect 611319 73695 611368 73697
rect 611461 73695 611492 73697
rect 611603 73695 611616 73697
rect 611176 73641 611244 73695
rect 611300 73641 611368 73695
rect 611424 73641 611492 73695
rect 611548 73641 611616 73695
rect 611672 73695 611689 73697
rect 611796 73695 611831 73697
rect 611920 73695 611973 73697
rect 611672 73641 611740 73695
rect 611796 73641 611864 73695
rect 611920 73641 611988 73695
rect 612044 73641 612112 73697
rect 612171 73695 612248 73751
rect 612168 73641 612248 73695
rect 610198 73609 612248 73641
rect 610198 73573 610269 73609
rect 610325 73573 610411 73609
rect 610467 73573 610553 73609
rect 610609 73573 610695 73609
rect 610751 73573 610837 73609
rect 610893 73573 610979 73609
rect 611035 73573 611121 73609
rect 611177 73573 611263 73609
rect 611319 73573 611405 73609
rect 611461 73573 611547 73609
rect 611603 73573 611689 73609
rect 611745 73573 611831 73609
rect 611887 73573 611973 73609
rect 612029 73573 612115 73609
rect 610198 73517 610252 73573
rect 610325 73553 610376 73573
rect 610467 73553 610500 73573
rect 610609 73553 610624 73573
rect 610308 73517 610376 73553
rect 610432 73517 610500 73553
rect 610556 73517 610624 73553
rect 610680 73553 610695 73573
rect 610804 73553 610837 73573
rect 610928 73553 610979 73573
rect 610680 73517 610748 73553
rect 610804 73517 610872 73553
rect 610928 73517 610996 73553
rect 611052 73517 611120 73573
rect 611177 73553 611244 73573
rect 611319 73553 611368 73573
rect 611461 73553 611492 73573
rect 611603 73553 611616 73573
rect 611176 73517 611244 73553
rect 611300 73517 611368 73553
rect 611424 73517 611492 73553
rect 611548 73517 611616 73553
rect 611672 73553 611689 73573
rect 611796 73553 611831 73573
rect 611920 73553 611973 73573
rect 611672 73517 611740 73553
rect 611796 73517 611864 73553
rect 611920 73517 611988 73553
rect 612044 73517 612112 73573
rect 612171 73553 612248 73609
rect 612168 73517 612248 73553
rect 610198 73467 612248 73517
rect 610198 73449 610269 73467
rect 610325 73449 610411 73467
rect 610467 73449 610553 73467
rect 610609 73449 610695 73467
rect 610751 73449 610837 73467
rect 610893 73449 610979 73467
rect 611035 73449 611121 73467
rect 611177 73449 611263 73467
rect 611319 73449 611405 73467
rect 611461 73449 611547 73467
rect 611603 73449 611689 73467
rect 611745 73449 611831 73467
rect 611887 73449 611973 73467
rect 612029 73449 612115 73467
rect 610198 73393 610252 73449
rect 610325 73411 610376 73449
rect 610467 73411 610500 73449
rect 610609 73411 610624 73449
rect 610308 73393 610376 73411
rect 610432 73393 610500 73411
rect 610556 73393 610624 73411
rect 610680 73411 610695 73449
rect 610804 73411 610837 73449
rect 610928 73411 610979 73449
rect 610680 73393 610748 73411
rect 610804 73393 610872 73411
rect 610928 73393 610996 73411
rect 611052 73393 611120 73449
rect 611177 73411 611244 73449
rect 611319 73411 611368 73449
rect 611461 73411 611492 73449
rect 611603 73411 611616 73449
rect 611176 73393 611244 73411
rect 611300 73393 611368 73411
rect 611424 73393 611492 73411
rect 611548 73393 611616 73411
rect 611672 73411 611689 73449
rect 611796 73411 611831 73449
rect 611920 73411 611973 73449
rect 611672 73393 611740 73411
rect 611796 73393 611864 73411
rect 611920 73393 611988 73411
rect 612044 73393 612112 73449
rect 612171 73411 612248 73467
rect 612168 73393 612248 73411
rect 610198 73325 612248 73393
rect 610198 73269 610252 73325
rect 610325 73269 610376 73325
rect 610467 73269 610500 73325
rect 610609 73269 610624 73325
rect 610680 73269 610695 73325
rect 610804 73269 610837 73325
rect 610928 73269 610979 73325
rect 611052 73269 611120 73325
rect 611177 73269 611244 73325
rect 611319 73269 611368 73325
rect 611461 73269 611492 73325
rect 611603 73269 611616 73325
rect 611672 73269 611689 73325
rect 611796 73269 611831 73325
rect 611920 73269 611973 73325
rect 612044 73269 612112 73325
rect 612171 73269 612248 73325
rect 610198 73201 612248 73269
rect 610198 73145 610252 73201
rect 610308 73183 610376 73201
rect 610432 73183 610500 73201
rect 610556 73183 610624 73201
rect 610325 73145 610376 73183
rect 610467 73145 610500 73183
rect 610609 73145 610624 73183
rect 610680 73183 610748 73201
rect 610804 73183 610872 73201
rect 610928 73183 610996 73201
rect 610680 73145 610695 73183
rect 610804 73145 610837 73183
rect 610928 73145 610979 73183
rect 611052 73145 611120 73201
rect 611176 73183 611244 73201
rect 611300 73183 611368 73201
rect 611424 73183 611492 73201
rect 611548 73183 611616 73201
rect 611177 73145 611244 73183
rect 611319 73145 611368 73183
rect 611461 73145 611492 73183
rect 611603 73145 611616 73183
rect 611672 73183 611740 73201
rect 611796 73183 611864 73201
rect 611920 73183 611988 73201
rect 611672 73145 611689 73183
rect 611796 73145 611831 73183
rect 611920 73145 611973 73183
rect 612044 73145 612112 73201
rect 612168 73183 612248 73201
rect 610198 73127 610269 73145
rect 610325 73127 610411 73145
rect 610467 73127 610553 73145
rect 610609 73127 610695 73145
rect 610751 73127 610837 73145
rect 610893 73127 610979 73145
rect 611035 73127 611121 73145
rect 611177 73127 611263 73145
rect 611319 73127 611405 73145
rect 611461 73127 611547 73145
rect 611603 73127 611689 73145
rect 611745 73127 611831 73145
rect 611887 73127 611973 73145
rect 612029 73127 612115 73145
rect 612171 73127 612248 73183
rect 610198 73077 612248 73127
rect 610198 73021 610252 73077
rect 610308 73041 610376 73077
rect 610432 73041 610500 73077
rect 610556 73041 610624 73077
rect 610325 73021 610376 73041
rect 610467 73021 610500 73041
rect 610609 73021 610624 73041
rect 610680 73041 610748 73077
rect 610804 73041 610872 73077
rect 610928 73041 610996 73077
rect 610680 73021 610695 73041
rect 610804 73021 610837 73041
rect 610928 73021 610979 73041
rect 611052 73021 611120 73077
rect 611176 73041 611244 73077
rect 611300 73041 611368 73077
rect 611424 73041 611492 73077
rect 611548 73041 611616 73077
rect 611177 73021 611244 73041
rect 611319 73021 611368 73041
rect 611461 73021 611492 73041
rect 611603 73021 611616 73041
rect 611672 73041 611740 73077
rect 611796 73041 611864 73077
rect 611920 73041 611988 73077
rect 611672 73021 611689 73041
rect 611796 73021 611831 73041
rect 611920 73021 611973 73041
rect 612044 73021 612112 73077
rect 612168 73041 612248 73077
rect 610198 72985 610269 73021
rect 610325 72985 610411 73021
rect 610467 72985 610553 73021
rect 610609 72985 610695 73021
rect 610751 72985 610837 73021
rect 610893 72985 610979 73021
rect 611035 72985 611121 73021
rect 611177 72985 611263 73021
rect 611319 72985 611405 73021
rect 611461 72985 611547 73021
rect 611603 72985 611689 73021
rect 611745 72985 611831 73021
rect 611887 72985 611973 73021
rect 612029 72985 612115 73021
rect 612171 72985 612248 73041
rect 610198 72953 612248 72985
rect 610198 72897 610252 72953
rect 610308 72899 610376 72953
rect 610432 72899 610500 72953
rect 610556 72899 610624 72953
rect 610325 72897 610376 72899
rect 610467 72897 610500 72899
rect 610609 72897 610624 72899
rect 610680 72899 610748 72953
rect 610804 72899 610872 72953
rect 610928 72899 610996 72953
rect 610680 72897 610695 72899
rect 610804 72897 610837 72899
rect 610928 72897 610979 72899
rect 611052 72897 611120 72953
rect 611176 72899 611244 72953
rect 611300 72899 611368 72953
rect 611424 72899 611492 72953
rect 611548 72899 611616 72953
rect 611177 72897 611244 72899
rect 611319 72897 611368 72899
rect 611461 72897 611492 72899
rect 611603 72897 611616 72899
rect 611672 72899 611740 72953
rect 611796 72899 611864 72953
rect 611920 72899 611988 72953
rect 611672 72897 611689 72899
rect 611796 72897 611831 72899
rect 611920 72897 611973 72899
rect 612044 72897 612112 72953
rect 612168 72899 612248 72953
rect 610198 72843 610269 72897
rect 610325 72843 610411 72897
rect 610467 72843 610553 72897
rect 610609 72843 610695 72897
rect 610751 72843 610837 72897
rect 610893 72843 610979 72897
rect 611035 72843 611121 72897
rect 611177 72843 611263 72897
rect 611319 72843 611405 72897
rect 611461 72843 611547 72897
rect 611603 72843 611689 72897
rect 611745 72843 611831 72897
rect 611887 72843 611973 72897
rect 612029 72843 612115 72897
rect 612171 72843 612248 72899
rect 610198 72829 612248 72843
rect 610198 72773 610252 72829
rect 610308 72773 610376 72829
rect 610432 72773 610500 72829
rect 610556 72773 610624 72829
rect 610680 72773 610748 72829
rect 610804 72773 610872 72829
rect 610928 72773 610996 72829
rect 611052 72773 611120 72829
rect 611176 72773 611244 72829
rect 611300 72773 611368 72829
rect 611424 72773 611492 72829
rect 611548 72773 611616 72829
rect 611672 72773 611740 72829
rect 611796 72773 611864 72829
rect 611920 72773 611988 72829
rect 612044 72773 612112 72829
rect 612168 72773 612248 72829
rect 610198 72757 612248 72773
rect 610198 72705 610269 72757
rect 610325 72705 610411 72757
rect 610467 72705 610553 72757
rect 610609 72705 610695 72757
rect 610751 72705 610837 72757
rect 610893 72705 610979 72757
rect 611035 72705 611121 72757
rect 611177 72705 611263 72757
rect 611319 72705 611405 72757
rect 611461 72705 611547 72757
rect 611603 72705 611689 72757
rect 611745 72705 611831 72757
rect 611887 72705 611973 72757
rect 612029 72705 612115 72757
rect 610198 72649 610252 72705
rect 610325 72701 610376 72705
rect 610467 72701 610500 72705
rect 610609 72701 610624 72705
rect 610308 72649 610376 72701
rect 610432 72649 610500 72701
rect 610556 72649 610624 72701
rect 610680 72701 610695 72705
rect 610804 72701 610837 72705
rect 610928 72701 610979 72705
rect 610680 72649 610748 72701
rect 610804 72649 610872 72701
rect 610928 72649 610996 72701
rect 611052 72649 611120 72705
rect 611177 72701 611244 72705
rect 611319 72701 611368 72705
rect 611461 72701 611492 72705
rect 611603 72701 611616 72705
rect 611176 72649 611244 72701
rect 611300 72649 611368 72701
rect 611424 72649 611492 72701
rect 611548 72649 611616 72701
rect 611672 72701 611689 72705
rect 611796 72701 611831 72705
rect 611920 72701 611973 72705
rect 611672 72649 611740 72701
rect 611796 72649 611864 72701
rect 611920 72649 611988 72701
rect 612044 72649 612112 72705
rect 612171 72701 612248 72757
rect 612168 72649 612248 72701
rect 610198 72615 612248 72649
rect 610198 72581 610269 72615
rect 610325 72581 610411 72615
rect 610467 72581 610553 72615
rect 610609 72581 610695 72615
rect 610751 72581 610837 72615
rect 610893 72581 610979 72615
rect 611035 72581 611121 72615
rect 611177 72581 611263 72615
rect 611319 72581 611405 72615
rect 611461 72581 611547 72615
rect 611603 72581 611689 72615
rect 611745 72581 611831 72615
rect 611887 72581 611973 72615
rect 612029 72581 612115 72615
rect 610198 72525 610252 72581
rect 610325 72559 610376 72581
rect 610467 72559 610500 72581
rect 610609 72559 610624 72581
rect 610308 72525 610376 72559
rect 610432 72525 610500 72559
rect 610556 72525 610624 72559
rect 610680 72559 610695 72581
rect 610804 72559 610837 72581
rect 610928 72559 610979 72581
rect 610680 72525 610748 72559
rect 610804 72525 610872 72559
rect 610928 72525 610996 72559
rect 611052 72525 611120 72581
rect 611177 72559 611244 72581
rect 611319 72559 611368 72581
rect 611461 72559 611492 72581
rect 611603 72559 611616 72581
rect 611176 72525 611244 72559
rect 611300 72525 611368 72559
rect 611424 72525 611492 72559
rect 611548 72525 611616 72559
rect 611672 72559 611689 72581
rect 611796 72559 611831 72581
rect 611920 72559 611973 72581
rect 611672 72525 611740 72559
rect 611796 72525 611864 72559
rect 611920 72525 611988 72559
rect 612044 72525 612112 72581
rect 612171 72559 612248 72615
rect 612168 72525 612248 72559
rect 610198 72473 612248 72525
rect 610198 72457 610269 72473
rect 610325 72457 610411 72473
rect 610467 72457 610553 72473
rect 610609 72457 610695 72473
rect 610751 72457 610837 72473
rect 610893 72457 610979 72473
rect 611035 72457 611121 72473
rect 611177 72457 611263 72473
rect 611319 72457 611405 72473
rect 611461 72457 611547 72473
rect 611603 72457 611689 72473
rect 611745 72457 611831 72473
rect 611887 72457 611973 72473
rect 612029 72457 612115 72473
rect 610198 72401 610252 72457
rect 610325 72417 610376 72457
rect 610467 72417 610500 72457
rect 610609 72417 610624 72457
rect 610308 72401 610376 72417
rect 610432 72401 610500 72417
rect 610556 72401 610624 72417
rect 610680 72417 610695 72457
rect 610804 72417 610837 72457
rect 610928 72417 610979 72457
rect 610680 72401 610748 72417
rect 610804 72401 610872 72417
rect 610928 72401 610996 72417
rect 611052 72401 611120 72457
rect 611177 72417 611244 72457
rect 611319 72417 611368 72457
rect 611461 72417 611492 72457
rect 611603 72417 611616 72457
rect 611176 72401 611244 72417
rect 611300 72401 611368 72417
rect 611424 72401 611492 72417
rect 611548 72401 611616 72417
rect 611672 72417 611689 72457
rect 611796 72417 611831 72457
rect 611920 72417 611973 72457
rect 611672 72401 611740 72417
rect 611796 72401 611864 72417
rect 611920 72401 611988 72417
rect 612044 72401 612112 72457
rect 612171 72417 612248 72473
rect 612168 72401 612248 72417
rect 610198 72333 612248 72401
rect 610198 72277 610252 72333
rect 610308 72331 610376 72333
rect 610432 72331 610500 72333
rect 610556 72331 610624 72333
rect 610325 72277 610376 72331
rect 610467 72277 610500 72331
rect 610609 72277 610624 72331
rect 610680 72331 610748 72333
rect 610804 72331 610872 72333
rect 610928 72331 610996 72333
rect 610680 72277 610695 72331
rect 610804 72277 610837 72331
rect 610928 72277 610979 72331
rect 611052 72277 611120 72333
rect 611176 72331 611244 72333
rect 611300 72331 611368 72333
rect 611424 72331 611492 72333
rect 611548 72331 611616 72333
rect 611177 72277 611244 72331
rect 611319 72277 611368 72331
rect 611461 72277 611492 72331
rect 611603 72277 611616 72331
rect 611672 72331 611740 72333
rect 611796 72331 611864 72333
rect 611920 72331 611988 72333
rect 611672 72277 611689 72331
rect 611796 72277 611831 72331
rect 611920 72277 611973 72331
rect 612044 72277 612112 72333
rect 612168 72331 612248 72333
rect 610198 72275 610269 72277
rect 610325 72275 610411 72277
rect 610467 72275 610553 72277
rect 610609 72275 610695 72277
rect 610751 72275 610837 72277
rect 610893 72275 610979 72277
rect 611035 72275 611121 72277
rect 611177 72275 611263 72277
rect 611319 72275 611405 72277
rect 611461 72275 611547 72277
rect 611603 72275 611689 72277
rect 611745 72275 611831 72277
rect 611887 72275 611973 72277
rect 612029 72275 612115 72277
rect 612171 72275 612248 72331
rect 610198 72209 612248 72275
rect 610198 72153 610252 72209
rect 610308 72189 610376 72209
rect 610432 72189 610500 72209
rect 610556 72189 610624 72209
rect 610325 72153 610376 72189
rect 610467 72153 610500 72189
rect 610609 72153 610624 72189
rect 610680 72189 610748 72209
rect 610804 72189 610872 72209
rect 610928 72189 610996 72209
rect 610680 72153 610695 72189
rect 610804 72153 610837 72189
rect 610928 72153 610979 72189
rect 611052 72153 611120 72209
rect 611176 72189 611244 72209
rect 611300 72189 611368 72209
rect 611424 72189 611492 72209
rect 611548 72189 611616 72209
rect 611177 72153 611244 72189
rect 611319 72153 611368 72189
rect 611461 72153 611492 72189
rect 611603 72153 611616 72189
rect 611672 72189 611740 72209
rect 611796 72189 611864 72209
rect 611920 72189 611988 72209
rect 611672 72153 611689 72189
rect 611796 72153 611831 72189
rect 611920 72153 611973 72189
rect 612044 72153 612112 72209
rect 612168 72189 612248 72209
rect 610198 72133 610269 72153
rect 610325 72133 610411 72153
rect 610467 72133 610553 72153
rect 610609 72133 610695 72153
rect 610751 72133 610837 72153
rect 610893 72133 610979 72153
rect 611035 72133 611121 72153
rect 611177 72133 611263 72153
rect 611319 72133 611405 72153
rect 611461 72133 611547 72153
rect 611603 72133 611689 72153
rect 611745 72133 611831 72153
rect 611887 72133 611973 72153
rect 612029 72133 612115 72153
rect 612171 72133 612248 72189
rect 610198 72088 612248 72133
rect 612828 74035 614728 74088
rect 612828 73979 612899 74035
rect 612955 73979 613041 74035
rect 613097 73979 613183 74035
rect 613239 73979 613325 74035
rect 613381 73979 613467 74035
rect 613523 73979 613609 74035
rect 613665 73979 613751 74035
rect 613807 73979 613893 74035
rect 613949 73979 614035 74035
rect 614091 73979 614177 74035
rect 614233 73979 614319 74035
rect 614375 73979 614461 74035
rect 614517 73979 614603 74035
rect 614659 73979 614728 74035
rect 612828 73945 614728 73979
rect 612828 73889 612882 73945
rect 612938 73893 613006 73945
rect 613062 73893 613130 73945
rect 613186 73893 613254 73945
rect 612955 73889 613006 73893
rect 613097 73889 613130 73893
rect 613239 73889 613254 73893
rect 613310 73893 613378 73945
rect 613434 73893 613502 73945
rect 613558 73893 613626 73945
rect 613310 73889 613325 73893
rect 613434 73889 613467 73893
rect 613558 73889 613609 73893
rect 613682 73889 613750 73945
rect 613806 73893 613874 73945
rect 613930 73893 613998 73945
rect 614054 73893 614122 73945
rect 614178 73893 614246 73945
rect 613807 73889 613874 73893
rect 613949 73889 613998 73893
rect 614091 73889 614122 73893
rect 614233 73889 614246 73893
rect 614302 73893 614370 73945
rect 614426 73893 614494 73945
rect 614550 73893 614618 73945
rect 614302 73889 614319 73893
rect 614426 73889 614461 73893
rect 614550 73889 614603 73893
rect 614674 73889 614728 73945
rect 612828 73837 612899 73889
rect 612955 73837 613041 73889
rect 613097 73837 613183 73889
rect 613239 73837 613325 73889
rect 613381 73837 613467 73889
rect 613523 73837 613609 73889
rect 613665 73837 613751 73889
rect 613807 73837 613893 73889
rect 613949 73837 614035 73889
rect 614091 73837 614177 73889
rect 614233 73837 614319 73889
rect 614375 73837 614461 73889
rect 614517 73837 614603 73889
rect 614659 73837 614728 73889
rect 612828 73821 614728 73837
rect 612828 73765 612882 73821
rect 612938 73765 613006 73821
rect 613062 73765 613130 73821
rect 613186 73765 613254 73821
rect 613310 73765 613378 73821
rect 613434 73765 613502 73821
rect 613558 73765 613626 73821
rect 613682 73765 613750 73821
rect 613806 73765 613874 73821
rect 613930 73765 613998 73821
rect 614054 73765 614122 73821
rect 614178 73765 614246 73821
rect 614302 73765 614370 73821
rect 614426 73765 614494 73821
rect 614550 73765 614618 73821
rect 614674 73765 614728 73821
rect 612828 73751 614728 73765
rect 612828 73697 612899 73751
rect 612955 73697 613041 73751
rect 613097 73697 613183 73751
rect 613239 73697 613325 73751
rect 613381 73697 613467 73751
rect 613523 73697 613609 73751
rect 613665 73697 613751 73751
rect 613807 73697 613893 73751
rect 613949 73697 614035 73751
rect 614091 73697 614177 73751
rect 614233 73697 614319 73751
rect 614375 73697 614461 73751
rect 614517 73697 614603 73751
rect 614659 73697 614728 73751
rect 612828 73641 612882 73697
rect 612955 73695 613006 73697
rect 613097 73695 613130 73697
rect 613239 73695 613254 73697
rect 612938 73641 613006 73695
rect 613062 73641 613130 73695
rect 613186 73641 613254 73695
rect 613310 73695 613325 73697
rect 613434 73695 613467 73697
rect 613558 73695 613609 73697
rect 613310 73641 613378 73695
rect 613434 73641 613502 73695
rect 613558 73641 613626 73695
rect 613682 73641 613750 73697
rect 613807 73695 613874 73697
rect 613949 73695 613998 73697
rect 614091 73695 614122 73697
rect 614233 73695 614246 73697
rect 613806 73641 613874 73695
rect 613930 73641 613998 73695
rect 614054 73641 614122 73695
rect 614178 73641 614246 73695
rect 614302 73695 614319 73697
rect 614426 73695 614461 73697
rect 614550 73695 614603 73697
rect 614302 73641 614370 73695
rect 614426 73641 614494 73695
rect 614550 73641 614618 73695
rect 614674 73641 614728 73697
rect 612828 73609 614728 73641
rect 612828 73573 612899 73609
rect 612955 73573 613041 73609
rect 613097 73573 613183 73609
rect 613239 73573 613325 73609
rect 613381 73573 613467 73609
rect 613523 73573 613609 73609
rect 613665 73573 613751 73609
rect 613807 73573 613893 73609
rect 613949 73573 614035 73609
rect 614091 73573 614177 73609
rect 614233 73573 614319 73609
rect 614375 73573 614461 73609
rect 614517 73573 614603 73609
rect 614659 73573 614728 73609
rect 612828 73517 612882 73573
rect 612955 73553 613006 73573
rect 613097 73553 613130 73573
rect 613239 73553 613254 73573
rect 612938 73517 613006 73553
rect 613062 73517 613130 73553
rect 613186 73517 613254 73553
rect 613310 73553 613325 73573
rect 613434 73553 613467 73573
rect 613558 73553 613609 73573
rect 613310 73517 613378 73553
rect 613434 73517 613502 73553
rect 613558 73517 613626 73553
rect 613682 73517 613750 73573
rect 613807 73553 613874 73573
rect 613949 73553 613998 73573
rect 614091 73553 614122 73573
rect 614233 73553 614246 73573
rect 613806 73517 613874 73553
rect 613930 73517 613998 73553
rect 614054 73517 614122 73553
rect 614178 73517 614246 73553
rect 614302 73553 614319 73573
rect 614426 73553 614461 73573
rect 614550 73553 614603 73573
rect 614302 73517 614370 73553
rect 614426 73517 614494 73553
rect 614550 73517 614618 73553
rect 614674 73517 614728 73573
rect 612828 73467 614728 73517
rect 612828 73449 612899 73467
rect 612955 73449 613041 73467
rect 613097 73449 613183 73467
rect 613239 73449 613325 73467
rect 613381 73449 613467 73467
rect 613523 73449 613609 73467
rect 613665 73449 613751 73467
rect 613807 73449 613893 73467
rect 613949 73449 614035 73467
rect 614091 73449 614177 73467
rect 614233 73449 614319 73467
rect 614375 73449 614461 73467
rect 614517 73449 614603 73467
rect 614659 73449 614728 73467
rect 612828 73393 612882 73449
rect 612955 73411 613006 73449
rect 613097 73411 613130 73449
rect 613239 73411 613254 73449
rect 612938 73393 613006 73411
rect 613062 73393 613130 73411
rect 613186 73393 613254 73411
rect 613310 73411 613325 73449
rect 613434 73411 613467 73449
rect 613558 73411 613609 73449
rect 613310 73393 613378 73411
rect 613434 73393 613502 73411
rect 613558 73393 613626 73411
rect 613682 73393 613750 73449
rect 613807 73411 613874 73449
rect 613949 73411 613998 73449
rect 614091 73411 614122 73449
rect 614233 73411 614246 73449
rect 613806 73393 613874 73411
rect 613930 73393 613998 73411
rect 614054 73393 614122 73411
rect 614178 73393 614246 73411
rect 614302 73411 614319 73449
rect 614426 73411 614461 73449
rect 614550 73411 614603 73449
rect 614302 73393 614370 73411
rect 614426 73393 614494 73411
rect 614550 73393 614618 73411
rect 614674 73393 614728 73449
rect 612828 73325 614728 73393
rect 612828 73269 612882 73325
rect 612955 73269 613006 73325
rect 613097 73269 613130 73325
rect 613239 73269 613254 73325
rect 613310 73269 613325 73325
rect 613434 73269 613467 73325
rect 613558 73269 613609 73325
rect 613682 73269 613750 73325
rect 613807 73269 613874 73325
rect 613949 73269 613998 73325
rect 614091 73269 614122 73325
rect 614233 73269 614246 73325
rect 614302 73269 614319 73325
rect 614426 73269 614461 73325
rect 614550 73269 614603 73325
rect 614674 73269 614728 73325
rect 612828 73201 614728 73269
rect 612828 73145 612882 73201
rect 612938 73183 613006 73201
rect 613062 73183 613130 73201
rect 613186 73183 613254 73201
rect 612955 73145 613006 73183
rect 613097 73145 613130 73183
rect 613239 73145 613254 73183
rect 613310 73183 613378 73201
rect 613434 73183 613502 73201
rect 613558 73183 613626 73201
rect 613310 73145 613325 73183
rect 613434 73145 613467 73183
rect 613558 73145 613609 73183
rect 613682 73145 613750 73201
rect 613806 73183 613874 73201
rect 613930 73183 613998 73201
rect 614054 73183 614122 73201
rect 614178 73183 614246 73201
rect 613807 73145 613874 73183
rect 613949 73145 613998 73183
rect 614091 73145 614122 73183
rect 614233 73145 614246 73183
rect 614302 73183 614370 73201
rect 614426 73183 614494 73201
rect 614550 73183 614618 73201
rect 614302 73145 614319 73183
rect 614426 73145 614461 73183
rect 614550 73145 614603 73183
rect 614674 73145 614728 73201
rect 612828 73127 612899 73145
rect 612955 73127 613041 73145
rect 613097 73127 613183 73145
rect 613239 73127 613325 73145
rect 613381 73127 613467 73145
rect 613523 73127 613609 73145
rect 613665 73127 613751 73145
rect 613807 73127 613893 73145
rect 613949 73127 614035 73145
rect 614091 73127 614177 73145
rect 614233 73127 614319 73145
rect 614375 73127 614461 73145
rect 614517 73127 614603 73145
rect 614659 73127 614728 73145
rect 612828 73077 614728 73127
rect 612828 73021 612882 73077
rect 612938 73041 613006 73077
rect 613062 73041 613130 73077
rect 613186 73041 613254 73077
rect 612955 73021 613006 73041
rect 613097 73021 613130 73041
rect 613239 73021 613254 73041
rect 613310 73041 613378 73077
rect 613434 73041 613502 73077
rect 613558 73041 613626 73077
rect 613310 73021 613325 73041
rect 613434 73021 613467 73041
rect 613558 73021 613609 73041
rect 613682 73021 613750 73077
rect 613806 73041 613874 73077
rect 613930 73041 613998 73077
rect 614054 73041 614122 73077
rect 614178 73041 614246 73077
rect 613807 73021 613874 73041
rect 613949 73021 613998 73041
rect 614091 73021 614122 73041
rect 614233 73021 614246 73041
rect 614302 73041 614370 73077
rect 614426 73041 614494 73077
rect 614550 73041 614618 73077
rect 614302 73021 614319 73041
rect 614426 73021 614461 73041
rect 614550 73021 614603 73041
rect 614674 73021 614728 73077
rect 612828 72985 612899 73021
rect 612955 72985 613041 73021
rect 613097 72985 613183 73021
rect 613239 72985 613325 73021
rect 613381 72985 613467 73021
rect 613523 72985 613609 73021
rect 613665 72985 613751 73021
rect 613807 72985 613893 73021
rect 613949 72985 614035 73021
rect 614091 72985 614177 73021
rect 614233 72985 614319 73021
rect 614375 72985 614461 73021
rect 614517 72985 614603 73021
rect 614659 72985 614728 73021
rect 612828 72953 614728 72985
rect 612828 72897 612882 72953
rect 612938 72899 613006 72953
rect 613062 72899 613130 72953
rect 613186 72899 613254 72953
rect 612955 72897 613006 72899
rect 613097 72897 613130 72899
rect 613239 72897 613254 72899
rect 613310 72899 613378 72953
rect 613434 72899 613502 72953
rect 613558 72899 613626 72953
rect 613310 72897 613325 72899
rect 613434 72897 613467 72899
rect 613558 72897 613609 72899
rect 613682 72897 613750 72953
rect 613806 72899 613874 72953
rect 613930 72899 613998 72953
rect 614054 72899 614122 72953
rect 614178 72899 614246 72953
rect 613807 72897 613874 72899
rect 613949 72897 613998 72899
rect 614091 72897 614122 72899
rect 614233 72897 614246 72899
rect 614302 72899 614370 72953
rect 614426 72899 614494 72953
rect 614550 72899 614618 72953
rect 614302 72897 614319 72899
rect 614426 72897 614461 72899
rect 614550 72897 614603 72899
rect 614674 72897 614728 72953
rect 612828 72843 612899 72897
rect 612955 72843 613041 72897
rect 613097 72843 613183 72897
rect 613239 72843 613325 72897
rect 613381 72843 613467 72897
rect 613523 72843 613609 72897
rect 613665 72843 613751 72897
rect 613807 72843 613893 72897
rect 613949 72843 614035 72897
rect 614091 72843 614177 72897
rect 614233 72843 614319 72897
rect 614375 72843 614461 72897
rect 614517 72843 614603 72897
rect 614659 72843 614728 72897
rect 612828 72829 614728 72843
rect 612828 72773 612882 72829
rect 612938 72773 613006 72829
rect 613062 72773 613130 72829
rect 613186 72773 613254 72829
rect 613310 72773 613378 72829
rect 613434 72773 613502 72829
rect 613558 72773 613626 72829
rect 613682 72773 613750 72829
rect 613806 72773 613874 72829
rect 613930 72773 613998 72829
rect 614054 72773 614122 72829
rect 614178 72773 614246 72829
rect 614302 72773 614370 72829
rect 614426 72773 614494 72829
rect 614550 72773 614618 72829
rect 614674 72773 614728 72829
rect 612828 72757 614728 72773
rect 612828 72705 612899 72757
rect 612955 72705 613041 72757
rect 613097 72705 613183 72757
rect 613239 72705 613325 72757
rect 613381 72705 613467 72757
rect 613523 72705 613609 72757
rect 613665 72705 613751 72757
rect 613807 72705 613893 72757
rect 613949 72705 614035 72757
rect 614091 72705 614177 72757
rect 614233 72705 614319 72757
rect 614375 72705 614461 72757
rect 614517 72705 614603 72757
rect 614659 72705 614728 72757
rect 612828 72649 612882 72705
rect 612955 72701 613006 72705
rect 613097 72701 613130 72705
rect 613239 72701 613254 72705
rect 612938 72649 613006 72701
rect 613062 72649 613130 72701
rect 613186 72649 613254 72701
rect 613310 72701 613325 72705
rect 613434 72701 613467 72705
rect 613558 72701 613609 72705
rect 613310 72649 613378 72701
rect 613434 72649 613502 72701
rect 613558 72649 613626 72701
rect 613682 72649 613750 72705
rect 613807 72701 613874 72705
rect 613949 72701 613998 72705
rect 614091 72701 614122 72705
rect 614233 72701 614246 72705
rect 613806 72649 613874 72701
rect 613930 72649 613998 72701
rect 614054 72649 614122 72701
rect 614178 72649 614246 72701
rect 614302 72701 614319 72705
rect 614426 72701 614461 72705
rect 614550 72701 614603 72705
rect 614302 72649 614370 72701
rect 614426 72649 614494 72701
rect 614550 72649 614618 72701
rect 614674 72649 614728 72705
rect 612828 72615 614728 72649
rect 612828 72581 612899 72615
rect 612955 72581 613041 72615
rect 613097 72581 613183 72615
rect 613239 72581 613325 72615
rect 613381 72581 613467 72615
rect 613523 72581 613609 72615
rect 613665 72581 613751 72615
rect 613807 72581 613893 72615
rect 613949 72581 614035 72615
rect 614091 72581 614177 72615
rect 614233 72581 614319 72615
rect 614375 72581 614461 72615
rect 614517 72581 614603 72615
rect 614659 72581 614728 72615
rect 612828 72525 612882 72581
rect 612955 72559 613006 72581
rect 613097 72559 613130 72581
rect 613239 72559 613254 72581
rect 612938 72525 613006 72559
rect 613062 72525 613130 72559
rect 613186 72525 613254 72559
rect 613310 72559 613325 72581
rect 613434 72559 613467 72581
rect 613558 72559 613609 72581
rect 613310 72525 613378 72559
rect 613434 72525 613502 72559
rect 613558 72525 613626 72559
rect 613682 72525 613750 72581
rect 613807 72559 613874 72581
rect 613949 72559 613998 72581
rect 614091 72559 614122 72581
rect 614233 72559 614246 72581
rect 613806 72525 613874 72559
rect 613930 72525 613998 72559
rect 614054 72525 614122 72559
rect 614178 72525 614246 72559
rect 614302 72559 614319 72581
rect 614426 72559 614461 72581
rect 614550 72559 614603 72581
rect 614302 72525 614370 72559
rect 614426 72525 614494 72559
rect 614550 72525 614618 72559
rect 614674 72525 614728 72581
rect 612828 72473 614728 72525
rect 612828 72457 612899 72473
rect 612955 72457 613041 72473
rect 613097 72457 613183 72473
rect 613239 72457 613325 72473
rect 613381 72457 613467 72473
rect 613523 72457 613609 72473
rect 613665 72457 613751 72473
rect 613807 72457 613893 72473
rect 613949 72457 614035 72473
rect 614091 72457 614177 72473
rect 614233 72457 614319 72473
rect 614375 72457 614461 72473
rect 614517 72457 614603 72473
rect 614659 72457 614728 72473
rect 612828 72401 612882 72457
rect 612955 72417 613006 72457
rect 613097 72417 613130 72457
rect 613239 72417 613254 72457
rect 612938 72401 613006 72417
rect 613062 72401 613130 72417
rect 613186 72401 613254 72417
rect 613310 72417 613325 72457
rect 613434 72417 613467 72457
rect 613558 72417 613609 72457
rect 613310 72401 613378 72417
rect 613434 72401 613502 72417
rect 613558 72401 613626 72417
rect 613682 72401 613750 72457
rect 613807 72417 613874 72457
rect 613949 72417 613998 72457
rect 614091 72417 614122 72457
rect 614233 72417 614246 72457
rect 613806 72401 613874 72417
rect 613930 72401 613998 72417
rect 614054 72401 614122 72417
rect 614178 72401 614246 72417
rect 614302 72417 614319 72457
rect 614426 72417 614461 72457
rect 614550 72417 614603 72457
rect 614302 72401 614370 72417
rect 614426 72401 614494 72417
rect 614550 72401 614618 72417
rect 614674 72401 614728 72457
rect 612828 72333 614728 72401
rect 612828 72277 612882 72333
rect 612938 72331 613006 72333
rect 613062 72331 613130 72333
rect 613186 72331 613254 72333
rect 612955 72277 613006 72331
rect 613097 72277 613130 72331
rect 613239 72277 613254 72331
rect 613310 72331 613378 72333
rect 613434 72331 613502 72333
rect 613558 72331 613626 72333
rect 613310 72277 613325 72331
rect 613434 72277 613467 72331
rect 613558 72277 613609 72331
rect 613682 72277 613750 72333
rect 613806 72331 613874 72333
rect 613930 72331 613998 72333
rect 614054 72331 614122 72333
rect 614178 72331 614246 72333
rect 613807 72277 613874 72331
rect 613949 72277 613998 72331
rect 614091 72277 614122 72331
rect 614233 72277 614246 72331
rect 614302 72331 614370 72333
rect 614426 72331 614494 72333
rect 614550 72331 614618 72333
rect 614302 72277 614319 72331
rect 614426 72277 614461 72331
rect 614550 72277 614603 72331
rect 614674 72277 614728 72333
rect 612828 72275 612899 72277
rect 612955 72275 613041 72277
rect 613097 72275 613183 72277
rect 613239 72275 613325 72277
rect 613381 72275 613467 72277
rect 613523 72275 613609 72277
rect 613665 72275 613751 72277
rect 613807 72275 613893 72277
rect 613949 72275 614035 72277
rect 614091 72275 614177 72277
rect 614233 72275 614319 72277
rect 614375 72275 614461 72277
rect 614517 72275 614603 72277
rect 614659 72275 614728 72277
rect 612828 72209 614728 72275
rect 612828 72153 612882 72209
rect 612938 72189 613006 72209
rect 613062 72189 613130 72209
rect 613186 72189 613254 72209
rect 612955 72153 613006 72189
rect 613097 72153 613130 72189
rect 613239 72153 613254 72189
rect 613310 72189 613378 72209
rect 613434 72189 613502 72209
rect 613558 72189 613626 72209
rect 613310 72153 613325 72189
rect 613434 72153 613467 72189
rect 613558 72153 613609 72189
rect 613682 72153 613750 72209
rect 613806 72189 613874 72209
rect 613930 72189 613998 72209
rect 614054 72189 614122 72209
rect 614178 72189 614246 72209
rect 613807 72153 613874 72189
rect 613949 72153 613998 72189
rect 614091 72153 614122 72189
rect 614233 72153 614246 72189
rect 614302 72189 614370 72209
rect 614426 72189 614494 72209
rect 614550 72189 614618 72209
rect 614302 72153 614319 72189
rect 614426 72153 614461 72189
rect 614550 72153 614603 72189
rect 614674 72153 614728 72209
rect 612828 72133 612899 72153
rect 612955 72133 613041 72153
rect 613097 72133 613183 72153
rect 613239 72133 613325 72153
rect 613381 72133 613467 72153
rect 613523 72133 613609 72153
rect 613665 72133 613751 72153
rect 613807 72133 613893 72153
rect 613949 72133 614035 72153
rect 614091 72133 614177 72153
rect 614233 72133 614319 72153
rect 614375 72133 614461 72153
rect 614517 72133 614603 72153
rect 614659 72133 614728 72153
rect 612828 72088 614728 72133
<< via3 >>
rect 379341 941655 379397 941675
rect 379483 941655 379539 941675
rect 379625 941655 379681 941675
rect 379767 941655 379823 941675
rect 379909 941655 379965 941675
rect 379341 941619 379382 941655
rect 379382 941619 379397 941655
rect 379483 941619 379506 941655
rect 379506 941619 379539 941655
rect 379625 941619 379630 941655
rect 379630 941619 379681 941655
rect 379767 941619 379822 941655
rect 379822 941619 379823 941655
rect 379909 941619 379946 941655
rect 379946 941619 379965 941655
rect 379341 941531 379397 941533
rect 379483 941531 379539 941533
rect 379625 941531 379681 941533
rect 379767 941531 379823 941533
rect 379909 941531 379965 941533
rect 379341 941477 379382 941531
rect 379382 941477 379397 941531
rect 379483 941477 379506 941531
rect 379506 941477 379539 941531
rect 379625 941477 379630 941531
rect 379630 941477 379681 941531
rect 379767 941477 379822 941531
rect 379822 941477 379823 941531
rect 379909 941477 379946 941531
rect 379946 941477 379965 941531
rect 379341 941351 379382 941391
rect 379382 941351 379397 941391
rect 379483 941351 379506 941391
rect 379506 941351 379539 941391
rect 379625 941351 379630 941391
rect 379630 941351 379681 941391
rect 379767 941351 379822 941391
rect 379822 941351 379823 941391
rect 379909 941351 379946 941391
rect 379946 941351 379965 941391
rect 379341 941335 379397 941351
rect 379483 941335 379539 941351
rect 379625 941335 379681 941351
rect 379767 941335 379823 941351
rect 379909 941335 379965 941351
rect 379341 941227 379382 941249
rect 379382 941227 379397 941249
rect 379483 941227 379506 941249
rect 379506 941227 379539 941249
rect 379625 941227 379630 941249
rect 379630 941227 379681 941249
rect 379767 941227 379822 941249
rect 379822 941227 379823 941249
rect 379909 941227 379946 941249
rect 379946 941227 379965 941249
rect 379341 941193 379397 941227
rect 379483 941193 379539 941227
rect 379625 941193 379681 941227
rect 379767 941193 379823 941227
rect 379909 941193 379965 941227
rect 379341 941103 379382 941107
rect 379382 941103 379397 941107
rect 379483 941103 379506 941107
rect 379506 941103 379539 941107
rect 379625 941103 379630 941107
rect 379630 941103 379681 941107
rect 379767 941103 379822 941107
rect 379822 941103 379823 941107
rect 379909 941103 379946 941107
rect 379946 941103 379965 941107
rect 379341 941051 379397 941103
rect 379483 941051 379539 941103
rect 379625 941051 379681 941103
rect 379767 941051 379823 941103
rect 379909 941051 379965 941103
rect 379341 940911 379397 940965
rect 379483 940911 379539 940965
rect 379625 940911 379681 940965
rect 379767 940911 379823 940965
rect 379909 940911 379965 940965
rect 379341 940909 379382 940911
rect 379382 940909 379397 940911
rect 379483 940909 379506 940911
rect 379506 940909 379539 940911
rect 379625 940909 379630 940911
rect 379630 940909 379681 940911
rect 379767 940909 379822 940911
rect 379822 940909 379823 940911
rect 379909 940909 379946 940911
rect 379946 940909 379965 940911
rect 379341 940787 379397 940823
rect 379483 940787 379539 940823
rect 379625 940787 379681 940823
rect 379767 940787 379823 940823
rect 379909 940787 379965 940823
rect 379341 940767 379382 940787
rect 379382 940767 379397 940787
rect 379483 940767 379506 940787
rect 379506 940767 379539 940787
rect 379625 940767 379630 940787
rect 379630 940767 379681 940787
rect 379767 940767 379822 940787
rect 379822 940767 379823 940787
rect 379909 940767 379946 940787
rect 379946 940767 379965 940787
rect 379341 940663 379397 940681
rect 379483 940663 379539 940681
rect 379625 940663 379681 940681
rect 379767 940663 379823 940681
rect 379909 940663 379965 940681
rect 379341 940625 379382 940663
rect 379382 940625 379397 940663
rect 379483 940625 379506 940663
rect 379506 940625 379539 940663
rect 379625 940625 379630 940663
rect 379630 940625 379681 940663
rect 379767 940625 379822 940663
rect 379822 940625 379823 940663
rect 379909 940625 379946 940663
rect 379946 940625 379965 940663
rect 379341 940483 379382 940539
rect 379382 940483 379397 940539
rect 379483 940483 379506 940539
rect 379506 940483 379539 940539
rect 379625 940483 379630 940539
rect 379630 940483 379681 940539
rect 379767 940483 379822 940539
rect 379822 940483 379823 940539
rect 379909 940483 379946 940539
rect 379946 940483 379965 940539
rect 379341 940359 379382 940397
rect 379382 940359 379397 940397
rect 379483 940359 379506 940397
rect 379506 940359 379539 940397
rect 379625 940359 379630 940397
rect 379630 940359 379681 940397
rect 379767 940359 379822 940397
rect 379822 940359 379823 940397
rect 379909 940359 379946 940397
rect 379946 940359 379965 940397
rect 379341 940341 379397 940359
rect 379483 940341 379539 940359
rect 379625 940341 379681 940359
rect 379767 940341 379823 940359
rect 379909 940341 379965 940359
rect 379341 940235 379382 940255
rect 379382 940235 379397 940255
rect 379483 940235 379506 940255
rect 379506 940235 379539 940255
rect 379625 940235 379630 940255
rect 379630 940235 379681 940255
rect 379767 940235 379822 940255
rect 379822 940235 379823 940255
rect 379909 940235 379946 940255
rect 379946 940235 379965 940255
rect 379341 940199 379397 940235
rect 379483 940199 379539 940235
rect 379625 940199 379681 940235
rect 379767 940199 379823 940235
rect 379909 940199 379965 940235
rect 379341 940111 379382 940113
rect 379382 940111 379397 940113
rect 379483 940111 379506 940113
rect 379506 940111 379539 940113
rect 379625 940111 379630 940113
rect 379630 940111 379681 940113
rect 379767 940111 379822 940113
rect 379822 940111 379823 940113
rect 379909 940111 379946 940113
rect 379946 940111 379965 940113
rect 379341 940057 379397 940111
rect 379483 940057 379539 940111
rect 379625 940057 379681 940111
rect 379767 940057 379823 940111
rect 379909 940057 379965 940111
rect 379341 939919 379397 939971
rect 379483 939919 379539 939971
rect 379625 939919 379681 939971
rect 379767 939919 379823 939971
rect 379909 939919 379965 939971
rect 379341 939915 379382 939919
rect 379382 939915 379397 939919
rect 379483 939915 379506 939919
rect 379506 939915 379539 939919
rect 379625 939915 379630 939919
rect 379630 939915 379681 939919
rect 379767 939915 379822 939919
rect 379822 939915 379823 939919
rect 379909 939915 379946 939919
rect 379946 939915 379965 939919
rect 379341 939773 379397 939829
rect 379483 939773 379539 939829
rect 379625 939773 379681 939829
rect 379767 939773 379823 939829
rect 379909 939773 379965 939829
rect 381829 941655 381885 941675
rect 381971 941655 382027 941675
rect 382113 941655 382169 941675
rect 382255 941655 382311 941675
rect 382397 941655 382453 941675
rect 382539 941655 382595 941675
rect 382681 941655 382737 941675
rect 382823 941655 382879 941675
rect 382965 941655 383021 941675
rect 383107 941655 383163 941675
rect 383249 941655 383305 941675
rect 383391 941655 383447 941675
rect 383533 941655 383589 941675
rect 383675 941655 383731 941675
rect 381829 941619 381832 941655
rect 381832 941619 381885 941655
rect 381971 941619 382012 941655
rect 382012 941619 382027 941655
rect 382113 941619 382136 941655
rect 382136 941619 382169 941655
rect 382255 941619 382260 941655
rect 382260 941619 382311 941655
rect 382397 941619 382452 941655
rect 382452 941619 382453 941655
rect 382539 941619 382576 941655
rect 382576 941619 382595 941655
rect 382681 941619 382700 941655
rect 382700 941619 382737 941655
rect 382823 941619 382824 941655
rect 382824 941619 382879 941655
rect 382965 941619 383004 941655
rect 383004 941619 383021 941655
rect 383107 941619 383128 941655
rect 383128 941619 383163 941655
rect 383249 941619 383252 941655
rect 383252 941619 383305 941655
rect 383391 941619 383444 941655
rect 383444 941619 383447 941655
rect 383533 941619 383568 941655
rect 383568 941619 383589 941655
rect 383675 941619 383692 941655
rect 383692 941619 383731 941655
rect 381829 941531 381885 941533
rect 381971 941531 382027 941533
rect 382113 941531 382169 941533
rect 382255 941531 382311 941533
rect 382397 941531 382453 941533
rect 382539 941531 382595 941533
rect 382681 941531 382737 941533
rect 382823 941531 382879 941533
rect 382965 941531 383021 941533
rect 383107 941531 383163 941533
rect 383249 941531 383305 941533
rect 383391 941531 383447 941533
rect 383533 941531 383589 941533
rect 383675 941531 383731 941533
rect 381829 941477 381832 941531
rect 381832 941477 381885 941531
rect 381971 941477 382012 941531
rect 382012 941477 382027 941531
rect 382113 941477 382136 941531
rect 382136 941477 382169 941531
rect 382255 941477 382260 941531
rect 382260 941477 382311 941531
rect 382397 941477 382452 941531
rect 382452 941477 382453 941531
rect 382539 941477 382576 941531
rect 382576 941477 382595 941531
rect 382681 941477 382700 941531
rect 382700 941477 382737 941531
rect 382823 941477 382824 941531
rect 382824 941477 382879 941531
rect 382965 941477 383004 941531
rect 383004 941477 383021 941531
rect 383107 941477 383128 941531
rect 383128 941477 383163 941531
rect 383249 941477 383252 941531
rect 383252 941477 383305 941531
rect 383391 941477 383444 941531
rect 383444 941477 383447 941531
rect 383533 941477 383568 941531
rect 383568 941477 383589 941531
rect 383675 941477 383692 941531
rect 383692 941477 383731 941531
rect 381829 941351 381832 941391
rect 381832 941351 381885 941391
rect 381971 941351 382012 941391
rect 382012 941351 382027 941391
rect 382113 941351 382136 941391
rect 382136 941351 382169 941391
rect 382255 941351 382260 941391
rect 382260 941351 382311 941391
rect 382397 941351 382452 941391
rect 382452 941351 382453 941391
rect 382539 941351 382576 941391
rect 382576 941351 382595 941391
rect 382681 941351 382700 941391
rect 382700 941351 382737 941391
rect 382823 941351 382824 941391
rect 382824 941351 382879 941391
rect 382965 941351 383004 941391
rect 383004 941351 383021 941391
rect 383107 941351 383128 941391
rect 383128 941351 383163 941391
rect 383249 941351 383252 941391
rect 383252 941351 383305 941391
rect 383391 941351 383444 941391
rect 383444 941351 383447 941391
rect 383533 941351 383568 941391
rect 383568 941351 383589 941391
rect 383675 941351 383692 941391
rect 383692 941351 383731 941391
rect 381829 941335 381885 941351
rect 381971 941335 382027 941351
rect 382113 941335 382169 941351
rect 382255 941335 382311 941351
rect 382397 941335 382453 941351
rect 382539 941335 382595 941351
rect 382681 941335 382737 941351
rect 382823 941335 382879 941351
rect 382965 941335 383021 941351
rect 383107 941335 383163 941351
rect 383249 941335 383305 941351
rect 383391 941335 383447 941351
rect 383533 941335 383589 941351
rect 383675 941335 383731 941351
rect 381829 941227 381832 941249
rect 381832 941227 381885 941249
rect 381971 941227 382012 941249
rect 382012 941227 382027 941249
rect 382113 941227 382136 941249
rect 382136 941227 382169 941249
rect 382255 941227 382260 941249
rect 382260 941227 382311 941249
rect 382397 941227 382452 941249
rect 382452 941227 382453 941249
rect 382539 941227 382576 941249
rect 382576 941227 382595 941249
rect 382681 941227 382700 941249
rect 382700 941227 382737 941249
rect 382823 941227 382824 941249
rect 382824 941227 382879 941249
rect 382965 941227 383004 941249
rect 383004 941227 383021 941249
rect 383107 941227 383128 941249
rect 383128 941227 383163 941249
rect 383249 941227 383252 941249
rect 383252 941227 383305 941249
rect 383391 941227 383444 941249
rect 383444 941227 383447 941249
rect 383533 941227 383568 941249
rect 383568 941227 383589 941249
rect 383675 941227 383692 941249
rect 383692 941227 383731 941249
rect 381829 941193 381885 941227
rect 381971 941193 382027 941227
rect 382113 941193 382169 941227
rect 382255 941193 382311 941227
rect 382397 941193 382453 941227
rect 382539 941193 382595 941227
rect 382681 941193 382737 941227
rect 382823 941193 382879 941227
rect 382965 941193 383021 941227
rect 383107 941193 383163 941227
rect 383249 941193 383305 941227
rect 383391 941193 383447 941227
rect 383533 941193 383589 941227
rect 383675 941193 383731 941227
rect 381829 941103 381832 941107
rect 381832 941103 381885 941107
rect 381971 941103 382012 941107
rect 382012 941103 382027 941107
rect 382113 941103 382136 941107
rect 382136 941103 382169 941107
rect 382255 941103 382260 941107
rect 382260 941103 382311 941107
rect 382397 941103 382452 941107
rect 382452 941103 382453 941107
rect 382539 941103 382576 941107
rect 382576 941103 382595 941107
rect 382681 941103 382700 941107
rect 382700 941103 382737 941107
rect 382823 941103 382824 941107
rect 382824 941103 382879 941107
rect 382965 941103 383004 941107
rect 383004 941103 383021 941107
rect 383107 941103 383128 941107
rect 383128 941103 383163 941107
rect 383249 941103 383252 941107
rect 383252 941103 383305 941107
rect 383391 941103 383444 941107
rect 383444 941103 383447 941107
rect 383533 941103 383568 941107
rect 383568 941103 383589 941107
rect 383675 941103 383692 941107
rect 383692 941103 383731 941107
rect 381829 941051 381885 941103
rect 381971 941051 382027 941103
rect 382113 941051 382169 941103
rect 382255 941051 382311 941103
rect 382397 941051 382453 941103
rect 382539 941051 382595 941103
rect 382681 941051 382737 941103
rect 382823 941051 382879 941103
rect 382965 941051 383021 941103
rect 383107 941051 383163 941103
rect 383249 941051 383305 941103
rect 383391 941051 383447 941103
rect 383533 941051 383589 941103
rect 383675 941051 383731 941103
rect 381829 940911 381885 940965
rect 381971 940911 382027 940965
rect 382113 940911 382169 940965
rect 382255 940911 382311 940965
rect 382397 940911 382453 940965
rect 382539 940911 382595 940965
rect 382681 940911 382737 940965
rect 382823 940911 382879 940965
rect 382965 940911 383021 940965
rect 383107 940911 383163 940965
rect 383249 940911 383305 940965
rect 383391 940911 383447 940965
rect 383533 940911 383589 940965
rect 383675 940911 383731 940965
rect 381829 940909 381832 940911
rect 381832 940909 381885 940911
rect 381971 940909 382012 940911
rect 382012 940909 382027 940911
rect 382113 940909 382136 940911
rect 382136 940909 382169 940911
rect 382255 940909 382260 940911
rect 382260 940909 382311 940911
rect 382397 940909 382452 940911
rect 382452 940909 382453 940911
rect 382539 940909 382576 940911
rect 382576 940909 382595 940911
rect 382681 940909 382700 940911
rect 382700 940909 382737 940911
rect 382823 940909 382824 940911
rect 382824 940909 382879 940911
rect 382965 940909 383004 940911
rect 383004 940909 383021 940911
rect 383107 940909 383128 940911
rect 383128 940909 383163 940911
rect 383249 940909 383252 940911
rect 383252 940909 383305 940911
rect 383391 940909 383444 940911
rect 383444 940909 383447 940911
rect 383533 940909 383568 940911
rect 383568 940909 383589 940911
rect 383675 940909 383692 940911
rect 383692 940909 383731 940911
rect 381829 940787 381885 940823
rect 381971 940787 382027 940823
rect 382113 940787 382169 940823
rect 382255 940787 382311 940823
rect 382397 940787 382453 940823
rect 382539 940787 382595 940823
rect 382681 940787 382737 940823
rect 382823 940787 382879 940823
rect 382965 940787 383021 940823
rect 383107 940787 383163 940823
rect 383249 940787 383305 940823
rect 383391 940787 383447 940823
rect 383533 940787 383589 940823
rect 383675 940787 383731 940823
rect 381829 940767 381832 940787
rect 381832 940767 381885 940787
rect 381971 940767 382012 940787
rect 382012 940767 382027 940787
rect 382113 940767 382136 940787
rect 382136 940767 382169 940787
rect 382255 940767 382260 940787
rect 382260 940767 382311 940787
rect 382397 940767 382452 940787
rect 382452 940767 382453 940787
rect 382539 940767 382576 940787
rect 382576 940767 382595 940787
rect 382681 940767 382700 940787
rect 382700 940767 382737 940787
rect 382823 940767 382824 940787
rect 382824 940767 382879 940787
rect 382965 940767 383004 940787
rect 383004 940767 383021 940787
rect 383107 940767 383128 940787
rect 383128 940767 383163 940787
rect 383249 940767 383252 940787
rect 383252 940767 383305 940787
rect 383391 940767 383444 940787
rect 383444 940767 383447 940787
rect 383533 940767 383568 940787
rect 383568 940767 383589 940787
rect 383675 940767 383692 940787
rect 383692 940767 383731 940787
rect 381829 940663 381885 940681
rect 381971 940663 382027 940681
rect 382113 940663 382169 940681
rect 382255 940663 382311 940681
rect 382397 940663 382453 940681
rect 382539 940663 382595 940681
rect 382681 940663 382737 940681
rect 382823 940663 382879 940681
rect 382965 940663 383021 940681
rect 383107 940663 383163 940681
rect 383249 940663 383305 940681
rect 383391 940663 383447 940681
rect 383533 940663 383589 940681
rect 383675 940663 383731 940681
rect 381829 940625 381832 940663
rect 381832 940625 381885 940663
rect 381971 940625 382012 940663
rect 382012 940625 382027 940663
rect 382113 940625 382136 940663
rect 382136 940625 382169 940663
rect 382255 940625 382260 940663
rect 382260 940625 382311 940663
rect 382397 940625 382452 940663
rect 382452 940625 382453 940663
rect 382539 940625 382576 940663
rect 382576 940625 382595 940663
rect 382681 940625 382700 940663
rect 382700 940625 382737 940663
rect 382823 940625 382824 940663
rect 382824 940625 382879 940663
rect 382965 940625 383004 940663
rect 383004 940625 383021 940663
rect 383107 940625 383128 940663
rect 383128 940625 383163 940663
rect 383249 940625 383252 940663
rect 383252 940625 383305 940663
rect 383391 940625 383444 940663
rect 383444 940625 383447 940663
rect 383533 940625 383568 940663
rect 383568 940625 383589 940663
rect 383675 940625 383692 940663
rect 383692 940625 383731 940663
rect 381829 940483 381832 940539
rect 381832 940483 381885 940539
rect 381971 940483 382012 940539
rect 382012 940483 382027 940539
rect 382113 940483 382136 940539
rect 382136 940483 382169 940539
rect 382255 940483 382260 940539
rect 382260 940483 382311 940539
rect 382397 940483 382452 940539
rect 382452 940483 382453 940539
rect 382539 940483 382576 940539
rect 382576 940483 382595 940539
rect 382681 940483 382700 940539
rect 382700 940483 382737 940539
rect 382823 940483 382824 940539
rect 382824 940483 382879 940539
rect 382965 940483 383004 940539
rect 383004 940483 383021 940539
rect 383107 940483 383128 940539
rect 383128 940483 383163 940539
rect 383249 940483 383252 940539
rect 383252 940483 383305 940539
rect 383391 940483 383444 940539
rect 383444 940483 383447 940539
rect 383533 940483 383568 940539
rect 383568 940483 383589 940539
rect 383675 940483 383692 940539
rect 383692 940483 383731 940539
rect 381829 940359 381832 940397
rect 381832 940359 381885 940397
rect 381971 940359 382012 940397
rect 382012 940359 382027 940397
rect 382113 940359 382136 940397
rect 382136 940359 382169 940397
rect 382255 940359 382260 940397
rect 382260 940359 382311 940397
rect 382397 940359 382452 940397
rect 382452 940359 382453 940397
rect 382539 940359 382576 940397
rect 382576 940359 382595 940397
rect 382681 940359 382700 940397
rect 382700 940359 382737 940397
rect 382823 940359 382824 940397
rect 382824 940359 382879 940397
rect 382965 940359 383004 940397
rect 383004 940359 383021 940397
rect 383107 940359 383128 940397
rect 383128 940359 383163 940397
rect 383249 940359 383252 940397
rect 383252 940359 383305 940397
rect 383391 940359 383444 940397
rect 383444 940359 383447 940397
rect 383533 940359 383568 940397
rect 383568 940359 383589 940397
rect 383675 940359 383692 940397
rect 383692 940359 383731 940397
rect 381829 940341 381885 940359
rect 381971 940341 382027 940359
rect 382113 940341 382169 940359
rect 382255 940341 382311 940359
rect 382397 940341 382453 940359
rect 382539 940341 382595 940359
rect 382681 940341 382737 940359
rect 382823 940341 382879 940359
rect 382965 940341 383021 940359
rect 383107 940341 383163 940359
rect 383249 940341 383305 940359
rect 383391 940341 383447 940359
rect 383533 940341 383589 940359
rect 383675 940341 383731 940359
rect 381829 940235 381832 940255
rect 381832 940235 381885 940255
rect 381971 940235 382012 940255
rect 382012 940235 382027 940255
rect 382113 940235 382136 940255
rect 382136 940235 382169 940255
rect 382255 940235 382260 940255
rect 382260 940235 382311 940255
rect 382397 940235 382452 940255
rect 382452 940235 382453 940255
rect 382539 940235 382576 940255
rect 382576 940235 382595 940255
rect 382681 940235 382700 940255
rect 382700 940235 382737 940255
rect 382823 940235 382824 940255
rect 382824 940235 382879 940255
rect 382965 940235 383004 940255
rect 383004 940235 383021 940255
rect 383107 940235 383128 940255
rect 383128 940235 383163 940255
rect 383249 940235 383252 940255
rect 383252 940235 383305 940255
rect 383391 940235 383444 940255
rect 383444 940235 383447 940255
rect 383533 940235 383568 940255
rect 383568 940235 383589 940255
rect 383675 940235 383692 940255
rect 383692 940235 383731 940255
rect 381829 940199 381885 940235
rect 381971 940199 382027 940235
rect 382113 940199 382169 940235
rect 382255 940199 382311 940235
rect 382397 940199 382453 940235
rect 382539 940199 382595 940235
rect 382681 940199 382737 940235
rect 382823 940199 382879 940235
rect 382965 940199 383021 940235
rect 383107 940199 383163 940235
rect 383249 940199 383305 940235
rect 383391 940199 383447 940235
rect 383533 940199 383589 940235
rect 383675 940199 383731 940235
rect 381829 940111 381832 940113
rect 381832 940111 381885 940113
rect 381971 940111 382012 940113
rect 382012 940111 382027 940113
rect 382113 940111 382136 940113
rect 382136 940111 382169 940113
rect 382255 940111 382260 940113
rect 382260 940111 382311 940113
rect 382397 940111 382452 940113
rect 382452 940111 382453 940113
rect 382539 940111 382576 940113
rect 382576 940111 382595 940113
rect 382681 940111 382700 940113
rect 382700 940111 382737 940113
rect 382823 940111 382824 940113
rect 382824 940111 382879 940113
rect 382965 940111 383004 940113
rect 383004 940111 383021 940113
rect 383107 940111 383128 940113
rect 383128 940111 383163 940113
rect 383249 940111 383252 940113
rect 383252 940111 383305 940113
rect 383391 940111 383444 940113
rect 383444 940111 383447 940113
rect 383533 940111 383568 940113
rect 383568 940111 383589 940113
rect 383675 940111 383692 940113
rect 383692 940111 383731 940113
rect 381829 940057 381885 940111
rect 381971 940057 382027 940111
rect 382113 940057 382169 940111
rect 382255 940057 382311 940111
rect 382397 940057 382453 940111
rect 382539 940057 382595 940111
rect 382681 940057 382737 940111
rect 382823 940057 382879 940111
rect 382965 940057 383021 940111
rect 383107 940057 383163 940111
rect 383249 940057 383305 940111
rect 383391 940057 383447 940111
rect 383533 940057 383589 940111
rect 383675 940057 383731 940111
rect 381829 939919 381885 939971
rect 381971 939919 382027 939971
rect 382113 939919 382169 939971
rect 382255 939919 382311 939971
rect 382397 939919 382453 939971
rect 382539 939919 382595 939971
rect 382681 939919 382737 939971
rect 382823 939919 382879 939971
rect 382965 939919 383021 939971
rect 383107 939919 383163 939971
rect 383249 939919 383305 939971
rect 383391 939919 383447 939971
rect 383533 939919 383589 939971
rect 383675 939919 383731 939971
rect 381829 939915 381832 939919
rect 381832 939915 381885 939919
rect 381971 939915 382012 939919
rect 382012 939915 382027 939919
rect 382113 939915 382136 939919
rect 382136 939915 382169 939919
rect 382255 939915 382260 939919
rect 382260 939915 382311 939919
rect 382397 939915 382452 939919
rect 382452 939915 382453 939919
rect 382539 939915 382576 939919
rect 382576 939915 382595 939919
rect 382681 939915 382700 939919
rect 382700 939915 382737 939919
rect 382823 939915 382824 939919
rect 382824 939915 382879 939919
rect 382965 939915 383004 939919
rect 383004 939915 383021 939919
rect 383107 939915 383128 939919
rect 383128 939915 383163 939919
rect 383249 939915 383252 939919
rect 383252 939915 383305 939919
rect 383391 939915 383444 939919
rect 383444 939915 383447 939919
rect 383533 939915 383568 939919
rect 383568 939915 383589 939919
rect 383675 939915 383692 939919
rect 383692 939915 383731 939919
rect 381829 939773 381885 939829
rect 381971 939773 382027 939829
rect 382113 939773 382169 939829
rect 382255 939773 382311 939829
rect 382397 939773 382453 939829
rect 382539 939773 382595 939829
rect 382681 939773 382737 939829
rect 382823 939773 382879 939829
rect 382965 939773 383021 939829
rect 383107 939773 383163 939829
rect 383249 939773 383305 939829
rect 383391 939773 383447 939829
rect 383533 939773 383589 939829
rect 383675 939773 383731 939829
rect 384199 941655 384255 941675
rect 384341 941655 384397 941675
rect 384483 941655 384539 941675
rect 384625 941655 384681 941675
rect 384767 941655 384823 941675
rect 384909 941655 384965 941675
rect 385051 941655 385107 941675
rect 385193 941655 385249 941675
rect 385335 941655 385391 941675
rect 385477 941655 385533 941675
rect 385619 941655 385675 941675
rect 385761 941655 385817 941675
rect 385903 941655 385959 941675
rect 386045 941655 386101 941675
rect 384199 941619 384202 941655
rect 384202 941619 384255 941655
rect 384341 941619 384382 941655
rect 384382 941619 384397 941655
rect 384483 941619 384506 941655
rect 384506 941619 384539 941655
rect 384625 941619 384630 941655
rect 384630 941619 384681 941655
rect 384767 941619 384822 941655
rect 384822 941619 384823 941655
rect 384909 941619 384946 941655
rect 384946 941619 384965 941655
rect 385051 941619 385070 941655
rect 385070 941619 385107 941655
rect 385193 941619 385194 941655
rect 385194 941619 385249 941655
rect 385335 941619 385374 941655
rect 385374 941619 385391 941655
rect 385477 941619 385498 941655
rect 385498 941619 385533 941655
rect 385619 941619 385622 941655
rect 385622 941619 385675 941655
rect 385761 941619 385814 941655
rect 385814 941619 385817 941655
rect 385903 941619 385938 941655
rect 385938 941619 385959 941655
rect 386045 941619 386062 941655
rect 386062 941619 386101 941655
rect 384199 941531 384255 941533
rect 384341 941531 384397 941533
rect 384483 941531 384539 941533
rect 384625 941531 384681 941533
rect 384767 941531 384823 941533
rect 384909 941531 384965 941533
rect 385051 941531 385107 941533
rect 385193 941531 385249 941533
rect 385335 941531 385391 941533
rect 385477 941531 385533 941533
rect 385619 941531 385675 941533
rect 385761 941531 385817 941533
rect 385903 941531 385959 941533
rect 386045 941531 386101 941533
rect 384199 941477 384202 941531
rect 384202 941477 384255 941531
rect 384341 941477 384382 941531
rect 384382 941477 384397 941531
rect 384483 941477 384506 941531
rect 384506 941477 384539 941531
rect 384625 941477 384630 941531
rect 384630 941477 384681 941531
rect 384767 941477 384822 941531
rect 384822 941477 384823 941531
rect 384909 941477 384946 941531
rect 384946 941477 384965 941531
rect 385051 941477 385070 941531
rect 385070 941477 385107 941531
rect 385193 941477 385194 941531
rect 385194 941477 385249 941531
rect 385335 941477 385374 941531
rect 385374 941477 385391 941531
rect 385477 941477 385498 941531
rect 385498 941477 385533 941531
rect 385619 941477 385622 941531
rect 385622 941477 385675 941531
rect 385761 941477 385814 941531
rect 385814 941477 385817 941531
rect 385903 941477 385938 941531
rect 385938 941477 385959 941531
rect 386045 941477 386062 941531
rect 386062 941477 386101 941531
rect 384199 941351 384202 941391
rect 384202 941351 384255 941391
rect 384341 941351 384382 941391
rect 384382 941351 384397 941391
rect 384483 941351 384506 941391
rect 384506 941351 384539 941391
rect 384625 941351 384630 941391
rect 384630 941351 384681 941391
rect 384767 941351 384822 941391
rect 384822 941351 384823 941391
rect 384909 941351 384946 941391
rect 384946 941351 384965 941391
rect 385051 941351 385070 941391
rect 385070 941351 385107 941391
rect 385193 941351 385194 941391
rect 385194 941351 385249 941391
rect 385335 941351 385374 941391
rect 385374 941351 385391 941391
rect 385477 941351 385498 941391
rect 385498 941351 385533 941391
rect 385619 941351 385622 941391
rect 385622 941351 385675 941391
rect 385761 941351 385814 941391
rect 385814 941351 385817 941391
rect 385903 941351 385938 941391
rect 385938 941351 385959 941391
rect 386045 941351 386062 941391
rect 386062 941351 386101 941391
rect 384199 941335 384255 941351
rect 384341 941335 384397 941351
rect 384483 941335 384539 941351
rect 384625 941335 384681 941351
rect 384767 941335 384823 941351
rect 384909 941335 384965 941351
rect 385051 941335 385107 941351
rect 385193 941335 385249 941351
rect 385335 941335 385391 941351
rect 385477 941335 385533 941351
rect 385619 941335 385675 941351
rect 385761 941335 385817 941351
rect 385903 941335 385959 941351
rect 386045 941335 386101 941351
rect 384199 941227 384202 941249
rect 384202 941227 384255 941249
rect 384341 941227 384382 941249
rect 384382 941227 384397 941249
rect 384483 941227 384506 941249
rect 384506 941227 384539 941249
rect 384625 941227 384630 941249
rect 384630 941227 384681 941249
rect 384767 941227 384822 941249
rect 384822 941227 384823 941249
rect 384909 941227 384946 941249
rect 384946 941227 384965 941249
rect 385051 941227 385070 941249
rect 385070 941227 385107 941249
rect 385193 941227 385194 941249
rect 385194 941227 385249 941249
rect 385335 941227 385374 941249
rect 385374 941227 385391 941249
rect 385477 941227 385498 941249
rect 385498 941227 385533 941249
rect 385619 941227 385622 941249
rect 385622 941227 385675 941249
rect 385761 941227 385814 941249
rect 385814 941227 385817 941249
rect 385903 941227 385938 941249
rect 385938 941227 385959 941249
rect 386045 941227 386062 941249
rect 386062 941227 386101 941249
rect 384199 941193 384255 941227
rect 384341 941193 384397 941227
rect 384483 941193 384539 941227
rect 384625 941193 384681 941227
rect 384767 941193 384823 941227
rect 384909 941193 384965 941227
rect 385051 941193 385107 941227
rect 385193 941193 385249 941227
rect 385335 941193 385391 941227
rect 385477 941193 385533 941227
rect 385619 941193 385675 941227
rect 385761 941193 385817 941227
rect 385903 941193 385959 941227
rect 386045 941193 386101 941227
rect 384199 941103 384202 941107
rect 384202 941103 384255 941107
rect 384341 941103 384382 941107
rect 384382 941103 384397 941107
rect 384483 941103 384506 941107
rect 384506 941103 384539 941107
rect 384625 941103 384630 941107
rect 384630 941103 384681 941107
rect 384767 941103 384822 941107
rect 384822 941103 384823 941107
rect 384909 941103 384946 941107
rect 384946 941103 384965 941107
rect 385051 941103 385070 941107
rect 385070 941103 385107 941107
rect 385193 941103 385194 941107
rect 385194 941103 385249 941107
rect 385335 941103 385374 941107
rect 385374 941103 385391 941107
rect 385477 941103 385498 941107
rect 385498 941103 385533 941107
rect 385619 941103 385622 941107
rect 385622 941103 385675 941107
rect 385761 941103 385814 941107
rect 385814 941103 385817 941107
rect 385903 941103 385938 941107
rect 385938 941103 385959 941107
rect 386045 941103 386062 941107
rect 386062 941103 386101 941107
rect 384199 941051 384255 941103
rect 384341 941051 384397 941103
rect 384483 941051 384539 941103
rect 384625 941051 384681 941103
rect 384767 941051 384823 941103
rect 384909 941051 384965 941103
rect 385051 941051 385107 941103
rect 385193 941051 385249 941103
rect 385335 941051 385391 941103
rect 385477 941051 385533 941103
rect 385619 941051 385675 941103
rect 385761 941051 385817 941103
rect 385903 941051 385959 941103
rect 386045 941051 386101 941103
rect 384199 940911 384255 940965
rect 384341 940911 384397 940965
rect 384483 940911 384539 940965
rect 384625 940911 384681 940965
rect 384767 940911 384823 940965
rect 384909 940911 384965 940965
rect 385051 940911 385107 940965
rect 385193 940911 385249 940965
rect 385335 940911 385391 940965
rect 385477 940911 385533 940965
rect 385619 940911 385675 940965
rect 385761 940911 385817 940965
rect 385903 940911 385959 940965
rect 386045 940911 386101 940965
rect 384199 940909 384202 940911
rect 384202 940909 384255 940911
rect 384341 940909 384382 940911
rect 384382 940909 384397 940911
rect 384483 940909 384506 940911
rect 384506 940909 384539 940911
rect 384625 940909 384630 940911
rect 384630 940909 384681 940911
rect 384767 940909 384822 940911
rect 384822 940909 384823 940911
rect 384909 940909 384946 940911
rect 384946 940909 384965 940911
rect 385051 940909 385070 940911
rect 385070 940909 385107 940911
rect 385193 940909 385194 940911
rect 385194 940909 385249 940911
rect 385335 940909 385374 940911
rect 385374 940909 385391 940911
rect 385477 940909 385498 940911
rect 385498 940909 385533 940911
rect 385619 940909 385622 940911
rect 385622 940909 385675 940911
rect 385761 940909 385814 940911
rect 385814 940909 385817 940911
rect 385903 940909 385938 940911
rect 385938 940909 385959 940911
rect 386045 940909 386062 940911
rect 386062 940909 386101 940911
rect 384199 940787 384255 940823
rect 384341 940787 384397 940823
rect 384483 940787 384539 940823
rect 384625 940787 384681 940823
rect 384767 940787 384823 940823
rect 384909 940787 384965 940823
rect 385051 940787 385107 940823
rect 385193 940787 385249 940823
rect 385335 940787 385391 940823
rect 385477 940787 385533 940823
rect 385619 940787 385675 940823
rect 385761 940787 385817 940823
rect 385903 940787 385959 940823
rect 386045 940787 386101 940823
rect 384199 940767 384202 940787
rect 384202 940767 384255 940787
rect 384341 940767 384382 940787
rect 384382 940767 384397 940787
rect 384483 940767 384506 940787
rect 384506 940767 384539 940787
rect 384625 940767 384630 940787
rect 384630 940767 384681 940787
rect 384767 940767 384822 940787
rect 384822 940767 384823 940787
rect 384909 940767 384946 940787
rect 384946 940767 384965 940787
rect 385051 940767 385070 940787
rect 385070 940767 385107 940787
rect 385193 940767 385194 940787
rect 385194 940767 385249 940787
rect 385335 940767 385374 940787
rect 385374 940767 385391 940787
rect 385477 940767 385498 940787
rect 385498 940767 385533 940787
rect 385619 940767 385622 940787
rect 385622 940767 385675 940787
rect 385761 940767 385814 940787
rect 385814 940767 385817 940787
rect 385903 940767 385938 940787
rect 385938 940767 385959 940787
rect 386045 940767 386062 940787
rect 386062 940767 386101 940787
rect 384199 940663 384255 940681
rect 384341 940663 384397 940681
rect 384483 940663 384539 940681
rect 384625 940663 384681 940681
rect 384767 940663 384823 940681
rect 384909 940663 384965 940681
rect 385051 940663 385107 940681
rect 385193 940663 385249 940681
rect 385335 940663 385391 940681
rect 385477 940663 385533 940681
rect 385619 940663 385675 940681
rect 385761 940663 385817 940681
rect 385903 940663 385959 940681
rect 386045 940663 386101 940681
rect 384199 940625 384202 940663
rect 384202 940625 384255 940663
rect 384341 940625 384382 940663
rect 384382 940625 384397 940663
rect 384483 940625 384506 940663
rect 384506 940625 384539 940663
rect 384625 940625 384630 940663
rect 384630 940625 384681 940663
rect 384767 940625 384822 940663
rect 384822 940625 384823 940663
rect 384909 940625 384946 940663
rect 384946 940625 384965 940663
rect 385051 940625 385070 940663
rect 385070 940625 385107 940663
rect 385193 940625 385194 940663
rect 385194 940625 385249 940663
rect 385335 940625 385374 940663
rect 385374 940625 385391 940663
rect 385477 940625 385498 940663
rect 385498 940625 385533 940663
rect 385619 940625 385622 940663
rect 385622 940625 385675 940663
rect 385761 940625 385814 940663
rect 385814 940625 385817 940663
rect 385903 940625 385938 940663
rect 385938 940625 385959 940663
rect 386045 940625 386062 940663
rect 386062 940625 386101 940663
rect 384199 940483 384202 940539
rect 384202 940483 384255 940539
rect 384341 940483 384382 940539
rect 384382 940483 384397 940539
rect 384483 940483 384506 940539
rect 384506 940483 384539 940539
rect 384625 940483 384630 940539
rect 384630 940483 384681 940539
rect 384767 940483 384822 940539
rect 384822 940483 384823 940539
rect 384909 940483 384946 940539
rect 384946 940483 384965 940539
rect 385051 940483 385070 940539
rect 385070 940483 385107 940539
rect 385193 940483 385194 940539
rect 385194 940483 385249 940539
rect 385335 940483 385374 940539
rect 385374 940483 385391 940539
rect 385477 940483 385498 940539
rect 385498 940483 385533 940539
rect 385619 940483 385622 940539
rect 385622 940483 385675 940539
rect 385761 940483 385814 940539
rect 385814 940483 385817 940539
rect 385903 940483 385938 940539
rect 385938 940483 385959 940539
rect 386045 940483 386062 940539
rect 386062 940483 386101 940539
rect 384199 940359 384202 940397
rect 384202 940359 384255 940397
rect 384341 940359 384382 940397
rect 384382 940359 384397 940397
rect 384483 940359 384506 940397
rect 384506 940359 384539 940397
rect 384625 940359 384630 940397
rect 384630 940359 384681 940397
rect 384767 940359 384822 940397
rect 384822 940359 384823 940397
rect 384909 940359 384946 940397
rect 384946 940359 384965 940397
rect 385051 940359 385070 940397
rect 385070 940359 385107 940397
rect 385193 940359 385194 940397
rect 385194 940359 385249 940397
rect 385335 940359 385374 940397
rect 385374 940359 385391 940397
rect 385477 940359 385498 940397
rect 385498 940359 385533 940397
rect 385619 940359 385622 940397
rect 385622 940359 385675 940397
rect 385761 940359 385814 940397
rect 385814 940359 385817 940397
rect 385903 940359 385938 940397
rect 385938 940359 385959 940397
rect 386045 940359 386062 940397
rect 386062 940359 386101 940397
rect 384199 940341 384255 940359
rect 384341 940341 384397 940359
rect 384483 940341 384539 940359
rect 384625 940341 384681 940359
rect 384767 940341 384823 940359
rect 384909 940341 384965 940359
rect 385051 940341 385107 940359
rect 385193 940341 385249 940359
rect 385335 940341 385391 940359
rect 385477 940341 385533 940359
rect 385619 940341 385675 940359
rect 385761 940341 385817 940359
rect 385903 940341 385959 940359
rect 386045 940341 386101 940359
rect 384199 940235 384202 940255
rect 384202 940235 384255 940255
rect 384341 940235 384382 940255
rect 384382 940235 384397 940255
rect 384483 940235 384506 940255
rect 384506 940235 384539 940255
rect 384625 940235 384630 940255
rect 384630 940235 384681 940255
rect 384767 940235 384822 940255
rect 384822 940235 384823 940255
rect 384909 940235 384946 940255
rect 384946 940235 384965 940255
rect 385051 940235 385070 940255
rect 385070 940235 385107 940255
rect 385193 940235 385194 940255
rect 385194 940235 385249 940255
rect 385335 940235 385374 940255
rect 385374 940235 385391 940255
rect 385477 940235 385498 940255
rect 385498 940235 385533 940255
rect 385619 940235 385622 940255
rect 385622 940235 385675 940255
rect 385761 940235 385814 940255
rect 385814 940235 385817 940255
rect 385903 940235 385938 940255
rect 385938 940235 385959 940255
rect 386045 940235 386062 940255
rect 386062 940235 386101 940255
rect 384199 940199 384255 940235
rect 384341 940199 384397 940235
rect 384483 940199 384539 940235
rect 384625 940199 384681 940235
rect 384767 940199 384823 940235
rect 384909 940199 384965 940235
rect 385051 940199 385107 940235
rect 385193 940199 385249 940235
rect 385335 940199 385391 940235
rect 385477 940199 385533 940235
rect 385619 940199 385675 940235
rect 385761 940199 385817 940235
rect 385903 940199 385959 940235
rect 386045 940199 386101 940235
rect 384199 940111 384202 940113
rect 384202 940111 384255 940113
rect 384341 940111 384382 940113
rect 384382 940111 384397 940113
rect 384483 940111 384506 940113
rect 384506 940111 384539 940113
rect 384625 940111 384630 940113
rect 384630 940111 384681 940113
rect 384767 940111 384822 940113
rect 384822 940111 384823 940113
rect 384909 940111 384946 940113
rect 384946 940111 384965 940113
rect 385051 940111 385070 940113
rect 385070 940111 385107 940113
rect 385193 940111 385194 940113
rect 385194 940111 385249 940113
rect 385335 940111 385374 940113
rect 385374 940111 385391 940113
rect 385477 940111 385498 940113
rect 385498 940111 385533 940113
rect 385619 940111 385622 940113
rect 385622 940111 385675 940113
rect 385761 940111 385814 940113
rect 385814 940111 385817 940113
rect 385903 940111 385938 940113
rect 385938 940111 385959 940113
rect 386045 940111 386062 940113
rect 386062 940111 386101 940113
rect 384199 940057 384255 940111
rect 384341 940057 384397 940111
rect 384483 940057 384539 940111
rect 384625 940057 384681 940111
rect 384767 940057 384823 940111
rect 384909 940057 384965 940111
rect 385051 940057 385107 940111
rect 385193 940057 385249 940111
rect 385335 940057 385391 940111
rect 385477 940057 385533 940111
rect 385619 940057 385675 940111
rect 385761 940057 385817 940111
rect 385903 940057 385959 940111
rect 386045 940057 386101 940111
rect 384199 939919 384255 939971
rect 384341 939919 384397 939971
rect 384483 939919 384539 939971
rect 384625 939919 384681 939971
rect 384767 939919 384823 939971
rect 384909 939919 384965 939971
rect 385051 939919 385107 939971
rect 385193 939919 385249 939971
rect 385335 939919 385391 939971
rect 385477 939919 385533 939971
rect 385619 939919 385675 939971
rect 385761 939919 385817 939971
rect 385903 939919 385959 939971
rect 386045 939919 386101 939971
rect 384199 939915 384202 939919
rect 384202 939915 384255 939919
rect 384341 939915 384382 939919
rect 384382 939915 384397 939919
rect 384483 939915 384506 939919
rect 384506 939915 384539 939919
rect 384625 939915 384630 939919
rect 384630 939915 384681 939919
rect 384767 939915 384822 939919
rect 384822 939915 384823 939919
rect 384909 939915 384946 939919
rect 384946 939915 384965 939919
rect 385051 939915 385070 939919
rect 385070 939915 385107 939919
rect 385193 939915 385194 939919
rect 385194 939915 385249 939919
rect 385335 939915 385374 939919
rect 385374 939915 385391 939919
rect 385477 939915 385498 939919
rect 385498 939915 385533 939919
rect 385619 939915 385622 939919
rect 385622 939915 385675 939919
rect 385761 939915 385814 939919
rect 385814 939915 385817 939919
rect 385903 939915 385938 939919
rect 385938 939915 385959 939919
rect 386045 939915 386062 939919
rect 386062 939915 386101 939919
rect 384199 939773 384255 939829
rect 384341 939773 384397 939829
rect 384483 939773 384539 939829
rect 384625 939773 384681 939829
rect 384767 939773 384823 939829
rect 384909 939773 384965 939829
rect 385051 939773 385107 939829
rect 385193 939773 385249 939829
rect 385335 939773 385391 939829
rect 385477 939773 385533 939829
rect 385619 939773 385675 939829
rect 385761 939773 385817 939829
rect 385903 939773 385959 939829
rect 386045 939773 386101 939829
rect 386905 941655 386961 941675
rect 387047 941655 387103 941675
rect 387189 941655 387245 941675
rect 387331 941655 387387 941675
rect 387473 941655 387529 941675
rect 387615 941655 387671 941675
rect 387757 941655 387813 941675
rect 387899 941655 387955 941675
rect 388041 941655 388097 941675
rect 388183 941655 388239 941675
rect 388325 941655 388381 941675
rect 388467 941655 388523 941675
rect 388609 941655 388665 941675
rect 388751 941655 388807 941675
rect 386905 941619 386908 941655
rect 386908 941619 386961 941655
rect 387047 941619 387088 941655
rect 387088 941619 387103 941655
rect 387189 941619 387212 941655
rect 387212 941619 387245 941655
rect 387331 941619 387336 941655
rect 387336 941619 387387 941655
rect 387473 941619 387528 941655
rect 387528 941619 387529 941655
rect 387615 941619 387652 941655
rect 387652 941619 387671 941655
rect 387757 941619 387776 941655
rect 387776 941619 387813 941655
rect 387899 941619 387900 941655
rect 387900 941619 387955 941655
rect 388041 941619 388080 941655
rect 388080 941619 388097 941655
rect 388183 941619 388204 941655
rect 388204 941619 388239 941655
rect 388325 941619 388328 941655
rect 388328 941619 388381 941655
rect 388467 941619 388520 941655
rect 388520 941619 388523 941655
rect 388609 941619 388644 941655
rect 388644 941619 388665 941655
rect 388751 941619 388768 941655
rect 388768 941619 388807 941655
rect 386905 941531 386961 941533
rect 387047 941531 387103 941533
rect 387189 941531 387245 941533
rect 387331 941531 387387 941533
rect 387473 941531 387529 941533
rect 387615 941531 387671 941533
rect 387757 941531 387813 941533
rect 387899 941531 387955 941533
rect 388041 941531 388097 941533
rect 388183 941531 388239 941533
rect 388325 941531 388381 941533
rect 388467 941531 388523 941533
rect 388609 941531 388665 941533
rect 388751 941531 388807 941533
rect 386905 941477 386908 941531
rect 386908 941477 386961 941531
rect 387047 941477 387088 941531
rect 387088 941477 387103 941531
rect 387189 941477 387212 941531
rect 387212 941477 387245 941531
rect 387331 941477 387336 941531
rect 387336 941477 387387 941531
rect 387473 941477 387528 941531
rect 387528 941477 387529 941531
rect 387615 941477 387652 941531
rect 387652 941477 387671 941531
rect 387757 941477 387776 941531
rect 387776 941477 387813 941531
rect 387899 941477 387900 941531
rect 387900 941477 387955 941531
rect 388041 941477 388080 941531
rect 388080 941477 388097 941531
rect 388183 941477 388204 941531
rect 388204 941477 388239 941531
rect 388325 941477 388328 941531
rect 388328 941477 388381 941531
rect 388467 941477 388520 941531
rect 388520 941477 388523 941531
rect 388609 941477 388644 941531
rect 388644 941477 388665 941531
rect 388751 941477 388768 941531
rect 388768 941477 388807 941531
rect 386905 941351 386908 941391
rect 386908 941351 386961 941391
rect 387047 941351 387088 941391
rect 387088 941351 387103 941391
rect 387189 941351 387212 941391
rect 387212 941351 387245 941391
rect 387331 941351 387336 941391
rect 387336 941351 387387 941391
rect 387473 941351 387528 941391
rect 387528 941351 387529 941391
rect 387615 941351 387652 941391
rect 387652 941351 387671 941391
rect 387757 941351 387776 941391
rect 387776 941351 387813 941391
rect 387899 941351 387900 941391
rect 387900 941351 387955 941391
rect 388041 941351 388080 941391
rect 388080 941351 388097 941391
rect 388183 941351 388204 941391
rect 388204 941351 388239 941391
rect 388325 941351 388328 941391
rect 388328 941351 388381 941391
rect 388467 941351 388520 941391
rect 388520 941351 388523 941391
rect 388609 941351 388644 941391
rect 388644 941351 388665 941391
rect 388751 941351 388768 941391
rect 388768 941351 388807 941391
rect 386905 941335 386961 941351
rect 387047 941335 387103 941351
rect 387189 941335 387245 941351
rect 387331 941335 387387 941351
rect 387473 941335 387529 941351
rect 387615 941335 387671 941351
rect 387757 941335 387813 941351
rect 387899 941335 387955 941351
rect 388041 941335 388097 941351
rect 388183 941335 388239 941351
rect 388325 941335 388381 941351
rect 388467 941335 388523 941351
rect 388609 941335 388665 941351
rect 388751 941335 388807 941351
rect 386905 941227 386908 941249
rect 386908 941227 386961 941249
rect 387047 941227 387088 941249
rect 387088 941227 387103 941249
rect 387189 941227 387212 941249
rect 387212 941227 387245 941249
rect 387331 941227 387336 941249
rect 387336 941227 387387 941249
rect 387473 941227 387528 941249
rect 387528 941227 387529 941249
rect 387615 941227 387652 941249
rect 387652 941227 387671 941249
rect 387757 941227 387776 941249
rect 387776 941227 387813 941249
rect 387899 941227 387900 941249
rect 387900 941227 387955 941249
rect 388041 941227 388080 941249
rect 388080 941227 388097 941249
rect 388183 941227 388204 941249
rect 388204 941227 388239 941249
rect 388325 941227 388328 941249
rect 388328 941227 388381 941249
rect 388467 941227 388520 941249
rect 388520 941227 388523 941249
rect 388609 941227 388644 941249
rect 388644 941227 388665 941249
rect 388751 941227 388768 941249
rect 388768 941227 388807 941249
rect 386905 941193 386961 941227
rect 387047 941193 387103 941227
rect 387189 941193 387245 941227
rect 387331 941193 387387 941227
rect 387473 941193 387529 941227
rect 387615 941193 387671 941227
rect 387757 941193 387813 941227
rect 387899 941193 387955 941227
rect 388041 941193 388097 941227
rect 388183 941193 388239 941227
rect 388325 941193 388381 941227
rect 388467 941193 388523 941227
rect 388609 941193 388665 941227
rect 388751 941193 388807 941227
rect 386905 941103 386908 941107
rect 386908 941103 386961 941107
rect 387047 941103 387088 941107
rect 387088 941103 387103 941107
rect 387189 941103 387212 941107
rect 387212 941103 387245 941107
rect 387331 941103 387336 941107
rect 387336 941103 387387 941107
rect 387473 941103 387528 941107
rect 387528 941103 387529 941107
rect 387615 941103 387652 941107
rect 387652 941103 387671 941107
rect 387757 941103 387776 941107
rect 387776 941103 387813 941107
rect 387899 941103 387900 941107
rect 387900 941103 387955 941107
rect 388041 941103 388080 941107
rect 388080 941103 388097 941107
rect 388183 941103 388204 941107
rect 388204 941103 388239 941107
rect 388325 941103 388328 941107
rect 388328 941103 388381 941107
rect 388467 941103 388520 941107
rect 388520 941103 388523 941107
rect 388609 941103 388644 941107
rect 388644 941103 388665 941107
rect 388751 941103 388768 941107
rect 388768 941103 388807 941107
rect 386905 941051 386961 941103
rect 387047 941051 387103 941103
rect 387189 941051 387245 941103
rect 387331 941051 387387 941103
rect 387473 941051 387529 941103
rect 387615 941051 387671 941103
rect 387757 941051 387813 941103
rect 387899 941051 387955 941103
rect 388041 941051 388097 941103
rect 388183 941051 388239 941103
rect 388325 941051 388381 941103
rect 388467 941051 388523 941103
rect 388609 941051 388665 941103
rect 388751 941051 388807 941103
rect 386905 940911 386961 940965
rect 387047 940911 387103 940965
rect 387189 940911 387245 940965
rect 387331 940911 387387 940965
rect 387473 940911 387529 940965
rect 387615 940911 387671 940965
rect 387757 940911 387813 940965
rect 387899 940911 387955 940965
rect 388041 940911 388097 940965
rect 388183 940911 388239 940965
rect 388325 940911 388381 940965
rect 388467 940911 388523 940965
rect 388609 940911 388665 940965
rect 388751 940911 388807 940965
rect 386905 940909 386908 940911
rect 386908 940909 386961 940911
rect 387047 940909 387088 940911
rect 387088 940909 387103 940911
rect 387189 940909 387212 940911
rect 387212 940909 387245 940911
rect 387331 940909 387336 940911
rect 387336 940909 387387 940911
rect 387473 940909 387528 940911
rect 387528 940909 387529 940911
rect 387615 940909 387652 940911
rect 387652 940909 387671 940911
rect 387757 940909 387776 940911
rect 387776 940909 387813 940911
rect 387899 940909 387900 940911
rect 387900 940909 387955 940911
rect 388041 940909 388080 940911
rect 388080 940909 388097 940911
rect 388183 940909 388204 940911
rect 388204 940909 388239 940911
rect 388325 940909 388328 940911
rect 388328 940909 388381 940911
rect 388467 940909 388520 940911
rect 388520 940909 388523 940911
rect 388609 940909 388644 940911
rect 388644 940909 388665 940911
rect 388751 940909 388768 940911
rect 388768 940909 388807 940911
rect 386905 940787 386961 940823
rect 387047 940787 387103 940823
rect 387189 940787 387245 940823
rect 387331 940787 387387 940823
rect 387473 940787 387529 940823
rect 387615 940787 387671 940823
rect 387757 940787 387813 940823
rect 387899 940787 387955 940823
rect 388041 940787 388097 940823
rect 388183 940787 388239 940823
rect 388325 940787 388381 940823
rect 388467 940787 388523 940823
rect 388609 940787 388665 940823
rect 388751 940787 388807 940823
rect 386905 940767 386908 940787
rect 386908 940767 386961 940787
rect 387047 940767 387088 940787
rect 387088 940767 387103 940787
rect 387189 940767 387212 940787
rect 387212 940767 387245 940787
rect 387331 940767 387336 940787
rect 387336 940767 387387 940787
rect 387473 940767 387528 940787
rect 387528 940767 387529 940787
rect 387615 940767 387652 940787
rect 387652 940767 387671 940787
rect 387757 940767 387776 940787
rect 387776 940767 387813 940787
rect 387899 940767 387900 940787
rect 387900 940767 387955 940787
rect 388041 940767 388080 940787
rect 388080 940767 388097 940787
rect 388183 940767 388204 940787
rect 388204 940767 388239 940787
rect 388325 940767 388328 940787
rect 388328 940767 388381 940787
rect 388467 940767 388520 940787
rect 388520 940767 388523 940787
rect 388609 940767 388644 940787
rect 388644 940767 388665 940787
rect 388751 940767 388768 940787
rect 388768 940767 388807 940787
rect 386905 940663 386961 940681
rect 387047 940663 387103 940681
rect 387189 940663 387245 940681
rect 387331 940663 387387 940681
rect 387473 940663 387529 940681
rect 387615 940663 387671 940681
rect 387757 940663 387813 940681
rect 387899 940663 387955 940681
rect 388041 940663 388097 940681
rect 388183 940663 388239 940681
rect 388325 940663 388381 940681
rect 388467 940663 388523 940681
rect 388609 940663 388665 940681
rect 388751 940663 388807 940681
rect 386905 940625 386908 940663
rect 386908 940625 386961 940663
rect 387047 940625 387088 940663
rect 387088 940625 387103 940663
rect 387189 940625 387212 940663
rect 387212 940625 387245 940663
rect 387331 940625 387336 940663
rect 387336 940625 387387 940663
rect 387473 940625 387528 940663
rect 387528 940625 387529 940663
rect 387615 940625 387652 940663
rect 387652 940625 387671 940663
rect 387757 940625 387776 940663
rect 387776 940625 387813 940663
rect 387899 940625 387900 940663
rect 387900 940625 387955 940663
rect 388041 940625 388080 940663
rect 388080 940625 388097 940663
rect 388183 940625 388204 940663
rect 388204 940625 388239 940663
rect 388325 940625 388328 940663
rect 388328 940625 388381 940663
rect 388467 940625 388520 940663
rect 388520 940625 388523 940663
rect 388609 940625 388644 940663
rect 388644 940625 388665 940663
rect 388751 940625 388768 940663
rect 388768 940625 388807 940663
rect 386905 940483 386908 940539
rect 386908 940483 386961 940539
rect 387047 940483 387088 940539
rect 387088 940483 387103 940539
rect 387189 940483 387212 940539
rect 387212 940483 387245 940539
rect 387331 940483 387336 940539
rect 387336 940483 387387 940539
rect 387473 940483 387528 940539
rect 387528 940483 387529 940539
rect 387615 940483 387652 940539
rect 387652 940483 387671 940539
rect 387757 940483 387776 940539
rect 387776 940483 387813 940539
rect 387899 940483 387900 940539
rect 387900 940483 387955 940539
rect 388041 940483 388080 940539
rect 388080 940483 388097 940539
rect 388183 940483 388204 940539
rect 388204 940483 388239 940539
rect 388325 940483 388328 940539
rect 388328 940483 388381 940539
rect 388467 940483 388520 940539
rect 388520 940483 388523 940539
rect 388609 940483 388644 940539
rect 388644 940483 388665 940539
rect 388751 940483 388768 940539
rect 388768 940483 388807 940539
rect 386905 940359 386908 940397
rect 386908 940359 386961 940397
rect 387047 940359 387088 940397
rect 387088 940359 387103 940397
rect 387189 940359 387212 940397
rect 387212 940359 387245 940397
rect 387331 940359 387336 940397
rect 387336 940359 387387 940397
rect 387473 940359 387528 940397
rect 387528 940359 387529 940397
rect 387615 940359 387652 940397
rect 387652 940359 387671 940397
rect 387757 940359 387776 940397
rect 387776 940359 387813 940397
rect 387899 940359 387900 940397
rect 387900 940359 387955 940397
rect 388041 940359 388080 940397
rect 388080 940359 388097 940397
rect 388183 940359 388204 940397
rect 388204 940359 388239 940397
rect 388325 940359 388328 940397
rect 388328 940359 388381 940397
rect 388467 940359 388520 940397
rect 388520 940359 388523 940397
rect 388609 940359 388644 940397
rect 388644 940359 388665 940397
rect 388751 940359 388768 940397
rect 388768 940359 388807 940397
rect 386905 940341 386961 940359
rect 387047 940341 387103 940359
rect 387189 940341 387245 940359
rect 387331 940341 387387 940359
rect 387473 940341 387529 940359
rect 387615 940341 387671 940359
rect 387757 940341 387813 940359
rect 387899 940341 387955 940359
rect 388041 940341 388097 940359
rect 388183 940341 388239 940359
rect 388325 940341 388381 940359
rect 388467 940341 388523 940359
rect 388609 940341 388665 940359
rect 388751 940341 388807 940359
rect 386905 940235 386908 940255
rect 386908 940235 386961 940255
rect 387047 940235 387088 940255
rect 387088 940235 387103 940255
rect 387189 940235 387212 940255
rect 387212 940235 387245 940255
rect 387331 940235 387336 940255
rect 387336 940235 387387 940255
rect 387473 940235 387528 940255
rect 387528 940235 387529 940255
rect 387615 940235 387652 940255
rect 387652 940235 387671 940255
rect 387757 940235 387776 940255
rect 387776 940235 387813 940255
rect 387899 940235 387900 940255
rect 387900 940235 387955 940255
rect 388041 940235 388080 940255
rect 388080 940235 388097 940255
rect 388183 940235 388204 940255
rect 388204 940235 388239 940255
rect 388325 940235 388328 940255
rect 388328 940235 388381 940255
rect 388467 940235 388520 940255
rect 388520 940235 388523 940255
rect 388609 940235 388644 940255
rect 388644 940235 388665 940255
rect 388751 940235 388768 940255
rect 388768 940235 388807 940255
rect 386905 940199 386961 940235
rect 387047 940199 387103 940235
rect 387189 940199 387245 940235
rect 387331 940199 387387 940235
rect 387473 940199 387529 940235
rect 387615 940199 387671 940235
rect 387757 940199 387813 940235
rect 387899 940199 387955 940235
rect 388041 940199 388097 940235
rect 388183 940199 388239 940235
rect 388325 940199 388381 940235
rect 388467 940199 388523 940235
rect 388609 940199 388665 940235
rect 388751 940199 388807 940235
rect 386905 940111 386908 940113
rect 386908 940111 386961 940113
rect 387047 940111 387088 940113
rect 387088 940111 387103 940113
rect 387189 940111 387212 940113
rect 387212 940111 387245 940113
rect 387331 940111 387336 940113
rect 387336 940111 387387 940113
rect 387473 940111 387528 940113
rect 387528 940111 387529 940113
rect 387615 940111 387652 940113
rect 387652 940111 387671 940113
rect 387757 940111 387776 940113
rect 387776 940111 387813 940113
rect 387899 940111 387900 940113
rect 387900 940111 387955 940113
rect 388041 940111 388080 940113
rect 388080 940111 388097 940113
rect 388183 940111 388204 940113
rect 388204 940111 388239 940113
rect 388325 940111 388328 940113
rect 388328 940111 388381 940113
rect 388467 940111 388520 940113
rect 388520 940111 388523 940113
rect 388609 940111 388644 940113
rect 388644 940111 388665 940113
rect 388751 940111 388768 940113
rect 388768 940111 388807 940113
rect 386905 940057 386961 940111
rect 387047 940057 387103 940111
rect 387189 940057 387245 940111
rect 387331 940057 387387 940111
rect 387473 940057 387529 940111
rect 387615 940057 387671 940111
rect 387757 940057 387813 940111
rect 387899 940057 387955 940111
rect 388041 940057 388097 940111
rect 388183 940057 388239 940111
rect 388325 940057 388381 940111
rect 388467 940057 388523 940111
rect 388609 940057 388665 940111
rect 388751 940057 388807 940111
rect 386905 939919 386961 939971
rect 387047 939919 387103 939971
rect 387189 939919 387245 939971
rect 387331 939919 387387 939971
rect 387473 939919 387529 939971
rect 387615 939919 387671 939971
rect 387757 939919 387813 939971
rect 387899 939919 387955 939971
rect 388041 939919 388097 939971
rect 388183 939919 388239 939971
rect 388325 939919 388381 939971
rect 388467 939919 388523 939971
rect 388609 939919 388665 939971
rect 388751 939919 388807 939971
rect 386905 939915 386908 939919
rect 386908 939915 386961 939919
rect 387047 939915 387088 939919
rect 387088 939915 387103 939919
rect 387189 939915 387212 939919
rect 387212 939915 387245 939919
rect 387331 939915 387336 939919
rect 387336 939915 387387 939919
rect 387473 939915 387528 939919
rect 387528 939915 387529 939919
rect 387615 939915 387652 939919
rect 387652 939915 387671 939919
rect 387757 939915 387776 939919
rect 387776 939915 387813 939919
rect 387899 939915 387900 939919
rect 387900 939915 387955 939919
rect 388041 939915 388080 939919
rect 388080 939915 388097 939919
rect 388183 939915 388204 939919
rect 388204 939915 388239 939919
rect 388325 939915 388328 939919
rect 388328 939915 388381 939919
rect 388467 939915 388520 939919
rect 388520 939915 388523 939919
rect 388609 939915 388644 939919
rect 388644 939915 388665 939919
rect 388751 939915 388768 939919
rect 388768 939915 388807 939919
rect 386905 939773 386961 939829
rect 387047 939773 387103 939829
rect 387189 939773 387245 939829
rect 387331 939773 387387 939829
rect 387473 939773 387529 939829
rect 387615 939773 387671 939829
rect 387757 939773 387813 939829
rect 387899 939773 387955 939829
rect 388041 939773 388097 939829
rect 388183 939773 388239 939829
rect 388325 939773 388381 939829
rect 388467 939773 388523 939829
rect 388609 939773 388665 939829
rect 388751 939773 388807 939829
rect 389275 941655 389331 941675
rect 389417 941655 389473 941675
rect 389559 941655 389615 941675
rect 389701 941655 389757 941675
rect 389843 941655 389899 941675
rect 389985 941655 390041 941675
rect 390127 941655 390183 941675
rect 390269 941655 390325 941675
rect 390411 941655 390467 941675
rect 390553 941655 390609 941675
rect 390695 941655 390751 941675
rect 390837 941655 390893 941675
rect 390979 941655 391035 941675
rect 391121 941655 391177 941675
rect 389275 941619 389278 941655
rect 389278 941619 389331 941655
rect 389417 941619 389458 941655
rect 389458 941619 389473 941655
rect 389559 941619 389582 941655
rect 389582 941619 389615 941655
rect 389701 941619 389706 941655
rect 389706 941619 389757 941655
rect 389843 941619 389898 941655
rect 389898 941619 389899 941655
rect 389985 941619 390022 941655
rect 390022 941619 390041 941655
rect 390127 941619 390146 941655
rect 390146 941619 390183 941655
rect 390269 941619 390270 941655
rect 390270 941619 390325 941655
rect 390411 941619 390450 941655
rect 390450 941619 390467 941655
rect 390553 941619 390574 941655
rect 390574 941619 390609 941655
rect 390695 941619 390698 941655
rect 390698 941619 390751 941655
rect 390837 941619 390890 941655
rect 390890 941619 390893 941655
rect 390979 941619 391014 941655
rect 391014 941619 391035 941655
rect 391121 941619 391138 941655
rect 391138 941619 391177 941655
rect 389275 941531 389331 941533
rect 389417 941531 389473 941533
rect 389559 941531 389615 941533
rect 389701 941531 389757 941533
rect 389843 941531 389899 941533
rect 389985 941531 390041 941533
rect 390127 941531 390183 941533
rect 390269 941531 390325 941533
rect 390411 941531 390467 941533
rect 390553 941531 390609 941533
rect 390695 941531 390751 941533
rect 390837 941531 390893 941533
rect 390979 941531 391035 941533
rect 391121 941531 391177 941533
rect 389275 941477 389278 941531
rect 389278 941477 389331 941531
rect 389417 941477 389458 941531
rect 389458 941477 389473 941531
rect 389559 941477 389582 941531
rect 389582 941477 389615 941531
rect 389701 941477 389706 941531
rect 389706 941477 389757 941531
rect 389843 941477 389898 941531
rect 389898 941477 389899 941531
rect 389985 941477 390022 941531
rect 390022 941477 390041 941531
rect 390127 941477 390146 941531
rect 390146 941477 390183 941531
rect 390269 941477 390270 941531
rect 390270 941477 390325 941531
rect 390411 941477 390450 941531
rect 390450 941477 390467 941531
rect 390553 941477 390574 941531
rect 390574 941477 390609 941531
rect 390695 941477 390698 941531
rect 390698 941477 390751 941531
rect 390837 941477 390890 941531
rect 390890 941477 390893 941531
rect 390979 941477 391014 941531
rect 391014 941477 391035 941531
rect 391121 941477 391138 941531
rect 391138 941477 391177 941531
rect 389275 941351 389278 941391
rect 389278 941351 389331 941391
rect 389417 941351 389458 941391
rect 389458 941351 389473 941391
rect 389559 941351 389582 941391
rect 389582 941351 389615 941391
rect 389701 941351 389706 941391
rect 389706 941351 389757 941391
rect 389843 941351 389898 941391
rect 389898 941351 389899 941391
rect 389985 941351 390022 941391
rect 390022 941351 390041 941391
rect 390127 941351 390146 941391
rect 390146 941351 390183 941391
rect 390269 941351 390270 941391
rect 390270 941351 390325 941391
rect 390411 941351 390450 941391
rect 390450 941351 390467 941391
rect 390553 941351 390574 941391
rect 390574 941351 390609 941391
rect 390695 941351 390698 941391
rect 390698 941351 390751 941391
rect 390837 941351 390890 941391
rect 390890 941351 390893 941391
rect 390979 941351 391014 941391
rect 391014 941351 391035 941391
rect 391121 941351 391138 941391
rect 391138 941351 391177 941391
rect 389275 941335 389331 941351
rect 389417 941335 389473 941351
rect 389559 941335 389615 941351
rect 389701 941335 389757 941351
rect 389843 941335 389899 941351
rect 389985 941335 390041 941351
rect 390127 941335 390183 941351
rect 390269 941335 390325 941351
rect 390411 941335 390467 941351
rect 390553 941335 390609 941351
rect 390695 941335 390751 941351
rect 390837 941335 390893 941351
rect 390979 941335 391035 941351
rect 391121 941335 391177 941351
rect 389275 941227 389278 941249
rect 389278 941227 389331 941249
rect 389417 941227 389458 941249
rect 389458 941227 389473 941249
rect 389559 941227 389582 941249
rect 389582 941227 389615 941249
rect 389701 941227 389706 941249
rect 389706 941227 389757 941249
rect 389843 941227 389898 941249
rect 389898 941227 389899 941249
rect 389985 941227 390022 941249
rect 390022 941227 390041 941249
rect 390127 941227 390146 941249
rect 390146 941227 390183 941249
rect 390269 941227 390270 941249
rect 390270 941227 390325 941249
rect 390411 941227 390450 941249
rect 390450 941227 390467 941249
rect 390553 941227 390574 941249
rect 390574 941227 390609 941249
rect 390695 941227 390698 941249
rect 390698 941227 390751 941249
rect 390837 941227 390890 941249
rect 390890 941227 390893 941249
rect 390979 941227 391014 941249
rect 391014 941227 391035 941249
rect 391121 941227 391138 941249
rect 391138 941227 391177 941249
rect 389275 941193 389331 941227
rect 389417 941193 389473 941227
rect 389559 941193 389615 941227
rect 389701 941193 389757 941227
rect 389843 941193 389899 941227
rect 389985 941193 390041 941227
rect 390127 941193 390183 941227
rect 390269 941193 390325 941227
rect 390411 941193 390467 941227
rect 390553 941193 390609 941227
rect 390695 941193 390751 941227
rect 390837 941193 390893 941227
rect 390979 941193 391035 941227
rect 391121 941193 391177 941227
rect 389275 941103 389278 941107
rect 389278 941103 389331 941107
rect 389417 941103 389458 941107
rect 389458 941103 389473 941107
rect 389559 941103 389582 941107
rect 389582 941103 389615 941107
rect 389701 941103 389706 941107
rect 389706 941103 389757 941107
rect 389843 941103 389898 941107
rect 389898 941103 389899 941107
rect 389985 941103 390022 941107
rect 390022 941103 390041 941107
rect 390127 941103 390146 941107
rect 390146 941103 390183 941107
rect 390269 941103 390270 941107
rect 390270 941103 390325 941107
rect 390411 941103 390450 941107
rect 390450 941103 390467 941107
rect 390553 941103 390574 941107
rect 390574 941103 390609 941107
rect 390695 941103 390698 941107
rect 390698 941103 390751 941107
rect 390837 941103 390890 941107
rect 390890 941103 390893 941107
rect 390979 941103 391014 941107
rect 391014 941103 391035 941107
rect 391121 941103 391138 941107
rect 391138 941103 391177 941107
rect 389275 941051 389331 941103
rect 389417 941051 389473 941103
rect 389559 941051 389615 941103
rect 389701 941051 389757 941103
rect 389843 941051 389899 941103
rect 389985 941051 390041 941103
rect 390127 941051 390183 941103
rect 390269 941051 390325 941103
rect 390411 941051 390467 941103
rect 390553 941051 390609 941103
rect 390695 941051 390751 941103
rect 390837 941051 390893 941103
rect 390979 941051 391035 941103
rect 391121 941051 391177 941103
rect 389275 940911 389331 940965
rect 389417 940911 389473 940965
rect 389559 940911 389615 940965
rect 389701 940911 389757 940965
rect 389843 940911 389899 940965
rect 389985 940911 390041 940965
rect 390127 940911 390183 940965
rect 390269 940911 390325 940965
rect 390411 940911 390467 940965
rect 390553 940911 390609 940965
rect 390695 940911 390751 940965
rect 390837 940911 390893 940965
rect 390979 940911 391035 940965
rect 391121 940911 391177 940965
rect 389275 940909 389278 940911
rect 389278 940909 389331 940911
rect 389417 940909 389458 940911
rect 389458 940909 389473 940911
rect 389559 940909 389582 940911
rect 389582 940909 389615 940911
rect 389701 940909 389706 940911
rect 389706 940909 389757 940911
rect 389843 940909 389898 940911
rect 389898 940909 389899 940911
rect 389985 940909 390022 940911
rect 390022 940909 390041 940911
rect 390127 940909 390146 940911
rect 390146 940909 390183 940911
rect 390269 940909 390270 940911
rect 390270 940909 390325 940911
rect 390411 940909 390450 940911
rect 390450 940909 390467 940911
rect 390553 940909 390574 940911
rect 390574 940909 390609 940911
rect 390695 940909 390698 940911
rect 390698 940909 390751 940911
rect 390837 940909 390890 940911
rect 390890 940909 390893 940911
rect 390979 940909 391014 940911
rect 391014 940909 391035 940911
rect 391121 940909 391138 940911
rect 391138 940909 391177 940911
rect 389275 940787 389331 940823
rect 389417 940787 389473 940823
rect 389559 940787 389615 940823
rect 389701 940787 389757 940823
rect 389843 940787 389899 940823
rect 389985 940787 390041 940823
rect 390127 940787 390183 940823
rect 390269 940787 390325 940823
rect 390411 940787 390467 940823
rect 390553 940787 390609 940823
rect 390695 940787 390751 940823
rect 390837 940787 390893 940823
rect 390979 940787 391035 940823
rect 391121 940787 391177 940823
rect 389275 940767 389278 940787
rect 389278 940767 389331 940787
rect 389417 940767 389458 940787
rect 389458 940767 389473 940787
rect 389559 940767 389582 940787
rect 389582 940767 389615 940787
rect 389701 940767 389706 940787
rect 389706 940767 389757 940787
rect 389843 940767 389898 940787
rect 389898 940767 389899 940787
rect 389985 940767 390022 940787
rect 390022 940767 390041 940787
rect 390127 940767 390146 940787
rect 390146 940767 390183 940787
rect 390269 940767 390270 940787
rect 390270 940767 390325 940787
rect 390411 940767 390450 940787
rect 390450 940767 390467 940787
rect 390553 940767 390574 940787
rect 390574 940767 390609 940787
rect 390695 940767 390698 940787
rect 390698 940767 390751 940787
rect 390837 940767 390890 940787
rect 390890 940767 390893 940787
rect 390979 940767 391014 940787
rect 391014 940767 391035 940787
rect 391121 940767 391138 940787
rect 391138 940767 391177 940787
rect 389275 940663 389331 940681
rect 389417 940663 389473 940681
rect 389559 940663 389615 940681
rect 389701 940663 389757 940681
rect 389843 940663 389899 940681
rect 389985 940663 390041 940681
rect 390127 940663 390183 940681
rect 390269 940663 390325 940681
rect 390411 940663 390467 940681
rect 390553 940663 390609 940681
rect 390695 940663 390751 940681
rect 390837 940663 390893 940681
rect 390979 940663 391035 940681
rect 391121 940663 391177 940681
rect 389275 940625 389278 940663
rect 389278 940625 389331 940663
rect 389417 940625 389458 940663
rect 389458 940625 389473 940663
rect 389559 940625 389582 940663
rect 389582 940625 389615 940663
rect 389701 940625 389706 940663
rect 389706 940625 389757 940663
rect 389843 940625 389898 940663
rect 389898 940625 389899 940663
rect 389985 940625 390022 940663
rect 390022 940625 390041 940663
rect 390127 940625 390146 940663
rect 390146 940625 390183 940663
rect 390269 940625 390270 940663
rect 390270 940625 390325 940663
rect 390411 940625 390450 940663
rect 390450 940625 390467 940663
rect 390553 940625 390574 940663
rect 390574 940625 390609 940663
rect 390695 940625 390698 940663
rect 390698 940625 390751 940663
rect 390837 940625 390890 940663
rect 390890 940625 390893 940663
rect 390979 940625 391014 940663
rect 391014 940625 391035 940663
rect 391121 940625 391138 940663
rect 391138 940625 391177 940663
rect 389275 940483 389278 940539
rect 389278 940483 389331 940539
rect 389417 940483 389458 940539
rect 389458 940483 389473 940539
rect 389559 940483 389582 940539
rect 389582 940483 389615 940539
rect 389701 940483 389706 940539
rect 389706 940483 389757 940539
rect 389843 940483 389898 940539
rect 389898 940483 389899 940539
rect 389985 940483 390022 940539
rect 390022 940483 390041 940539
rect 390127 940483 390146 940539
rect 390146 940483 390183 940539
rect 390269 940483 390270 940539
rect 390270 940483 390325 940539
rect 390411 940483 390450 940539
rect 390450 940483 390467 940539
rect 390553 940483 390574 940539
rect 390574 940483 390609 940539
rect 390695 940483 390698 940539
rect 390698 940483 390751 940539
rect 390837 940483 390890 940539
rect 390890 940483 390893 940539
rect 390979 940483 391014 940539
rect 391014 940483 391035 940539
rect 391121 940483 391138 940539
rect 391138 940483 391177 940539
rect 389275 940359 389278 940397
rect 389278 940359 389331 940397
rect 389417 940359 389458 940397
rect 389458 940359 389473 940397
rect 389559 940359 389582 940397
rect 389582 940359 389615 940397
rect 389701 940359 389706 940397
rect 389706 940359 389757 940397
rect 389843 940359 389898 940397
rect 389898 940359 389899 940397
rect 389985 940359 390022 940397
rect 390022 940359 390041 940397
rect 390127 940359 390146 940397
rect 390146 940359 390183 940397
rect 390269 940359 390270 940397
rect 390270 940359 390325 940397
rect 390411 940359 390450 940397
rect 390450 940359 390467 940397
rect 390553 940359 390574 940397
rect 390574 940359 390609 940397
rect 390695 940359 390698 940397
rect 390698 940359 390751 940397
rect 390837 940359 390890 940397
rect 390890 940359 390893 940397
rect 390979 940359 391014 940397
rect 391014 940359 391035 940397
rect 391121 940359 391138 940397
rect 391138 940359 391177 940397
rect 389275 940341 389331 940359
rect 389417 940341 389473 940359
rect 389559 940341 389615 940359
rect 389701 940341 389757 940359
rect 389843 940341 389899 940359
rect 389985 940341 390041 940359
rect 390127 940341 390183 940359
rect 390269 940341 390325 940359
rect 390411 940341 390467 940359
rect 390553 940341 390609 940359
rect 390695 940341 390751 940359
rect 390837 940341 390893 940359
rect 390979 940341 391035 940359
rect 391121 940341 391177 940359
rect 389275 940235 389278 940255
rect 389278 940235 389331 940255
rect 389417 940235 389458 940255
rect 389458 940235 389473 940255
rect 389559 940235 389582 940255
rect 389582 940235 389615 940255
rect 389701 940235 389706 940255
rect 389706 940235 389757 940255
rect 389843 940235 389898 940255
rect 389898 940235 389899 940255
rect 389985 940235 390022 940255
rect 390022 940235 390041 940255
rect 390127 940235 390146 940255
rect 390146 940235 390183 940255
rect 390269 940235 390270 940255
rect 390270 940235 390325 940255
rect 390411 940235 390450 940255
rect 390450 940235 390467 940255
rect 390553 940235 390574 940255
rect 390574 940235 390609 940255
rect 390695 940235 390698 940255
rect 390698 940235 390751 940255
rect 390837 940235 390890 940255
rect 390890 940235 390893 940255
rect 390979 940235 391014 940255
rect 391014 940235 391035 940255
rect 391121 940235 391138 940255
rect 391138 940235 391177 940255
rect 389275 940199 389331 940235
rect 389417 940199 389473 940235
rect 389559 940199 389615 940235
rect 389701 940199 389757 940235
rect 389843 940199 389899 940235
rect 389985 940199 390041 940235
rect 390127 940199 390183 940235
rect 390269 940199 390325 940235
rect 390411 940199 390467 940235
rect 390553 940199 390609 940235
rect 390695 940199 390751 940235
rect 390837 940199 390893 940235
rect 390979 940199 391035 940235
rect 391121 940199 391177 940235
rect 389275 940111 389278 940113
rect 389278 940111 389331 940113
rect 389417 940111 389458 940113
rect 389458 940111 389473 940113
rect 389559 940111 389582 940113
rect 389582 940111 389615 940113
rect 389701 940111 389706 940113
rect 389706 940111 389757 940113
rect 389843 940111 389898 940113
rect 389898 940111 389899 940113
rect 389985 940111 390022 940113
rect 390022 940111 390041 940113
rect 390127 940111 390146 940113
rect 390146 940111 390183 940113
rect 390269 940111 390270 940113
rect 390270 940111 390325 940113
rect 390411 940111 390450 940113
rect 390450 940111 390467 940113
rect 390553 940111 390574 940113
rect 390574 940111 390609 940113
rect 390695 940111 390698 940113
rect 390698 940111 390751 940113
rect 390837 940111 390890 940113
rect 390890 940111 390893 940113
rect 390979 940111 391014 940113
rect 391014 940111 391035 940113
rect 391121 940111 391138 940113
rect 391138 940111 391177 940113
rect 389275 940057 389331 940111
rect 389417 940057 389473 940111
rect 389559 940057 389615 940111
rect 389701 940057 389757 940111
rect 389843 940057 389899 940111
rect 389985 940057 390041 940111
rect 390127 940057 390183 940111
rect 390269 940057 390325 940111
rect 390411 940057 390467 940111
rect 390553 940057 390609 940111
rect 390695 940057 390751 940111
rect 390837 940057 390893 940111
rect 390979 940057 391035 940111
rect 391121 940057 391177 940111
rect 389275 939919 389331 939971
rect 389417 939919 389473 939971
rect 389559 939919 389615 939971
rect 389701 939919 389757 939971
rect 389843 939919 389899 939971
rect 389985 939919 390041 939971
rect 390127 939919 390183 939971
rect 390269 939919 390325 939971
rect 390411 939919 390467 939971
rect 390553 939919 390609 939971
rect 390695 939919 390751 939971
rect 390837 939919 390893 939971
rect 390979 939919 391035 939971
rect 391121 939919 391177 939971
rect 389275 939915 389278 939919
rect 389278 939915 389331 939919
rect 389417 939915 389458 939919
rect 389458 939915 389473 939919
rect 389559 939915 389582 939919
rect 389582 939915 389615 939919
rect 389701 939915 389706 939919
rect 389706 939915 389757 939919
rect 389843 939915 389898 939919
rect 389898 939915 389899 939919
rect 389985 939915 390022 939919
rect 390022 939915 390041 939919
rect 390127 939915 390146 939919
rect 390146 939915 390183 939919
rect 390269 939915 390270 939919
rect 390270 939915 390325 939919
rect 390411 939915 390450 939919
rect 390450 939915 390467 939919
rect 390553 939915 390574 939919
rect 390574 939915 390609 939919
rect 390695 939915 390698 939919
rect 390698 939915 390751 939919
rect 390837 939915 390890 939919
rect 390890 939915 390893 939919
rect 390979 939915 391014 939919
rect 391014 939915 391035 939919
rect 391121 939915 391138 939919
rect 391138 939915 391177 939919
rect 389275 939773 389331 939829
rect 389417 939773 389473 939829
rect 389559 939773 389615 939829
rect 389701 939773 389757 939829
rect 389843 939773 389899 939829
rect 389985 939773 390041 939829
rect 390127 939773 390183 939829
rect 390269 939773 390325 939829
rect 390411 939773 390467 939829
rect 390553 939773 390609 939829
rect 390695 939773 390751 939829
rect 390837 939773 390893 939829
rect 390979 939773 391035 939829
rect 391121 939773 391177 939829
rect 391897 941655 391953 941675
rect 392039 941655 392095 941675
rect 392181 941655 392237 941675
rect 392323 941655 392379 941675
rect 392465 941655 392521 941675
rect 392607 941655 392663 941675
rect 392749 941655 392805 941675
rect 392891 941655 392947 941675
rect 393033 941655 393089 941675
rect 393175 941655 393231 941675
rect 393317 941655 393373 941675
rect 393459 941655 393515 941675
rect 393601 941655 393657 941675
rect 391897 941619 391938 941655
rect 391938 941619 391953 941655
rect 392039 941619 392062 941655
rect 392062 941619 392095 941655
rect 392181 941619 392186 941655
rect 392186 941619 392237 941655
rect 392323 941619 392378 941655
rect 392378 941619 392379 941655
rect 392465 941619 392502 941655
rect 392502 941619 392521 941655
rect 392607 941619 392626 941655
rect 392626 941619 392663 941655
rect 392749 941619 392750 941655
rect 392750 941619 392805 941655
rect 392891 941619 392930 941655
rect 392930 941619 392947 941655
rect 393033 941619 393054 941655
rect 393054 941619 393089 941655
rect 393175 941619 393178 941655
rect 393178 941619 393231 941655
rect 393317 941619 393370 941655
rect 393370 941619 393373 941655
rect 393459 941619 393494 941655
rect 393494 941619 393515 941655
rect 393601 941619 393618 941655
rect 393618 941619 393657 941655
rect 391897 941531 391953 941533
rect 392039 941531 392095 941533
rect 392181 941531 392237 941533
rect 392323 941531 392379 941533
rect 392465 941531 392521 941533
rect 392607 941531 392663 941533
rect 392749 941531 392805 941533
rect 392891 941531 392947 941533
rect 393033 941531 393089 941533
rect 393175 941531 393231 941533
rect 393317 941531 393373 941533
rect 393459 941531 393515 941533
rect 393601 941531 393657 941533
rect 391897 941477 391938 941531
rect 391938 941477 391953 941531
rect 392039 941477 392062 941531
rect 392062 941477 392095 941531
rect 392181 941477 392186 941531
rect 392186 941477 392237 941531
rect 392323 941477 392378 941531
rect 392378 941477 392379 941531
rect 392465 941477 392502 941531
rect 392502 941477 392521 941531
rect 392607 941477 392626 941531
rect 392626 941477 392663 941531
rect 392749 941477 392750 941531
rect 392750 941477 392805 941531
rect 392891 941477 392930 941531
rect 392930 941477 392947 941531
rect 393033 941477 393054 941531
rect 393054 941477 393089 941531
rect 393175 941477 393178 941531
rect 393178 941477 393231 941531
rect 393317 941477 393370 941531
rect 393370 941477 393373 941531
rect 393459 941477 393494 941531
rect 393494 941477 393515 941531
rect 393601 941477 393618 941531
rect 393618 941477 393657 941531
rect 391897 941351 391938 941391
rect 391938 941351 391953 941391
rect 392039 941351 392062 941391
rect 392062 941351 392095 941391
rect 392181 941351 392186 941391
rect 392186 941351 392237 941391
rect 392323 941351 392378 941391
rect 392378 941351 392379 941391
rect 392465 941351 392502 941391
rect 392502 941351 392521 941391
rect 392607 941351 392626 941391
rect 392626 941351 392663 941391
rect 392749 941351 392750 941391
rect 392750 941351 392805 941391
rect 392891 941351 392930 941391
rect 392930 941351 392947 941391
rect 393033 941351 393054 941391
rect 393054 941351 393089 941391
rect 393175 941351 393178 941391
rect 393178 941351 393231 941391
rect 393317 941351 393370 941391
rect 393370 941351 393373 941391
rect 393459 941351 393494 941391
rect 393494 941351 393515 941391
rect 393601 941351 393618 941391
rect 393618 941351 393657 941391
rect 391897 941335 391953 941351
rect 392039 941335 392095 941351
rect 392181 941335 392237 941351
rect 392323 941335 392379 941351
rect 392465 941335 392521 941351
rect 392607 941335 392663 941351
rect 392749 941335 392805 941351
rect 392891 941335 392947 941351
rect 393033 941335 393089 941351
rect 393175 941335 393231 941351
rect 393317 941335 393373 941351
rect 393459 941335 393515 941351
rect 393601 941335 393657 941351
rect 391897 941227 391938 941249
rect 391938 941227 391953 941249
rect 392039 941227 392062 941249
rect 392062 941227 392095 941249
rect 392181 941227 392186 941249
rect 392186 941227 392237 941249
rect 392323 941227 392378 941249
rect 392378 941227 392379 941249
rect 392465 941227 392502 941249
rect 392502 941227 392521 941249
rect 392607 941227 392626 941249
rect 392626 941227 392663 941249
rect 392749 941227 392750 941249
rect 392750 941227 392805 941249
rect 392891 941227 392930 941249
rect 392930 941227 392947 941249
rect 393033 941227 393054 941249
rect 393054 941227 393089 941249
rect 393175 941227 393178 941249
rect 393178 941227 393231 941249
rect 393317 941227 393370 941249
rect 393370 941227 393373 941249
rect 393459 941227 393494 941249
rect 393494 941227 393515 941249
rect 393601 941227 393618 941249
rect 393618 941227 393657 941249
rect 391897 941193 391953 941227
rect 392039 941193 392095 941227
rect 392181 941193 392237 941227
rect 392323 941193 392379 941227
rect 392465 941193 392521 941227
rect 392607 941193 392663 941227
rect 392749 941193 392805 941227
rect 392891 941193 392947 941227
rect 393033 941193 393089 941227
rect 393175 941193 393231 941227
rect 393317 941193 393373 941227
rect 393459 941193 393515 941227
rect 393601 941193 393657 941227
rect 391897 941103 391938 941107
rect 391938 941103 391953 941107
rect 392039 941103 392062 941107
rect 392062 941103 392095 941107
rect 392181 941103 392186 941107
rect 392186 941103 392237 941107
rect 392323 941103 392378 941107
rect 392378 941103 392379 941107
rect 392465 941103 392502 941107
rect 392502 941103 392521 941107
rect 392607 941103 392626 941107
rect 392626 941103 392663 941107
rect 392749 941103 392750 941107
rect 392750 941103 392805 941107
rect 392891 941103 392930 941107
rect 392930 941103 392947 941107
rect 393033 941103 393054 941107
rect 393054 941103 393089 941107
rect 393175 941103 393178 941107
rect 393178 941103 393231 941107
rect 393317 941103 393370 941107
rect 393370 941103 393373 941107
rect 393459 941103 393494 941107
rect 393494 941103 393515 941107
rect 393601 941103 393618 941107
rect 393618 941103 393657 941107
rect 391897 941051 391953 941103
rect 392039 941051 392095 941103
rect 392181 941051 392237 941103
rect 392323 941051 392379 941103
rect 392465 941051 392521 941103
rect 392607 941051 392663 941103
rect 392749 941051 392805 941103
rect 392891 941051 392947 941103
rect 393033 941051 393089 941103
rect 393175 941051 393231 941103
rect 393317 941051 393373 941103
rect 393459 941051 393515 941103
rect 393601 941051 393657 941103
rect 391897 940911 391953 940965
rect 392039 940911 392095 940965
rect 392181 940911 392237 940965
rect 392323 940911 392379 940965
rect 392465 940911 392521 940965
rect 392607 940911 392663 940965
rect 392749 940911 392805 940965
rect 392891 940911 392947 940965
rect 393033 940911 393089 940965
rect 393175 940911 393231 940965
rect 393317 940911 393373 940965
rect 393459 940911 393515 940965
rect 393601 940911 393657 940965
rect 391897 940909 391938 940911
rect 391938 940909 391953 940911
rect 392039 940909 392062 940911
rect 392062 940909 392095 940911
rect 392181 940909 392186 940911
rect 392186 940909 392237 940911
rect 392323 940909 392378 940911
rect 392378 940909 392379 940911
rect 392465 940909 392502 940911
rect 392502 940909 392521 940911
rect 392607 940909 392626 940911
rect 392626 940909 392663 940911
rect 392749 940909 392750 940911
rect 392750 940909 392805 940911
rect 392891 940909 392930 940911
rect 392930 940909 392947 940911
rect 393033 940909 393054 940911
rect 393054 940909 393089 940911
rect 393175 940909 393178 940911
rect 393178 940909 393231 940911
rect 393317 940909 393370 940911
rect 393370 940909 393373 940911
rect 393459 940909 393494 940911
rect 393494 940909 393515 940911
rect 393601 940909 393618 940911
rect 393618 940909 393657 940911
rect 391897 940787 391953 940823
rect 392039 940787 392095 940823
rect 392181 940787 392237 940823
rect 392323 940787 392379 940823
rect 392465 940787 392521 940823
rect 392607 940787 392663 940823
rect 392749 940787 392805 940823
rect 392891 940787 392947 940823
rect 393033 940787 393089 940823
rect 393175 940787 393231 940823
rect 393317 940787 393373 940823
rect 393459 940787 393515 940823
rect 393601 940787 393657 940823
rect 391897 940767 391938 940787
rect 391938 940767 391953 940787
rect 392039 940767 392062 940787
rect 392062 940767 392095 940787
rect 392181 940767 392186 940787
rect 392186 940767 392237 940787
rect 392323 940767 392378 940787
rect 392378 940767 392379 940787
rect 392465 940767 392502 940787
rect 392502 940767 392521 940787
rect 392607 940767 392626 940787
rect 392626 940767 392663 940787
rect 392749 940767 392750 940787
rect 392750 940767 392805 940787
rect 392891 940767 392930 940787
rect 392930 940767 392947 940787
rect 393033 940767 393054 940787
rect 393054 940767 393089 940787
rect 393175 940767 393178 940787
rect 393178 940767 393231 940787
rect 393317 940767 393370 940787
rect 393370 940767 393373 940787
rect 393459 940767 393494 940787
rect 393494 940767 393515 940787
rect 393601 940767 393618 940787
rect 393618 940767 393657 940787
rect 391897 940663 391953 940681
rect 392039 940663 392095 940681
rect 392181 940663 392237 940681
rect 392323 940663 392379 940681
rect 392465 940663 392521 940681
rect 392607 940663 392663 940681
rect 392749 940663 392805 940681
rect 392891 940663 392947 940681
rect 393033 940663 393089 940681
rect 393175 940663 393231 940681
rect 393317 940663 393373 940681
rect 393459 940663 393515 940681
rect 393601 940663 393657 940681
rect 391897 940625 391938 940663
rect 391938 940625 391953 940663
rect 392039 940625 392062 940663
rect 392062 940625 392095 940663
rect 392181 940625 392186 940663
rect 392186 940625 392237 940663
rect 392323 940625 392378 940663
rect 392378 940625 392379 940663
rect 392465 940625 392502 940663
rect 392502 940625 392521 940663
rect 392607 940625 392626 940663
rect 392626 940625 392663 940663
rect 392749 940625 392750 940663
rect 392750 940625 392805 940663
rect 392891 940625 392930 940663
rect 392930 940625 392947 940663
rect 393033 940625 393054 940663
rect 393054 940625 393089 940663
rect 393175 940625 393178 940663
rect 393178 940625 393231 940663
rect 393317 940625 393370 940663
rect 393370 940625 393373 940663
rect 393459 940625 393494 940663
rect 393494 940625 393515 940663
rect 393601 940625 393618 940663
rect 393618 940625 393657 940663
rect 391897 940483 391938 940539
rect 391938 940483 391953 940539
rect 392039 940483 392062 940539
rect 392062 940483 392095 940539
rect 392181 940483 392186 940539
rect 392186 940483 392237 940539
rect 392323 940483 392378 940539
rect 392378 940483 392379 940539
rect 392465 940483 392502 940539
rect 392502 940483 392521 940539
rect 392607 940483 392626 940539
rect 392626 940483 392663 940539
rect 392749 940483 392750 940539
rect 392750 940483 392805 940539
rect 392891 940483 392930 940539
rect 392930 940483 392947 940539
rect 393033 940483 393054 940539
rect 393054 940483 393089 940539
rect 393175 940483 393178 940539
rect 393178 940483 393231 940539
rect 393317 940483 393370 940539
rect 393370 940483 393373 940539
rect 393459 940483 393494 940539
rect 393494 940483 393515 940539
rect 393601 940483 393618 940539
rect 393618 940483 393657 940539
rect 391897 940359 391938 940397
rect 391938 940359 391953 940397
rect 392039 940359 392062 940397
rect 392062 940359 392095 940397
rect 392181 940359 392186 940397
rect 392186 940359 392237 940397
rect 392323 940359 392378 940397
rect 392378 940359 392379 940397
rect 392465 940359 392502 940397
rect 392502 940359 392521 940397
rect 392607 940359 392626 940397
rect 392626 940359 392663 940397
rect 392749 940359 392750 940397
rect 392750 940359 392805 940397
rect 392891 940359 392930 940397
rect 392930 940359 392947 940397
rect 393033 940359 393054 940397
rect 393054 940359 393089 940397
rect 393175 940359 393178 940397
rect 393178 940359 393231 940397
rect 393317 940359 393370 940397
rect 393370 940359 393373 940397
rect 393459 940359 393494 940397
rect 393494 940359 393515 940397
rect 393601 940359 393618 940397
rect 393618 940359 393657 940397
rect 391897 940341 391953 940359
rect 392039 940341 392095 940359
rect 392181 940341 392237 940359
rect 392323 940341 392379 940359
rect 392465 940341 392521 940359
rect 392607 940341 392663 940359
rect 392749 940341 392805 940359
rect 392891 940341 392947 940359
rect 393033 940341 393089 940359
rect 393175 940341 393231 940359
rect 393317 940341 393373 940359
rect 393459 940341 393515 940359
rect 393601 940341 393657 940359
rect 391897 940235 391938 940255
rect 391938 940235 391953 940255
rect 392039 940235 392062 940255
rect 392062 940235 392095 940255
rect 392181 940235 392186 940255
rect 392186 940235 392237 940255
rect 392323 940235 392378 940255
rect 392378 940235 392379 940255
rect 392465 940235 392502 940255
rect 392502 940235 392521 940255
rect 392607 940235 392626 940255
rect 392626 940235 392663 940255
rect 392749 940235 392750 940255
rect 392750 940235 392805 940255
rect 392891 940235 392930 940255
rect 392930 940235 392947 940255
rect 393033 940235 393054 940255
rect 393054 940235 393089 940255
rect 393175 940235 393178 940255
rect 393178 940235 393231 940255
rect 393317 940235 393370 940255
rect 393370 940235 393373 940255
rect 393459 940235 393494 940255
rect 393494 940235 393515 940255
rect 393601 940235 393618 940255
rect 393618 940235 393657 940255
rect 391897 940199 391953 940235
rect 392039 940199 392095 940235
rect 392181 940199 392237 940235
rect 392323 940199 392379 940235
rect 392465 940199 392521 940235
rect 392607 940199 392663 940235
rect 392749 940199 392805 940235
rect 392891 940199 392947 940235
rect 393033 940199 393089 940235
rect 393175 940199 393231 940235
rect 393317 940199 393373 940235
rect 393459 940199 393515 940235
rect 393601 940199 393657 940235
rect 391897 940111 391938 940113
rect 391938 940111 391953 940113
rect 392039 940111 392062 940113
rect 392062 940111 392095 940113
rect 392181 940111 392186 940113
rect 392186 940111 392237 940113
rect 392323 940111 392378 940113
rect 392378 940111 392379 940113
rect 392465 940111 392502 940113
rect 392502 940111 392521 940113
rect 392607 940111 392626 940113
rect 392626 940111 392663 940113
rect 392749 940111 392750 940113
rect 392750 940111 392805 940113
rect 392891 940111 392930 940113
rect 392930 940111 392947 940113
rect 393033 940111 393054 940113
rect 393054 940111 393089 940113
rect 393175 940111 393178 940113
rect 393178 940111 393231 940113
rect 393317 940111 393370 940113
rect 393370 940111 393373 940113
rect 393459 940111 393494 940113
rect 393494 940111 393515 940113
rect 393601 940111 393618 940113
rect 393618 940111 393657 940113
rect 391897 940057 391953 940111
rect 392039 940057 392095 940111
rect 392181 940057 392237 940111
rect 392323 940057 392379 940111
rect 392465 940057 392521 940111
rect 392607 940057 392663 940111
rect 392749 940057 392805 940111
rect 392891 940057 392947 940111
rect 393033 940057 393089 940111
rect 393175 940057 393231 940111
rect 393317 940057 393373 940111
rect 393459 940057 393515 940111
rect 393601 940057 393657 940111
rect 391897 939919 391953 939971
rect 392039 939919 392095 939971
rect 392181 939919 392237 939971
rect 392323 939919 392379 939971
rect 392465 939919 392521 939971
rect 392607 939919 392663 939971
rect 392749 939919 392805 939971
rect 392891 939919 392947 939971
rect 393033 939919 393089 939971
rect 393175 939919 393231 939971
rect 393317 939919 393373 939971
rect 393459 939919 393515 939971
rect 393601 939919 393657 939971
rect 391897 939915 391938 939919
rect 391938 939915 391953 939919
rect 392039 939915 392062 939919
rect 392062 939915 392095 939919
rect 392181 939915 392186 939919
rect 392186 939915 392237 939919
rect 392323 939915 392378 939919
rect 392378 939915 392379 939919
rect 392465 939915 392502 939919
rect 392502 939915 392521 939919
rect 392607 939915 392626 939919
rect 392626 939915 392663 939919
rect 392749 939915 392750 939919
rect 392750 939915 392805 939919
rect 392891 939915 392930 939919
rect 392930 939915 392947 939919
rect 393033 939915 393054 939919
rect 393054 939915 393089 939919
rect 393175 939915 393178 939919
rect 393178 939915 393231 939919
rect 393317 939915 393370 939919
rect 393370 939915 393373 939919
rect 393459 939915 393494 939919
rect 393494 939915 393515 939919
rect 393601 939915 393618 939919
rect 393618 939915 393657 939919
rect 391897 939773 391953 939829
rect 392039 939773 392095 939829
rect 392181 939773 392237 939829
rect 392323 939773 392379 939829
rect 392465 939773 392521 939829
rect 392607 939773 392663 939829
rect 392749 939773 392805 939829
rect 392891 939773 392947 939829
rect 393033 939773 393089 939829
rect 393175 939773 393231 939829
rect 393317 939773 393373 939829
rect 393459 939773 393515 939829
rect 393601 939773 393657 939829
rect 599341 941655 599397 941675
rect 599483 941655 599539 941675
rect 599625 941655 599681 941675
rect 599767 941655 599823 941675
rect 599909 941655 599965 941675
rect 600051 941655 600107 941675
rect 600193 941655 600249 941675
rect 600335 941655 600391 941675
rect 600477 941655 600533 941675
rect 600619 941655 600675 941675
rect 600761 941655 600817 941675
rect 600903 941655 600959 941675
rect 601045 941655 601101 941675
rect 599341 941619 599382 941655
rect 599382 941619 599397 941655
rect 599483 941619 599506 941655
rect 599506 941619 599539 941655
rect 599625 941619 599630 941655
rect 599630 941619 599681 941655
rect 599767 941619 599822 941655
rect 599822 941619 599823 941655
rect 599909 941619 599946 941655
rect 599946 941619 599965 941655
rect 600051 941619 600070 941655
rect 600070 941619 600107 941655
rect 600193 941619 600194 941655
rect 600194 941619 600249 941655
rect 600335 941619 600374 941655
rect 600374 941619 600391 941655
rect 600477 941619 600498 941655
rect 600498 941619 600533 941655
rect 600619 941619 600622 941655
rect 600622 941619 600675 941655
rect 600761 941619 600814 941655
rect 600814 941619 600817 941655
rect 600903 941619 600938 941655
rect 600938 941619 600959 941655
rect 601045 941619 601062 941655
rect 601062 941619 601101 941655
rect 599341 941531 599397 941533
rect 599483 941531 599539 941533
rect 599625 941531 599681 941533
rect 599767 941531 599823 941533
rect 599909 941531 599965 941533
rect 600051 941531 600107 941533
rect 600193 941531 600249 941533
rect 600335 941531 600391 941533
rect 600477 941531 600533 941533
rect 600619 941531 600675 941533
rect 600761 941531 600817 941533
rect 600903 941531 600959 941533
rect 601045 941531 601101 941533
rect 599341 941477 599382 941531
rect 599382 941477 599397 941531
rect 599483 941477 599506 941531
rect 599506 941477 599539 941531
rect 599625 941477 599630 941531
rect 599630 941477 599681 941531
rect 599767 941477 599822 941531
rect 599822 941477 599823 941531
rect 599909 941477 599946 941531
rect 599946 941477 599965 941531
rect 600051 941477 600070 941531
rect 600070 941477 600107 941531
rect 600193 941477 600194 941531
rect 600194 941477 600249 941531
rect 600335 941477 600374 941531
rect 600374 941477 600391 941531
rect 600477 941477 600498 941531
rect 600498 941477 600533 941531
rect 600619 941477 600622 941531
rect 600622 941477 600675 941531
rect 600761 941477 600814 941531
rect 600814 941477 600817 941531
rect 600903 941477 600938 941531
rect 600938 941477 600959 941531
rect 601045 941477 601062 941531
rect 601062 941477 601101 941531
rect 599341 941351 599382 941391
rect 599382 941351 599397 941391
rect 599483 941351 599506 941391
rect 599506 941351 599539 941391
rect 599625 941351 599630 941391
rect 599630 941351 599681 941391
rect 599767 941351 599822 941391
rect 599822 941351 599823 941391
rect 599909 941351 599946 941391
rect 599946 941351 599965 941391
rect 600051 941351 600070 941391
rect 600070 941351 600107 941391
rect 600193 941351 600194 941391
rect 600194 941351 600249 941391
rect 600335 941351 600374 941391
rect 600374 941351 600391 941391
rect 600477 941351 600498 941391
rect 600498 941351 600533 941391
rect 600619 941351 600622 941391
rect 600622 941351 600675 941391
rect 600761 941351 600814 941391
rect 600814 941351 600817 941391
rect 600903 941351 600938 941391
rect 600938 941351 600959 941391
rect 601045 941351 601062 941391
rect 601062 941351 601101 941391
rect 599341 941335 599397 941351
rect 599483 941335 599539 941351
rect 599625 941335 599681 941351
rect 599767 941335 599823 941351
rect 599909 941335 599965 941351
rect 600051 941335 600107 941351
rect 600193 941335 600249 941351
rect 600335 941335 600391 941351
rect 600477 941335 600533 941351
rect 600619 941335 600675 941351
rect 600761 941335 600817 941351
rect 600903 941335 600959 941351
rect 601045 941335 601101 941351
rect 599341 941227 599382 941249
rect 599382 941227 599397 941249
rect 599483 941227 599506 941249
rect 599506 941227 599539 941249
rect 599625 941227 599630 941249
rect 599630 941227 599681 941249
rect 599767 941227 599822 941249
rect 599822 941227 599823 941249
rect 599909 941227 599946 941249
rect 599946 941227 599965 941249
rect 600051 941227 600070 941249
rect 600070 941227 600107 941249
rect 600193 941227 600194 941249
rect 600194 941227 600249 941249
rect 600335 941227 600374 941249
rect 600374 941227 600391 941249
rect 600477 941227 600498 941249
rect 600498 941227 600533 941249
rect 600619 941227 600622 941249
rect 600622 941227 600675 941249
rect 600761 941227 600814 941249
rect 600814 941227 600817 941249
rect 600903 941227 600938 941249
rect 600938 941227 600959 941249
rect 601045 941227 601062 941249
rect 601062 941227 601101 941249
rect 599341 941193 599397 941227
rect 599483 941193 599539 941227
rect 599625 941193 599681 941227
rect 599767 941193 599823 941227
rect 599909 941193 599965 941227
rect 600051 941193 600107 941227
rect 600193 941193 600249 941227
rect 600335 941193 600391 941227
rect 600477 941193 600533 941227
rect 600619 941193 600675 941227
rect 600761 941193 600817 941227
rect 600903 941193 600959 941227
rect 601045 941193 601101 941227
rect 599341 941103 599382 941107
rect 599382 941103 599397 941107
rect 599483 941103 599506 941107
rect 599506 941103 599539 941107
rect 599625 941103 599630 941107
rect 599630 941103 599681 941107
rect 599767 941103 599822 941107
rect 599822 941103 599823 941107
rect 599909 941103 599946 941107
rect 599946 941103 599965 941107
rect 600051 941103 600070 941107
rect 600070 941103 600107 941107
rect 600193 941103 600194 941107
rect 600194 941103 600249 941107
rect 600335 941103 600374 941107
rect 600374 941103 600391 941107
rect 600477 941103 600498 941107
rect 600498 941103 600533 941107
rect 600619 941103 600622 941107
rect 600622 941103 600675 941107
rect 600761 941103 600814 941107
rect 600814 941103 600817 941107
rect 600903 941103 600938 941107
rect 600938 941103 600959 941107
rect 601045 941103 601062 941107
rect 601062 941103 601101 941107
rect 599341 941051 599397 941103
rect 599483 941051 599539 941103
rect 599625 941051 599681 941103
rect 599767 941051 599823 941103
rect 599909 941051 599965 941103
rect 600051 941051 600107 941103
rect 600193 941051 600249 941103
rect 600335 941051 600391 941103
rect 600477 941051 600533 941103
rect 600619 941051 600675 941103
rect 600761 941051 600817 941103
rect 600903 941051 600959 941103
rect 601045 941051 601101 941103
rect 599341 940911 599397 940965
rect 599483 940911 599539 940965
rect 599625 940911 599681 940965
rect 599767 940911 599823 940965
rect 599909 940911 599965 940965
rect 600051 940911 600107 940965
rect 600193 940911 600249 940965
rect 600335 940911 600391 940965
rect 600477 940911 600533 940965
rect 600619 940911 600675 940965
rect 600761 940911 600817 940965
rect 600903 940911 600959 940965
rect 601045 940911 601101 940965
rect 599341 940909 599382 940911
rect 599382 940909 599397 940911
rect 599483 940909 599506 940911
rect 599506 940909 599539 940911
rect 599625 940909 599630 940911
rect 599630 940909 599681 940911
rect 599767 940909 599822 940911
rect 599822 940909 599823 940911
rect 599909 940909 599946 940911
rect 599946 940909 599965 940911
rect 600051 940909 600070 940911
rect 600070 940909 600107 940911
rect 600193 940909 600194 940911
rect 600194 940909 600249 940911
rect 600335 940909 600374 940911
rect 600374 940909 600391 940911
rect 600477 940909 600498 940911
rect 600498 940909 600533 940911
rect 600619 940909 600622 940911
rect 600622 940909 600675 940911
rect 600761 940909 600814 940911
rect 600814 940909 600817 940911
rect 600903 940909 600938 940911
rect 600938 940909 600959 940911
rect 601045 940909 601062 940911
rect 601062 940909 601101 940911
rect 599341 940787 599397 940823
rect 599483 940787 599539 940823
rect 599625 940787 599681 940823
rect 599767 940787 599823 940823
rect 599909 940787 599965 940823
rect 600051 940787 600107 940823
rect 600193 940787 600249 940823
rect 600335 940787 600391 940823
rect 600477 940787 600533 940823
rect 600619 940787 600675 940823
rect 600761 940787 600817 940823
rect 600903 940787 600959 940823
rect 601045 940787 601101 940823
rect 599341 940767 599382 940787
rect 599382 940767 599397 940787
rect 599483 940767 599506 940787
rect 599506 940767 599539 940787
rect 599625 940767 599630 940787
rect 599630 940767 599681 940787
rect 599767 940767 599822 940787
rect 599822 940767 599823 940787
rect 599909 940767 599946 940787
rect 599946 940767 599965 940787
rect 600051 940767 600070 940787
rect 600070 940767 600107 940787
rect 600193 940767 600194 940787
rect 600194 940767 600249 940787
rect 600335 940767 600374 940787
rect 600374 940767 600391 940787
rect 600477 940767 600498 940787
rect 600498 940767 600533 940787
rect 600619 940767 600622 940787
rect 600622 940767 600675 940787
rect 600761 940767 600814 940787
rect 600814 940767 600817 940787
rect 600903 940767 600938 940787
rect 600938 940767 600959 940787
rect 601045 940767 601062 940787
rect 601062 940767 601101 940787
rect 599341 940663 599397 940681
rect 599483 940663 599539 940681
rect 599625 940663 599681 940681
rect 599767 940663 599823 940681
rect 599909 940663 599965 940681
rect 600051 940663 600107 940681
rect 600193 940663 600249 940681
rect 600335 940663 600391 940681
rect 600477 940663 600533 940681
rect 600619 940663 600675 940681
rect 600761 940663 600817 940681
rect 600903 940663 600959 940681
rect 601045 940663 601101 940681
rect 599341 940625 599382 940663
rect 599382 940625 599397 940663
rect 599483 940625 599506 940663
rect 599506 940625 599539 940663
rect 599625 940625 599630 940663
rect 599630 940625 599681 940663
rect 599767 940625 599822 940663
rect 599822 940625 599823 940663
rect 599909 940625 599946 940663
rect 599946 940625 599965 940663
rect 600051 940625 600070 940663
rect 600070 940625 600107 940663
rect 600193 940625 600194 940663
rect 600194 940625 600249 940663
rect 600335 940625 600374 940663
rect 600374 940625 600391 940663
rect 600477 940625 600498 940663
rect 600498 940625 600533 940663
rect 600619 940625 600622 940663
rect 600622 940625 600675 940663
rect 600761 940625 600814 940663
rect 600814 940625 600817 940663
rect 600903 940625 600938 940663
rect 600938 940625 600959 940663
rect 601045 940625 601062 940663
rect 601062 940625 601101 940663
rect 599341 940483 599382 940539
rect 599382 940483 599397 940539
rect 599483 940483 599506 940539
rect 599506 940483 599539 940539
rect 599625 940483 599630 940539
rect 599630 940483 599681 940539
rect 599767 940483 599822 940539
rect 599822 940483 599823 940539
rect 599909 940483 599946 940539
rect 599946 940483 599965 940539
rect 600051 940483 600070 940539
rect 600070 940483 600107 940539
rect 600193 940483 600194 940539
rect 600194 940483 600249 940539
rect 600335 940483 600374 940539
rect 600374 940483 600391 940539
rect 600477 940483 600498 940539
rect 600498 940483 600533 940539
rect 600619 940483 600622 940539
rect 600622 940483 600675 940539
rect 600761 940483 600814 940539
rect 600814 940483 600817 940539
rect 600903 940483 600938 940539
rect 600938 940483 600959 940539
rect 601045 940483 601062 940539
rect 601062 940483 601101 940539
rect 599341 940359 599382 940397
rect 599382 940359 599397 940397
rect 599483 940359 599506 940397
rect 599506 940359 599539 940397
rect 599625 940359 599630 940397
rect 599630 940359 599681 940397
rect 599767 940359 599822 940397
rect 599822 940359 599823 940397
rect 599909 940359 599946 940397
rect 599946 940359 599965 940397
rect 600051 940359 600070 940397
rect 600070 940359 600107 940397
rect 600193 940359 600194 940397
rect 600194 940359 600249 940397
rect 600335 940359 600374 940397
rect 600374 940359 600391 940397
rect 600477 940359 600498 940397
rect 600498 940359 600533 940397
rect 600619 940359 600622 940397
rect 600622 940359 600675 940397
rect 600761 940359 600814 940397
rect 600814 940359 600817 940397
rect 600903 940359 600938 940397
rect 600938 940359 600959 940397
rect 601045 940359 601062 940397
rect 601062 940359 601101 940397
rect 599341 940341 599397 940359
rect 599483 940341 599539 940359
rect 599625 940341 599681 940359
rect 599767 940341 599823 940359
rect 599909 940341 599965 940359
rect 600051 940341 600107 940359
rect 600193 940341 600249 940359
rect 600335 940341 600391 940359
rect 600477 940341 600533 940359
rect 600619 940341 600675 940359
rect 600761 940341 600817 940359
rect 600903 940341 600959 940359
rect 601045 940341 601101 940359
rect 599341 940235 599382 940255
rect 599382 940235 599397 940255
rect 599483 940235 599506 940255
rect 599506 940235 599539 940255
rect 599625 940235 599630 940255
rect 599630 940235 599681 940255
rect 599767 940235 599822 940255
rect 599822 940235 599823 940255
rect 599909 940235 599946 940255
rect 599946 940235 599965 940255
rect 600051 940235 600070 940255
rect 600070 940235 600107 940255
rect 600193 940235 600194 940255
rect 600194 940235 600249 940255
rect 600335 940235 600374 940255
rect 600374 940235 600391 940255
rect 600477 940235 600498 940255
rect 600498 940235 600533 940255
rect 600619 940235 600622 940255
rect 600622 940235 600675 940255
rect 600761 940235 600814 940255
rect 600814 940235 600817 940255
rect 600903 940235 600938 940255
rect 600938 940235 600959 940255
rect 601045 940235 601062 940255
rect 601062 940235 601101 940255
rect 599341 940199 599397 940235
rect 599483 940199 599539 940235
rect 599625 940199 599681 940235
rect 599767 940199 599823 940235
rect 599909 940199 599965 940235
rect 600051 940199 600107 940235
rect 600193 940199 600249 940235
rect 600335 940199 600391 940235
rect 600477 940199 600533 940235
rect 600619 940199 600675 940235
rect 600761 940199 600817 940235
rect 600903 940199 600959 940235
rect 601045 940199 601101 940235
rect 599341 940111 599382 940113
rect 599382 940111 599397 940113
rect 599483 940111 599506 940113
rect 599506 940111 599539 940113
rect 599625 940111 599630 940113
rect 599630 940111 599681 940113
rect 599767 940111 599822 940113
rect 599822 940111 599823 940113
rect 599909 940111 599946 940113
rect 599946 940111 599965 940113
rect 600051 940111 600070 940113
rect 600070 940111 600107 940113
rect 600193 940111 600194 940113
rect 600194 940111 600249 940113
rect 600335 940111 600374 940113
rect 600374 940111 600391 940113
rect 600477 940111 600498 940113
rect 600498 940111 600533 940113
rect 600619 940111 600622 940113
rect 600622 940111 600675 940113
rect 600761 940111 600814 940113
rect 600814 940111 600817 940113
rect 600903 940111 600938 940113
rect 600938 940111 600959 940113
rect 601045 940111 601062 940113
rect 601062 940111 601101 940113
rect 599341 940057 599397 940111
rect 599483 940057 599539 940111
rect 599625 940057 599681 940111
rect 599767 940057 599823 940111
rect 599909 940057 599965 940111
rect 600051 940057 600107 940111
rect 600193 940057 600249 940111
rect 600335 940057 600391 940111
rect 600477 940057 600533 940111
rect 600619 940057 600675 940111
rect 600761 940057 600817 940111
rect 600903 940057 600959 940111
rect 601045 940057 601101 940111
rect 599341 939919 599397 939971
rect 599483 939919 599539 939971
rect 599625 939919 599681 939971
rect 599767 939919 599823 939971
rect 599909 939919 599965 939971
rect 600051 939919 600107 939971
rect 600193 939919 600249 939971
rect 600335 939919 600391 939971
rect 600477 939919 600533 939971
rect 600619 939919 600675 939971
rect 600761 939919 600817 939971
rect 600903 939919 600959 939971
rect 601045 939919 601101 939971
rect 599341 939915 599382 939919
rect 599382 939915 599397 939919
rect 599483 939915 599506 939919
rect 599506 939915 599539 939919
rect 599625 939915 599630 939919
rect 599630 939915 599681 939919
rect 599767 939915 599822 939919
rect 599822 939915 599823 939919
rect 599909 939915 599946 939919
rect 599946 939915 599965 939919
rect 600051 939915 600070 939919
rect 600070 939915 600107 939919
rect 600193 939915 600194 939919
rect 600194 939915 600249 939919
rect 600335 939915 600374 939919
rect 600374 939915 600391 939919
rect 600477 939915 600498 939919
rect 600498 939915 600533 939919
rect 600619 939915 600622 939919
rect 600622 939915 600675 939919
rect 600761 939915 600814 939919
rect 600814 939915 600817 939919
rect 600903 939915 600938 939919
rect 600938 939915 600959 939919
rect 601045 939915 601062 939919
rect 601062 939915 601101 939919
rect 599341 939773 599397 939829
rect 599483 939773 599539 939829
rect 599625 939773 599681 939829
rect 599767 939773 599823 939829
rect 599909 939773 599965 939829
rect 600051 939773 600107 939829
rect 600193 939773 600249 939829
rect 600335 939773 600391 939829
rect 600477 939773 600533 939829
rect 600619 939773 600675 939829
rect 600761 939773 600817 939829
rect 600903 939773 600959 939829
rect 601045 939773 601101 939829
rect 601829 941655 601885 941675
rect 601971 941655 602027 941675
rect 602113 941655 602169 941675
rect 602255 941655 602311 941675
rect 602397 941655 602453 941675
rect 602539 941655 602595 941675
rect 602681 941655 602737 941675
rect 602823 941655 602879 941675
rect 602965 941655 603021 941675
rect 603107 941655 603163 941675
rect 603249 941655 603305 941675
rect 603391 941655 603447 941675
rect 603533 941655 603589 941675
rect 603675 941655 603731 941675
rect 601829 941619 601832 941655
rect 601832 941619 601885 941655
rect 601971 941619 602012 941655
rect 602012 941619 602027 941655
rect 602113 941619 602136 941655
rect 602136 941619 602169 941655
rect 602255 941619 602260 941655
rect 602260 941619 602311 941655
rect 602397 941619 602452 941655
rect 602452 941619 602453 941655
rect 602539 941619 602576 941655
rect 602576 941619 602595 941655
rect 602681 941619 602700 941655
rect 602700 941619 602737 941655
rect 602823 941619 602824 941655
rect 602824 941619 602879 941655
rect 602965 941619 603004 941655
rect 603004 941619 603021 941655
rect 603107 941619 603128 941655
rect 603128 941619 603163 941655
rect 603249 941619 603252 941655
rect 603252 941619 603305 941655
rect 603391 941619 603444 941655
rect 603444 941619 603447 941655
rect 603533 941619 603568 941655
rect 603568 941619 603589 941655
rect 603675 941619 603692 941655
rect 603692 941619 603731 941655
rect 601829 941531 601885 941533
rect 601971 941531 602027 941533
rect 602113 941531 602169 941533
rect 602255 941531 602311 941533
rect 602397 941531 602453 941533
rect 602539 941531 602595 941533
rect 602681 941531 602737 941533
rect 602823 941531 602879 941533
rect 602965 941531 603021 941533
rect 603107 941531 603163 941533
rect 603249 941531 603305 941533
rect 603391 941531 603447 941533
rect 603533 941531 603589 941533
rect 603675 941531 603731 941533
rect 601829 941477 601832 941531
rect 601832 941477 601885 941531
rect 601971 941477 602012 941531
rect 602012 941477 602027 941531
rect 602113 941477 602136 941531
rect 602136 941477 602169 941531
rect 602255 941477 602260 941531
rect 602260 941477 602311 941531
rect 602397 941477 602452 941531
rect 602452 941477 602453 941531
rect 602539 941477 602576 941531
rect 602576 941477 602595 941531
rect 602681 941477 602700 941531
rect 602700 941477 602737 941531
rect 602823 941477 602824 941531
rect 602824 941477 602879 941531
rect 602965 941477 603004 941531
rect 603004 941477 603021 941531
rect 603107 941477 603128 941531
rect 603128 941477 603163 941531
rect 603249 941477 603252 941531
rect 603252 941477 603305 941531
rect 603391 941477 603444 941531
rect 603444 941477 603447 941531
rect 603533 941477 603568 941531
rect 603568 941477 603589 941531
rect 603675 941477 603692 941531
rect 603692 941477 603731 941531
rect 601829 941351 601832 941391
rect 601832 941351 601885 941391
rect 601971 941351 602012 941391
rect 602012 941351 602027 941391
rect 602113 941351 602136 941391
rect 602136 941351 602169 941391
rect 602255 941351 602260 941391
rect 602260 941351 602311 941391
rect 602397 941351 602452 941391
rect 602452 941351 602453 941391
rect 602539 941351 602576 941391
rect 602576 941351 602595 941391
rect 602681 941351 602700 941391
rect 602700 941351 602737 941391
rect 602823 941351 602824 941391
rect 602824 941351 602879 941391
rect 602965 941351 603004 941391
rect 603004 941351 603021 941391
rect 603107 941351 603128 941391
rect 603128 941351 603163 941391
rect 603249 941351 603252 941391
rect 603252 941351 603305 941391
rect 603391 941351 603444 941391
rect 603444 941351 603447 941391
rect 603533 941351 603568 941391
rect 603568 941351 603589 941391
rect 603675 941351 603692 941391
rect 603692 941351 603731 941391
rect 601829 941335 601885 941351
rect 601971 941335 602027 941351
rect 602113 941335 602169 941351
rect 602255 941335 602311 941351
rect 602397 941335 602453 941351
rect 602539 941335 602595 941351
rect 602681 941335 602737 941351
rect 602823 941335 602879 941351
rect 602965 941335 603021 941351
rect 603107 941335 603163 941351
rect 603249 941335 603305 941351
rect 603391 941335 603447 941351
rect 603533 941335 603589 941351
rect 603675 941335 603731 941351
rect 601829 941227 601832 941249
rect 601832 941227 601885 941249
rect 601971 941227 602012 941249
rect 602012 941227 602027 941249
rect 602113 941227 602136 941249
rect 602136 941227 602169 941249
rect 602255 941227 602260 941249
rect 602260 941227 602311 941249
rect 602397 941227 602452 941249
rect 602452 941227 602453 941249
rect 602539 941227 602576 941249
rect 602576 941227 602595 941249
rect 602681 941227 602700 941249
rect 602700 941227 602737 941249
rect 602823 941227 602824 941249
rect 602824 941227 602879 941249
rect 602965 941227 603004 941249
rect 603004 941227 603021 941249
rect 603107 941227 603128 941249
rect 603128 941227 603163 941249
rect 603249 941227 603252 941249
rect 603252 941227 603305 941249
rect 603391 941227 603444 941249
rect 603444 941227 603447 941249
rect 603533 941227 603568 941249
rect 603568 941227 603589 941249
rect 603675 941227 603692 941249
rect 603692 941227 603731 941249
rect 601829 941193 601885 941227
rect 601971 941193 602027 941227
rect 602113 941193 602169 941227
rect 602255 941193 602311 941227
rect 602397 941193 602453 941227
rect 602539 941193 602595 941227
rect 602681 941193 602737 941227
rect 602823 941193 602879 941227
rect 602965 941193 603021 941227
rect 603107 941193 603163 941227
rect 603249 941193 603305 941227
rect 603391 941193 603447 941227
rect 603533 941193 603589 941227
rect 603675 941193 603731 941227
rect 601829 941103 601832 941107
rect 601832 941103 601885 941107
rect 601971 941103 602012 941107
rect 602012 941103 602027 941107
rect 602113 941103 602136 941107
rect 602136 941103 602169 941107
rect 602255 941103 602260 941107
rect 602260 941103 602311 941107
rect 602397 941103 602452 941107
rect 602452 941103 602453 941107
rect 602539 941103 602576 941107
rect 602576 941103 602595 941107
rect 602681 941103 602700 941107
rect 602700 941103 602737 941107
rect 602823 941103 602824 941107
rect 602824 941103 602879 941107
rect 602965 941103 603004 941107
rect 603004 941103 603021 941107
rect 603107 941103 603128 941107
rect 603128 941103 603163 941107
rect 603249 941103 603252 941107
rect 603252 941103 603305 941107
rect 603391 941103 603444 941107
rect 603444 941103 603447 941107
rect 603533 941103 603568 941107
rect 603568 941103 603589 941107
rect 603675 941103 603692 941107
rect 603692 941103 603731 941107
rect 601829 941051 601885 941103
rect 601971 941051 602027 941103
rect 602113 941051 602169 941103
rect 602255 941051 602311 941103
rect 602397 941051 602453 941103
rect 602539 941051 602595 941103
rect 602681 941051 602737 941103
rect 602823 941051 602879 941103
rect 602965 941051 603021 941103
rect 603107 941051 603163 941103
rect 603249 941051 603305 941103
rect 603391 941051 603447 941103
rect 603533 941051 603589 941103
rect 603675 941051 603731 941103
rect 601829 940911 601885 940965
rect 601971 940911 602027 940965
rect 602113 940911 602169 940965
rect 602255 940911 602311 940965
rect 602397 940911 602453 940965
rect 602539 940911 602595 940965
rect 602681 940911 602737 940965
rect 602823 940911 602879 940965
rect 602965 940911 603021 940965
rect 603107 940911 603163 940965
rect 603249 940911 603305 940965
rect 603391 940911 603447 940965
rect 603533 940911 603589 940965
rect 603675 940911 603731 940965
rect 601829 940909 601832 940911
rect 601832 940909 601885 940911
rect 601971 940909 602012 940911
rect 602012 940909 602027 940911
rect 602113 940909 602136 940911
rect 602136 940909 602169 940911
rect 602255 940909 602260 940911
rect 602260 940909 602311 940911
rect 602397 940909 602452 940911
rect 602452 940909 602453 940911
rect 602539 940909 602576 940911
rect 602576 940909 602595 940911
rect 602681 940909 602700 940911
rect 602700 940909 602737 940911
rect 602823 940909 602824 940911
rect 602824 940909 602879 940911
rect 602965 940909 603004 940911
rect 603004 940909 603021 940911
rect 603107 940909 603128 940911
rect 603128 940909 603163 940911
rect 603249 940909 603252 940911
rect 603252 940909 603305 940911
rect 603391 940909 603444 940911
rect 603444 940909 603447 940911
rect 603533 940909 603568 940911
rect 603568 940909 603589 940911
rect 603675 940909 603692 940911
rect 603692 940909 603731 940911
rect 601829 940787 601885 940823
rect 601971 940787 602027 940823
rect 602113 940787 602169 940823
rect 602255 940787 602311 940823
rect 602397 940787 602453 940823
rect 602539 940787 602595 940823
rect 602681 940787 602737 940823
rect 602823 940787 602879 940823
rect 602965 940787 603021 940823
rect 603107 940787 603163 940823
rect 603249 940787 603305 940823
rect 603391 940787 603447 940823
rect 603533 940787 603589 940823
rect 603675 940787 603731 940823
rect 601829 940767 601832 940787
rect 601832 940767 601885 940787
rect 601971 940767 602012 940787
rect 602012 940767 602027 940787
rect 602113 940767 602136 940787
rect 602136 940767 602169 940787
rect 602255 940767 602260 940787
rect 602260 940767 602311 940787
rect 602397 940767 602452 940787
rect 602452 940767 602453 940787
rect 602539 940767 602576 940787
rect 602576 940767 602595 940787
rect 602681 940767 602700 940787
rect 602700 940767 602737 940787
rect 602823 940767 602824 940787
rect 602824 940767 602879 940787
rect 602965 940767 603004 940787
rect 603004 940767 603021 940787
rect 603107 940767 603128 940787
rect 603128 940767 603163 940787
rect 603249 940767 603252 940787
rect 603252 940767 603305 940787
rect 603391 940767 603444 940787
rect 603444 940767 603447 940787
rect 603533 940767 603568 940787
rect 603568 940767 603589 940787
rect 603675 940767 603692 940787
rect 603692 940767 603731 940787
rect 601829 940663 601885 940681
rect 601971 940663 602027 940681
rect 602113 940663 602169 940681
rect 602255 940663 602311 940681
rect 602397 940663 602453 940681
rect 602539 940663 602595 940681
rect 602681 940663 602737 940681
rect 602823 940663 602879 940681
rect 602965 940663 603021 940681
rect 603107 940663 603163 940681
rect 603249 940663 603305 940681
rect 603391 940663 603447 940681
rect 603533 940663 603589 940681
rect 603675 940663 603731 940681
rect 601829 940625 601832 940663
rect 601832 940625 601885 940663
rect 601971 940625 602012 940663
rect 602012 940625 602027 940663
rect 602113 940625 602136 940663
rect 602136 940625 602169 940663
rect 602255 940625 602260 940663
rect 602260 940625 602311 940663
rect 602397 940625 602452 940663
rect 602452 940625 602453 940663
rect 602539 940625 602576 940663
rect 602576 940625 602595 940663
rect 602681 940625 602700 940663
rect 602700 940625 602737 940663
rect 602823 940625 602824 940663
rect 602824 940625 602879 940663
rect 602965 940625 603004 940663
rect 603004 940625 603021 940663
rect 603107 940625 603128 940663
rect 603128 940625 603163 940663
rect 603249 940625 603252 940663
rect 603252 940625 603305 940663
rect 603391 940625 603444 940663
rect 603444 940625 603447 940663
rect 603533 940625 603568 940663
rect 603568 940625 603589 940663
rect 603675 940625 603692 940663
rect 603692 940625 603731 940663
rect 601829 940483 601832 940539
rect 601832 940483 601885 940539
rect 601971 940483 602012 940539
rect 602012 940483 602027 940539
rect 602113 940483 602136 940539
rect 602136 940483 602169 940539
rect 602255 940483 602260 940539
rect 602260 940483 602311 940539
rect 602397 940483 602452 940539
rect 602452 940483 602453 940539
rect 602539 940483 602576 940539
rect 602576 940483 602595 940539
rect 602681 940483 602700 940539
rect 602700 940483 602737 940539
rect 602823 940483 602824 940539
rect 602824 940483 602879 940539
rect 602965 940483 603004 940539
rect 603004 940483 603021 940539
rect 603107 940483 603128 940539
rect 603128 940483 603163 940539
rect 603249 940483 603252 940539
rect 603252 940483 603305 940539
rect 603391 940483 603444 940539
rect 603444 940483 603447 940539
rect 603533 940483 603568 940539
rect 603568 940483 603589 940539
rect 603675 940483 603692 940539
rect 603692 940483 603731 940539
rect 601829 940359 601832 940397
rect 601832 940359 601885 940397
rect 601971 940359 602012 940397
rect 602012 940359 602027 940397
rect 602113 940359 602136 940397
rect 602136 940359 602169 940397
rect 602255 940359 602260 940397
rect 602260 940359 602311 940397
rect 602397 940359 602452 940397
rect 602452 940359 602453 940397
rect 602539 940359 602576 940397
rect 602576 940359 602595 940397
rect 602681 940359 602700 940397
rect 602700 940359 602737 940397
rect 602823 940359 602824 940397
rect 602824 940359 602879 940397
rect 602965 940359 603004 940397
rect 603004 940359 603021 940397
rect 603107 940359 603128 940397
rect 603128 940359 603163 940397
rect 603249 940359 603252 940397
rect 603252 940359 603305 940397
rect 603391 940359 603444 940397
rect 603444 940359 603447 940397
rect 603533 940359 603568 940397
rect 603568 940359 603589 940397
rect 603675 940359 603692 940397
rect 603692 940359 603731 940397
rect 601829 940341 601885 940359
rect 601971 940341 602027 940359
rect 602113 940341 602169 940359
rect 602255 940341 602311 940359
rect 602397 940341 602453 940359
rect 602539 940341 602595 940359
rect 602681 940341 602737 940359
rect 602823 940341 602879 940359
rect 602965 940341 603021 940359
rect 603107 940341 603163 940359
rect 603249 940341 603305 940359
rect 603391 940341 603447 940359
rect 603533 940341 603589 940359
rect 603675 940341 603731 940359
rect 601829 940235 601832 940255
rect 601832 940235 601885 940255
rect 601971 940235 602012 940255
rect 602012 940235 602027 940255
rect 602113 940235 602136 940255
rect 602136 940235 602169 940255
rect 602255 940235 602260 940255
rect 602260 940235 602311 940255
rect 602397 940235 602452 940255
rect 602452 940235 602453 940255
rect 602539 940235 602576 940255
rect 602576 940235 602595 940255
rect 602681 940235 602700 940255
rect 602700 940235 602737 940255
rect 602823 940235 602824 940255
rect 602824 940235 602879 940255
rect 602965 940235 603004 940255
rect 603004 940235 603021 940255
rect 603107 940235 603128 940255
rect 603128 940235 603163 940255
rect 603249 940235 603252 940255
rect 603252 940235 603305 940255
rect 603391 940235 603444 940255
rect 603444 940235 603447 940255
rect 603533 940235 603568 940255
rect 603568 940235 603589 940255
rect 603675 940235 603692 940255
rect 603692 940235 603731 940255
rect 601829 940199 601885 940235
rect 601971 940199 602027 940235
rect 602113 940199 602169 940235
rect 602255 940199 602311 940235
rect 602397 940199 602453 940235
rect 602539 940199 602595 940235
rect 602681 940199 602737 940235
rect 602823 940199 602879 940235
rect 602965 940199 603021 940235
rect 603107 940199 603163 940235
rect 603249 940199 603305 940235
rect 603391 940199 603447 940235
rect 603533 940199 603589 940235
rect 603675 940199 603731 940235
rect 601829 940111 601832 940113
rect 601832 940111 601885 940113
rect 601971 940111 602012 940113
rect 602012 940111 602027 940113
rect 602113 940111 602136 940113
rect 602136 940111 602169 940113
rect 602255 940111 602260 940113
rect 602260 940111 602311 940113
rect 602397 940111 602452 940113
rect 602452 940111 602453 940113
rect 602539 940111 602576 940113
rect 602576 940111 602595 940113
rect 602681 940111 602700 940113
rect 602700 940111 602737 940113
rect 602823 940111 602824 940113
rect 602824 940111 602879 940113
rect 602965 940111 603004 940113
rect 603004 940111 603021 940113
rect 603107 940111 603128 940113
rect 603128 940111 603163 940113
rect 603249 940111 603252 940113
rect 603252 940111 603305 940113
rect 603391 940111 603444 940113
rect 603444 940111 603447 940113
rect 603533 940111 603568 940113
rect 603568 940111 603589 940113
rect 603675 940111 603692 940113
rect 603692 940111 603731 940113
rect 601829 940057 601885 940111
rect 601971 940057 602027 940111
rect 602113 940057 602169 940111
rect 602255 940057 602311 940111
rect 602397 940057 602453 940111
rect 602539 940057 602595 940111
rect 602681 940057 602737 940111
rect 602823 940057 602879 940111
rect 602965 940057 603021 940111
rect 603107 940057 603163 940111
rect 603249 940057 603305 940111
rect 603391 940057 603447 940111
rect 603533 940057 603589 940111
rect 603675 940057 603731 940111
rect 601829 939919 601885 939971
rect 601971 939919 602027 939971
rect 602113 939919 602169 939971
rect 602255 939919 602311 939971
rect 602397 939919 602453 939971
rect 602539 939919 602595 939971
rect 602681 939919 602737 939971
rect 602823 939919 602879 939971
rect 602965 939919 603021 939971
rect 603107 939919 603163 939971
rect 603249 939919 603305 939971
rect 603391 939919 603447 939971
rect 603533 939919 603589 939971
rect 603675 939919 603731 939971
rect 601829 939915 601832 939919
rect 601832 939915 601885 939919
rect 601971 939915 602012 939919
rect 602012 939915 602027 939919
rect 602113 939915 602136 939919
rect 602136 939915 602169 939919
rect 602255 939915 602260 939919
rect 602260 939915 602311 939919
rect 602397 939915 602452 939919
rect 602452 939915 602453 939919
rect 602539 939915 602576 939919
rect 602576 939915 602595 939919
rect 602681 939915 602700 939919
rect 602700 939915 602737 939919
rect 602823 939915 602824 939919
rect 602824 939915 602879 939919
rect 602965 939915 603004 939919
rect 603004 939915 603021 939919
rect 603107 939915 603128 939919
rect 603128 939915 603163 939919
rect 603249 939915 603252 939919
rect 603252 939915 603305 939919
rect 603391 939915 603444 939919
rect 603444 939915 603447 939919
rect 603533 939915 603568 939919
rect 603568 939915 603589 939919
rect 603675 939915 603692 939919
rect 603692 939915 603731 939919
rect 601829 939773 601885 939829
rect 601971 939773 602027 939829
rect 602113 939773 602169 939829
rect 602255 939773 602311 939829
rect 602397 939773 602453 939829
rect 602539 939773 602595 939829
rect 602681 939773 602737 939829
rect 602823 939773 602879 939829
rect 602965 939773 603021 939829
rect 603107 939773 603163 939829
rect 603249 939773 603305 939829
rect 603391 939773 603447 939829
rect 603533 939773 603589 939829
rect 603675 939773 603731 939829
rect 605051 941655 605107 941675
rect 605193 941655 605249 941675
rect 605335 941655 605391 941675
rect 605477 941655 605533 941675
rect 605619 941655 605675 941675
rect 605761 941655 605817 941675
rect 605903 941655 605959 941675
rect 606045 941655 606101 941675
rect 605051 941619 605070 941655
rect 605070 941619 605107 941655
rect 605193 941619 605194 941655
rect 605194 941619 605249 941655
rect 605335 941619 605374 941655
rect 605374 941619 605391 941655
rect 605477 941619 605498 941655
rect 605498 941619 605533 941655
rect 605619 941619 605622 941655
rect 605622 941619 605675 941655
rect 605761 941619 605814 941655
rect 605814 941619 605817 941655
rect 605903 941619 605938 941655
rect 605938 941619 605959 941655
rect 606045 941619 606062 941655
rect 606062 941619 606101 941655
rect 605051 941531 605107 941533
rect 605193 941531 605249 941533
rect 605335 941531 605391 941533
rect 605477 941531 605533 941533
rect 605619 941531 605675 941533
rect 605761 941531 605817 941533
rect 605903 941531 605959 941533
rect 606045 941531 606101 941533
rect 605051 941477 605070 941531
rect 605070 941477 605107 941531
rect 605193 941477 605194 941531
rect 605194 941477 605249 941531
rect 605335 941477 605374 941531
rect 605374 941477 605391 941531
rect 605477 941477 605498 941531
rect 605498 941477 605533 941531
rect 605619 941477 605622 941531
rect 605622 941477 605675 941531
rect 605761 941477 605814 941531
rect 605814 941477 605817 941531
rect 605903 941477 605938 941531
rect 605938 941477 605959 941531
rect 606045 941477 606062 941531
rect 606062 941477 606101 941531
rect 605051 941351 605070 941391
rect 605070 941351 605107 941391
rect 605193 941351 605194 941391
rect 605194 941351 605249 941391
rect 605335 941351 605374 941391
rect 605374 941351 605391 941391
rect 605477 941351 605498 941391
rect 605498 941351 605533 941391
rect 605619 941351 605622 941391
rect 605622 941351 605675 941391
rect 605761 941351 605814 941391
rect 605814 941351 605817 941391
rect 605903 941351 605938 941391
rect 605938 941351 605959 941391
rect 606045 941351 606062 941391
rect 606062 941351 606101 941391
rect 605051 941335 605107 941351
rect 605193 941335 605249 941351
rect 605335 941335 605391 941351
rect 605477 941335 605533 941351
rect 605619 941335 605675 941351
rect 605761 941335 605817 941351
rect 605903 941335 605959 941351
rect 606045 941335 606101 941351
rect 605051 941227 605070 941249
rect 605070 941227 605107 941249
rect 605193 941227 605194 941249
rect 605194 941227 605249 941249
rect 605335 941227 605374 941249
rect 605374 941227 605391 941249
rect 605477 941227 605498 941249
rect 605498 941227 605533 941249
rect 605619 941227 605622 941249
rect 605622 941227 605675 941249
rect 605761 941227 605814 941249
rect 605814 941227 605817 941249
rect 605903 941227 605938 941249
rect 605938 941227 605959 941249
rect 606045 941227 606062 941249
rect 606062 941227 606101 941249
rect 605051 941193 605107 941227
rect 605193 941193 605249 941227
rect 605335 941193 605391 941227
rect 605477 941193 605533 941227
rect 605619 941193 605675 941227
rect 605761 941193 605817 941227
rect 605903 941193 605959 941227
rect 606045 941193 606101 941227
rect 605051 941103 605070 941107
rect 605070 941103 605107 941107
rect 605193 941103 605194 941107
rect 605194 941103 605249 941107
rect 605335 941103 605374 941107
rect 605374 941103 605391 941107
rect 605477 941103 605498 941107
rect 605498 941103 605533 941107
rect 605619 941103 605622 941107
rect 605622 941103 605675 941107
rect 605761 941103 605814 941107
rect 605814 941103 605817 941107
rect 605903 941103 605938 941107
rect 605938 941103 605959 941107
rect 606045 941103 606062 941107
rect 606062 941103 606101 941107
rect 605051 941051 605107 941103
rect 605193 941051 605249 941103
rect 605335 941051 605391 941103
rect 605477 941051 605533 941103
rect 605619 941051 605675 941103
rect 605761 941051 605817 941103
rect 605903 941051 605959 941103
rect 606045 941051 606101 941103
rect 605051 940911 605107 940965
rect 605193 940911 605249 940965
rect 605335 940911 605391 940965
rect 605477 940911 605533 940965
rect 605619 940911 605675 940965
rect 605761 940911 605817 940965
rect 605903 940911 605959 940965
rect 606045 940911 606101 940965
rect 605051 940909 605070 940911
rect 605070 940909 605107 940911
rect 605193 940909 605194 940911
rect 605194 940909 605249 940911
rect 605335 940909 605374 940911
rect 605374 940909 605391 940911
rect 605477 940909 605498 940911
rect 605498 940909 605533 940911
rect 605619 940909 605622 940911
rect 605622 940909 605675 940911
rect 605761 940909 605814 940911
rect 605814 940909 605817 940911
rect 605903 940909 605938 940911
rect 605938 940909 605959 940911
rect 606045 940909 606062 940911
rect 606062 940909 606101 940911
rect 605051 940787 605107 940823
rect 605193 940787 605249 940823
rect 605335 940787 605391 940823
rect 605477 940787 605533 940823
rect 605619 940787 605675 940823
rect 605761 940787 605817 940823
rect 605903 940787 605959 940823
rect 606045 940787 606101 940823
rect 605051 940767 605070 940787
rect 605070 940767 605107 940787
rect 605193 940767 605194 940787
rect 605194 940767 605249 940787
rect 605335 940767 605374 940787
rect 605374 940767 605391 940787
rect 605477 940767 605498 940787
rect 605498 940767 605533 940787
rect 605619 940767 605622 940787
rect 605622 940767 605675 940787
rect 605761 940767 605814 940787
rect 605814 940767 605817 940787
rect 605903 940767 605938 940787
rect 605938 940767 605959 940787
rect 606045 940767 606062 940787
rect 606062 940767 606101 940787
rect 605051 940663 605107 940681
rect 605193 940663 605249 940681
rect 605335 940663 605391 940681
rect 605477 940663 605533 940681
rect 605619 940663 605675 940681
rect 605761 940663 605817 940681
rect 605903 940663 605959 940681
rect 606045 940663 606101 940681
rect 605051 940625 605070 940663
rect 605070 940625 605107 940663
rect 605193 940625 605194 940663
rect 605194 940625 605249 940663
rect 605335 940625 605374 940663
rect 605374 940625 605391 940663
rect 605477 940625 605498 940663
rect 605498 940625 605533 940663
rect 605619 940625 605622 940663
rect 605622 940625 605675 940663
rect 605761 940625 605814 940663
rect 605814 940625 605817 940663
rect 605903 940625 605938 940663
rect 605938 940625 605959 940663
rect 606045 940625 606062 940663
rect 606062 940625 606101 940663
rect 605051 940483 605070 940539
rect 605070 940483 605107 940539
rect 605193 940483 605194 940539
rect 605194 940483 605249 940539
rect 605335 940483 605374 940539
rect 605374 940483 605391 940539
rect 605477 940483 605498 940539
rect 605498 940483 605533 940539
rect 605619 940483 605622 940539
rect 605622 940483 605675 940539
rect 605761 940483 605814 940539
rect 605814 940483 605817 940539
rect 605903 940483 605938 940539
rect 605938 940483 605959 940539
rect 606045 940483 606062 940539
rect 606062 940483 606101 940539
rect 605051 940359 605070 940397
rect 605070 940359 605107 940397
rect 605193 940359 605194 940397
rect 605194 940359 605249 940397
rect 605335 940359 605374 940397
rect 605374 940359 605391 940397
rect 605477 940359 605498 940397
rect 605498 940359 605533 940397
rect 605619 940359 605622 940397
rect 605622 940359 605675 940397
rect 605761 940359 605814 940397
rect 605814 940359 605817 940397
rect 605903 940359 605938 940397
rect 605938 940359 605959 940397
rect 606045 940359 606062 940397
rect 606062 940359 606101 940397
rect 605051 940341 605107 940359
rect 605193 940341 605249 940359
rect 605335 940341 605391 940359
rect 605477 940341 605533 940359
rect 605619 940341 605675 940359
rect 605761 940341 605817 940359
rect 605903 940341 605959 940359
rect 606045 940341 606101 940359
rect 605051 940235 605070 940255
rect 605070 940235 605107 940255
rect 605193 940235 605194 940255
rect 605194 940235 605249 940255
rect 605335 940235 605374 940255
rect 605374 940235 605391 940255
rect 605477 940235 605498 940255
rect 605498 940235 605533 940255
rect 605619 940235 605622 940255
rect 605622 940235 605675 940255
rect 605761 940235 605814 940255
rect 605814 940235 605817 940255
rect 605903 940235 605938 940255
rect 605938 940235 605959 940255
rect 606045 940235 606062 940255
rect 606062 940235 606101 940255
rect 605051 940199 605107 940235
rect 605193 940199 605249 940235
rect 605335 940199 605391 940235
rect 605477 940199 605533 940235
rect 605619 940199 605675 940235
rect 605761 940199 605817 940235
rect 605903 940199 605959 940235
rect 606045 940199 606101 940235
rect 605051 940111 605070 940113
rect 605070 940111 605107 940113
rect 605193 940111 605194 940113
rect 605194 940111 605249 940113
rect 605335 940111 605374 940113
rect 605374 940111 605391 940113
rect 605477 940111 605498 940113
rect 605498 940111 605533 940113
rect 605619 940111 605622 940113
rect 605622 940111 605675 940113
rect 605761 940111 605814 940113
rect 605814 940111 605817 940113
rect 605903 940111 605938 940113
rect 605938 940111 605959 940113
rect 606045 940111 606062 940113
rect 606062 940111 606101 940113
rect 605051 940057 605107 940111
rect 605193 940057 605249 940111
rect 605335 940057 605391 940111
rect 605477 940057 605533 940111
rect 605619 940057 605675 940111
rect 605761 940057 605817 940111
rect 605903 940057 605959 940111
rect 606045 940057 606101 940111
rect 605051 939919 605107 939971
rect 605193 939919 605249 939971
rect 605335 939919 605391 939971
rect 605477 939919 605533 939971
rect 605619 939919 605675 939971
rect 605761 939919 605817 939971
rect 605903 939919 605959 939971
rect 606045 939919 606101 939971
rect 605051 939915 605070 939919
rect 605070 939915 605107 939919
rect 605193 939915 605194 939919
rect 605194 939915 605249 939919
rect 605335 939915 605374 939919
rect 605374 939915 605391 939919
rect 605477 939915 605498 939919
rect 605498 939915 605533 939919
rect 605619 939915 605622 939919
rect 605622 939915 605675 939919
rect 605761 939915 605814 939919
rect 605814 939915 605817 939919
rect 605903 939915 605938 939919
rect 605938 939915 605959 939919
rect 606045 939915 606062 939919
rect 606062 939915 606101 939919
rect 605051 939773 605107 939829
rect 605193 939773 605249 939829
rect 605335 939773 605391 939829
rect 605477 939773 605533 939829
rect 605619 939773 605675 939829
rect 605761 939773 605817 939829
rect 605903 939773 605959 939829
rect 606045 939773 606101 939829
rect 606905 941655 606961 941675
rect 607047 941655 607103 941675
rect 607189 941655 607245 941675
rect 607331 941655 607387 941675
rect 607473 941655 607529 941675
rect 607615 941655 607671 941675
rect 607757 941655 607813 941675
rect 607899 941655 607955 941675
rect 608041 941655 608097 941675
rect 608183 941655 608239 941675
rect 608325 941655 608381 941675
rect 608467 941655 608523 941675
rect 608609 941655 608665 941675
rect 608751 941655 608807 941675
rect 606905 941619 606908 941655
rect 606908 941619 606961 941655
rect 607047 941619 607088 941655
rect 607088 941619 607103 941655
rect 607189 941619 607212 941655
rect 607212 941619 607245 941655
rect 607331 941619 607336 941655
rect 607336 941619 607387 941655
rect 607473 941619 607528 941655
rect 607528 941619 607529 941655
rect 607615 941619 607652 941655
rect 607652 941619 607671 941655
rect 607757 941619 607776 941655
rect 607776 941619 607813 941655
rect 607899 941619 607900 941655
rect 607900 941619 607955 941655
rect 608041 941619 608080 941655
rect 608080 941619 608097 941655
rect 608183 941619 608204 941655
rect 608204 941619 608239 941655
rect 608325 941619 608328 941655
rect 608328 941619 608381 941655
rect 608467 941619 608520 941655
rect 608520 941619 608523 941655
rect 608609 941619 608644 941655
rect 608644 941619 608665 941655
rect 608751 941619 608768 941655
rect 608768 941619 608807 941655
rect 606905 941531 606961 941533
rect 607047 941531 607103 941533
rect 607189 941531 607245 941533
rect 607331 941531 607387 941533
rect 607473 941531 607529 941533
rect 607615 941531 607671 941533
rect 607757 941531 607813 941533
rect 607899 941531 607955 941533
rect 608041 941531 608097 941533
rect 608183 941531 608239 941533
rect 608325 941531 608381 941533
rect 608467 941531 608523 941533
rect 608609 941531 608665 941533
rect 608751 941531 608807 941533
rect 606905 941477 606908 941531
rect 606908 941477 606961 941531
rect 607047 941477 607088 941531
rect 607088 941477 607103 941531
rect 607189 941477 607212 941531
rect 607212 941477 607245 941531
rect 607331 941477 607336 941531
rect 607336 941477 607387 941531
rect 607473 941477 607528 941531
rect 607528 941477 607529 941531
rect 607615 941477 607652 941531
rect 607652 941477 607671 941531
rect 607757 941477 607776 941531
rect 607776 941477 607813 941531
rect 607899 941477 607900 941531
rect 607900 941477 607955 941531
rect 608041 941477 608080 941531
rect 608080 941477 608097 941531
rect 608183 941477 608204 941531
rect 608204 941477 608239 941531
rect 608325 941477 608328 941531
rect 608328 941477 608381 941531
rect 608467 941477 608520 941531
rect 608520 941477 608523 941531
rect 608609 941477 608644 941531
rect 608644 941477 608665 941531
rect 608751 941477 608768 941531
rect 608768 941477 608807 941531
rect 606905 941351 606908 941391
rect 606908 941351 606961 941391
rect 607047 941351 607088 941391
rect 607088 941351 607103 941391
rect 607189 941351 607212 941391
rect 607212 941351 607245 941391
rect 607331 941351 607336 941391
rect 607336 941351 607387 941391
rect 607473 941351 607528 941391
rect 607528 941351 607529 941391
rect 607615 941351 607652 941391
rect 607652 941351 607671 941391
rect 607757 941351 607776 941391
rect 607776 941351 607813 941391
rect 607899 941351 607900 941391
rect 607900 941351 607955 941391
rect 608041 941351 608080 941391
rect 608080 941351 608097 941391
rect 608183 941351 608204 941391
rect 608204 941351 608239 941391
rect 608325 941351 608328 941391
rect 608328 941351 608381 941391
rect 608467 941351 608520 941391
rect 608520 941351 608523 941391
rect 608609 941351 608644 941391
rect 608644 941351 608665 941391
rect 608751 941351 608768 941391
rect 608768 941351 608807 941391
rect 606905 941335 606961 941351
rect 607047 941335 607103 941351
rect 607189 941335 607245 941351
rect 607331 941335 607387 941351
rect 607473 941335 607529 941351
rect 607615 941335 607671 941351
rect 607757 941335 607813 941351
rect 607899 941335 607955 941351
rect 608041 941335 608097 941351
rect 608183 941335 608239 941351
rect 608325 941335 608381 941351
rect 608467 941335 608523 941351
rect 608609 941335 608665 941351
rect 608751 941335 608807 941351
rect 606905 941227 606908 941249
rect 606908 941227 606961 941249
rect 607047 941227 607088 941249
rect 607088 941227 607103 941249
rect 607189 941227 607212 941249
rect 607212 941227 607245 941249
rect 607331 941227 607336 941249
rect 607336 941227 607387 941249
rect 607473 941227 607528 941249
rect 607528 941227 607529 941249
rect 607615 941227 607652 941249
rect 607652 941227 607671 941249
rect 607757 941227 607776 941249
rect 607776 941227 607813 941249
rect 607899 941227 607900 941249
rect 607900 941227 607955 941249
rect 608041 941227 608080 941249
rect 608080 941227 608097 941249
rect 608183 941227 608204 941249
rect 608204 941227 608239 941249
rect 608325 941227 608328 941249
rect 608328 941227 608381 941249
rect 608467 941227 608520 941249
rect 608520 941227 608523 941249
rect 608609 941227 608644 941249
rect 608644 941227 608665 941249
rect 608751 941227 608768 941249
rect 608768 941227 608807 941249
rect 606905 941193 606961 941227
rect 607047 941193 607103 941227
rect 607189 941193 607245 941227
rect 607331 941193 607387 941227
rect 607473 941193 607529 941227
rect 607615 941193 607671 941227
rect 607757 941193 607813 941227
rect 607899 941193 607955 941227
rect 608041 941193 608097 941227
rect 608183 941193 608239 941227
rect 608325 941193 608381 941227
rect 608467 941193 608523 941227
rect 608609 941193 608665 941227
rect 608751 941193 608807 941227
rect 606905 941103 606908 941107
rect 606908 941103 606961 941107
rect 607047 941103 607088 941107
rect 607088 941103 607103 941107
rect 607189 941103 607212 941107
rect 607212 941103 607245 941107
rect 607331 941103 607336 941107
rect 607336 941103 607387 941107
rect 607473 941103 607528 941107
rect 607528 941103 607529 941107
rect 607615 941103 607652 941107
rect 607652 941103 607671 941107
rect 607757 941103 607776 941107
rect 607776 941103 607813 941107
rect 607899 941103 607900 941107
rect 607900 941103 607955 941107
rect 608041 941103 608080 941107
rect 608080 941103 608097 941107
rect 608183 941103 608204 941107
rect 608204 941103 608239 941107
rect 608325 941103 608328 941107
rect 608328 941103 608381 941107
rect 608467 941103 608520 941107
rect 608520 941103 608523 941107
rect 608609 941103 608644 941107
rect 608644 941103 608665 941107
rect 608751 941103 608768 941107
rect 608768 941103 608807 941107
rect 606905 941051 606961 941103
rect 607047 941051 607103 941103
rect 607189 941051 607245 941103
rect 607331 941051 607387 941103
rect 607473 941051 607529 941103
rect 607615 941051 607671 941103
rect 607757 941051 607813 941103
rect 607899 941051 607955 941103
rect 608041 941051 608097 941103
rect 608183 941051 608239 941103
rect 608325 941051 608381 941103
rect 608467 941051 608523 941103
rect 608609 941051 608665 941103
rect 608751 941051 608807 941103
rect 606905 940911 606961 940965
rect 607047 940911 607103 940965
rect 607189 940911 607245 940965
rect 607331 940911 607387 940965
rect 607473 940911 607529 940965
rect 607615 940911 607671 940965
rect 607757 940911 607813 940965
rect 607899 940911 607955 940965
rect 608041 940911 608097 940965
rect 608183 940911 608239 940965
rect 608325 940911 608381 940965
rect 608467 940911 608523 940965
rect 608609 940911 608665 940965
rect 608751 940911 608807 940965
rect 606905 940909 606908 940911
rect 606908 940909 606961 940911
rect 607047 940909 607088 940911
rect 607088 940909 607103 940911
rect 607189 940909 607212 940911
rect 607212 940909 607245 940911
rect 607331 940909 607336 940911
rect 607336 940909 607387 940911
rect 607473 940909 607528 940911
rect 607528 940909 607529 940911
rect 607615 940909 607652 940911
rect 607652 940909 607671 940911
rect 607757 940909 607776 940911
rect 607776 940909 607813 940911
rect 607899 940909 607900 940911
rect 607900 940909 607955 940911
rect 608041 940909 608080 940911
rect 608080 940909 608097 940911
rect 608183 940909 608204 940911
rect 608204 940909 608239 940911
rect 608325 940909 608328 940911
rect 608328 940909 608381 940911
rect 608467 940909 608520 940911
rect 608520 940909 608523 940911
rect 608609 940909 608644 940911
rect 608644 940909 608665 940911
rect 608751 940909 608768 940911
rect 608768 940909 608807 940911
rect 606905 940787 606961 940823
rect 607047 940787 607103 940823
rect 607189 940787 607245 940823
rect 607331 940787 607387 940823
rect 607473 940787 607529 940823
rect 607615 940787 607671 940823
rect 607757 940787 607813 940823
rect 607899 940787 607955 940823
rect 608041 940787 608097 940823
rect 608183 940787 608239 940823
rect 608325 940787 608381 940823
rect 608467 940787 608523 940823
rect 608609 940787 608665 940823
rect 608751 940787 608807 940823
rect 606905 940767 606908 940787
rect 606908 940767 606961 940787
rect 607047 940767 607088 940787
rect 607088 940767 607103 940787
rect 607189 940767 607212 940787
rect 607212 940767 607245 940787
rect 607331 940767 607336 940787
rect 607336 940767 607387 940787
rect 607473 940767 607528 940787
rect 607528 940767 607529 940787
rect 607615 940767 607652 940787
rect 607652 940767 607671 940787
rect 607757 940767 607776 940787
rect 607776 940767 607813 940787
rect 607899 940767 607900 940787
rect 607900 940767 607955 940787
rect 608041 940767 608080 940787
rect 608080 940767 608097 940787
rect 608183 940767 608204 940787
rect 608204 940767 608239 940787
rect 608325 940767 608328 940787
rect 608328 940767 608381 940787
rect 608467 940767 608520 940787
rect 608520 940767 608523 940787
rect 608609 940767 608644 940787
rect 608644 940767 608665 940787
rect 608751 940767 608768 940787
rect 608768 940767 608807 940787
rect 606905 940663 606961 940681
rect 607047 940663 607103 940681
rect 607189 940663 607245 940681
rect 607331 940663 607387 940681
rect 607473 940663 607529 940681
rect 607615 940663 607671 940681
rect 607757 940663 607813 940681
rect 607899 940663 607955 940681
rect 608041 940663 608097 940681
rect 608183 940663 608239 940681
rect 608325 940663 608381 940681
rect 608467 940663 608523 940681
rect 608609 940663 608665 940681
rect 608751 940663 608807 940681
rect 606905 940625 606908 940663
rect 606908 940625 606961 940663
rect 607047 940625 607088 940663
rect 607088 940625 607103 940663
rect 607189 940625 607212 940663
rect 607212 940625 607245 940663
rect 607331 940625 607336 940663
rect 607336 940625 607387 940663
rect 607473 940625 607528 940663
rect 607528 940625 607529 940663
rect 607615 940625 607652 940663
rect 607652 940625 607671 940663
rect 607757 940625 607776 940663
rect 607776 940625 607813 940663
rect 607899 940625 607900 940663
rect 607900 940625 607955 940663
rect 608041 940625 608080 940663
rect 608080 940625 608097 940663
rect 608183 940625 608204 940663
rect 608204 940625 608239 940663
rect 608325 940625 608328 940663
rect 608328 940625 608381 940663
rect 608467 940625 608520 940663
rect 608520 940625 608523 940663
rect 608609 940625 608644 940663
rect 608644 940625 608665 940663
rect 608751 940625 608768 940663
rect 608768 940625 608807 940663
rect 606905 940483 606908 940539
rect 606908 940483 606961 940539
rect 607047 940483 607088 940539
rect 607088 940483 607103 940539
rect 607189 940483 607212 940539
rect 607212 940483 607245 940539
rect 607331 940483 607336 940539
rect 607336 940483 607387 940539
rect 607473 940483 607528 940539
rect 607528 940483 607529 940539
rect 607615 940483 607652 940539
rect 607652 940483 607671 940539
rect 607757 940483 607776 940539
rect 607776 940483 607813 940539
rect 607899 940483 607900 940539
rect 607900 940483 607955 940539
rect 608041 940483 608080 940539
rect 608080 940483 608097 940539
rect 608183 940483 608204 940539
rect 608204 940483 608239 940539
rect 608325 940483 608328 940539
rect 608328 940483 608381 940539
rect 608467 940483 608520 940539
rect 608520 940483 608523 940539
rect 608609 940483 608644 940539
rect 608644 940483 608665 940539
rect 608751 940483 608768 940539
rect 608768 940483 608807 940539
rect 606905 940359 606908 940397
rect 606908 940359 606961 940397
rect 607047 940359 607088 940397
rect 607088 940359 607103 940397
rect 607189 940359 607212 940397
rect 607212 940359 607245 940397
rect 607331 940359 607336 940397
rect 607336 940359 607387 940397
rect 607473 940359 607528 940397
rect 607528 940359 607529 940397
rect 607615 940359 607652 940397
rect 607652 940359 607671 940397
rect 607757 940359 607776 940397
rect 607776 940359 607813 940397
rect 607899 940359 607900 940397
rect 607900 940359 607955 940397
rect 608041 940359 608080 940397
rect 608080 940359 608097 940397
rect 608183 940359 608204 940397
rect 608204 940359 608239 940397
rect 608325 940359 608328 940397
rect 608328 940359 608381 940397
rect 608467 940359 608520 940397
rect 608520 940359 608523 940397
rect 608609 940359 608644 940397
rect 608644 940359 608665 940397
rect 608751 940359 608768 940397
rect 608768 940359 608807 940397
rect 606905 940341 606961 940359
rect 607047 940341 607103 940359
rect 607189 940341 607245 940359
rect 607331 940341 607387 940359
rect 607473 940341 607529 940359
rect 607615 940341 607671 940359
rect 607757 940341 607813 940359
rect 607899 940341 607955 940359
rect 608041 940341 608097 940359
rect 608183 940341 608239 940359
rect 608325 940341 608381 940359
rect 608467 940341 608523 940359
rect 608609 940341 608665 940359
rect 608751 940341 608807 940359
rect 606905 940235 606908 940255
rect 606908 940235 606961 940255
rect 607047 940235 607088 940255
rect 607088 940235 607103 940255
rect 607189 940235 607212 940255
rect 607212 940235 607245 940255
rect 607331 940235 607336 940255
rect 607336 940235 607387 940255
rect 607473 940235 607528 940255
rect 607528 940235 607529 940255
rect 607615 940235 607652 940255
rect 607652 940235 607671 940255
rect 607757 940235 607776 940255
rect 607776 940235 607813 940255
rect 607899 940235 607900 940255
rect 607900 940235 607955 940255
rect 608041 940235 608080 940255
rect 608080 940235 608097 940255
rect 608183 940235 608204 940255
rect 608204 940235 608239 940255
rect 608325 940235 608328 940255
rect 608328 940235 608381 940255
rect 608467 940235 608520 940255
rect 608520 940235 608523 940255
rect 608609 940235 608644 940255
rect 608644 940235 608665 940255
rect 608751 940235 608768 940255
rect 608768 940235 608807 940255
rect 606905 940199 606961 940235
rect 607047 940199 607103 940235
rect 607189 940199 607245 940235
rect 607331 940199 607387 940235
rect 607473 940199 607529 940235
rect 607615 940199 607671 940235
rect 607757 940199 607813 940235
rect 607899 940199 607955 940235
rect 608041 940199 608097 940235
rect 608183 940199 608239 940235
rect 608325 940199 608381 940235
rect 608467 940199 608523 940235
rect 608609 940199 608665 940235
rect 608751 940199 608807 940235
rect 606905 940111 606908 940113
rect 606908 940111 606961 940113
rect 607047 940111 607088 940113
rect 607088 940111 607103 940113
rect 607189 940111 607212 940113
rect 607212 940111 607245 940113
rect 607331 940111 607336 940113
rect 607336 940111 607387 940113
rect 607473 940111 607528 940113
rect 607528 940111 607529 940113
rect 607615 940111 607652 940113
rect 607652 940111 607671 940113
rect 607757 940111 607776 940113
rect 607776 940111 607813 940113
rect 607899 940111 607900 940113
rect 607900 940111 607955 940113
rect 608041 940111 608080 940113
rect 608080 940111 608097 940113
rect 608183 940111 608204 940113
rect 608204 940111 608239 940113
rect 608325 940111 608328 940113
rect 608328 940111 608381 940113
rect 608467 940111 608520 940113
rect 608520 940111 608523 940113
rect 608609 940111 608644 940113
rect 608644 940111 608665 940113
rect 608751 940111 608768 940113
rect 608768 940111 608807 940113
rect 606905 940057 606961 940111
rect 607047 940057 607103 940111
rect 607189 940057 607245 940111
rect 607331 940057 607387 940111
rect 607473 940057 607529 940111
rect 607615 940057 607671 940111
rect 607757 940057 607813 940111
rect 607899 940057 607955 940111
rect 608041 940057 608097 940111
rect 608183 940057 608239 940111
rect 608325 940057 608381 940111
rect 608467 940057 608523 940111
rect 608609 940057 608665 940111
rect 608751 940057 608807 940111
rect 606905 939919 606961 939971
rect 607047 939919 607103 939971
rect 607189 939919 607245 939971
rect 607331 939919 607387 939971
rect 607473 939919 607529 939971
rect 607615 939919 607671 939971
rect 607757 939919 607813 939971
rect 607899 939919 607955 939971
rect 608041 939919 608097 939971
rect 608183 939919 608239 939971
rect 608325 939919 608381 939971
rect 608467 939919 608523 939971
rect 608609 939919 608665 939971
rect 608751 939919 608807 939971
rect 606905 939915 606908 939919
rect 606908 939915 606961 939919
rect 607047 939915 607088 939919
rect 607088 939915 607103 939919
rect 607189 939915 607212 939919
rect 607212 939915 607245 939919
rect 607331 939915 607336 939919
rect 607336 939915 607387 939919
rect 607473 939915 607528 939919
rect 607528 939915 607529 939919
rect 607615 939915 607652 939919
rect 607652 939915 607671 939919
rect 607757 939915 607776 939919
rect 607776 939915 607813 939919
rect 607899 939915 607900 939919
rect 607900 939915 607955 939919
rect 608041 939915 608080 939919
rect 608080 939915 608097 939919
rect 608183 939915 608204 939919
rect 608204 939915 608239 939919
rect 608325 939915 608328 939919
rect 608328 939915 608381 939919
rect 608467 939915 608520 939919
rect 608520 939915 608523 939919
rect 608609 939915 608644 939919
rect 608644 939915 608665 939919
rect 608751 939915 608768 939919
rect 608768 939915 608807 939919
rect 606905 939773 606961 939829
rect 607047 939773 607103 939829
rect 607189 939773 607245 939829
rect 607331 939773 607387 939829
rect 607473 939773 607529 939829
rect 607615 939773 607671 939829
rect 607757 939773 607813 939829
rect 607899 939773 607955 939829
rect 608041 939773 608097 939829
rect 608183 939773 608239 939829
rect 608325 939773 608381 939829
rect 608467 939773 608523 939829
rect 608609 939773 608665 939829
rect 608751 939773 608807 939829
rect 609275 941655 609331 941675
rect 609417 941655 609473 941675
rect 609559 941655 609615 941675
rect 609701 941655 609757 941675
rect 609843 941655 609899 941675
rect 609985 941655 610041 941675
rect 610127 941655 610183 941675
rect 610269 941655 610325 941675
rect 610411 941655 610467 941675
rect 610553 941655 610609 941675
rect 610695 941655 610751 941675
rect 610837 941655 610893 941675
rect 610979 941655 611035 941675
rect 611121 941655 611177 941675
rect 609275 941619 609278 941655
rect 609278 941619 609331 941655
rect 609417 941619 609458 941655
rect 609458 941619 609473 941655
rect 609559 941619 609582 941655
rect 609582 941619 609615 941655
rect 609701 941619 609706 941655
rect 609706 941619 609757 941655
rect 609843 941619 609898 941655
rect 609898 941619 609899 941655
rect 609985 941619 610022 941655
rect 610022 941619 610041 941655
rect 610127 941619 610146 941655
rect 610146 941619 610183 941655
rect 610269 941619 610270 941655
rect 610270 941619 610325 941655
rect 610411 941619 610450 941655
rect 610450 941619 610467 941655
rect 610553 941619 610574 941655
rect 610574 941619 610609 941655
rect 610695 941619 610698 941655
rect 610698 941619 610751 941655
rect 610837 941619 610890 941655
rect 610890 941619 610893 941655
rect 610979 941619 611014 941655
rect 611014 941619 611035 941655
rect 611121 941619 611138 941655
rect 611138 941619 611177 941655
rect 609275 941531 609331 941533
rect 609417 941531 609473 941533
rect 609559 941531 609615 941533
rect 609701 941531 609757 941533
rect 609843 941531 609899 941533
rect 609985 941531 610041 941533
rect 610127 941531 610183 941533
rect 610269 941531 610325 941533
rect 610411 941531 610467 941533
rect 610553 941531 610609 941533
rect 610695 941531 610751 941533
rect 610837 941531 610893 941533
rect 610979 941531 611035 941533
rect 611121 941531 611177 941533
rect 609275 941477 609278 941531
rect 609278 941477 609331 941531
rect 609417 941477 609458 941531
rect 609458 941477 609473 941531
rect 609559 941477 609582 941531
rect 609582 941477 609615 941531
rect 609701 941477 609706 941531
rect 609706 941477 609757 941531
rect 609843 941477 609898 941531
rect 609898 941477 609899 941531
rect 609985 941477 610022 941531
rect 610022 941477 610041 941531
rect 610127 941477 610146 941531
rect 610146 941477 610183 941531
rect 610269 941477 610270 941531
rect 610270 941477 610325 941531
rect 610411 941477 610450 941531
rect 610450 941477 610467 941531
rect 610553 941477 610574 941531
rect 610574 941477 610609 941531
rect 610695 941477 610698 941531
rect 610698 941477 610751 941531
rect 610837 941477 610890 941531
rect 610890 941477 610893 941531
rect 610979 941477 611014 941531
rect 611014 941477 611035 941531
rect 611121 941477 611138 941531
rect 611138 941477 611177 941531
rect 609275 941351 609278 941391
rect 609278 941351 609331 941391
rect 609417 941351 609458 941391
rect 609458 941351 609473 941391
rect 609559 941351 609582 941391
rect 609582 941351 609615 941391
rect 609701 941351 609706 941391
rect 609706 941351 609757 941391
rect 609843 941351 609898 941391
rect 609898 941351 609899 941391
rect 609985 941351 610022 941391
rect 610022 941351 610041 941391
rect 610127 941351 610146 941391
rect 610146 941351 610183 941391
rect 610269 941351 610270 941391
rect 610270 941351 610325 941391
rect 610411 941351 610450 941391
rect 610450 941351 610467 941391
rect 610553 941351 610574 941391
rect 610574 941351 610609 941391
rect 610695 941351 610698 941391
rect 610698 941351 610751 941391
rect 610837 941351 610890 941391
rect 610890 941351 610893 941391
rect 610979 941351 611014 941391
rect 611014 941351 611035 941391
rect 611121 941351 611138 941391
rect 611138 941351 611177 941391
rect 609275 941335 609331 941351
rect 609417 941335 609473 941351
rect 609559 941335 609615 941351
rect 609701 941335 609757 941351
rect 609843 941335 609899 941351
rect 609985 941335 610041 941351
rect 610127 941335 610183 941351
rect 610269 941335 610325 941351
rect 610411 941335 610467 941351
rect 610553 941335 610609 941351
rect 610695 941335 610751 941351
rect 610837 941335 610893 941351
rect 610979 941335 611035 941351
rect 611121 941335 611177 941351
rect 609275 941227 609278 941249
rect 609278 941227 609331 941249
rect 609417 941227 609458 941249
rect 609458 941227 609473 941249
rect 609559 941227 609582 941249
rect 609582 941227 609615 941249
rect 609701 941227 609706 941249
rect 609706 941227 609757 941249
rect 609843 941227 609898 941249
rect 609898 941227 609899 941249
rect 609985 941227 610022 941249
rect 610022 941227 610041 941249
rect 610127 941227 610146 941249
rect 610146 941227 610183 941249
rect 610269 941227 610270 941249
rect 610270 941227 610325 941249
rect 610411 941227 610450 941249
rect 610450 941227 610467 941249
rect 610553 941227 610574 941249
rect 610574 941227 610609 941249
rect 610695 941227 610698 941249
rect 610698 941227 610751 941249
rect 610837 941227 610890 941249
rect 610890 941227 610893 941249
rect 610979 941227 611014 941249
rect 611014 941227 611035 941249
rect 611121 941227 611138 941249
rect 611138 941227 611177 941249
rect 609275 941193 609331 941227
rect 609417 941193 609473 941227
rect 609559 941193 609615 941227
rect 609701 941193 609757 941227
rect 609843 941193 609899 941227
rect 609985 941193 610041 941227
rect 610127 941193 610183 941227
rect 610269 941193 610325 941227
rect 610411 941193 610467 941227
rect 610553 941193 610609 941227
rect 610695 941193 610751 941227
rect 610837 941193 610893 941227
rect 610979 941193 611035 941227
rect 611121 941193 611177 941227
rect 609275 941103 609278 941107
rect 609278 941103 609331 941107
rect 609417 941103 609458 941107
rect 609458 941103 609473 941107
rect 609559 941103 609582 941107
rect 609582 941103 609615 941107
rect 609701 941103 609706 941107
rect 609706 941103 609757 941107
rect 609843 941103 609898 941107
rect 609898 941103 609899 941107
rect 609985 941103 610022 941107
rect 610022 941103 610041 941107
rect 610127 941103 610146 941107
rect 610146 941103 610183 941107
rect 610269 941103 610270 941107
rect 610270 941103 610325 941107
rect 610411 941103 610450 941107
rect 610450 941103 610467 941107
rect 610553 941103 610574 941107
rect 610574 941103 610609 941107
rect 610695 941103 610698 941107
rect 610698 941103 610751 941107
rect 610837 941103 610890 941107
rect 610890 941103 610893 941107
rect 610979 941103 611014 941107
rect 611014 941103 611035 941107
rect 611121 941103 611138 941107
rect 611138 941103 611177 941107
rect 609275 941051 609331 941103
rect 609417 941051 609473 941103
rect 609559 941051 609615 941103
rect 609701 941051 609757 941103
rect 609843 941051 609899 941103
rect 609985 941051 610041 941103
rect 610127 941051 610183 941103
rect 610269 941051 610325 941103
rect 610411 941051 610467 941103
rect 610553 941051 610609 941103
rect 610695 941051 610751 941103
rect 610837 941051 610893 941103
rect 610979 941051 611035 941103
rect 611121 941051 611177 941103
rect 609275 940911 609331 940965
rect 609417 940911 609473 940965
rect 609559 940911 609615 940965
rect 609701 940911 609757 940965
rect 609843 940911 609899 940965
rect 609985 940911 610041 940965
rect 610127 940911 610183 940965
rect 610269 940911 610325 940965
rect 610411 940911 610467 940965
rect 610553 940911 610609 940965
rect 610695 940911 610751 940965
rect 610837 940911 610893 940965
rect 610979 940911 611035 940965
rect 611121 940911 611177 940965
rect 609275 940909 609278 940911
rect 609278 940909 609331 940911
rect 609417 940909 609458 940911
rect 609458 940909 609473 940911
rect 609559 940909 609582 940911
rect 609582 940909 609615 940911
rect 609701 940909 609706 940911
rect 609706 940909 609757 940911
rect 609843 940909 609898 940911
rect 609898 940909 609899 940911
rect 609985 940909 610022 940911
rect 610022 940909 610041 940911
rect 610127 940909 610146 940911
rect 610146 940909 610183 940911
rect 610269 940909 610270 940911
rect 610270 940909 610325 940911
rect 610411 940909 610450 940911
rect 610450 940909 610467 940911
rect 610553 940909 610574 940911
rect 610574 940909 610609 940911
rect 610695 940909 610698 940911
rect 610698 940909 610751 940911
rect 610837 940909 610890 940911
rect 610890 940909 610893 940911
rect 610979 940909 611014 940911
rect 611014 940909 611035 940911
rect 611121 940909 611138 940911
rect 611138 940909 611177 940911
rect 609275 940787 609331 940823
rect 609417 940787 609473 940823
rect 609559 940787 609615 940823
rect 609701 940787 609757 940823
rect 609843 940787 609899 940823
rect 609985 940787 610041 940823
rect 610127 940787 610183 940823
rect 610269 940787 610325 940823
rect 610411 940787 610467 940823
rect 610553 940787 610609 940823
rect 610695 940787 610751 940823
rect 610837 940787 610893 940823
rect 610979 940787 611035 940823
rect 611121 940787 611177 940823
rect 609275 940767 609278 940787
rect 609278 940767 609331 940787
rect 609417 940767 609458 940787
rect 609458 940767 609473 940787
rect 609559 940767 609582 940787
rect 609582 940767 609615 940787
rect 609701 940767 609706 940787
rect 609706 940767 609757 940787
rect 609843 940767 609898 940787
rect 609898 940767 609899 940787
rect 609985 940767 610022 940787
rect 610022 940767 610041 940787
rect 610127 940767 610146 940787
rect 610146 940767 610183 940787
rect 610269 940767 610270 940787
rect 610270 940767 610325 940787
rect 610411 940767 610450 940787
rect 610450 940767 610467 940787
rect 610553 940767 610574 940787
rect 610574 940767 610609 940787
rect 610695 940767 610698 940787
rect 610698 940767 610751 940787
rect 610837 940767 610890 940787
rect 610890 940767 610893 940787
rect 610979 940767 611014 940787
rect 611014 940767 611035 940787
rect 611121 940767 611138 940787
rect 611138 940767 611177 940787
rect 609275 940663 609331 940681
rect 609417 940663 609473 940681
rect 609559 940663 609615 940681
rect 609701 940663 609757 940681
rect 609843 940663 609899 940681
rect 609985 940663 610041 940681
rect 610127 940663 610183 940681
rect 610269 940663 610325 940681
rect 610411 940663 610467 940681
rect 610553 940663 610609 940681
rect 610695 940663 610751 940681
rect 610837 940663 610893 940681
rect 610979 940663 611035 940681
rect 611121 940663 611177 940681
rect 609275 940625 609278 940663
rect 609278 940625 609331 940663
rect 609417 940625 609458 940663
rect 609458 940625 609473 940663
rect 609559 940625 609582 940663
rect 609582 940625 609615 940663
rect 609701 940625 609706 940663
rect 609706 940625 609757 940663
rect 609843 940625 609898 940663
rect 609898 940625 609899 940663
rect 609985 940625 610022 940663
rect 610022 940625 610041 940663
rect 610127 940625 610146 940663
rect 610146 940625 610183 940663
rect 610269 940625 610270 940663
rect 610270 940625 610325 940663
rect 610411 940625 610450 940663
rect 610450 940625 610467 940663
rect 610553 940625 610574 940663
rect 610574 940625 610609 940663
rect 610695 940625 610698 940663
rect 610698 940625 610751 940663
rect 610837 940625 610890 940663
rect 610890 940625 610893 940663
rect 610979 940625 611014 940663
rect 611014 940625 611035 940663
rect 611121 940625 611138 940663
rect 611138 940625 611177 940663
rect 609275 940483 609278 940539
rect 609278 940483 609331 940539
rect 609417 940483 609458 940539
rect 609458 940483 609473 940539
rect 609559 940483 609582 940539
rect 609582 940483 609615 940539
rect 609701 940483 609706 940539
rect 609706 940483 609757 940539
rect 609843 940483 609898 940539
rect 609898 940483 609899 940539
rect 609985 940483 610022 940539
rect 610022 940483 610041 940539
rect 610127 940483 610146 940539
rect 610146 940483 610183 940539
rect 610269 940483 610270 940539
rect 610270 940483 610325 940539
rect 610411 940483 610450 940539
rect 610450 940483 610467 940539
rect 610553 940483 610574 940539
rect 610574 940483 610609 940539
rect 610695 940483 610698 940539
rect 610698 940483 610751 940539
rect 610837 940483 610890 940539
rect 610890 940483 610893 940539
rect 610979 940483 611014 940539
rect 611014 940483 611035 940539
rect 611121 940483 611138 940539
rect 611138 940483 611177 940539
rect 609275 940359 609278 940397
rect 609278 940359 609331 940397
rect 609417 940359 609458 940397
rect 609458 940359 609473 940397
rect 609559 940359 609582 940397
rect 609582 940359 609615 940397
rect 609701 940359 609706 940397
rect 609706 940359 609757 940397
rect 609843 940359 609898 940397
rect 609898 940359 609899 940397
rect 609985 940359 610022 940397
rect 610022 940359 610041 940397
rect 610127 940359 610146 940397
rect 610146 940359 610183 940397
rect 610269 940359 610270 940397
rect 610270 940359 610325 940397
rect 610411 940359 610450 940397
rect 610450 940359 610467 940397
rect 610553 940359 610574 940397
rect 610574 940359 610609 940397
rect 610695 940359 610698 940397
rect 610698 940359 610751 940397
rect 610837 940359 610890 940397
rect 610890 940359 610893 940397
rect 610979 940359 611014 940397
rect 611014 940359 611035 940397
rect 611121 940359 611138 940397
rect 611138 940359 611177 940397
rect 609275 940341 609331 940359
rect 609417 940341 609473 940359
rect 609559 940341 609615 940359
rect 609701 940341 609757 940359
rect 609843 940341 609899 940359
rect 609985 940341 610041 940359
rect 610127 940341 610183 940359
rect 610269 940341 610325 940359
rect 610411 940341 610467 940359
rect 610553 940341 610609 940359
rect 610695 940341 610751 940359
rect 610837 940341 610893 940359
rect 610979 940341 611035 940359
rect 611121 940341 611177 940359
rect 609275 940235 609278 940255
rect 609278 940235 609331 940255
rect 609417 940235 609458 940255
rect 609458 940235 609473 940255
rect 609559 940235 609582 940255
rect 609582 940235 609615 940255
rect 609701 940235 609706 940255
rect 609706 940235 609757 940255
rect 609843 940235 609898 940255
rect 609898 940235 609899 940255
rect 609985 940235 610022 940255
rect 610022 940235 610041 940255
rect 610127 940235 610146 940255
rect 610146 940235 610183 940255
rect 610269 940235 610270 940255
rect 610270 940235 610325 940255
rect 610411 940235 610450 940255
rect 610450 940235 610467 940255
rect 610553 940235 610574 940255
rect 610574 940235 610609 940255
rect 610695 940235 610698 940255
rect 610698 940235 610751 940255
rect 610837 940235 610890 940255
rect 610890 940235 610893 940255
rect 610979 940235 611014 940255
rect 611014 940235 611035 940255
rect 611121 940235 611138 940255
rect 611138 940235 611177 940255
rect 609275 940199 609331 940235
rect 609417 940199 609473 940235
rect 609559 940199 609615 940235
rect 609701 940199 609757 940235
rect 609843 940199 609899 940235
rect 609985 940199 610041 940235
rect 610127 940199 610183 940235
rect 610269 940199 610325 940235
rect 610411 940199 610467 940235
rect 610553 940199 610609 940235
rect 610695 940199 610751 940235
rect 610837 940199 610893 940235
rect 610979 940199 611035 940235
rect 611121 940199 611177 940235
rect 609275 940111 609278 940113
rect 609278 940111 609331 940113
rect 609417 940111 609458 940113
rect 609458 940111 609473 940113
rect 609559 940111 609582 940113
rect 609582 940111 609615 940113
rect 609701 940111 609706 940113
rect 609706 940111 609757 940113
rect 609843 940111 609898 940113
rect 609898 940111 609899 940113
rect 609985 940111 610022 940113
rect 610022 940111 610041 940113
rect 610127 940111 610146 940113
rect 610146 940111 610183 940113
rect 610269 940111 610270 940113
rect 610270 940111 610325 940113
rect 610411 940111 610450 940113
rect 610450 940111 610467 940113
rect 610553 940111 610574 940113
rect 610574 940111 610609 940113
rect 610695 940111 610698 940113
rect 610698 940111 610751 940113
rect 610837 940111 610890 940113
rect 610890 940111 610893 940113
rect 610979 940111 611014 940113
rect 611014 940111 611035 940113
rect 611121 940111 611138 940113
rect 611138 940111 611177 940113
rect 609275 940057 609331 940111
rect 609417 940057 609473 940111
rect 609559 940057 609615 940111
rect 609701 940057 609757 940111
rect 609843 940057 609899 940111
rect 609985 940057 610041 940111
rect 610127 940057 610183 940111
rect 610269 940057 610325 940111
rect 610411 940057 610467 940111
rect 610553 940057 610609 940111
rect 610695 940057 610751 940111
rect 610837 940057 610893 940111
rect 610979 940057 611035 940111
rect 611121 940057 611177 940111
rect 609275 939919 609331 939971
rect 609417 939919 609473 939971
rect 609559 939919 609615 939971
rect 609701 939919 609757 939971
rect 609843 939919 609899 939971
rect 609985 939919 610041 939971
rect 610127 939919 610183 939971
rect 610269 939919 610325 939971
rect 610411 939919 610467 939971
rect 610553 939919 610609 939971
rect 610695 939919 610751 939971
rect 610837 939919 610893 939971
rect 610979 939919 611035 939971
rect 611121 939919 611177 939971
rect 609275 939915 609278 939919
rect 609278 939915 609331 939919
rect 609417 939915 609458 939919
rect 609458 939915 609473 939919
rect 609559 939915 609582 939919
rect 609582 939915 609615 939919
rect 609701 939915 609706 939919
rect 609706 939915 609757 939919
rect 609843 939915 609898 939919
rect 609898 939915 609899 939919
rect 609985 939915 610022 939919
rect 610022 939915 610041 939919
rect 610127 939915 610146 939919
rect 610146 939915 610183 939919
rect 610269 939915 610270 939919
rect 610270 939915 610325 939919
rect 610411 939915 610450 939919
rect 610450 939915 610467 939919
rect 610553 939915 610574 939919
rect 610574 939915 610609 939919
rect 610695 939915 610698 939919
rect 610698 939915 610751 939919
rect 610837 939915 610890 939919
rect 610890 939915 610893 939919
rect 610979 939915 611014 939919
rect 611014 939915 611035 939919
rect 611121 939915 611138 939919
rect 611138 939915 611177 939919
rect 609275 939773 609331 939829
rect 609417 939773 609473 939829
rect 609559 939773 609615 939829
rect 609701 939773 609757 939829
rect 609843 939773 609899 939829
rect 609985 939773 610041 939829
rect 610127 939773 610183 939829
rect 610269 939773 610325 939829
rect 610411 939773 610467 939829
rect 610553 939773 610609 939829
rect 610695 939773 610751 939829
rect 610837 939773 610893 939829
rect 610979 939773 611035 939829
rect 611121 939773 611177 939829
rect 611897 941655 611953 941675
rect 612039 941655 612095 941675
rect 612181 941655 612237 941675
rect 612323 941655 612379 941675
rect 612465 941655 612521 941675
rect 612607 941655 612663 941675
rect 612749 941655 612805 941675
rect 612891 941655 612947 941675
rect 613033 941655 613089 941675
rect 613175 941655 613231 941675
rect 613317 941655 613373 941675
rect 613459 941655 613515 941675
rect 613601 941655 613657 941675
rect 611897 941619 611938 941655
rect 611938 941619 611953 941655
rect 612039 941619 612062 941655
rect 612062 941619 612095 941655
rect 612181 941619 612186 941655
rect 612186 941619 612237 941655
rect 612323 941619 612378 941655
rect 612378 941619 612379 941655
rect 612465 941619 612502 941655
rect 612502 941619 612521 941655
rect 612607 941619 612626 941655
rect 612626 941619 612663 941655
rect 612749 941619 612750 941655
rect 612750 941619 612805 941655
rect 612891 941619 612930 941655
rect 612930 941619 612947 941655
rect 613033 941619 613054 941655
rect 613054 941619 613089 941655
rect 613175 941619 613178 941655
rect 613178 941619 613231 941655
rect 613317 941619 613370 941655
rect 613370 941619 613373 941655
rect 613459 941619 613494 941655
rect 613494 941619 613515 941655
rect 613601 941619 613618 941655
rect 613618 941619 613657 941655
rect 611897 941531 611953 941533
rect 612039 941531 612095 941533
rect 612181 941531 612237 941533
rect 612323 941531 612379 941533
rect 612465 941531 612521 941533
rect 612607 941531 612663 941533
rect 612749 941531 612805 941533
rect 612891 941531 612947 941533
rect 613033 941531 613089 941533
rect 613175 941531 613231 941533
rect 613317 941531 613373 941533
rect 613459 941531 613515 941533
rect 613601 941531 613657 941533
rect 611897 941477 611938 941531
rect 611938 941477 611953 941531
rect 612039 941477 612062 941531
rect 612062 941477 612095 941531
rect 612181 941477 612186 941531
rect 612186 941477 612237 941531
rect 612323 941477 612378 941531
rect 612378 941477 612379 941531
rect 612465 941477 612502 941531
rect 612502 941477 612521 941531
rect 612607 941477 612626 941531
rect 612626 941477 612663 941531
rect 612749 941477 612750 941531
rect 612750 941477 612805 941531
rect 612891 941477 612930 941531
rect 612930 941477 612947 941531
rect 613033 941477 613054 941531
rect 613054 941477 613089 941531
rect 613175 941477 613178 941531
rect 613178 941477 613231 941531
rect 613317 941477 613370 941531
rect 613370 941477 613373 941531
rect 613459 941477 613494 941531
rect 613494 941477 613515 941531
rect 613601 941477 613618 941531
rect 613618 941477 613657 941531
rect 611897 941351 611938 941391
rect 611938 941351 611953 941391
rect 612039 941351 612062 941391
rect 612062 941351 612095 941391
rect 612181 941351 612186 941391
rect 612186 941351 612237 941391
rect 612323 941351 612378 941391
rect 612378 941351 612379 941391
rect 612465 941351 612502 941391
rect 612502 941351 612521 941391
rect 612607 941351 612626 941391
rect 612626 941351 612663 941391
rect 612749 941351 612750 941391
rect 612750 941351 612805 941391
rect 612891 941351 612930 941391
rect 612930 941351 612947 941391
rect 613033 941351 613054 941391
rect 613054 941351 613089 941391
rect 613175 941351 613178 941391
rect 613178 941351 613231 941391
rect 613317 941351 613370 941391
rect 613370 941351 613373 941391
rect 613459 941351 613494 941391
rect 613494 941351 613515 941391
rect 613601 941351 613618 941391
rect 613618 941351 613657 941391
rect 611897 941335 611953 941351
rect 612039 941335 612095 941351
rect 612181 941335 612237 941351
rect 612323 941335 612379 941351
rect 612465 941335 612521 941351
rect 612607 941335 612663 941351
rect 612749 941335 612805 941351
rect 612891 941335 612947 941351
rect 613033 941335 613089 941351
rect 613175 941335 613231 941351
rect 613317 941335 613373 941351
rect 613459 941335 613515 941351
rect 613601 941335 613657 941351
rect 611897 941227 611938 941249
rect 611938 941227 611953 941249
rect 612039 941227 612062 941249
rect 612062 941227 612095 941249
rect 612181 941227 612186 941249
rect 612186 941227 612237 941249
rect 612323 941227 612378 941249
rect 612378 941227 612379 941249
rect 612465 941227 612502 941249
rect 612502 941227 612521 941249
rect 612607 941227 612626 941249
rect 612626 941227 612663 941249
rect 612749 941227 612750 941249
rect 612750 941227 612805 941249
rect 612891 941227 612930 941249
rect 612930 941227 612947 941249
rect 613033 941227 613054 941249
rect 613054 941227 613089 941249
rect 613175 941227 613178 941249
rect 613178 941227 613231 941249
rect 613317 941227 613370 941249
rect 613370 941227 613373 941249
rect 613459 941227 613494 941249
rect 613494 941227 613515 941249
rect 613601 941227 613618 941249
rect 613618 941227 613657 941249
rect 611897 941193 611953 941227
rect 612039 941193 612095 941227
rect 612181 941193 612237 941227
rect 612323 941193 612379 941227
rect 612465 941193 612521 941227
rect 612607 941193 612663 941227
rect 612749 941193 612805 941227
rect 612891 941193 612947 941227
rect 613033 941193 613089 941227
rect 613175 941193 613231 941227
rect 613317 941193 613373 941227
rect 613459 941193 613515 941227
rect 613601 941193 613657 941227
rect 611897 941103 611938 941107
rect 611938 941103 611953 941107
rect 612039 941103 612062 941107
rect 612062 941103 612095 941107
rect 612181 941103 612186 941107
rect 612186 941103 612237 941107
rect 612323 941103 612378 941107
rect 612378 941103 612379 941107
rect 612465 941103 612502 941107
rect 612502 941103 612521 941107
rect 612607 941103 612626 941107
rect 612626 941103 612663 941107
rect 612749 941103 612750 941107
rect 612750 941103 612805 941107
rect 612891 941103 612930 941107
rect 612930 941103 612947 941107
rect 613033 941103 613054 941107
rect 613054 941103 613089 941107
rect 613175 941103 613178 941107
rect 613178 941103 613231 941107
rect 613317 941103 613370 941107
rect 613370 941103 613373 941107
rect 613459 941103 613494 941107
rect 613494 941103 613515 941107
rect 613601 941103 613618 941107
rect 613618 941103 613657 941107
rect 611897 941051 611953 941103
rect 612039 941051 612095 941103
rect 612181 941051 612237 941103
rect 612323 941051 612379 941103
rect 612465 941051 612521 941103
rect 612607 941051 612663 941103
rect 612749 941051 612805 941103
rect 612891 941051 612947 941103
rect 613033 941051 613089 941103
rect 613175 941051 613231 941103
rect 613317 941051 613373 941103
rect 613459 941051 613515 941103
rect 613601 941051 613657 941103
rect 611897 940911 611953 940965
rect 612039 940911 612095 940965
rect 612181 940911 612237 940965
rect 612323 940911 612379 940965
rect 612465 940911 612521 940965
rect 612607 940911 612663 940965
rect 612749 940911 612805 940965
rect 612891 940911 612947 940965
rect 613033 940911 613089 940965
rect 613175 940911 613231 940965
rect 613317 940911 613373 940965
rect 613459 940911 613515 940965
rect 613601 940911 613657 940965
rect 611897 940909 611938 940911
rect 611938 940909 611953 940911
rect 612039 940909 612062 940911
rect 612062 940909 612095 940911
rect 612181 940909 612186 940911
rect 612186 940909 612237 940911
rect 612323 940909 612378 940911
rect 612378 940909 612379 940911
rect 612465 940909 612502 940911
rect 612502 940909 612521 940911
rect 612607 940909 612626 940911
rect 612626 940909 612663 940911
rect 612749 940909 612750 940911
rect 612750 940909 612805 940911
rect 612891 940909 612930 940911
rect 612930 940909 612947 940911
rect 613033 940909 613054 940911
rect 613054 940909 613089 940911
rect 613175 940909 613178 940911
rect 613178 940909 613231 940911
rect 613317 940909 613370 940911
rect 613370 940909 613373 940911
rect 613459 940909 613494 940911
rect 613494 940909 613515 940911
rect 613601 940909 613618 940911
rect 613618 940909 613657 940911
rect 611897 940787 611953 940823
rect 612039 940787 612095 940823
rect 612181 940787 612237 940823
rect 612323 940787 612379 940823
rect 612465 940787 612521 940823
rect 612607 940787 612663 940823
rect 612749 940787 612805 940823
rect 612891 940787 612947 940823
rect 613033 940787 613089 940823
rect 613175 940787 613231 940823
rect 613317 940787 613373 940823
rect 613459 940787 613515 940823
rect 613601 940787 613657 940823
rect 611897 940767 611938 940787
rect 611938 940767 611953 940787
rect 612039 940767 612062 940787
rect 612062 940767 612095 940787
rect 612181 940767 612186 940787
rect 612186 940767 612237 940787
rect 612323 940767 612378 940787
rect 612378 940767 612379 940787
rect 612465 940767 612502 940787
rect 612502 940767 612521 940787
rect 612607 940767 612626 940787
rect 612626 940767 612663 940787
rect 612749 940767 612750 940787
rect 612750 940767 612805 940787
rect 612891 940767 612930 940787
rect 612930 940767 612947 940787
rect 613033 940767 613054 940787
rect 613054 940767 613089 940787
rect 613175 940767 613178 940787
rect 613178 940767 613231 940787
rect 613317 940767 613370 940787
rect 613370 940767 613373 940787
rect 613459 940767 613494 940787
rect 613494 940767 613515 940787
rect 613601 940767 613618 940787
rect 613618 940767 613657 940787
rect 611897 940663 611953 940681
rect 612039 940663 612095 940681
rect 612181 940663 612237 940681
rect 612323 940663 612379 940681
rect 612465 940663 612521 940681
rect 612607 940663 612663 940681
rect 612749 940663 612805 940681
rect 612891 940663 612947 940681
rect 613033 940663 613089 940681
rect 613175 940663 613231 940681
rect 613317 940663 613373 940681
rect 613459 940663 613515 940681
rect 613601 940663 613657 940681
rect 611897 940625 611938 940663
rect 611938 940625 611953 940663
rect 612039 940625 612062 940663
rect 612062 940625 612095 940663
rect 612181 940625 612186 940663
rect 612186 940625 612237 940663
rect 612323 940625 612378 940663
rect 612378 940625 612379 940663
rect 612465 940625 612502 940663
rect 612502 940625 612521 940663
rect 612607 940625 612626 940663
rect 612626 940625 612663 940663
rect 612749 940625 612750 940663
rect 612750 940625 612805 940663
rect 612891 940625 612930 940663
rect 612930 940625 612947 940663
rect 613033 940625 613054 940663
rect 613054 940625 613089 940663
rect 613175 940625 613178 940663
rect 613178 940625 613231 940663
rect 613317 940625 613370 940663
rect 613370 940625 613373 940663
rect 613459 940625 613494 940663
rect 613494 940625 613515 940663
rect 613601 940625 613618 940663
rect 613618 940625 613657 940663
rect 611897 940483 611938 940539
rect 611938 940483 611953 940539
rect 612039 940483 612062 940539
rect 612062 940483 612095 940539
rect 612181 940483 612186 940539
rect 612186 940483 612237 940539
rect 612323 940483 612378 940539
rect 612378 940483 612379 940539
rect 612465 940483 612502 940539
rect 612502 940483 612521 940539
rect 612607 940483 612626 940539
rect 612626 940483 612663 940539
rect 612749 940483 612750 940539
rect 612750 940483 612805 940539
rect 612891 940483 612930 940539
rect 612930 940483 612947 940539
rect 613033 940483 613054 940539
rect 613054 940483 613089 940539
rect 613175 940483 613178 940539
rect 613178 940483 613231 940539
rect 613317 940483 613370 940539
rect 613370 940483 613373 940539
rect 613459 940483 613494 940539
rect 613494 940483 613515 940539
rect 613601 940483 613618 940539
rect 613618 940483 613657 940539
rect 611897 940359 611938 940397
rect 611938 940359 611953 940397
rect 612039 940359 612062 940397
rect 612062 940359 612095 940397
rect 612181 940359 612186 940397
rect 612186 940359 612237 940397
rect 612323 940359 612378 940397
rect 612378 940359 612379 940397
rect 612465 940359 612502 940397
rect 612502 940359 612521 940397
rect 612607 940359 612626 940397
rect 612626 940359 612663 940397
rect 612749 940359 612750 940397
rect 612750 940359 612805 940397
rect 612891 940359 612930 940397
rect 612930 940359 612947 940397
rect 613033 940359 613054 940397
rect 613054 940359 613089 940397
rect 613175 940359 613178 940397
rect 613178 940359 613231 940397
rect 613317 940359 613370 940397
rect 613370 940359 613373 940397
rect 613459 940359 613494 940397
rect 613494 940359 613515 940397
rect 613601 940359 613618 940397
rect 613618 940359 613657 940397
rect 611897 940341 611953 940359
rect 612039 940341 612095 940359
rect 612181 940341 612237 940359
rect 612323 940341 612379 940359
rect 612465 940341 612521 940359
rect 612607 940341 612663 940359
rect 612749 940341 612805 940359
rect 612891 940341 612947 940359
rect 613033 940341 613089 940359
rect 613175 940341 613231 940359
rect 613317 940341 613373 940359
rect 613459 940341 613515 940359
rect 613601 940341 613657 940359
rect 611897 940235 611938 940255
rect 611938 940235 611953 940255
rect 612039 940235 612062 940255
rect 612062 940235 612095 940255
rect 612181 940235 612186 940255
rect 612186 940235 612237 940255
rect 612323 940235 612378 940255
rect 612378 940235 612379 940255
rect 612465 940235 612502 940255
rect 612502 940235 612521 940255
rect 612607 940235 612626 940255
rect 612626 940235 612663 940255
rect 612749 940235 612750 940255
rect 612750 940235 612805 940255
rect 612891 940235 612930 940255
rect 612930 940235 612947 940255
rect 613033 940235 613054 940255
rect 613054 940235 613089 940255
rect 613175 940235 613178 940255
rect 613178 940235 613231 940255
rect 613317 940235 613370 940255
rect 613370 940235 613373 940255
rect 613459 940235 613494 940255
rect 613494 940235 613515 940255
rect 613601 940235 613618 940255
rect 613618 940235 613657 940255
rect 611897 940199 611953 940235
rect 612039 940199 612095 940235
rect 612181 940199 612237 940235
rect 612323 940199 612379 940235
rect 612465 940199 612521 940235
rect 612607 940199 612663 940235
rect 612749 940199 612805 940235
rect 612891 940199 612947 940235
rect 613033 940199 613089 940235
rect 613175 940199 613231 940235
rect 613317 940199 613373 940235
rect 613459 940199 613515 940235
rect 613601 940199 613657 940235
rect 611897 940111 611938 940113
rect 611938 940111 611953 940113
rect 612039 940111 612062 940113
rect 612062 940111 612095 940113
rect 612181 940111 612186 940113
rect 612186 940111 612237 940113
rect 612323 940111 612378 940113
rect 612378 940111 612379 940113
rect 612465 940111 612502 940113
rect 612502 940111 612521 940113
rect 612607 940111 612626 940113
rect 612626 940111 612663 940113
rect 612749 940111 612750 940113
rect 612750 940111 612805 940113
rect 612891 940111 612930 940113
rect 612930 940111 612947 940113
rect 613033 940111 613054 940113
rect 613054 940111 613089 940113
rect 613175 940111 613178 940113
rect 613178 940111 613231 940113
rect 613317 940111 613370 940113
rect 613370 940111 613373 940113
rect 613459 940111 613494 940113
rect 613494 940111 613515 940113
rect 613601 940111 613618 940113
rect 613618 940111 613657 940113
rect 611897 940057 611953 940111
rect 612039 940057 612095 940111
rect 612181 940057 612237 940111
rect 612323 940057 612379 940111
rect 612465 940057 612521 940111
rect 612607 940057 612663 940111
rect 612749 940057 612805 940111
rect 612891 940057 612947 940111
rect 613033 940057 613089 940111
rect 613175 940057 613231 940111
rect 613317 940057 613373 940111
rect 613459 940057 613515 940111
rect 613601 940057 613657 940111
rect 611897 939919 611953 939971
rect 612039 939919 612095 939971
rect 612181 939919 612237 939971
rect 612323 939919 612379 939971
rect 612465 939919 612521 939971
rect 612607 939919 612663 939971
rect 612749 939919 612805 939971
rect 612891 939919 612947 939971
rect 613033 939919 613089 939971
rect 613175 939919 613231 939971
rect 613317 939919 613373 939971
rect 613459 939919 613515 939971
rect 613601 939919 613657 939971
rect 611897 939915 611938 939919
rect 611938 939915 611953 939919
rect 612039 939915 612062 939919
rect 612062 939915 612095 939919
rect 612181 939915 612186 939919
rect 612186 939915 612237 939919
rect 612323 939915 612378 939919
rect 612378 939915 612379 939919
rect 612465 939915 612502 939919
rect 612502 939915 612521 939919
rect 612607 939915 612626 939919
rect 612626 939915 612663 939919
rect 612749 939915 612750 939919
rect 612750 939915 612805 939919
rect 612891 939915 612930 939919
rect 612930 939915 612947 939919
rect 613033 939915 613054 939919
rect 613054 939915 613089 939919
rect 613175 939915 613178 939919
rect 613178 939915 613231 939919
rect 613317 939915 613370 939919
rect 613370 939915 613373 939919
rect 613459 939915 613494 939919
rect 613494 939915 613515 939919
rect 613601 939915 613618 939919
rect 613618 939915 613657 939919
rect 611897 939773 611953 939829
rect 612039 939773 612095 939829
rect 612181 939773 612237 939829
rect 612323 939773 612379 939829
rect 612465 939773 612521 939829
rect 612607 939773 612663 939829
rect 612749 939773 612805 939829
rect 612891 939773 612947 939829
rect 613033 939773 613089 939829
rect 613175 939773 613231 939829
rect 613317 939773 613373 939829
rect 613459 939773 613515 939829
rect 613601 939773 613657 939829
rect 73866 878594 73922 878650
rect 74008 878594 74064 878650
rect 74150 878594 74206 878650
rect 74292 878594 74348 878650
rect 74434 878594 74490 878650
rect 74576 878594 74632 878650
rect 74718 878594 74774 878650
rect 74860 878594 74916 878650
rect 75002 878594 75058 878650
rect 75144 878594 75200 878650
rect 75286 878594 75342 878650
rect 75428 878594 75484 878650
rect 75570 878594 75626 878650
rect 75712 878594 75768 878650
rect 73866 878452 73922 878508
rect 74008 878452 74064 878508
rect 74150 878452 74206 878508
rect 74292 878452 74348 878508
rect 74434 878452 74490 878508
rect 74576 878452 74632 878508
rect 74718 878452 74774 878508
rect 74860 878452 74916 878508
rect 75002 878452 75058 878508
rect 75144 878452 75200 878508
rect 75286 878452 75342 878508
rect 75428 878452 75484 878508
rect 75570 878452 75626 878508
rect 75712 878452 75768 878508
rect 73866 878310 73922 878366
rect 74008 878310 74064 878366
rect 74150 878310 74206 878366
rect 74292 878310 74348 878366
rect 74434 878310 74490 878366
rect 74576 878310 74632 878366
rect 74718 878310 74774 878366
rect 74860 878310 74916 878366
rect 75002 878310 75058 878366
rect 75144 878310 75200 878366
rect 75286 878310 75342 878366
rect 75428 878310 75484 878366
rect 75570 878310 75626 878366
rect 75712 878310 75768 878366
rect 73866 878168 73922 878224
rect 74008 878168 74064 878224
rect 74150 878168 74206 878224
rect 74292 878168 74348 878224
rect 74434 878168 74490 878224
rect 74576 878168 74632 878224
rect 74718 878168 74774 878224
rect 74860 878168 74916 878224
rect 75002 878168 75058 878224
rect 75144 878168 75200 878224
rect 75286 878168 75342 878224
rect 75428 878168 75484 878224
rect 75570 878168 75626 878224
rect 75712 878168 75768 878224
rect 73866 878026 73922 878082
rect 74008 878026 74064 878082
rect 74150 878026 74206 878082
rect 74292 878026 74348 878082
rect 74434 878026 74490 878082
rect 74576 878026 74632 878082
rect 74718 878026 74774 878082
rect 74860 878026 74916 878082
rect 75002 878026 75058 878082
rect 75144 878026 75200 878082
rect 75286 878026 75342 878082
rect 75428 878026 75484 878082
rect 75570 878026 75626 878082
rect 75712 878026 75768 878082
rect 73866 877884 73922 877940
rect 74008 877884 74064 877940
rect 74150 877884 74206 877940
rect 74292 877884 74348 877940
rect 74434 877884 74490 877940
rect 74576 877884 74632 877940
rect 74718 877884 74774 877940
rect 74860 877884 74916 877940
rect 75002 877884 75058 877940
rect 75144 877884 75200 877940
rect 75286 877884 75342 877940
rect 75428 877884 75484 877940
rect 75570 877884 75626 877940
rect 75712 877884 75768 877940
rect 73866 877742 73922 877798
rect 74008 877742 74064 877798
rect 74150 877742 74206 877798
rect 74292 877742 74348 877798
rect 74434 877742 74490 877798
rect 74576 877742 74632 877798
rect 74718 877742 74774 877798
rect 74860 877742 74916 877798
rect 75002 877742 75058 877798
rect 75144 877742 75200 877798
rect 75286 877742 75342 877798
rect 75428 877742 75484 877798
rect 75570 877742 75626 877798
rect 75712 877742 75768 877798
rect 73866 877600 73922 877656
rect 74008 877600 74064 877656
rect 74150 877600 74206 877656
rect 74292 877600 74348 877656
rect 74434 877600 74490 877656
rect 74576 877600 74632 877656
rect 74718 877600 74774 877656
rect 74860 877600 74916 877656
rect 75002 877600 75058 877656
rect 75144 877600 75200 877656
rect 75286 877600 75342 877656
rect 75428 877600 75484 877656
rect 75570 877600 75626 877656
rect 75712 877600 75768 877656
rect 73866 877458 73922 877514
rect 74008 877458 74064 877514
rect 74150 877458 74206 877514
rect 74292 877458 74348 877514
rect 74434 877458 74490 877514
rect 74576 877458 74632 877514
rect 74718 877458 74774 877514
rect 74860 877458 74916 877514
rect 75002 877458 75058 877514
rect 75144 877458 75200 877514
rect 75286 877458 75342 877514
rect 75428 877458 75484 877514
rect 75570 877458 75626 877514
rect 75712 877458 75768 877514
rect 73866 877316 73922 877372
rect 74008 877316 74064 877372
rect 74150 877316 74206 877372
rect 74292 877316 74348 877372
rect 74434 877316 74490 877372
rect 74576 877316 74632 877372
rect 74718 877316 74774 877372
rect 74860 877316 74916 877372
rect 75002 877316 75058 877372
rect 75144 877316 75200 877372
rect 75286 877316 75342 877372
rect 75428 877316 75484 877372
rect 75570 877316 75626 877372
rect 75712 877316 75768 877372
rect 73866 877174 73922 877230
rect 74008 877174 74064 877230
rect 74150 877174 74206 877230
rect 74292 877174 74348 877230
rect 74434 877174 74490 877230
rect 74576 877174 74632 877230
rect 74718 877174 74774 877230
rect 74860 877174 74916 877230
rect 75002 877174 75058 877230
rect 75144 877174 75200 877230
rect 75286 877174 75342 877230
rect 75428 877174 75484 877230
rect 75570 877174 75626 877230
rect 75712 877174 75768 877230
rect 73866 877032 73922 877088
rect 74008 877032 74064 877088
rect 74150 877032 74206 877088
rect 74292 877032 74348 877088
rect 74434 877032 74490 877088
rect 74576 877032 74632 877088
rect 74718 877032 74774 877088
rect 74860 877032 74916 877088
rect 75002 877032 75058 877088
rect 75144 877032 75200 877088
rect 75286 877032 75342 877088
rect 75428 877032 75484 877088
rect 75570 877032 75626 877088
rect 75712 877032 75768 877088
rect 73866 876890 73922 876946
rect 74008 876890 74064 876946
rect 74150 876890 74206 876946
rect 74292 876890 74348 876946
rect 74434 876890 74490 876946
rect 74576 876890 74632 876946
rect 74718 876890 74774 876946
rect 74860 876890 74916 876946
rect 75002 876890 75058 876946
rect 75144 876890 75200 876946
rect 75286 876890 75342 876946
rect 75428 876890 75484 876946
rect 75570 876890 75626 876946
rect 75712 876890 75768 876946
rect 700040 877610 700096 877666
rect 700182 877610 700238 877666
rect 700324 877610 700380 877666
rect 700466 877610 700522 877666
rect 700608 877610 700664 877666
rect 700750 877610 700806 877666
rect 700892 877610 700948 877666
rect 701034 877610 701090 877666
rect 701176 877610 701232 877666
rect 701318 877610 701374 877666
rect 701460 877610 701516 877666
rect 701602 877610 701658 877666
rect 701744 877610 701800 877666
rect 701886 877610 701942 877666
rect 700040 877468 700096 877524
rect 700182 877468 700238 877524
rect 700324 877468 700380 877524
rect 700466 877468 700522 877524
rect 700608 877468 700664 877524
rect 700750 877468 700806 877524
rect 700892 877468 700948 877524
rect 701034 877468 701090 877524
rect 701176 877468 701232 877524
rect 701318 877468 701374 877524
rect 701460 877468 701516 877524
rect 701602 877468 701658 877524
rect 701744 877468 701800 877524
rect 701886 877468 701942 877524
rect 700040 877326 700096 877382
rect 700182 877326 700238 877382
rect 700324 877326 700380 877382
rect 700466 877326 700522 877382
rect 700608 877326 700664 877382
rect 700750 877326 700806 877382
rect 700892 877326 700948 877382
rect 701034 877326 701090 877382
rect 701176 877326 701232 877382
rect 701318 877326 701374 877382
rect 701460 877326 701516 877382
rect 701602 877326 701658 877382
rect 701744 877326 701800 877382
rect 701886 877326 701942 877382
rect 700040 877184 700096 877240
rect 700182 877184 700238 877240
rect 700324 877184 700380 877240
rect 700466 877184 700522 877240
rect 700608 877184 700664 877240
rect 700750 877184 700806 877240
rect 700892 877184 700948 877240
rect 701034 877184 701090 877240
rect 701176 877184 701232 877240
rect 701318 877184 701374 877240
rect 701460 877184 701516 877240
rect 701602 877184 701658 877240
rect 701744 877184 701800 877240
rect 701886 877184 701942 877240
rect 700040 877042 700096 877098
rect 700182 877042 700238 877098
rect 700324 877042 700380 877098
rect 700466 877042 700522 877098
rect 700608 877042 700664 877098
rect 700750 877042 700806 877098
rect 700892 877042 700948 877098
rect 701034 877042 701090 877098
rect 701176 877042 701232 877098
rect 701318 877042 701374 877098
rect 701460 877042 701516 877098
rect 701602 877042 701658 877098
rect 701744 877042 701800 877098
rect 701886 877042 701942 877098
rect 700040 876900 700096 876956
rect 700182 876900 700238 876956
rect 700324 876900 700380 876956
rect 700466 876900 700522 876956
rect 700608 876900 700664 876956
rect 700750 876900 700806 876956
rect 700892 876900 700948 876956
rect 701034 876900 701090 876956
rect 701176 876900 701232 876956
rect 701318 876900 701374 876956
rect 701460 876900 701516 876956
rect 701602 876900 701658 876956
rect 701744 876900 701800 876956
rect 701886 876900 701942 876956
rect 700040 876758 700096 876814
rect 700182 876758 700238 876814
rect 700324 876758 700380 876814
rect 700466 876758 700522 876814
rect 700608 876758 700664 876814
rect 700750 876758 700806 876814
rect 700892 876758 700948 876814
rect 701034 876758 701090 876814
rect 701176 876758 701232 876814
rect 701318 876758 701374 876814
rect 701460 876758 701516 876814
rect 701602 876758 701658 876814
rect 701744 876758 701800 876814
rect 701886 876758 701942 876814
rect 700040 876616 700096 876672
rect 700182 876616 700238 876672
rect 700324 876616 700380 876672
rect 700466 876616 700522 876672
rect 700608 876616 700664 876672
rect 700750 876616 700806 876672
rect 700892 876616 700948 876672
rect 701034 876616 701090 876672
rect 701176 876616 701232 876672
rect 701318 876616 701374 876672
rect 701460 876616 701516 876672
rect 701602 876616 701658 876672
rect 701744 876616 701800 876672
rect 701886 876616 701942 876672
rect 700040 876474 700096 876530
rect 700182 876474 700238 876530
rect 700324 876474 700380 876530
rect 700466 876474 700522 876530
rect 700608 876474 700664 876530
rect 700750 876474 700806 876530
rect 700892 876474 700948 876530
rect 701034 876474 701090 876530
rect 701176 876474 701232 876530
rect 701318 876474 701374 876530
rect 701460 876474 701516 876530
rect 701602 876474 701658 876530
rect 701744 876474 701800 876530
rect 701886 876474 701942 876530
rect 700040 876332 700096 876388
rect 700182 876332 700238 876388
rect 700324 876332 700380 876388
rect 700466 876332 700522 876388
rect 700608 876332 700664 876388
rect 700750 876332 700806 876388
rect 700892 876332 700948 876388
rect 701034 876332 701090 876388
rect 701176 876332 701232 876388
rect 701318 876332 701374 876388
rect 701460 876332 701516 876388
rect 701602 876332 701658 876388
rect 701744 876332 701800 876388
rect 701886 876332 701942 876388
rect 73855 876113 73911 876169
rect 73997 876113 74053 876169
rect 74139 876113 74195 876169
rect 74281 876113 74337 876169
rect 74423 876113 74479 876169
rect 74565 876113 74621 876169
rect 74707 876113 74763 876169
rect 74849 876113 74905 876169
rect 74991 876113 75047 876169
rect 75133 876113 75189 876169
rect 75275 876113 75331 876169
rect 75417 876113 75473 876169
rect 75559 876113 75615 876169
rect 75701 876113 75757 876169
rect 73855 875971 73911 876027
rect 73997 875971 74053 876027
rect 74139 875971 74195 876027
rect 74281 875971 74337 876027
rect 74423 875971 74479 876027
rect 74565 875971 74621 876027
rect 74707 875971 74763 876027
rect 74849 875971 74905 876027
rect 74991 875971 75047 876027
rect 75133 875971 75189 876027
rect 75275 875971 75331 876027
rect 75417 875971 75473 876027
rect 75559 875971 75615 876027
rect 75701 875971 75757 876027
rect 73855 875829 73911 875885
rect 73997 875829 74053 875885
rect 74139 875829 74195 875885
rect 74281 875829 74337 875885
rect 74423 875829 74479 875885
rect 74565 875829 74621 875885
rect 74707 875829 74763 875885
rect 74849 875829 74905 875885
rect 74991 875829 75047 875885
rect 75133 875829 75189 875885
rect 75275 875829 75331 875885
rect 75417 875829 75473 875885
rect 75559 875829 75615 875885
rect 75701 875829 75757 875885
rect 700040 876190 700096 876246
rect 700182 876190 700238 876246
rect 700324 876190 700380 876246
rect 700466 876190 700522 876246
rect 700608 876190 700664 876246
rect 700750 876190 700806 876246
rect 700892 876190 700948 876246
rect 701034 876190 701090 876246
rect 701176 876190 701232 876246
rect 701318 876190 701374 876246
rect 701460 876190 701516 876246
rect 701602 876190 701658 876246
rect 701744 876190 701800 876246
rect 701886 876190 701942 876246
rect 700040 876048 700096 876104
rect 700182 876048 700238 876104
rect 700324 876048 700380 876104
rect 700466 876048 700522 876104
rect 700608 876048 700664 876104
rect 700750 876048 700806 876104
rect 700892 876048 700948 876104
rect 701034 876048 701090 876104
rect 701176 876048 701232 876104
rect 701318 876048 701374 876104
rect 701460 876048 701516 876104
rect 701602 876048 701658 876104
rect 701744 876048 701800 876104
rect 701886 876048 701942 876104
rect 700040 875906 700096 875962
rect 700182 875906 700238 875962
rect 700324 875906 700380 875962
rect 700466 875906 700522 875962
rect 700608 875906 700664 875962
rect 700750 875906 700806 875962
rect 700892 875906 700948 875962
rect 701034 875906 701090 875962
rect 701176 875906 701232 875962
rect 701318 875906 701374 875962
rect 701460 875906 701516 875962
rect 701602 875906 701658 875962
rect 701744 875906 701800 875962
rect 701886 875906 701942 875962
rect 73855 875687 73911 875743
rect 73997 875687 74053 875743
rect 74139 875687 74195 875743
rect 74281 875687 74337 875743
rect 74423 875687 74479 875743
rect 74565 875687 74621 875743
rect 74707 875687 74763 875743
rect 74849 875687 74905 875743
rect 74991 875687 75047 875743
rect 75133 875687 75189 875743
rect 75275 875687 75331 875743
rect 75417 875687 75473 875743
rect 75559 875687 75615 875743
rect 75701 875687 75757 875743
rect 73855 875545 73911 875601
rect 73997 875545 74053 875601
rect 74139 875545 74195 875601
rect 74281 875545 74337 875601
rect 74423 875545 74479 875601
rect 74565 875545 74621 875601
rect 74707 875545 74763 875601
rect 74849 875545 74905 875601
rect 74991 875545 75047 875601
rect 75133 875545 75189 875601
rect 75275 875545 75331 875601
rect 75417 875545 75473 875601
rect 75559 875545 75615 875601
rect 75701 875545 75757 875601
rect 73855 875403 73911 875459
rect 73997 875403 74053 875459
rect 74139 875403 74195 875459
rect 74281 875403 74337 875459
rect 74423 875403 74479 875459
rect 74565 875403 74621 875459
rect 74707 875403 74763 875459
rect 74849 875403 74905 875459
rect 74991 875403 75047 875459
rect 75133 875403 75189 875459
rect 75275 875403 75331 875459
rect 75417 875403 75473 875459
rect 75559 875403 75615 875459
rect 75701 875403 75757 875459
rect 73855 875261 73911 875317
rect 73997 875261 74053 875317
rect 74139 875261 74195 875317
rect 74281 875261 74337 875317
rect 74423 875261 74479 875317
rect 74565 875261 74621 875317
rect 74707 875261 74763 875317
rect 74849 875261 74905 875317
rect 74991 875261 75047 875317
rect 75133 875261 75189 875317
rect 75275 875261 75331 875317
rect 75417 875261 75473 875317
rect 75559 875261 75615 875317
rect 75701 875261 75757 875317
rect 73855 875119 73911 875175
rect 73997 875119 74053 875175
rect 74139 875119 74195 875175
rect 74281 875119 74337 875175
rect 74423 875119 74479 875175
rect 74565 875119 74621 875175
rect 74707 875119 74763 875175
rect 74849 875119 74905 875175
rect 74991 875119 75047 875175
rect 75133 875119 75189 875175
rect 75275 875119 75331 875175
rect 75417 875119 75473 875175
rect 75559 875119 75615 875175
rect 75701 875119 75757 875175
rect 73855 874977 73911 875033
rect 73997 874977 74053 875033
rect 74139 874977 74195 875033
rect 74281 874977 74337 875033
rect 74423 874977 74479 875033
rect 74565 874977 74621 875033
rect 74707 874977 74763 875033
rect 74849 874977 74905 875033
rect 74991 874977 75047 875033
rect 75133 874977 75189 875033
rect 75275 874977 75331 875033
rect 75417 874977 75473 875033
rect 75559 874977 75615 875033
rect 75701 874977 75757 875033
rect 73855 874835 73911 874891
rect 73997 874835 74053 874891
rect 74139 874835 74195 874891
rect 74281 874835 74337 874891
rect 74423 874835 74479 874891
rect 74565 874835 74621 874891
rect 74707 874835 74763 874891
rect 74849 874835 74905 874891
rect 74991 874835 75047 874891
rect 75133 874835 75189 874891
rect 75275 874835 75331 874891
rect 75417 874835 75473 874891
rect 75559 874835 75615 874891
rect 75701 874835 75757 874891
rect 73855 874693 73911 874749
rect 73997 874693 74053 874749
rect 74139 874693 74195 874749
rect 74281 874693 74337 874749
rect 74423 874693 74479 874749
rect 74565 874693 74621 874749
rect 74707 874693 74763 874749
rect 74849 874693 74905 874749
rect 74991 874693 75047 874749
rect 75133 874693 75189 874749
rect 75275 874693 75331 874749
rect 75417 874693 75473 874749
rect 75559 874693 75615 874749
rect 75701 874693 75757 874749
rect 73855 874551 73911 874607
rect 73997 874551 74053 874607
rect 74139 874551 74195 874607
rect 74281 874551 74337 874607
rect 74423 874551 74479 874607
rect 74565 874551 74621 874607
rect 74707 874551 74763 874607
rect 74849 874551 74905 874607
rect 74991 874551 75047 874607
rect 75133 874551 75189 874607
rect 75275 874551 75331 874607
rect 75417 874551 75473 874607
rect 75559 874551 75615 874607
rect 75701 874551 75757 874607
rect 73855 874409 73911 874465
rect 73997 874409 74053 874465
rect 74139 874409 74195 874465
rect 74281 874409 74337 874465
rect 74423 874409 74479 874465
rect 74565 874409 74621 874465
rect 74707 874409 74763 874465
rect 74849 874409 74905 874465
rect 74991 874409 75047 874465
rect 75133 874409 75189 874465
rect 75275 874409 75331 874465
rect 75417 874409 75473 874465
rect 75559 874409 75615 874465
rect 75701 874409 75757 874465
rect 73855 874267 73911 874323
rect 73997 874267 74053 874323
rect 74139 874267 74195 874323
rect 74281 874267 74337 874323
rect 74423 874267 74479 874323
rect 74565 874267 74621 874323
rect 74707 874267 74763 874323
rect 74849 874267 74905 874323
rect 74991 874267 75047 874323
rect 75133 874267 75189 874323
rect 75275 874267 75331 874323
rect 75417 874267 75473 874323
rect 75559 874267 75615 874323
rect 75701 874267 75757 874323
rect 700051 875123 700107 875179
rect 700193 875123 700249 875179
rect 700335 875123 700391 875179
rect 700477 875123 700533 875179
rect 700619 875123 700675 875179
rect 700761 875123 700817 875179
rect 700903 875123 700959 875179
rect 701045 875123 701101 875179
rect 701187 875123 701243 875179
rect 701329 875123 701385 875179
rect 701471 875123 701527 875179
rect 701613 875123 701669 875179
rect 701755 875123 701811 875179
rect 701897 875123 701953 875179
rect 700051 874981 700107 875037
rect 700193 874981 700249 875037
rect 700335 874981 700391 875037
rect 700477 874981 700533 875037
rect 700619 874981 700675 875037
rect 700761 874981 700817 875037
rect 700903 874981 700959 875037
rect 701045 874981 701101 875037
rect 701187 874981 701243 875037
rect 701329 874981 701385 875037
rect 701471 874981 701527 875037
rect 701613 874981 701669 875037
rect 701755 874981 701811 875037
rect 701897 874981 701953 875037
rect 700051 874839 700107 874895
rect 700193 874839 700249 874895
rect 700335 874839 700391 874895
rect 700477 874839 700533 874895
rect 700619 874839 700675 874895
rect 700761 874839 700817 874895
rect 700903 874839 700959 874895
rect 701045 874839 701101 874895
rect 701187 874839 701243 874895
rect 701329 874839 701385 874895
rect 701471 874839 701527 874895
rect 701613 874839 701669 874895
rect 701755 874839 701811 874895
rect 701897 874839 701953 874895
rect 700051 874697 700107 874753
rect 700193 874697 700249 874753
rect 700335 874697 700391 874753
rect 700477 874697 700533 874753
rect 700619 874697 700675 874753
rect 700761 874697 700817 874753
rect 700903 874697 700959 874753
rect 701045 874697 701101 874753
rect 701187 874697 701243 874753
rect 701329 874697 701385 874753
rect 701471 874697 701527 874753
rect 701613 874697 701669 874753
rect 701755 874697 701811 874753
rect 701897 874697 701953 874753
rect 700051 874555 700107 874611
rect 700193 874555 700249 874611
rect 700335 874555 700391 874611
rect 700477 874555 700533 874611
rect 700619 874555 700675 874611
rect 700761 874555 700817 874611
rect 700903 874555 700959 874611
rect 701045 874555 701101 874611
rect 701187 874555 701243 874611
rect 701329 874555 701385 874611
rect 701471 874555 701527 874611
rect 701613 874555 701669 874611
rect 701755 874555 701811 874611
rect 701897 874555 701953 874611
rect 700051 874413 700107 874469
rect 700193 874413 700249 874469
rect 700335 874413 700391 874469
rect 700477 874413 700533 874469
rect 700619 874413 700675 874469
rect 700761 874413 700817 874469
rect 700903 874413 700959 874469
rect 701045 874413 701101 874469
rect 701187 874413 701243 874469
rect 701329 874413 701385 874469
rect 701471 874413 701527 874469
rect 701613 874413 701669 874469
rect 701755 874413 701811 874469
rect 701897 874413 701953 874469
rect 700051 874271 700107 874327
rect 700193 874271 700249 874327
rect 700335 874271 700391 874327
rect 700477 874271 700533 874327
rect 700619 874271 700675 874327
rect 700761 874271 700817 874327
rect 700903 874271 700959 874327
rect 701045 874271 701101 874327
rect 701187 874271 701243 874327
rect 701329 874271 701385 874327
rect 701471 874271 701527 874327
rect 701613 874271 701669 874327
rect 701755 874271 701811 874327
rect 701897 874271 701953 874327
rect 700051 874129 700107 874185
rect 700193 874129 700249 874185
rect 700335 874129 700391 874185
rect 700477 874129 700533 874185
rect 700619 874129 700675 874185
rect 700761 874129 700817 874185
rect 700903 874129 700959 874185
rect 701045 874129 701101 874185
rect 701187 874129 701243 874185
rect 701329 874129 701385 874185
rect 701471 874129 701527 874185
rect 701613 874129 701669 874185
rect 701755 874129 701811 874185
rect 701897 874129 701953 874185
rect 700051 873987 700107 874043
rect 700193 873987 700249 874043
rect 700335 873987 700391 874043
rect 700477 873987 700533 874043
rect 700619 873987 700675 874043
rect 700761 873987 700817 874043
rect 700903 873987 700959 874043
rect 701045 873987 701101 874043
rect 701187 873987 701243 874043
rect 701329 873987 701385 874043
rect 701471 873987 701527 874043
rect 701613 873987 701669 874043
rect 701755 873987 701811 874043
rect 701897 873987 701953 874043
rect 73855 873743 73911 873799
rect 73997 873743 74053 873799
rect 74139 873743 74195 873799
rect 74281 873743 74337 873799
rect 74423 873743 74479 873799
rect 74565 873743 74621 873799
rect 74707 873743 74763 873799
rect 74849 873743 74905 873799
rect 74991 873743 75047 873799
rect 75133 873743 75189 873799
rect 75275 873743 75331 873799
rect 75417 873743 75473 873799
rect 75559 873743 75615 873799
rect 75701 873743 75757 873799
rect 73855 873601 73911 873657
rect 73997 873601 74053 873657
rect 74139 873601 74195 873657
rect 74281 873601 74337 873657
rect 74423 873601 74479 873657
rect 74565 873601 74621 873657
rect 74707 873601 74763 873657
rect 74849 873601 74905 873657
rect 74991 873601 75047 873657
rect 75133 873601 75189 873657
rect 75275 873601 75331 873657
rect 75417 873601 75473 873657
rect 75559 873601 75615 873657
rect 75701 873601 75757 873657
rect 73855 873459 73911 873515
rect 73997 873459 74053 873515
rect 74139 873459 74195 873515
rect 74281 873459 74337 873515
rect 74423 873459 74479 873515
rect 74565 873459 74621 873515
rect 74707 873459 74763 873515
rect 74849 873459 74905 873515
rect 74991 873459 75047 873515
rect 75133 873459 75189 873515
rect 75275 873459 75331 873515
rect 75417 873459 75473 873515
rect 75559 873459 75615 873515
rect 75701 873459 75757 873515
rect 73855 873317 73911 873373
rect 73997 873317 74053 873373
rect 74139 873317 74195 873373
rect 74281 873317 74337 873373
rect 74423 873317 74479 873373
rect 74565 873317 74621 873373
rect 74707 873317 74763 873373
rect 74849 873317 74905 873373
rect 74991 873317 75047 873373
rect 75133 873317 75189 873373
rect 75275 873317 75331 873373
rect 75417 873317 75473 873373
rect 75559 873317 75615 873373
rect 75701 873317 75757 873373
rect 73855 873175 73911 873231
rect 73997 873175 74053 873231
rect 74139 873175 74195 873231
rect 74281 873175 74337 873231
rect 74423 873175 74479 873231
rect 74565 873175 74621 873231
rect 74707 873175 74763 873231
rect 74849 873175 74905 873231
rect 74991 873175 75047 873231
rect 75133 873175 75189 873231
rect 75275 873175 75331 873231
rect 75417 873175 75473 873231
rect 75559 873175 75615 873231
rect 75701 873175 75757 873231
rect 700051 873845 700107 873901
rect 700193 873845 700249 873901
rect 700335 873845 700391 873901
rect 700477 873845 700533 873901
rect 700619 873845 700675 873901
rect 700761 873845 700817 873901
rect 700903 873845 700959 873901
rect 701045 873845 701101 873901
rect 701187 873845 701243 873901
rect 701329 873845 701385 873901
rect 701471 873845 701527 873901
rect 701613 873845 701669 873901
rect 701755 873845 701811 873901
rect 701897 873845 701953 873901
rect 700051 873703 700107 873759
rect 700193 873703 700249 873759
rect 700335 873703 700391 873759
rect 700477 873703 700533 873759
rect 700619 873703 700675 873759
rect 700761 873703 700817 873759
rect 700903 873703 700959 873759
rect 701045 873703 701101 873759
rect 701187 873703 701243 873759
rect 701329 873703 701385 873759
rect 701471 873703 701527 873759
rect 701613 873703 701669 873759
rect 701755 873703 701811 873759
rect 701897 873703 701953 873759
rect 700051 873561 700107 873617
rect 700193 873561 700249 873617
rect 700335 873561 700391 873617
rect 700477 873561 700533 873617
rect 700619 873561 700675 873617
rect 700761 873561 700817 873617
rect 700903 873561 700959 873617
rect 701045 873561 701101 873617
rect 701187 873561 701243 873617
rect 701329 873561 701385 873617
rect 701471 873561 701527 873617
rect 701613 873561 701669 873617
rect 701755 873561 701811 873617
rect 701897 873561 701953 873617
rect 700051 873419 700107 873475
rect 700193 873419 700249 873475
rect 700335 873419 700391 873475
rect 700477 873419 700533 873475
rect 700619 873419 700675 873475
rect 700761 873419 700817 873475
rect 700903 873419 700959 873475
rect 701045 873419 701101 873475
rect 701187 873419 701243 873475
rect 701329 873419 701385 873475
rect 701471 873419 701527 873475
rect 701613 873419 701669 873475
rect 701755 873419 701811 873475
rect 701897 873419 701953 873475
rect 700051 873277 700107 873333
rect 700193 873277 700249 873333
rect 700335 873277 700391 873333
rect 700477 873277 700533 873333
rect 700619 873277 700675 873333
rect 700761 873277 700817 873333
rect 700903 873277 700959 873333
rect 701045 873277 701101 873333
rect 701187 873277 701243 873333
rect 701329 873277 701385 873333
rect 701471 873277 701527 873333
rect 701613 873277 701669 873333
rect 701755 873277 701811 873333
rect 701897 873277 701953 873333
rect 73855 873033 73911 873089
rect 73997 873033 74053 873089
rect 74139 873033 74195 873089
rect 74281 873033 74337 873089
rect 74423 873033 74479 873089
rect 74565 873033 74621 873089
rect 74707 873033 74763 873089
rect 74849 873033 74905 873089
rect 74991 873033 75047 873089
rect 75133 873033 75189 873089
rect 75275 873033 75331 873089
rect 75417 873033 75473 873089
rect 75559 873033 75615 873089
rect 75701 873033 75757 873089
rect 73855 872891 73911 872947
rect 73997 872891 74053 872947
rect 74139 872891 74195 872947
rect 74281 872891 74337 872947
rect 74423 872891 74479 872947
rect 74565 872891 74621 872947
rect 74707 872891 74763 872947
rect 74849 872891 74905 872947
rect 74991 872891 75047 872947
rect 75133 872891 75189 872947
rect 75275 872891 75331 872947
rect 75417 872891 75473 872947
rect 75559 872891 75615 872947
rect 75701 872891 75757 872947
rect 73855 872749 73911 872805
rect 73997 872749 74053 872805
rect 74139 872749 74195 872805
rect 74281 872749 74337 872805
rect 74423 872749 74479 872805
rect 74565 872749 74621 872805
rect 74707 872749 74763 872805
rect 74849 872749 74905 872805
rect 74991 872749 75047 872805
rect 75133 872749 75189 872805
rect 75275 872749 75331 872805
rect 75417 872749 75473 872805
rect 75559 872749 75615 872805
rect 75701 872749 75757 872805
rect 73855 872607 73911 872663
rect 73997 872607 74053 872663
rect 74139 872607 74195 872663
rect 74281 872607 74337 872663
rect 74423 872607 74479 872663
rect 74565 872607 74621 872663
rect 74707 872607 74763 872663
rect 74849 872607 74905 872663
rect 74991 872607 75047 872663
rect 75133 872607 75189 872663
rect 75275 872607 75331 872663
rect 75417 872607 75473 872663
rect 75559 872607 75615 872663
rect 75701 872607 75757 872663
rect 73855 872465 73911 872521
rect 73997 872465 74053 872521
rect 74139 872465 74195 872521
rect 74281 872465 74337 872521
rect 74423 872465 74479 872521
rect 74565 872465 74621 872521
rect 74707 872465 74763 872521
rect 74849 872465 74905 872521
rect 74991 872465 75047 872521
rect 75133 872465 75189 872521
rect 75275 872465 75331 872521
rect 75417 872465 75473 872521
rect 75559 872465 75615 872521
rect 75701 872465 75757 872521
rect 73855 872323 73911 872379
rect 73997 872323 74053 872379
rect 74139 872323 74195 872379
rect 74281 872323 74337 872379
rect 74423 872323 74479 872379
rect 74565 872323 74621 872379
rect 74707 872323 74763 872379
rect 74849 872323 74905 872379
rect 74991 872323 75047 872379
rect 75133 872323 75189 872379
rect 75275 872323 75331 872379
rect 75417 872323 75473 872379
rect 75559 872323 75615 872379
rect 75701 872323 75757 872379
rect 73855 872181 73911 872237
rect 73997 872181 74053 872237
rect 74139 872181 74195 872237
rect 74281 872181 74337 872237
rect 74423 872181 74479 872237
rect 74565 872181 74621 872237
rect 74707 872181 74763 872237
rect 74849 872181 74905 872237
rect 74991 872181 75047 872237
rect 75133 872181 75189 872237
rect 75275 872181 75331 872237
rect 75417 872181 75473 872237
rect 75559 872181 75615 872237
rect 75701 872181 75757 872237
rect 73855 872039 73911 872095
rect 73997 872039 74053 872095
rect 74139 872039 74195 872095
rect 74281 872039 74337 872095
rect 74423 872039 74479 872095
rect 74565 872039 74621 872095
rect 74707 872039 74763 872095
rect 74849 872039 74905 872095
rect 74991 872039 75047 872095
rect 75133 872039 75189 872095
rect 75275 872039 75331 872095
rect 75417 872039 75473 872095
rect 75559 872039 75615 872095
rect 75701 872039 75757 872095
rect 73855 871897 73911 871953
rect 73997 871897 74053 871953
rect 74139 871897 74195 871953
rect 74281 871897 74337 871953
rect 74423 871897 74479 871953
rect 74565 871897 74621 871953
rect 74707 871897 74763 871953
rect 74849 871897 74905 871953
rect 74991 871897 75047 871953
rect 75133 871897 75189 871953
rect 75275 871897 75331 871953
rect 75417 871897 75473 871953
rect 75559 871897 75615 871953
rect 75701 871897 75757 871953
rect 700051 872753 700107 872809
rect 700193 872753 700249 872809
rect 700335 872753 700391 872809
rect 700477 872753 700533 872809
rect 700619 872753 700675 872809
rect 700761 872753 700817 872809
rect 700903 872753 700959 872809
rect 701045 872753 701101 872809
rect 701187 872753 701243 872809
rect 701329 872753 701385 872809
rect 701471 872753 701527 872809
rect 701613 872753 701669 872809
rect 701755 872753 701811 872809
rect 701897 872753 701953 872809
rect 700051 872611 700107 872667
rect 700193 872611 700249 872667
rect 700335 872611 700391 872667
rect 700477 872611 700533 872667
rect 700619 872611 700675 872667
rect 700761 872611 700817 872667
rect 700903 872611 700959 872667
rect 701045 872611 701101 872667
rect 701187 872611 701243 872667
rect 701329 872611 701385 872667
rect 701471 872611 701527 872667
rect 701613 872611 701669 872667
rect 701755 872611 701811 872667
rect 701897 872611 701953 872667
rect 700051 872469 700107 872525
rect 700193 872469 700249 872525
rect 700335 872469 700391 872525
rect 700477 872469 700533 872525
rect 700619 872469 700675 872525
rect 700761 872469 700817 872525
rect 700903 872469 700959 872525
rect 701045 872469 701101 872525
rect 701187 872469 701243 872525
rect 701329 872469 701385 872525
rect 701471 872469 701527 872525
rect 701613 872469 701669 872525
rect 701755 872469 701811 872525
rect 701897 872469 701953 872525
rect 700051 872327 700107 872383
rect 700193 872327 700249 872383
rect 700335 872327 700391 872383
rect 700477 872327 700533 872383
rect 700619 872327 700675 872383
rect 700761 872327 700817 872383
rect 700903 872327 700959 872383
rect 701045 872327 701101 872383
rect 701187 872327 701243 872383
rect 701329 872327 701385 872383
rect 701471 872327 701527 872383
rect 701613 872327 701669 872383
rect 701755 872327 701811 872383
rect 701897 872327 701953 872383
rect 700051 872185 700107 872241
rect 700193 872185 700249 872241
rect 700335 872185 700391 872241
rect 700477 872185 700533 872241
rect 700619 872185 700675 872241
rect 700761 872185 700817 872241
rect 700903 872185 700959 872241
rect 701045 872185 701101 872241
rect 701187 872185 701243 872241
rect 701329 872185 701385 872241
rect 701471 872185 701527 872241
rect 701613 872185 701669 872241
rect 701755 872185 701811 872241
rect 701897 872185 701953 872241
rect 700051 872043 700107 872099
rect 700193 872043 700249 872099
rect 700335 872043 700391 872099
rect 700477 872043 700533 872099
rect 700619 872043 700675 872099
rect 700761 872043 700817 872099
rect 700903 872043 700959 872099
rect 701045 872043 701101 872099
rect 701187 872043 701243 872099
rect 701329 872043 701385 872099
rect 701471 872043 701527 872099
rect 701613 872043 701669 872099
rect 701755 872043 701811 872099
rect 701897 872043 701953 872099
rect 700051 871901 700107 871957
rect 700193 871901 700249 871957
rect 700335 871901 700391 871957
rect 700477 871901 700533 871957
rect 700619 871901 700675 871957
rect 700761 871901 700817 871957
rect 700903 871901 700959 871957
rect 701045 871901 701101 871957
rect 701187 871901 701243 871957
rect 701329 871901 701385 871957
rect 701471 871901 701527 871957
rect 701613 871901 701669 871957
rect 701755 871901 701811 871957
rect 701897 871901 701953 871957
rect 700051 871759 700107 871815
rect 700193 871759 700249 871815
rect 700335 871759 700391 871815
rect 700477 871759 700533 871815
rect 700619 871759 700675 871815
rect 700761 871759 700817 871815
rect 700903 871759 700959 871815
rect 701045 871759 701101 871815
rect 701187 871759 701243 871815
rect 701329 871759 701385 871815
rect 701471 871759 701527 871815
rect 701613 871759 701669 871815
rect 701755 871759 701811 871815
rect 701897 871759 701953 871815
rect 700051 871617 700107 871673
rect 700193 871617 700249 871673
rect 700335 871617 700391 871673
rect 700477 871617 700533 871673
rect 700619 871617 700675 871673
rect 700761 871617 700817 871673
rect 700903 871617 700959 871673
rect 701045 871617 701101 871673
rect 701187 871617 701243 871673
rect 701329 871617 701385 871673
rect 701471 871617 701527 871673
rect 701613 871617 701669 871673
rect 701755 871617 701811 871673
rect 701897 871617 701953 871673
rect 700051 871475 700107 871531
rect 700193 871475 700249 871531
rect 700335 871475 700391 871531
rect 700477 871475 700533 871531
rect 700619 871475 700675 871531
rect 700761 871475 700817 871531
rect 700903 871475 700959 871531
rect 701045 871475 701101 871531
rect 701187 871475 701243 871531
rect 701329 871475 701385 871531
rect 701471 871475 701527 871531
rect 701613 871475 701669 871531
rect 701755 871475 701811 871531
rect 701897 871475 701953 871531
rect 700051 871333 700107 871389
rect 700193 871333 700249 871389
rect 700335 871333 700391 871389
rect 700477 871333 700533 871389
rect 700619 871333 700675 871389
rect 700761 871333 700817 871389
rect 700903 871333 700959 871389
rect 701045 871333 701101 871389
rect 701187 871333 701243 871389
rect 701329 871333 701385 871389
rect 701471 871333 701527 871389
rect 701613 871333 701669 871389
rect 701755 871333 701811 871389
rect 701897 871333 701953 871389
rect 700051 871191 700107 871247
rect 700193 871191 700249 871247
rect 700335 871191 700391 871247
rect 700477 871191 700533 871247
rect 700619 871191 700675 871247
rect 700761 871191 700817 871247
rect 700903 871191 700959 871247
rect 701045 871191 701101 871247
rect 701187 871191 701243 871247
rect 701329 871191 701385 871247
rect 701471 871191 701527 871247
rect 701613 871191 701669 871247
rect 701755 871191 701811 871247
rect 701897 871191 701953 871247
rect 73855 871037 73911 871093
rect 73997 871037 74053 871093
rect 74139 871037 74195 871093
rect 74281 871037 74337 871093
rect 74423 871037 74479 871093
rect 74565 871037 74621 871093
rect 74707 871037 74763 871093
rect 74849 871037 74905 871093
rect 74991 871037 75047 871093
rect 75133 871037 75189 871093
rect 75275 871037 75331 871093
rect 75417 871037 75473 871093
rect 75559 871037 75615 871093
rect 75701 871037 75757 871093
rect 73855 870895 73911 870951
rect 73997 870895 74053 870951
rect 74139 870895 74195 870951
rect 74281 870895 74337 870951
rect 74423 870895 74479 870951
rect 74565 870895 74621 870951
rect 74707 870895 74763 870951
rect 74849 870895 74905 870951
rect 74991 870895 75047 870951
rect 75133 870895 75189 870951
rect 75275 870895 75331 870951
rect 75417 870895 75473 870951
rect 75559 870895 75615 870951
rect 75701 870895 75757 870951
rect 700051 871049 700107 871105
rect 700193 871049 700249 871105
rect 700335 871049 700391 871105
rect 700477 871049 700533 871105
rect 700619 871049 700675 871105
rect 700761 871049 700817 871105
rect 700903 871049 700959 871105
rect 701045 871049 701101 871105
rect 701187 871049 701243 871105
rect 701329 871049 701385 871105
rect 701471 871049 701527 871105
rect 701613 871049 701669 871105
rect 701755 871049 701811 871105
rect 701897 871049 701953 871105
rect 700051 870907 700107 870963
rect 700193 870907 700249 870963
rect 700335 870907 700391 870963
rect 700477 870907 700533 870963
rect 700619 870907 700675 870963
rect 700761 870907 700817 870963
rect 700903 870907 700959 870963
rect 701045 870907 701101 870963
rect 701187 870907 701243 870963
rect 701329 870907 701385 870963
rect 701471 870907 701527 870963
rect 701613 870907 701669 870963
rect 701755 870907 701811 870963
rect 701897 870907 701953 870963
rect 73855 870753 73911 870809
rect 73997 870753 74053 870809
rect 74139 870753 74195 870809
rect 74281 870753 74337 870809
rect 74423 870753 74479 870809
rect 74565 870753 74621 870809
rect 74707 870753 74763 870809
rect 74849 870753 74905 870809
rect 74991 870753 75047 870809
rect 75133 870753 75189 870809
rect 75275 870753 75331 870809
rect 75417 870753 75473 870809
rect 75559 870753 75615 870809
rect 75701 870753 75757 870809
rect 73855 870611 73911 870667
rect 73997 870611 74053 870667
rect 74139 870611 74195 870667
rect 74281 870611 74337 870667
rect 74423 870611 74479 870667
rect 74565 870611 74621 870667
rect 74707 870611 74763 870667
rect 74849 870611 74905 870667
rect 74991 870611 75047 870667
rect 75133 870611 75189 870667
rect 75275 870611 75331 870667
rect 75417 870611 75473 870667
rect 75559 870611 75615 870667
rect 75701 870611 75757 870667
rect 73855 870469 73911 870525
rect 73997 870469 74053 870525
rect 74139 870469 74195 870525
rect 74281 870469 74337 870525
rect 74423 870469 74479 870525
rect 74565 870469 74621 870525
rect 74707 870469 74763 870525
rect 74849 870469 74905 870525
rect 74991 870469 75047 870525
rect 75133 870469 75189 870525
rect 75275 870469 75331 870525
rect 75417 870469 75473 870525
rect 75559 870469 75615 870525
rect 75701 870469 75757 870525
rect 73855 870327 73911 870383
rect 73997 870327 74053 870383
rect 74139 870327 74195 870383
rect 74281 870327 74337 870383
rect 74423 870327 74479 870383
rect 74565 870327 74621 870383
rect 74707 870327 74763 870383
rect 74849 870327 74905 870383
rect 74991 870327 75047 870383
rect 75133 870327 75189 870383
rect 75275 870327 75331 870383
rect 75417 870327 75473 870383
rect 75559 870327 75615 870383
rect 75701 870327 75757 870383
rect 73855 870185 73911 870241
rect 73997 870185 74053 870241
rect 74139 870185 74195 870241
rect 74281 870185 74337 870241
rect 74423 870185 74479 870241
rect 74565 870185 74621 870241
rect 74707 870185 74763 870241
rect 74849 870185 74905 870241
rect 74991 870185 75047 870241
rect 75133 870185 75189 870241
rect 75275 870185 75331 870241
rect 75417 870185 75473 870241
rect 75559 870185 75615 870241
rect 75701 870185 75757 870241
rect 73855 870043 73911 870099
rect 73997 870043 74053 870099
rect 74139 870043 74195 870099
rect 74281 870043 74337 870099
rect 74423 870043 74479 870099
rect 74565 870043 74621 870099
rect 74707 870043 74763 870099
rect 74849 870043 74905 870099
rect 74991 870043 75047 870099
rect 75133 870043 75189 870099
rect 75275 870043 75331 870099
rect 75417 870043 75473 870099
rect 75559 870043 75615 870099
rect 75701 870043 75757 870099
rect 73855 869901 73911 869957
rect 73997 869901 74053 869957
rect 74139 869901 74195 869957
rect 74281 869901 74337 869957
rect 74423 869901 74479 869957
rect 74565 869901 74621 869957
rect 74707 869901 74763 869957
rect 74849 869901 74905 869957
rect 74991 869901 75047 869957
rect 75133 869901 75189 869957
rect 75275 869901 75331 869957
rect 75417 869901 75473 869957
rect 75559 869901 75615 869957
rect 75701 869901 75757 869957
rect 73855 869759 73911 869815
rect 73997 869759 74053 869815
rect 74139 869759 74195 869815
rect 74281 869759 74337 869815
rect 74423 869759 74479 869815
rect 74565 869759 74621 869815
rect 74707 869759 74763 869815
rect 74849 869759 74905 869815
rect 74991 869759 75047 869815
rect 75133 869759 75189 869815
rect 75275 869759 75331 869815
rect 75417 869759 75473 869815
rect 75559 869759 75615 869815
rect 75701 869759 75757 869815
rect 73855 869617 73911 869673
rect 73997 869617 74053 869673
rect 74139 869617 74195 869673
rect 74281 869617 74337 869673
rect 74423 869617 74479 869673
rect 74565 869617 74621 869673
rect 74707 869617 74763 869673
rect 74849 869617 74905 869673
rect 74991 869617 75047 869673
rect 75133 869617 75189 869673
rect 75275 869617 75331 869673
rect 75417 869617 75473 869673
rect 75559 869617 75615 869673
rect 75701 869617 75757 869673
rect 73855 869475 73911 869531
rect 73997 869475 74053 869531
rect 74139 869475 74195 869531
rect 74281 869475 74337 869531
rect 74423 869475 74479 869531
rect 74565 869475 74621 869531
rect 74707 869475 74763 869531
rect 74849 869475 74905 869531
rect 74991 869475 75047 869531
rect 75133 869475 75189 869531
rect 75275 869475 75331 869531
rect 75417 869475 75473 869531
rect 75559 869475 75615 869531
rect 75701 869475 75757 869531
rect 73855 869333 73911 869389
rect 73997 869333 74053 869389
rect 74139 869333 74195 869389
rect 74281 869333 74337 869389
rect 74423 869333 74479 869389
rect 74565 869333 74621 869389
rect 74707 869333 74763 869389
rect 74849 869333 74905 869389
rect 74991 869333 75047 869389
rect 75133 869333 75189 869389
rect 75275 869333 75331 869389
rect 75417 869333 75473 869389
rect 75559 869333 75615 869389
rect 75701 869333 75757 869389
rect 73855 869191 73911 869247
rect 73997 869191 74053 869247
rect 74139 869191 74195 869247
rect 74281 869191 74337 869247
rect 74423 869191 74479 869247
rect 74565 869191 74621 869247
rect 74707 869191 74763 869247
rect 74849 869191 74905 869247
rect 74991 869191 75047 869247
rect 75133 869191 75189 869247
rect 75275 869191 75331 869247
rect 75417 869191 75473 869247
rect 75559 869191 75615 869247
rect 75701 869191 75757 869247
rect 700051 870047 700107 870103
rect 700193 870047 700249 870103
rect 700335 870047 700391 870103
rect 700477 870047 700533 870103
rect 700619 870047 700675 870103
rect 700761 870047 700817 870103
rect 700903 870047 700959 870103
rect 701045 870047 701101 870103
rect 701187 870047 701243 870103
rect 701329 870047 701385 870103
rect 701471 870047 701527 870103
rect 701613 870047 701669 870103
rect 701755 870047 701811 870103
rect 701897 870047 701953 870103
rect 700051 869905 700107 869961
rect 700193 869905 700249 869961
rect 700335 869905 700391 869961
rect 700477 869905 700533 869961
rect 700619 869905 700675 869961
rect 700761 869905 700817 869961
rect 700903 869905 700959 869961
rect 701045 869905 701101 869961
rect 701187 869905 701243 869961
rect 701329 869905 701385 869961
rect 701471 869905 701527 869961
rect 701613 869905 701669 869961
rect 701755 869905 701811 869961
rect 701897 869905 701953 869961
rect 700051 869763 700107 869819
rect 700193 869763 700249 869819
rect 700335 869763 700391 869819
rect 700477 869763 700533 869819
rect 700619 869763 700675 869819
rect 700761 869763 700817 869819
rect 700903 869763 700959 869819
rect 701045 869763 701101 869819
rect 701187 869763 701243 869819
rect 701329 869763 701385 869819
rect 701471 869763 701527 869819
rect 701613 869763 701669 869819
rect 701755 869763 701811 869819
rect 701897 869763 701953 869819
rect 700051 869621 700107 869677
rect 700193 869621 700249 869677
rect 700335 869621 700391 869677
rect 700477 869621 700533 869677
rect 700619 869621 700675 869677
rect 700761 869621 700817 869677
rect 700903 869621 700959 869677
rect 701045 869621 701101 869677
rect 701187 869621 701243 869677
rect 701329 869621 701385 869677
rect 701471 869621 701527 869677
rect 701613 869621 701669 869677
rect 701755 869621 701811 869677
rect 701897 869621 701953 869677
rect 700051 869479 700107 869535
rect 700193 869479 700249 869535
rect 700335 869479 700391 869535
rect 700477 869479 700533 869535
rect 700619 869479 700675 869535
rect 700761 869479 700817 869535
rect 700903 869479 700959 869535
rect 701045 869479 701101 869535
rect 701187 869479 701243 869535
rect 701329 869479 701385 869535
rect 701471 869479 701527 869535
rect 701613 869479 701669 869535
rect 701755 869479 701811 869535
rect 701897 869479 701953 869535
rect 700051 869337 700107 869393
rect 700193 869337 700249 869393
rect 700335 869337 700391 869393
rect 700477 869337 700533 869393
rect 700619 869337 700675 869393
rect 700761 869337 700817 869393
rect 700903 869337 700959 869393
rect 701045 869337 701101 869393
rect 701187 869337 701243 869393
rect 701329 869337 701385 869393
rect 701471 869337 701527 869393
rect 701613 869337 701669 869393
rect 701755 869337 701811 869393
rect 701897 869337 701953 869393
rect 700051 869195 700107 869251
rect 700193 869195 700249 869251
rect 700335 869195 700391 869251
rect 700477 869195 700533 869251
rect 700619 869195 700675 869251
rect 700761 869195 700817 869251
rect 700903 869195 700959 869251
rect 701045 869195 701101 869251
rect 701187 869195 701243 869251
rect 701329 869195 701385 869251
rect 701471 869195 701527 869251
rect 701613 869195 701669 869251
rect 701755 869195 701811 869251
rect 701897 869195 701953 869251
rect 700051 869053 700107 869109
rect 700193 869053 700249 869109
rect 700335 869053 700391 869109
rect 700477 869053 700533 869109
rect 700619 869053 700675 869109
rect 700761 869053 700817 869109
rect 700903 869053 700959 869109
rect 701045 869053 701101 869109
rect 701187 869053 701243 869109
rect 701329 869053 701385 869109
rect 701471 869053 701527 869109
rect 701613 869053 701669 869109
rect 701755 869053 701811 869109
rect 701897 869053 701953 869109
rect 700051 868911 700107 868967
rect 700193 868911 700249 868967
rect 700335 868911 700391 868967
rect 700477 868911 700533 868967
rect 700619 868911 700675 868967
rect 700761 868911 700817 868967
rect 700903 868911 700959 868967
rect 701045 868911 701101 868967
rect 701187 868911 701243 868967
rect 701329 868911 701385 868967
rect 701471 868911 701527 868967
rect 701613 868911 701669 868967
rect 701755 868911 701811 868967
rect 701897 868911 701953 868967
rect 73855 868667 73911 868723
rect 73997 868667 74053 868723
rect 74139 868667 74195 868723
rect 74281 868667 74337 868723
rect 74423 868667 74479 868723
rect 74565 868667 74621 868723
rect 74707 868667 74763 868723
rect 74849 868667 74905 868723
rect 74991 868667 75047 868723
rect 75133 868667 75189 868723
rect 75275 868667 75331 868723
rect 75417 868667 75473 868723
rect 75559 868667 75615 868723
rect 75701 868667 75757 868723
rect 73855 868525 73911 868581
rect 73997 868525 74053 868581
rect 74139 868525 74195 868581
rect 74281 868525 74337 868581
rect 74423 868525 74479 868581
rect 74565 868525 74621 868581
rect 74707 868525 74763 868581
rect 74849 868525 74905 868581
rect 74991 868525 75047 868581
rect 75133 868525 75189 868581
rect 75275 868525 75331 868581
rect 75417 868525 75473 868581
rect 75559 868525 75615 868581
rect 75701 868525 75757 868581
rect 73855 868383 73911 868439
rect 73997 868383 74053 868439
rect 74139 868383 74195 868439
rect 74281 868383 74337 868439
rect 74423 868383 74479 868439
rect 74565 868383 74621 868439
rect 74707 868383 74763 868439
rect 74849 868383 74905 868439
rect 74991 868383 75047 868439
rect 75133 868383 75189 868439
rect 75275 868383 75331 868439
rect 75417 868383 75473 868439
rect 75559 868383 75615 868439
rect 75701 868383 75757 868439
rect 73855 868241 73911 868297
rect 73997 868241 74053 868297
rect 74139 868241 74195 868297
rect 74281 868241 74337 868297
rect 74423 868241 74479 868297
rect 74565 868241 74621 868297
rect 74707 868241 74763 868297
rect 74849 868241 74905 868297
rect 74991 868241 75047 868297
rect 75133 868241 75189 868297
rect 75275 868241 75331 868297
rect 75417 868241 75473 868297
rect 75559 868241 75615 868297
rect 75701 868241 75757 868297
rect 73855 868099 73911 868155
rect 73997 868099 74053 868155
rect 74139 868099 74195 868155
rect 74281 868099 74337 868155
rect 74423 868099 74479 868155
rect 74565 868099 74621 868155
rect 74707 868099 74763 868155
rect 74849 868099 74905 868155
rect 74991 868099 75047 868155
rect 75133 868099 75189 868155
rect 75275 868099 75331 868155
rect 75417 868099 75473 868155
rect 75559 868099 75615 868155
rect 75701 868099 75757 868155
rect 700051 868769 700107 868825
rect 700193 868769 700249 868825
rect 700335 868769 700391 868825
rect 700477 868769 700533 868825
rect 700619 868769 700675 868825
rect 700761 868769 700817 868825
rect 700903 868769 700959 868825
rect 701045 868769 701101 868825
rect 701187 868769 701243 868825
rect 701329 868769 701385 868825
rect 701471 868769 701527 868825
rect 701613 868769 701669 868825
rect 701755 868769 701811 868825
rect 701897 868769 701953 868825
rect 700051 868627 700107 868683
rect 700193 868627 700249 868683
rect 700335 868627 700391 868683
rect 700477 868627 700533 868683
rect 700619 868627 700675 868683
rect 700761 868627 700817 868683
rect 700903 868627 700959 868683
rect 701045 868627 701101 868683
rect 701187 868627 701243 868683
rect 701329 868627 701385 868683
rect 701471 868627 701527 868683
rect 701613 868627 701669 868683
rect 701755 868627 701811 868683
rect 701897 868627 701953 868683
rect 700051 868485 700107 868541
rect 700193 868485 700249 868541
rect 700335 868485 700391 868541
rect 700477 868485 700533 868541
rect 700619 868485 700675 868541
rect 700761 868485 700817 868541
rect 700903 868485 700959 868541
rect 701045 868485 701101 868541
rect 701187 868485 701243 868541
rect 701329 868485 701385 868541
rect 701471 868485 701527 868541
rect 701613 868485 701669 868541
rect 701755 868485 701811 868541
rect 701897 868485 701953 868541
rect 700051 868343 700107 868399
rect 700193 868343 700249 868399
rect 700335 868343 700391 868399
rect 700477 868343 700533 868399
rect 700619 868343 700675 868399
rect 700761 868343 700817 868399
rect 700903 868343 700959 868399
rect 701045 868343 701101 868399
rect 701187 868343 701243 868399
rect 701329 868343 701385 868399
rect 701471 868343 701527 868399
rect 701613 868343 701669 868399
rect 701755 868343 701811 868399
rect 701897 868343 701953 868399
rect 700051 868201 700107 868257
rect 700193 868201 700249 868257
rect 700335 868201 700391 868257
rect 700477 868201 700533 868257
rect 700619 868201 700675 868257
rect 700761 868201 700817 868257
rect 700903 868201 700959 868257
rect 701045 868201 701101 868257
rect 701187 868201 701243 868257
rect 701329 868201 701385 868257
rect 701471 868201 701527 868257
rect 701613 868201 701669 868257
rect 701755 868201 701811 868257
rect 701897 868201 701953 868257
rect 73855 867957 73911 868013
rect 73997 867957 74053 868013
rect 74139 867957 74195 868013
rect 74281 867957 74337 868013
rect 74423 867957 74479 868013
rect 74565 867957 74621 868013
rect 74707 867957 74763 868013
rect 74849 867957 74905 868013
rect 74991 867957 75047 868013
rect 75133 867957 75189 868013
rect 75275 867957 75331 868013
rect 75417 867957 75473 868013
rect 75559 867957 75615 868013
rect 75701 867957 75757 868013
rect 73855 867815 73911 867871
rect 73997 867815 74053 867871
rect 74139 867815 74195 867871
rect 74281 867815 74337 867871
rect 74423 867815 74479 867871
rect 74565 867815 74621 867871
rect 74707 867815 74763 867871
rect 74849 867815 74905 867871
rect 74991 867815 75047 867871
rect 75133 867815 75189 867871
rect 75275 867815 75331 867871
rect 75417 867815 75473 867871
rect 75559 867815 75615 867871
rect 75701 867815 75757 867871
rect 73855 867673 73911 867729
rect 73997 867673 74053 867729
rect 74139 867673 74195 867729
rect 74281 867673 74337 867729
rect 74423 867673 74479 867729
rect 74565 867673 74621 867729
rect 74707 867673 74763 867729
rect 74849 867673 74905 867729
rect 74991 867673 75047 867729
rect 75133 867673 75189 867729
rect 75275 867673 75331 867729
rect 75417 867673 75473 867729
rect 75559 867673 75615 867729
rect 75701 867673 75757 867729
rect 73855 867531 73911 867587
rect 73997 867531 74053 867587
rect 74139 867531 74195 867587
rect 74281 867531 74337 867587
rect 74423 867531 74479 867587
rect 74565 867531 74621 867587
rect 74707 867531 74763 867587
rect 74849 867531 74905 867587
rect 74991 867531 75047 867587
rect 75133 867531 75189 867587
rect 75275 867531 75331 867587
rect 75417 867531 75473 867587
rect 75559 867531 75615 867587
rect 75701 867531 75757 867587
rect 73855 867389 73911 867445
rect 73997 867389 74053 867445
rect 74139 867389 74195 867445
rect 74281 867389 74337 867445
rect 74423 867389 74479 867445
rect 74565 867389 74621 867445
rect 74707 867389 74763 867445
rect 74849 867389 74905 867445
rect 74991 867389 75047 867445
rect 75133 867389 75189 867445
rect 75275 867389 75331 867445
rect 75417 867389 75473 867445
rect 75559 867389 75615 867445
rect 75701 867389 75757 867445
rect 73855 867247 73911 867303
rect 73997 867247 74053 867303
rect 74139 867247 74195 867303
rect 74281 867247 74337 867303
rect 74423 867247 74479 867303
rect 74565 867247 74621 867303
rect 74707 867247 74763 867303
rect 74849 867247 74905 867303
rect 74991 867247 75047 867303
rect 75133 867247 75189 867303
rect 75275 867247 75331 867303
rect 75417 867247 75473 867303
rect 75559 867247 75615 867303
rect 75701 867247 75757 867303
rect 73855 867105 73911 867161
rect 73997 867105 74053 867161
rect 74139 867105 74195 867161
rect 74281 867105 74337 867161
rect 74423 867105 74479 867161
rect 74565 867105 74621 867161
rect 74707 867105 74763 867161
rect 74849 867105 74905 867161
rect 74991 867105 75047 867161
rect 75133 867105 75189 867161
rect 75275 867105 75331 867161
rect 75417 867105 75473 867161
rect 75559 867105 75615 867161
rect 75701 867105 75757 867161
rect 73855 866963 73911 867019
rect 73997 866963 74053 867019
rect 74139 866963 74195 867019
rect 74281 866963 74337 867019
rect 74423 866963 74479 867019
rect 74565 866963 74621 867019
rect 74707 866963 74763 867019
rect 74849 866963 74905 867019
rect 74991 866963 75047 867019
rect 75133 866963 75189 867019
rect 75275 866963 75331 867019
rect 75417 866963 75473 867019
rect 75559 866963 75615 867019
rect 75701 866963 75757 867019
rect 73855 866821 73911 866877
rect 73997 866821 74053 866877
rect 74139 866821 74195 866877
rect 74281 866821 74337 866877
rect 74423 866821 74479 866877
rect 74565 866821 74621 866877
rect 74707 866821 74763 866877
rect 74849 866821 74905 866877
rect 74991 866821 75047 866877
rect 75133 866821 75189 866877
rect 75275 866821 75331 866877
rect 75417 866821 75473 866877
rect 75559 866821 75615 866877
rect 75701 866821 75757 866877
rect 700051 867677 700107 867733
rect 700193 867677 700249 867733
rect 700335 867677 700391 867733
rect 700477 867677 700533 867733
rect 700619 867677 700675 867733
rect 700761 867677 700817 867733
rect 700903 867677 700959 867733
rect 701045 867677 701101 867733
rect 701187 867677 701243 867733
rect 701329 867677 701385 867733
rect 701471 867677 701527 867733
rect 701613 867677 701669 867733
rect 701755 867677 701811 867733
rect 701897 867677 701953 867733
rect 700051 867535 700107 867591
rect 700193 867535 700249 867591
rect 700335 867535 700391 867591
rect 700477 867535 700533 867591
rect 700619 867535 700675 867591
rect 700761 867535 700817 867591
rect 700903 867535 700959 867591
rect 701045 867535 701101 867591
rect 701187 867535 701243 867591
rect 701329 867535 701385 867591
rect 701471 867535 701527 867591
rect 701613 867535 701669 867591
rect 701755 867535 701811 867591
rect 701897 867535 701953 867591
rect 700051 867393 700107 867449
rect 700193 867393 700249 867449
rect 700335 867393 700391 867449
rect 700477 867393 700533 867449
rect 700619 867393 700675 867449
rect 700761 867393 700817 867449
rect 700903 867393 700959 867449
rect 701045 867393 701101 867449
rect 701187 867393 701243 867449
rect 701329 867393 701385 867449
rect 701471 867393 701527 867449
rect 701613 867393 701669 867449
rect 701755 867393 701811 867449
rect 701897 867393 701953 867449
rect 700051 867251 700107 867307
rect 700193 867251 700249 867307
rect 700335 867251 700391 867307
rect 700477 867251 700533 867307
rect 700619 867251 700675 867307
rect 700761 867251 700817 867307
rect 700903 867251 700959 867307
rect 701045 867251 701101 867307
rect 701187 867251 701243 867307
rect 701329 867251 701385 867307
rect 701471 867251 701527 867307
rect 701613 867251 701669 867307
rect 701755 867251 701811 867307
rect 701897 867251 701953 867307
rect 700051 867109 700107 867165
rect 700193 867109 700249 867165
rect 700335 867109 700391 867165
rect 700477 867109 700533 867165
rect 700619 867109 700675 867165
rect 700761 867109 700817 867165
rect 700903 867109 700959 867165
rect 701045 867109 701101 867165
rect 701187 867109 701243 867165
rect 701329 867109 701385 867165
rect 701471 867109 701527 867165
rect 701613 867109 701669 867165
rect 701755 867109 701811 867165
rect 701897 867109 701953 867165
rect 700051 866967 700107 867023
rect 700193 866967 700249 867023
rect 700335 866967 700391 867023
rect 700477 866967 700533 867023
rect 700619 866967 700675 867023
rect 700761 866967 700817 867023
rect 700903 866967 700959 867023
rect 701045 866967 701101 867023
rect 701187 866967 701243 867023
rect 701329 866967 701385 867023
rect 701471 866967 701527 867023
rect 701613 866967 701669 867023
rect 701755 866967 701811 867023
rect 701897 866967 701953 867023
rect 700051 866825 700107 866881
rect 700193 866825 700249 866881
rect 700335 866825 700391 866881
rect 700477 866825 700533 866881
rect 700619 866825 700675 866881
rect 700761 866825 700817 866881
rect 700903 866825 700959 866881
rect 701045 866825 701101 866881
rect 701187 866825 701243 866881
rect 701329 866825 701385 866881
rect 701471 866825 701527 866881
rect 701613 866825 701669 866881
rect 701755 866825 701811 866881
rect 701897 866825 701953 866881
rect 700051 866683 700107 866739
rect 700193 866683 700249 866739
rect 700335 866683 700391 866739
rect 700477 866683 700533 866739
rect 700619 866683 700675 866739
rect 700761 866683 700817 866739
rect 700903 866683 700959 866739
rect 701045 866683 701101 866739
rect 701187 866683 701243 866739
rect 701329 866683 701385 866739
rect 701471 866683 701527 866739
rect 701613 866683 701669 866739
rect 701755 866683 701811 866739
rect 701897 866683 701953 866739
rect 700051 866541 700107 866597
rect 700193 866541 700249 866597
rect 700335 866541 700391 866597
rect 700477 866541 700533 866597
rect 700619 866541 700675 866597
rect 700761 866541 700817 866597
rect 700903 866541 700959 866597
rect 701045 866541 701101 866597
rect 701187 866541 701243 866597
rect 701329 866541 701385 866597
rect 701471 866541 701527 866597
rect 701613 866541 701669 866597
rect 701755 866541 701811 866597
rect 701897 866541 701953 866597
rect 700051 866399 700107 866455
rect 700193 866399 700249 866455
rect 700335 866399 700391 866455
rect 700477 866399 700533 866455
rect 700619 866399 700675 866455
rect 700761 866399 700817 866455
rect 700903 866399 700959 866455
rect 701045 866399 701101 866455
rect 701187 866399 701243 866455
rect 701329 866399 701385 866455
rect 701471 866399 701527 866455
rect 701613 866399 701669 866455
rect 701755 866399 701811 866455
rect 701897 866399 701953 866455
rect 700051 866257 700107 866313
rect 700193 866257 700249 866313
rect 700335 866257 700391 866313
rect 700477 866257 700533 866313
rect 700619 866257 700675 866313
rect 700761 866257 700817 866313
rect 700903 866257 700959 866313
rect 701045 866257 701101 866313
rect 701187 866257 701243 866313
rect 701329 866257 701385 866313
rect 701471 866257 701527 866313
rect 701613 866257 701669 866313
rect 701755 866257 701811 866313
rect 701897 866257 701953 866313
rect 73866 866038 73922 866094
rect 74008 866038 74064 866094
rect 74150 866038 74206 866094
rect 74292 866038 74348 866094
rect 74434 866038 74490 866094
rect 74576 866038 74632 866094
rect 74718 866038 74774 866094
rect 74860 866038 74916 866094
rect 75002 866038 75058 866094
rect 75144 866038 75200 866094
rect 75286 866038 75342 866094
rect 75428 866038 75484 866094
rect 75570 866038 75626 866094
rect 75712 866038 75768 866094
rect 73866 865896 73922 865952
rect 74008 865896 74064 865952
rect 74150 865896 74206 865952
rect 74292 865896 74348 865952
rect 74434 865896 74490 865952
rect 74576 865896 74632 865952
rect 74718 865896 74774 865952
rect 74860 865896 74916 865952
rect 75002 865896 75058 865952
rect 75144 865896 75200 865952
rect 75286 865896 75342 865952
rect 75428 865896 75484 865952
rect 75570 865896 75626 865952
rect 75712 865896 75768 865952
rect 73866 865754 73922 865810
rect 74008 865754 74064 865810
rect 74150 865754 74206 865810
rect 74292 865754 74348 865810
rect 74434 865754 74490 865810
rect 74576 865754 74632 865810
rect 74718 865754 74774 865810
rect 74860 865754 74916 865810
rect 75002 865754 75058 865810
rect 75144 865754 75200 865810
rect 75286 865754 75342 865810
rect 75428 865754 75484 865810
rect 75570 865754 75626 865810
rect 75712 865754 75768 865810
rect 700051 866115 700107 866171
rect 700193 866115 700249 866171
rect 700335 866115 700391 866171
rect 700477 866115 700533 866171
rect 700619 866115 700675 866171
rect 700761 866115 700817 866171
rect 700903 866115 700959 866171
rect 701045 866115 701101 866171
rect 701187 866115 701243 866171
rect 701329 866115 701385 866171
rect 701471 866115 701527 866171
rect 701613 866115 701669 866171
rect 701755 866115 701811 866171
rect 701897 866115 701953 866171
rect 700051 865973 700107 866029
rect 700193 865973 700249 866029
rect 700335 865973 700391 866029
rect 700477 865973 700533 866029
rect 700619 865973 700675 866029
rect 700761 865973 700817 866029
rect 700903 865973 700959 866029
rect 701045 865973 701101 866029
rect 701187 865973 701243 866029
rect 701329 865973 701385 866029
rect 701471 865973 701527 866029
rect 701613 865973 701669 866029
rect 701755 865973 701811 866029
rect 701897 865973 701953 866029
rect 700051 865831 700107 865887
rect 700193 865831 700249 865887
rect 700335 865831 700391 865887
rect 700477 865831 700533 865887
rect 700619 865831 700675 865887
rect 700761 865831 700817 865887
rect 700903 865831 700959 865887
rect 701045 865831 701101 865887
rect 701187 865831 701243 865887
rect 701329 865831 701385 865887
rect 701471 865831 701527 865887
rect 701613 865831 701669 865887
rect 701755 865831 701811 865887
rect 701897 865831 701953 865887
rect 73866 865612 73922 865668
rect 74008 865612 74064 865668
rect 74150 865612 74206 865668
rect 74292 865612 74348 865668
rect 74434 865612 74490 865668
rect 74576 865612 74632 865668
rect 74718 865612 74774 865668
rect 74860 865612 74916 865668
rect 75002 865612 75058 865668
rect 75144 865612 75200 865668
rect 75286 865612 75342 865668
rect 75428 865612 75484 865668
rect 75570 865612 75626 865668
rect 75712 865612 75768 865668
rect 73866 865470 73922 865526
rect 74008 865470 74064 865526
rect 74150 865470 74206 865526
rect 74292 865470 74348 865526
rect 74434 865470 74490 865526
rect 74576 865470 74632 865526
rect 74718 865470 74774 865526
rect 74860 865470 74916 865526
rect 75002 865470 75058 865526
rect 75144 865470 75200 865526
rect 75286 865470 75342 865526
rect 75428 865470 75484 865526
rect 75570 865470 75626 865526
rect 75712 865470 75768 865526
rect 73866 865328 73922 865384
rect 74008 865328 74064 865384
rect 74150 865328 74206 865384
rect 74292 865328 74348 865384
rect 74434 865328 74490 865384
rect 74576 865328 74632 865384
rect 74718 865328 74774 865384
rect 74860 865328 74916 865384
rect 75002 865328 75058 865384
rect 75144 865328 75200 865384
rect 75286 865328 75342 865384
rect 75428 865328 75484 865384
rect 75570 865328 75626 865384
rect 75712 865328 75768 865384
rect 73866 865186 73922 865242
rect 74008 865186 74064 865242
rect 74150 865186 74206 865242
rect 74292 865186 74348 865242
rect 74434 865186 74490 865242
rect 74576 865186 74632 865242
rect 74718 865186 74774 865242
rect 74860 865186 74916 865242
rect 75002 865186 75058 865242
rect 75144 865186 75200 865242
rect 75286 865186 75342 865242
rect 75428 865186 75484 865242
rect 75570 865186 75626 865242
rect 75712 865186 75768 865242
rect 73866 865044 73922 865100
rect 74008 865044 74064 865100
rect 74150 865044 74206 865100
rect 74292 865044 74348 865100
rect 74434 865044 74490 865100
rect 74576 865044 74632 865100
rect 74718 865044 74774 865100
rect 74860 865044 74916 865100
rect 75002 865044 75058 865100
rect 75144 865044 75200 865100
rect 75286 865044 75342 865100
rect 75428 865044 75484 865100
rect 75570 865044 75626 865100
rect 75712 865044 75768 865100
rect 73866 864902 73922 864958
rect 74008 864902 74064 864958
rect 74150 864902 74206 864958
rect 74292 864902 74348 864958
rect 74434 864902 74490 864958
rect 74576 864902 74632 864958
rect 74718 864902 74774 864958
rect 74860 864902 74916 864958
rect 75002 864902 75058 864958
rect 75144 864902 75200 864958
rect 75286 864902 75342 864958
rect 75428 864902 75484 864958
rect 75570 864902 75626 864958
rect 75712 864902 75768 864958
rect 73866 864760 73922 864816
rect 74008 864760 74064 864816
rect 74150 864760 74206 864816
rect 74292 864760 74348 864816
rect 74434 864760 74490 864816
rect 74576 864760 74632 864816
rect 74718 864760 74774 864816
rect 74860 864760 74916 864816
rect 75002 864760 75058 864816
rect 75144 864760 75200 864816
rect 75286 864760 75342 864816
rect 75428 864760 75484 864816
rect 75570 864760 75626 864816
rect 75712 864760 75768 864816
rect 73866 864618 73922 864674
rect 74008 864618 74064 864674
rect 74150 864618 74206 864674
rect 74292 864618 74348 864674
rect 74434 864618 74490 864674
rect 74576 864618 74632 864674
rect 74718 864618 74774 864674
rect 74860 864618 74916 864674
rect 75002 864618 75058 864674
rect 75144 864618 75200 864674
rect 75286 864618 75342 864674
rect 75428 864618 75484 864674
rect 75570 864618 75626 864674
rect 75712 864618 75768 864674
rect 73866 864476 73922 864532
rect 74008 864476 74064 864532
rect 74150 864476 74206 864532
rect 74292 864476 74348 864532
rect 74434 864476 74490 864532
rect 74576 864476 74632 864532
rect 74718 864476 74774 864532
rect 74860 864476 74916 864532
rect 75002 864476 75058 864532
rect 75144 864476 75200 864532
rect 75286 864476 75342 864532
rect 75428 864476 75484 864532
rect 75570 864476 75626 864532
rect 75712 864476 75768 864532
rect 73866 864334 73922 864390
rect 74008 864334 74064 864390
rect 74150 864334 74206 864390
rect 74292 864334 74348 864390
rect 74434 864334 74490 864390
rect 74576 864334 74632 864390
rect 74718 864334 74774 864390
rect 74860 864334 74916 864390
rect 75002 864334 75058 864390
rect 75144 864334 75200 864390
rect 75286 864334 75342 864390
rect 75428 864334 75484 864390
rect 75570 864334 75626 864390
rect 75712 864334 75768 864390
rect 700040 865054 700096 865110
rect 700182 865054 700238 865110
rect 700324 865054 700380 865110
rect 700466 865054 700522 865110
rect 700608 865054 700664 865110
rect 700750 865054 700806 865110
rect 700892 865054 700948 865110
rect 701034 865054 701090 865110
rect 701176 865054 701232 865110
rect 701318 865054 701374 865110
rect 701460 865054 701516 865110
rect 701602 865054 701658 865110
rect 701744 865054 701800 865110
rect 701886 865054 701942 865110
rect 700040 864912 700096 864968
rect 700182 864912 700238 864968
rect 700324 864912 700380 864968
rect 700466 864912 700522 864968
rect 700608 864912 700664 864968
rect 700750 864912 700806 864968
rect 700892 864912 700948 864968
rect 701034 864912 701090 864968
rect 701176 864912 701232 864968
rect 701318 864912 701374 864968
rect 701460 864912 701516 864968
rect 701602 864912 701658 864968
rect 701744 864912 701800 864968
rect 701886 864912 701942 864968
rect 700040 864770 700096 864826
rect 700182 864770 700238 864826
rect 700324 864770 700380 864826
rect 700466 864770 700522 864826
rect 700608 864770 700664 864826
rect 700750 864770 700806 864826
rect 700892 864770 700948 864826
rect 701034 864770 701090 864826
rect 701176 864770 701232 864826
rect 701318 864770 701374 864826
rect 701460 864770 701516 864826
rect 701602 864770 701658 864826
rect 701744 864770 701800 864826
rect 701886 864770 701942 864826
rect 700040 864628 700096 864684
rect 700182 864628 700238 864684
rect 700324 864628 700380 864684
rect 700466 864628 700522 864684
rect 700608 864628 700664 864684
rect 700750 864628 700806 864684
rect 700892 864628 700948 864684
rect 701034 864628 701090 864684
rect 701176 864628 701232 864684
rect 701318 864628 701374 864684
rect 701460 864628 701516 864684
rect 701602 864628 701658 864684
rect 701744 864628 701800 864684
rect 701886 864628 701942 864684
rect 700040 864486 700096 864542
rect 700182 864486 700238 864542
rect 700324 864486 700380 864542
rect 700466 864486 700522 864542
rect 700608 864486 700664 864542
rect 700750 864486 700806 864542
rect 700892 864486 700948 864542
rect 701034 864486 701090 864542
rect 701176 864486 701232 864542
rect 701318 864486 701374 864542
rect 701460 864486 701516 864542
rect 701602 864486 701658 864542
rect 701744 864486 701800 864542
rect 701886 864486 701942 864542
rect 700040 864344 700096 864400
rect 700182 864344 700238 864400
rect 700324 864344 700380 864400
rect 700466 864344 700522 864400
rect 700608 864344 700664 864400
rect 700750 864344 700806 864400
rect 700892 864344 700948 864400
rect 701034 864344 701090 864400
rect 701176 864344 701232 864400
rect 701318 864344 701374 864400
rect 701460 864344 701516 864400
rect 701602 864344 701658 864400
rect 701744 864344 701800 864400
rect 701886 864344 701942 864400
rect 700040 864202 700096 864258
rect 700182 864202 700238 864258
rect 700324 864202 700380 864258
rect 700466 864202 700522 864258
rect 700608 864202 700664 864258
rect 700750 864202 700806 864258
rect 700892 864202 700948 864258
rect 701034 864202 701090 864258
rect 701176 864202 701232 864258
rect 701318 864202 701374 864258
rect 701460 864202 701516 864258
rect 701602 864202 701658 864258
rect 701744 864202 701800 864258
rect 701886 864202 701942 864258
rect 700040 864060 700096 864116
rect 700182 864060 700238 864116
rect 700324 864060 700380 864116
rect 700466 864060 700522 864116
rect 700608 864060 700664 864116
rect 700750 864060 700806 864116
rect 700892 864060 700948 864116
rect 701034 864060 701090 864116
rect 701176 864060 701232 864116
rect 701318 864060 701374 864116
rect 701460 864060 701516 864116
rect 701602 864060 701658 864116
rect 701744 864060 701800 864116
rect 701886 864060 701942 864116
rect 700040 863918 700096 863974
rect 700182 863918 700238 863974
rect 700324 863918 700380 863974
rect 700466 863918 700522 863974
rect 700608 863918 700664 863974
rect 700750 863918 700806 863974
rect 700892 863918 700948 863974
rect 701034 863918 701090 863974
rect 701176 863918 701232 863974
rect 701318 863918 701374 863974
rect 701460 863918 701516 863974
rect 701602 863918 701658 863974
rect 701744 863918 701800 863974
rect 701886 863918 701942 863974
rect 700040 863776 700096 863832
rect 700182 863776 700238 863832
rect 700324 863776 700380 863832
rect 700466 863776 700522 863832
rect 700608 863776 700664 863832
rect 700750 863776 700806 863832
rect 700892 863776 700948 863832
rect 701034 863776 701090 863832
rect 701176 863776 701232 863832
rect 701318 863776 701374 863832
rect 701460 863776 701516 863832
rect 701602 863776 701658 863832
rect 701744 863776 701800 863832
rect 701886 863776 701942 863832
rect 700040 863634 700096 863690
rect 700182 863634 700238 863690
rect 700324 863634 700380 863690
rect 700466 863634 700522 863690
rect 700608 863634 700664 863690
rect 700750 863634 700806 863690
rect 700892 863634 700948 863690
rect 701034 863634 701090 863690
rect 701176 863634 701232 863690
rect 701318 863634 701374 863690
rect 701460 863634 701516 863690
rect 701602 863634 701658 863690
rect 701744 863634 701800 863690
rect 701886 863634 701942 863690
rect 700040 863492 700096 863548
rect 700182 863492 700238 863548
rect 700324 863492 700380 863548
rect 700466 863492 700522 863548
rect 700608 863492 700664 863548
rect 700750 863492 700806 863548
rect 700892 863492 700948 863548
rect 701034 863492 701090 863548
rect 701176 863492 701232 863548
rect 701318 863492 701374 863548
rect 701460 863492 701516 863548
rect 701602 863492 701658 863548
rect 701744 863492 701800 863548
rect 701886 863492 701942 863548
rect 700040 863350 700096 863406
rect 700182 863350 700238 863406
rect 700324 863350 700380 863406
rect 700466 863350 700522 863406
rect 700608 863350 700664 863406
rect 700750 863350 700806 863406
rect 700892 863350 700948 863406
rect 701034 863350 701090 863406
rect 701176 863350 701232 863406
rect 701318 863350 701374 863406
rect 701460 863350 701516 863406
rect 701602 863350 701658 863406
rect 701744 863350 701800 863406
rect 701886 863350 701942 863406
rect 73866 837594 73922 837650
rect 74008 837594 74064 837650
rect 74150 837594 74206 837650
rect 74292 837594 74348 837650
rect 74434 837594 74490 837650
rect 74576 837594 74632 837650
rect 74718 837594 74774 837650
rect 74860 837594 74916 837650
rect 75002 837594 75058 837650
rect 75144 837594 75200 837650
rect 75286 837594 75342 837650
rect 73866 837452 73922 837508
rect 74008 837452 74064 837508
rect 74150 837452 74206 837508
rect 74292 837452 74348 837508
rect 74434 837452 74490 837508
rect 74576 837452 74632 837508
rect 74718 837452 74774 837508
rect 74860 837452 74916 837508
rect 75002 837452 75058 837508
rect 75144 837452 75200 837508
rect 75286 837452 75342 837508
rect 73866 837310 73922 837366
rect 74008 837310 74064 837366
rect 74150 837310 74206 837366
rect 74292 837310 74348 837366
rect 74434 837310 74490 837366
rect 74576 837310 74632 837366
rect 74718 837310 74774 837366
rect 74860 837310 74916 837366
rect 75002 837310 75058 837366
rect 75144 837310 75200 837366
rect 75286 837310 75342 837366
rect 73866 837168 73922 837224
rect 74008 837168 74064 837224
rect 74150 837168 74206 837224
rect 74292 837168 74348 837224
rect 74434 837168 74490 837224
rect 74576 837168 74632 837224
rect 74718 837168 74774 837224
rect 74860 837168 74916 837224
rect 75002 837168 75058 837224
rect 75144 837168 75200 837224
rect 75286 837168 75342 837224
rect 73866 837026 73922 837082
rect 74008 837026 74064 837082
rect 74150 837026 74206 837082
rect 74292 837026 74348 837082
rect 74434 837026 74490 837082
rect 74576 837026 74632 837082
rect 74718 837026 74774 837082
rect 74860 837026 74916 837082
rect 75002 837026 75058 837082
rect 75144 837026 75200 837082
rect 75286 837026 75342 837082
rect 73866 836884 73922 836940
rect 74008 836884 74064 836940
rect 74150 836884 74206 836940
rect 74292 836884 74348 836940
rect 74434 836884 74490 836940
rect 74576 836884 74632 836940
rect 74718 836884 74774 836940
rect 74860 836884 74916 836940
rect 75002 836884 75058 836940
rect 75144 836884 75200 836940
rect 75286 836884 75342 836940
rect 73866 836742 73922 836798
rect 74008 836742 74064 836798
rect 74150 836742 74206 836798
rect 74292 836742 74348 836798
rect 74434 836742 74490 836798
rect 74576 836742 74632 836798
rect 74718 836742 74774 836798
rect 74860 836742 74916 836798
rect 75002 836742 75058 836798
rect 75144 836742 75200 836798
rect 75286 836742 75342 836798
rect 73866 836600 73922 836656
rect 74008 836600 74064 836656
rect 74150 836600 74206 836656
rect 74292 836600 74348 836656
rect 74434 836600 74490 836656
rect 74576 836600 74632 836656
rect 74718 836600 74774 836656
rect 74860 836600 74916 836656
rect 75002 836600 75058 836656
rect 75144 836600 75200 836656
rect 75286 836600 75342 836656
rect 73866 836458 73922 836514
rect 74008 836458 74064 836514
rect 74150 836458 74206 836514
rect 74292 836458 74348 836514
rect 74434 836458 74490 836514
rect 74576 836458 74632 836514
rect 74718 836458 74774 836514
rect 74860 836458 74916 836514
rect 75002 836458 75058 836514
rect 75144 836458 75200 836514
rect 75286 836458 75342 836514
rect 73866 836316 73922 836372
rect 74008 836316 74064 836372
rect 74150 836316 74206 836372
rect 74292 836316 74348 836372
rect 74434 836316 74490 836372
rect 74576 836316 74632 836372
rect 74718 836316 74774 836372
rect 74860 836316 74916 836372
rect 75002 836316 75058 836372
rect 75144 836316 75200 836372
rect 75286 836316 75342 836372
rect 73866 836174 73922 836230
rect 74008 836174 74064 836230
rect 74150 836174 74206 836230
rect 74292 836174 74348 836230
rect 74434 836174 74490 836230
rect 74576 836174 74632 836230
rect 74718 836174 74774 836230
rect 74860 836174 74916 836230
rect 75002 836174 75058 836230
rect 75144 836174 75200 836230
rect 75286 836174 75342 836230
rect 73866 836032 73922 836088
rect 74008 836032 74064 836088
rect 74150 836032 74206 836088
rect 74292 836032 74348 836088
rect 74434 836032 74490 836088
rect 74576 836032 74632 836088
rect 74718 836032 74774 836088
rect 74860 836032 74916 836088
rect 75002 836032 75058 836088
rect 75144 836032 75200 836088
rect 75286 836032 75342 836088
rect 73866 835890 73922 835946
rect 74008 835890 74064 835946
rect 74150 835890 74206 835946
rect 74292 835890 74348 835946
rect 74434 835890 74490 835946
rect 74576 835890 74632 835946
rect 74718 835890 74774 835946
rect 74860 835890 74916 835946
rect 75002 835890 75058 835946
rect 75144 835890 75200 835946
rect 75286 835890 75342 835946
rect 73855 835113 73911 835169
rect 73997 835113 74053 835169
rect 74139 835113 74195 835169
rect 74281 835113 74337 835169
rect 74423 835113 74479 835169
rect 74565 835113 74621 835169
rect 74707 835113 74763 835169
rect 74849 835113 74905 835169
rect 74991 835113 75047 835169
rect 75133 835113 75189 835169
rect 75275 835113 75331 835169
rect 73855 834971 73911 835027
rect 73997 834971 74053 835027
rect 74139 834971 74195 835027
rect 74281 834971 74337 835027
rect 74423 834971 74479 835027
rect 74565 834971 74621 835027
rect 74707 834971 74763 835027
rect 74849 834971 74905 835027
rect 74991 834971 75047 835027
rect 75133 834971 75189 835027
rect 75275 834971 75331 835027
rect 73855 834829 73911 834885
rect 73997 834829 74053 834885
rect 74139 834829 74195 834885
rect 74281 834829 74337 834885
rect 74423 834829 74479 834885
rect 74565 834829 74621 834885
rect 74707 834829 74763 834885
rect 74849 834829 74905 834885
rect 74991 834829 75047 834885
rect 75133 834829 75189 834885
rect 75275 834829 75331 834885
rect 73855 834687 73911 834743
rect 73997 834687 74053 834743
rect 74139 834687 74195 834743
rect 74281 834687 74337 834743
rect 74423 834687 74479 834743
rect 74565 834687 74621 834743
rect 74707 834687 74763 834743
rect 74849 834687 74905 834743
rect 74991 834687 75047 834743
rect 75133 834687 75189 834743
rect 75275 834687 75331 834743
rect 73855 834545 73911 834601
rect 73997 834545 74053 834601
rect 74139 834545 74195 834601
rect 74281 834545 74337 834601
rect 74423 834545 74479 834601
rect 74565 834545 74621 834601
rect 74707 834545 74763 834601
rect 74849 834545 74905 834601
rect 74991 834545 75047 834601
rect 75133 834545 75189 834601
rect 75275 834545 75331 834601
rect 73855 834403 73911 834459
rect 73997 834403 74053 834459
rect 74139 834403 74195 834459
rect 74281 834403 74337 834459
rect 74423 834403 74479 834459
rect 74565 834403 74621 834459
rect 74707 834403 74763 834459
rect 74849 834403 74905 834459
rect 74991 834403 75047 834459
rect 75133 834403 75189 834459
rect 75275 834403 75331 834459
rect 73855 834261 73911 834317
rect 73997 834261 74053 834317
rect 74139 834261 74195 834317
rect 74281 834261 74337 834317
rect 74423 834261 74479 834317
rect 74565 834261 74621 834317
rect 74707 834261 74763 834317
rect 74849 834261 74905 834317
rect 74991 834261 75047 834317
rect 75133 834261 75189 834317
rect 75275 834261 75331 834317
rect 73855 834119 73911 834175
rect 73997 834119 74053 834175
rect 74139 834119 74195 834175
rect 74281 834119 74337 834175
rect 74423 834119 74479 834175
rect 74565 834119 74621 834175
rect 74707 834119 74763 834175
rect 74849 834119 74905 834175
rect 74991 834119 75047 834175
rect 75133 834119 75189 834175
rect 75275 834119 75331 834175
rect 73855 833977 73911 834033
rect 73997 833977 74053 834033
rect 74139 833977 74195 834033
rect 74281 833977 74337 834033
rect 74423 833977 74479 834033
rect 74565 833977 74621 834033
rect 74707 833977 74763 834033
rect 74849 833977 74905 834033
rect 74991 833977 75047 834033
rect 75133 833977 75189 834033
rect 75275 833977 75331 834033
rect 73855 833835 73911 833891
rect 73997 833835 74053 833891
rect 74139 833835 74195 833891
rect 74281 833835 74337 833891
rect 74423 833835 74479 833891
rect 74565 833835 74621 833891
rect 74707 833835 74763 833891
rect 74849 833835 74905 833891
rect 74991 833835 75047 833891
rect 75133 833835 75189 833891
rect 75275 833835 75331 833891
rect 73855 833693 73911 833749
rect 73997 833693 74053 833749
rect 74139 833693 74195 833749
rect 74281 833693 74337 833749
rect 74423 833693 74479 833749
rect 74565 833693 74621 833749
rect 74707 833693 74763 833749
rect 74849 833693 74905 833749
rect 74991 833693 75047 833749
rect 75133 833693 75189 833749
rect 75275 833693 75331 833749
rect 73855 833551 73911 833607
rect 73997 833551 74053 833607
rect 74139 833551 74195 833607
rect 74281 833551 74337 833607
rect 74423 833551 74479 833607
rect 74565 833551 74621 833607
rect 74707 833551 74763 833607
rect 74849 833551 74905 833607
rect 74991 833551 75047 833607
rect 75133 833551 75189 833607
rect 75275 833551 75331 833607
rect 73855 833409 73911 833465
rect 73997 833409 74053 833465
rect 74139 833409 74195 833465
rect 74281 833409 74337 833465
rect 74423 833409 74479 833465
rect 74565 833409 74621 833465
rect 74707 833409 74763 833465
rect 74849 833409 74905 833465
rect 74991 833409 75047 833465
rect 75133 833409 75189 833465
rect 75275 833409 75331 833465
rect 73855 833267 73911 833323
rect 73997 833267 74053 833323
rect 74139 833267 74195 833323
rect 74281 833267 74337 833323
rect 74423 833267 74479 833323
rect 74565 833267 74621 833323
rect 74707 833267 74763 833323
rect 74849 833267 74905 833323
rect 74991 833267 75047 833323
rect 75133 833267 75189 833323
rect 75275 833267 75331 833323
rect 73855 832743 73911 832799
rect 73997 832743 74053 832799
rect 74139 832743 74195 832799
rect 74281 832743 74337 832799
rect 74423 832743 74479 832799
rect 74565 832743 74621 832799
rect 74707 832743 74763 832799
rect 74849 832743 74905 832799
rect 74991 832743 75047 832799
rect 75133 832743 75189 832799
rect 75275 832743 75331 832799
rect 73855 832601 73911 832657
rect 73997 832601 74053 832657
rect 74139 832601 74195 832657
rect 74281 832601 74337 832657
rect 74423 832601 74479 832657
rect 74565 832601 74621 832657
rect 74707 832601 74763 832657
rect 74849 832601 74905 832657
rect 74991 832601 75047 832657
rect 75133 832601 75189 832657
rect 75275 832601 75331 832657
rect 73855 832459 73911 832515
rect 73997 832459 74053 832515
rect 74139 832459 74195 832515
rect 74281 832459 74337 832515
rect 74423 832459 74479 832515
rect 74565 832459 74621 832515
rect 74707 832459 74763 832515
rect 74849 832459 74905 832515
rect 74991 832459 75047 832515
rect 75133 832459 75189 832515
rect 75275 832459 75331 832515
rect 73855 832317 73911 832373
rect 73997 832317 74053 832373
rect 74139 832317 74195 832373
rect 74281 832317 74337 832373
rect 74423 832317 74479 832373
rect 74565 832317 74621 832373
rect 74707 832317 74763 832373
rect 74849 832317 74905 832373
rect 74991 832317 75047 832373
rect 75133 832317 75189 832373
rect 75275 832317 75331 832373
rect 73855 832175 73911 832231
rect 73997 832175 74053 832231
rect 74139 832175 74195 832231
rect 74281 832175 74337 832231
rect 74423 832175 74479 832231
rect 74565 832175 74621 832231
rect 74707 832175 74763 832231
rect 74849 832175 74905 832231
rect 74991 832175 75047 832231
rect 75133 832175 75189 832231
rect 75275 832175 75331 832231
rect 73855 832033 73911 832089
rect 73997 832033 74053 832089
rect 74139 832033 74195 832089
rect 74281 832033 74337 832089
rect 74423 832033 74479 832089
rect 74565 832033 74621 832089
rect 74707 832033 74763 832089
rect 74849 832033 74905 832089
rect 74991 832033 75047 832089
rect 75133 832033 75189 832089
rect 75275 832033 75331 832089
rect 73855 831891 73911 831947
rect 73997 831891 74053 831947
rect 74139 831891 74195 831947
rect 74281 831891 74337 831947
rect 74423 831891 74479 831947
rect 74565 831891 74621 831947
rect 74707 831891 74763 831947
rect 74849 831891 74905 831947
rect 74991 831891 75047 831947
rect 75133 831891 75189 831947
rect 75275 831891 75331 831947
rect 73855 831749 73911 831805
rect 73997 831749 74053 831805
rect 74139 831749 74195 831805
rect 74281 831749 74337 831805
rect 74423 831749 74479 831805
rect 74565 831749 74621 831805
rect 74707 831749 74763 831805
rect 74849 831749 74905 831805
rect 74991 831749 75047 831805
rect 75133 831749 75189 831805
rect 75275 831749 75331 831805
rect 73855 831607 73911 831663
rect 73997 831607 74053 831663
rect 74139 831607 74195 831663
rect 74281 831607 74337 831663
rect 74423 831607 74479 831663
rect 74565 831607 74621 831663
rect 74707 831607 74763 831663
rect 74849 831607 74905 831663
rect 74991 831607 75047 831663
rect 75133 831607 75189 831663
rect 75275 831607 75331 831663
rect 73855 831465 73911 831521
rect 73997 831465 74053 831521
rect 74139 831465 74195 831521
rect 74281 831465 74337 831521
rect 74423 831465 74479 831521
rect 74565 831465 74621 831521
rect 74707 831465 74763 831521
rect 74849 831465 74905 831521
rect 74991 831465 75047 831521
rect 75133 831465 75189 831521
rect 75275 831465 75331 831521
rect 73855 831323 73911 831379
rect 73997 831323 74053 831379
rect 74139 831323 74195 831379
rect 74281 831323 74337 831379
rect 74423 831323 74479 831379
rect 74565 831323 74621 831379
rect 74707 831323 74763 831379
rect 74849 831323 74905 831379
rect 74991 831323 75047 831379
rect 75133 831323 75189 831379
rect 75275 831323 75331 831379
rect 73855 831181 73911 831237
rect 73997 831181 74053 831237
rect 74139 831181 74195 831237
rect 74281 831181 74337 831237
rect 74423 831181 74479 831237
rect 74565 831181 74621 831237
rect 74707 831181 74763 831237
rect 74849 831181 74905 831237
rect 74991 831181 75047 831237
rect 75133 831181 75189 831237
rect 75275 831181 75331 831237
rect 73855 831039 73911 831095
rect 73997 831039 74053 831095
rect 74139 831039 74195 831095
rect 74281 831039 74337 831095
rect 74423 831039 74479 831095
rect 74565 831039 74621 831095
rect 74707 831039 74763 831095
rect 74849 831039 74905 831095
rect 74991 831039 75047 831095
rect 75133 831039 75189 831095
rect 75275 831039 75331 831095
rect 73855 830897 73911 830953
rect 73997 830897 74053 830953
rect 74139 830897 74195 830953
rect 74281 830897 74337 830953
rect 74423 830897 74479 830953
rect 74565 830897 74621 830953
rect 74707 830897 74763 830953
rect 74849 830897 74905 830953
rect 74991 830897 75047 830953
rect 75133 830897 75189 830953
rect 75275 830897 75331 830953
rect 73855 830037 73911 830093
rect 73997 830037 74053 830093
rect 74139 830037 74195 830093
rect 74281 830037 74337 830093
rect 74423 830037 74479 830093
rect 74565 830037 74621 830093
rect 74707 830037 74763 830093
rect 74849 830037 74905 830093
rect 74991 830037 75047 830093
rect 75133 830037 75189 830093
rect 75275 830037 75331 830093
rect 73855 829895 73911 829951
rect 73997 829895 74053 829951
rect 74139 829895 74195 829951
rect 74281 829895 74337 829951
rect 74423 829895 74479 829951
rect 74565 829895 74621 829951
rect 74707 829895 74763 829951
rect 74849 829895 74905 829951
rect 74991 829895 75047 829951
rect 75133 829895 75189 829951
rect 75275 829895 75331 829951
rect 73855 829753 73911 829809
rect 73997 829753 74053 829809
rect 74139 829753 74195 829809
rect 74281 829753 74337 829809
rect 74423 829753 74479 829809
rect 74565 829753 74621 829809
rect 74707 829753 74763 829809
rect 74849 829753 74905 829809
rect 74991 829753 75047 829809
rect 75133 829753 75189 829809
rect 75275 829753 75331 829809
rect 73855 829611 73911 829667
rect 73997 829611 74053 829667
rect 74139 829611 74195 829667
rect 74281 829611 74337 829667
rect 74423 829611 74479 829667
rect 74565 829611 74621 829667
rect 74707 829611 74763 829667
rect 74849 829611 74905 829667
rect 74991 829611 75047 829667
rect 75133 829611 75189 829667
rect 75275 829611 75331 829667
rect 73855 829469 73911 829525
rect 73997 829469 74053 829525
rect 74139 829469 74195 829525
rect 74281 829469 74337 829525
rect 74423 829469 74479 829525
rect 74565 829469 74621 829525
rect 74707 829469 74763 829525
rect 74849 829469 74905 829525
rect 74991 829469 75047 829525
rect 75133 829469 75189 829525
rect 75275 829469 75331 829525
rect 73855 829327 73911 829383
rect 73997 829327 74053 829383
rect 74139 829327 74195 829383
rect 74281 829327 74337 829383
rect 74423 829327 74479 829383
rect 74565 829327 74621 829383
rect 74707 829327 74763 829383
rect 74849 829327 74905 829383
rect 74991 829327 75047 829383
rect 75133 829327 75189 829383
rect 75275 829327 75331 829383
rect 73855 829185 73911 829241
rect 73997 829185 74053 829241
rect 74139 829185 74195 829241
rect 74281 829185 74337 829241
rect 74423 829185 74479 829241
rect 74565 829185 74621 829241
rect 74707 829185 74763 829241
rect 74849 829185 74905 829241
rect 74991 829185 75047 829241
rect 75133 829185 75189 829241
rect 75275 829185 75331 829241
rect 73855 829043 73911 829099
rect 73997 829043 74053 829099
rect 74139 829043 74195 829099
rect 74281 829043 74337 829099
rect 74423 829043 74479 829099
rect 74565 829043 74621 829099
rect 74707 829043 74763 829099
rect 74849 829043 74905 829099
rect 74991 829043 75047 829099
rect 75133 829043 75189 829099
rect 75275 829043 75331 829099
rect 73855 828901 73911 828957
rect 73997 828901 74053 828957
rect 74139 828901 74195 828957
rect 74281 828901 74337 828957
rect 74423 828901 74479 828957
rect 74565 828901 74621 828957
rect 74707 828901 74763 828957
rect 74849 828901 74905 828957
rect 74991 828901 75047 828957
rect 75133 828901 75189 828957
rect 75275 828901 75331 828957
rect 73855 828759 73911 828815
rect 73997 828759 74053 828815
rect 74139 828759 74195 828815
rect 74281 828759 74337 828815
rect 74423 828759 74479 828815
rect 74565 828759 74621 828815
rect 74707 828759 74763 828815
rect 74849 828759 74905 828815
rect 74991 828759 75047 828815
rect 75133 828759 75189 828815
rect 75275 828759 75331 828815
rect 73855 828617 73911 828673
rect 73997 828617 74053 828673
rect 74139 828617 74195 828673
rect 74281 828617 74337 828673
rect 74423 828617 74479 828673
rect 74565 828617 74621 828673
rect 74707 828617 74763 828673
rect 74849 828617 74905 828673
rect 74991 828617 75047 828673
rect 75133 828617 75189 828673
rect 75275 828617 75331 828673
rect 73855 828475 73911 828531
rect 73997 828475 74053 828531
rect 74139 828475 74195 828531
rect 74281 828475 74337 828531
rect 74423 828475 74479 828531
rect 74565 828475 74621 828531
rect 74707 828475 74763 828531
rect 74849 828475 74905 828531
rect 74991 828475 75047 828531
rect 75133 828475 75189 828531
rect 75275 828475 75331 828531
rect 73855 828333 73911 828389
rect 73997 828333 74053 828389
rect 74139 828333 74195 828389
rect 74281 828333 74337 828389
rect 74423 828333 74479 828389
rect 74565 828333 74621 828389
rect 74707 828333 74763 828389
rect 74849 828333 74905 828389
rect 74991 828333 75047 828389
rect 75133 828333 75189 828389
rect 75275 828333 75331 828389
rect 73855 828191 73911 828247
rect 73997 828191 74053 828247
rect 74139 828191 74195 828247
rect 74281 828191 74337 828247
rect 74423 828191 74479 828247
rect 74565 828191 74621 828247
rect 74707 828191 74763 828247
rect 74849 828191 74905 828247
rect 74991 828191 75047 828247
rect 75133 828191 75189 828247
rect 75275 828191 75331 828247
rect 73855 827667 73911 827723
rect 73997 827667 74053 827723
rect 74139 827667 74195 827723
rect 74281 827667 74337 827723
rect 74423 827667 74479 827723
rect 74565 827667 74621 827723
rect 74707 827667 74763 827723
rect 74849 827667 74905 827723
rect 74991 827667 75047 827723
rect 75133 827667 75189 827723
rect 75275 827667 75331 827723
rect 73855 827525 73911 827581
rect 73997 827525 74053 827581
rect 74139 827525 74195 827581
rect 74281 827525 74337 827581
rect 74423 827525 74479 827581
rect 74565 827525 74621 827581
rect 74707 827525 74763 827581
rect 74849 827525 74905 827581
rect 74991 827525 75047 827581
rect 75133 827525 75189 827581
rect 75275 827525 75331 827581
rect 73855 827383 73911 827439
rect 73997 827383 74053 827439
rect 74139 827383 74195 827439
rect 74281 827383 74337 827439
rect 74423 827383 74479 827439
rect 74565 827383 74621 827439
rect 74707 827383 74763 827439
rect 74849 827383 74905 827439
rect 74991 827383 75047 827439
rect 75133 827383 75189 827439
rect 75275 827383 75331 827439
rect 73855 827241 73911 827297
rect 73997 827241 74053 827297
rect 74139 827241 74195 827297
rect 74281 827241 74337 827297
rect 74423 827241 74479 827297
rect 74565 827241 74621 827297
rect 74707 827241 74763 827297
rect 74849 827241 74905 827297
rect 74991 827241 75047 827297
rect 75133 827241 75189 827297
rect 75275 827241 75331 827297
rect 73855 827099 73911 827155
rect 73997 827099 74053 827155
rect 74139 827099 74195 827155
rect 74281 827099 74337 827155
rect 74423 827099 74479 827155
rect 74565 827099 74621 827155
rect 74707 827099 74763 827155
rect 74849 827099 74905 827155
rect 74991 827099 75047 827155
rect 75133 827099 75189 827155
rect 75275 827099 75331 827155
rect 73855 826957 73911 827013
rect 73997 826957 74053 827013
rect 74139 826957 74195 827013
rect 74281 826957 74337 827013
rect 74423 826957 74479 827013
rect 74565 826957 74621 827013
rect 74707 826957 74763 827013
rect 74849 826957 74905 827013
rect 74991 826957 75047 827013
rect 75133 826957 75189 827013
rect 75275 826957 75331 827013
rect 73855 826815 73911 826871
rect 73997 826815 74053 826871
rect 74139 826815 74195 826871
rect 74281 826815 74337 826871
rect 74423 826815 74479 826871
rect 74565 826815 74621 826871
rect 74707 826815 74763 826871
rect 74849 826815 74905 826871
rect 74991 826815 75047 826871
rect 75133 826815 75189 826871
rect 75275 826815 75331 826871
rect 73855 826673 73911 826729
rect 73997 826673 74053 826729
rect 74139 826673 74195 826729
rect 74281 826673 74337 826729
rect 74423 826673 74479 826729
rect 74565 826673 74621 826729
rect 74707 826673 74763 826729
rect 74849 826673 74905 826729
rect 74991 826673 75047 826729
rect 75133 826673 75189 826729
rect 75275 826673 75331 826729
rect 73855 826531 73911 826587
rect 73997 826531 74053 826587
rect 74139 826531 74195 826587
rect 74281 826531 74337 826587
rect 74423 826531 74479 826587
rect 74565 826531 74621 826587
rect 74707 826531 74763 826587
rect 74849 826531 74905 826587
rect 74991 826531 75047 826587
rect 75133 826531 75189 826587
rect 75275 826531 75331 826587
rect 73855 826389 73911 826445
rect 73997 826389 74053 826445
rect 74139 826389 74195 826445
rect 74281 826389 74337 826445
rect 74423 826389 74479 826445
rect 74565 826389 74621 826445
rect 74707 826389 74763 826445
rect 74849 826389 74905 826445
rect 74991 826389 75047 826445
rect 75133 826389 75189 826445
rect 75275 826389 75331 826445
rect 73855 826247 73911 826303
rect 73997 826247 74053 826303
rect 74139 826247 74195 826303
rect 74281 826247 74337 826303
rect 74423 826247 74479 826303
rect 74565 826247 74621 826303
rect 74707 826247 74763 826303
rect 74849 826247 74905 826303
rect 74991 826247 75047 826303
rect 75133 826247 75189 826303
rect 75275 826247 75331 826303
rect 73855 826105 73911 826161
rect 73997 826105 74053 826161
rect 74139 826105 74195 826161
rect 74281 826105 74337 826161
rect 74423 826105 74479 826161
rect 74565 826105 74621 826161
rect 74707 826105 74763 826161
rect 74849 826105 74905 826161
rect 74991 826105 75047 826161
rect 75133 826105 75189 826161
rect 75275 826105 75331 826161
rect 73855 825963 73911 826019
rect 73997 825963 74053 826019
rect 74139 825963 74195 826019
rect 74281 825963 74337 826019
rect 74423 825963 74479 826019
rect 74565 825963 74621 826019
rect 74707 825963 74763 826019
rect 74849 825963 74905 826019
rect 74991 825963 75047 826019
rect 75133 825963 75189 826019
rect 75275 825963 75331 826019
rect 73855 825821 73911 825877
rect 73997 825821 74053 825877
rect 74139 825821 74195 825877
rect 74281 825821 74337 825877
rect 74423 825821 74479 825877
rect 74565 825821 74621 825877
rect 74707 825821 74763 825877
rect 74849 825821 74905 825877
rect 74991 825821 75047 825877
rect 75133 825821 75189 825877
rect 75275 825821 75331 825877
rect 73866 825038 73922 825094
rect 74008 825038 74064 825094
rect 74150 825038 74206 825094
rect 74292 825038 74348 825094
rect 74434 825038 74490 825094
rect 74576 825038 74632 825094
rect 74718 825038 74774 825094
rect 74860 825038 74916 825094
rect 75002 825038 75058 825094
rect 75144 825038 75200 825094
rect 75286 825038 75342 825094
rect 73866 824896 73922 824952
rect 74008 824896 74064 824952
rect 74150 824896 74206 824952
rect 74292 824896 74348 824952
rect 74434 824896 74490 824952
rect 74576 824896 74632 824952
rect 74718 824896 74774 824952
rect 74860 824896 74916 824952
rect 75002 824896 75058 824952
rect 75144 824896 75200 824952
rect 75286 824896 75342 824952
rect 73866 824754 73922 824810
rect 74008 824754 74064 824810
rect 74150 824754 74206 824810
rect 74292 824754 74348 824810
rect 74434 824754 74490 824810
rect 74576 824754 74632 824810
rect 74718 824754 74774 824810
rect 74860 824754 74916 824810
rect 75002 824754 75058 824810
rect 75144 824754 75200 824810
rect 75286 824754 75342 824810
rect 73866 824612 73922 824668
rect 74008 824612 74064 824668
rect 74150 824612 74206 824668
rect 74292 824612 74348 824668
rect 74434 824612 74490 824668
rect 74576 824612 74632 824668
rect 74718 824612 74774 824668
rect 74860 824612 74916 824668
rect 75002 824612 75058 824668
rect 75144 824612 75200 824668
rect 75286 824612 75342 824668
rect 73866 824470 73922 824526
rect 74008 824470 74064 824526
rect 74150 824470 74206 824526
rect 74292 824470 74348 824526
rect 74434 824470 74490 824526
rect 74576 824470 74632 824526
rect 74718 824470 74774 824526
rect 74860 824470 74916 824526
rect 75002 824470 75058 824526
rect 75144 824470 75200 824526
rect 75286 824470 75342 824526
rect 73866 824328 73922 824384
rect 74008 824328 74064 824384
rect 74150 824328 74206 824384
rect 74292 824328 74348 824384
rect 74434 824328 74490 824384
rect 74576 824328 74632 824384
rect 74718 824328 74774 824384
rect 74860 824328 74916 824384
rect 75002 824328 75058 824384
rect 75144 824328 75200 824384
rect 75286 824328 75342 824384
rect 73866 824186 73922 824242
rect 74008 824186 74064 824242
rect 74150 824186 74206 824242
rect 74292 824186 74348 824242
rect 74434 824186 74490 824242
rect 74576 824186 74632 824242
rect 74718 824186 74774 824242
rect 74860 824186 74916 824242
rect 75002 824186 75058 824242
rect 75144 824186 75200 824242
rect 75286 824186 75342 824242
rect 73866 824044 73922 824100
rect 74008 824044 74064 824100
rect 74150 824044 74206 824100
rect 74292 824044 74348 824100
rect 74434 824044 74490 824100
rect 74576 824044 74632 824100
rect 74718 824044 74774 824100
rect 74860 824044 74916 824100
rect 75002 824044 75058 824100
rect 75144 824044 75200 824100
rect 75286 824044 75342 824100
rect 73866 823902 73922 823958
rect 74008 823902 74064 823958
rect 74150 823902 74206 823958
rect 74292 823902 74348 823958
rect 74434 823902 74490 823958
rect 74576 823902 74632 823958
rect 74718 823902 74774 823958
rect 74860 823902 74916 823958
rect 75002 823902 75058 823958
rect 75144 823902 75200 823958
rect 75286 823902 75342 823958
rect 73866 823760 73922 823816
rect 74008 823760 74064 823816
rect 74150 823760 74206 823816
rect 74292 823760 74348 823816
rect 74434 823760 74490 823816
rect 74576 823760 74632 823816
rect 74718 823760 74774 823816
rect 74860 823760 74916 823816
rect 75002 823760 75058 823816
rect 75144 823760 75200 823816
rect 75286 823760 75342 823816
rect 73866 823618 73922 823674
rect 74008 823618 74064 823674
rect 74150 823618 74206 823674
rect 74292 823618 74348 823674
rect 74434 823618 74490 823674
rect 74576 823618 74632 823674
rect 74718 823618 74774 823674
rect 74860 823618 74916 823674
rect 75002 823618 75058 823674
rect 75144 823618 75200 823674
rect 75286 823618 75342 823674
rect 73866 823476 73922 823532
rect 74008 823476 74064 823532
rect 74150 823476 74206 823532
rect 74292 823476 74348 823532
rect 74434 823476 74490 823532
rect 74576 823476 74632 823532
rect 74718 823476 74774 823532
rect 74860 823476 74916 823532
rect 75002 823476 75058 823532
rect 75144 823476 75200 823532
rect 75286 823476 75342 823532
rect 73866 823334 73922 823390
rect 74008 823334 74064 823390
rect 74150 823334 74206 823390
rect 74292 823334 74348 823390
rect 74434 823334 74490 823390
rect 74576 823334 74632 823390
rect 74718 823334 74774 823390
rect 74860 823334 74916 823390
rect 75002 823334 75058 823390
rect 75144 823334 75200 823390
rect 75286 823334 75342 823390
rect 71466 796594 71522 796650
rect 71608 796594 71664 796650
rect 71750 796594 71806 796650
rect 71892 796594 71948 796650
rect 72034 796594 72090 796650
rect 72176 796594 72232 796650
rect 72318 796594 72374 796650
rect 72460 796594 72516 796650
rect 72602 796594 72658 796650
rect 72744 796594 72800 796650
rect 72886 796594 72942 796650
rect 73028 796594 73084 796650
rect 73170 796594 73226 796650
rect 73312 796594 73368 796650
rect 71466 796452 71522 796508
rect 71608 796452 71664 796508
rect 71750 796452 71806 796508
rect 71892 796452 71948 796508
rect 72034 796452 72090 796508
rect 72176 796452 72232 796508
rect 72318 796452 72374 796508
rect 72460 796452 72516 796508
rect 72602 796452 72658 796508
rect 72744 796452 72800 796508
rect 72886 796452 72942 796508
rect 73028 796452 73084 796508
rect 73170 796452 73226 796508
rect 73312 796452 73368 796508
rect 71466 796310 71522 796366
rect 71608 796310 71664 796366
rect 71750 796310 71806 796366
rect 71892 796310 71948 796366
rect 72034 796310 72090 796366
rect 72176 796310 72232 796366
rect 72318 796310 72374 796366
rect 72460 796310 72516 796366
rect 72602 796310 72658 796366
rect 72744 796310 72800 796366
rect 72886 796310 72942 796366
rect 73028 796310 73084 796366
rect 73170 796310 73226 796366
rect 73312 796310 73368 796366
rect 71466 796168 71522 796224
rect 71608 796168 71664 796224
rect 71750 796168 71806 796224
rect 71892 796168 71948 796224
rect 72034 796168 72090 796224
rect 72176 796168 72232 796224
rect 72318 796168 72374 796224
rect 72460 796168 72516 796224
rect 72602 796168 72658 796224
rect 72744 796168 72800 796224
rect 72886 796168 72942 796224
rect 73028 796168 73084 796224
rect 73170 796168 73226 796224
rect 73312 796168 73368 796224
rect 71466 796026 71522 796082
rect 71608 796026 71664 796082
rect 71750 796026 71806 796082
rect 71892 796026 71948 796082
rect 72034 796026 72090 796082
rect 72176 796026 72232 796082
rect 72318 796026 72374 796082
rect 72460 796026 72516 796082
rect 72602 796026 72658 796082
rect 72744 796026 72800 796082
rect 72886 796026 72942 796082
rect 73028 796026 73084 796082
rect 73170 796026 73226 796082
rect 73312 796026 73368 796082
rect 71466 795884 71522 795940
rect 71608 795884 71664 795940
rect 71750 795884 71806 795940
rect 71892 795884 71948 795940
rect 72034 795884 72090 795940
rect 72176 795884 72232 795940
rect 72318 795884 72374 795940
rect 72460 795884 72516 795940
rect 72602 795884 72658 795940
rect 72744 795884 72800 795940
rect 72886 795884 72942 795940
rect 73028 795884 73084 795940
rect 73170 795884 73226 795940
rect 73312 795884 73368 795940
rect 71466 795742 71522 795798
rect 71608 795742 71664 795798
rect 71750 795742 71806 795798
rect 71892 795742 71948 795798
rect 72034 795742 72090 795798
rect 72176 795742 72232 795798
rect 72318 795742 72374 795798
rect 72460 795742 72516 795798
rect 72602 795742 72658 795798
rect 72744 795742 72800 795798
rect 72886 795742 72942 795798
rect 73028 795742 73084 795798
rect 73170 795742 73226 795798
rect 73312 795742 73368 795798
rect 71466 795600 71522 795656
rect 71608 795600 71664 795656
rect 71750 795600 71806 795656
rect 71892 795600 71948 795656
rect 72034 795600 72090 795656
rect 72176 795600 72232 795656
rect 72318 795600 72374 795656
rect 72460 795600 72516 795656
rect 72602 795600 72658 795656
rect 72744 795600 72800 795656
rect 72886 795600 72942 795656
rect 73028 795600 73084 795656
rect 73170 795600 73226 795656
rect 73312 795600 73368 795656
rect 71466 795458 71522 795514
rect 71608 795458 71664 795514
rect 71750 795458 71806 795514
rect 71892 795458 71948 795514
rect 72034 795458 72090 795514
rect 72176 795458 72232 795514
rect 72318 795458 72374 795514
rect 72460 795458 72516 795514
rect 72602 795458 72658 795514
rect 72744 795458 72800 795514
rect 72886 795458 72942 795514
rect 73028 795458 73084 795514
rect 73170 795458 73226 795514
rect 73312 795458 73368 795514
rect 71466 795316 71522 795372
rect 71608 795316 71664 795372
rect 71750 795316 71806 795372
rect 71892 795316 71948 795372
rect 72034 795316 72090 795372
rect 72176 795316 72232 795372
rect 72318 795316 72374 795372
rect 72460 795316 72516 795372
rect 72602 795316 72658 795372
rect 72744 795316 72800 795372
rect 72886 795316 72942 795372
rect 73028 795316 73084 795372
rect 73170 795316 73226 795372
rect 73312 795316 73368 795372
rect 71466 795174 71522 795230
rect 71608 795174 71664 795230
rect 71750 795174 71806 795230
rect 71892 795174 71948 795230
rect 72034 795174 72090 795230
rect 72176 795174 72232 795230
rect 72318 795174 72374 795230
rect 72460 795174 72516 795230
rect 72602 795174 72658 795230
rect 72744 795174 72800 795230
rect 72886 795174 72942 795230
rect 73028 795174 73084 795230
rect 73170 795174 73226 795230
rect 73312 795174 73368 795230
rect 71466 795032 71522 795088
rect 71608 795032 71664 795088
rect 71750 795032 71806 795088
rect 71892 795032 71948 795088
rect 72034 795032 72090 795088
rect 72176 795032 72232 795088
rect 72318 795032 72374 795088
rect 72460 795032 72516 795088
rect 72602 795032 72658 795088
rect 72744 795032 72800 795088
rect 72886 795032 72942 795088
rect 73028 795032 73084 795088
rect 73170 795032 73226 795088
rect 73312 795032 73368 795088
rect 71466 794890 71522 794946
rect 71608 794890 71664 794946
rect 71750 794890 71806 794946
rect 71892 794890 71948 794946
rect 72034 794890 72090 794946
rect 72176 794890 72232 794946
rect 72318 794890 72374 794946
rect 72460 794890 72516 794946
rect 72602 794890 72658 794946
rect 72744 794890 72800 794946
rect 72886 794890 72942 794946
rect 73028 794890 73084 794946
rect 73170 794890 73226 794946
rect 73312 794890 73368 794946
rect 71455 794113 71511 794169
rect 71597 794113 71653 794169
rect 71739 794113 71795 794169
rect 71881 794113 71937 794169
rect 72023 794113 72079 794169
rect 72165 794113 72221 794169
rect 72307 794113 72363 794169
rect 72449 794113 72505 794169
rect 72591 794113 72647 794169
rect 72733 794113 72789 794169
rect 72875 794113 72931 794169
rect 73017 794113 73073 794169
rect 73159 794113 73215 794169
rect 73301 794113 73357 794169
rect 71455 793971 71511 794027
rect 71597 793971 71653 794027
rect 71739 793971 71795 794027
rect 71881 793971 71937 794027
rect 72023 793971 72079 794027
rect 72165 793971 72221 794027
rect 72307 793971 72363 794027
rect 72449 793971 72505 794027
rect 72591 793971 72647 794027
rect 72733 793971 72789 794027
rect 72875 793971 72931 794027
rect 73017 793971 73073 794027
rect 73159 793971 73215 794027
rect 73301 793971 73357 794027
rect 71455 793829 71511 793885
rect 71597 793829 71653 793885
rect 71739 793829 71795 793885
rect 71881 793829 71937 793885
rect 72023 793829 72079 793885
rect 72165 793829 72221 793885
rect 72307 793829 72363 793885
rect 72449 793829 72505 793885
rect 72591 793829 72647 793885
rect 72733 793829 72789 793885
rect 72875 793829 72931 793885
rect 73017 793829 73073 793885
rect 73159 793829 73215 793885
rect 73301 793829 73357 793885
rect 71455 793687 71511 793743
rect 71597 793687 71653 793743
rect 71739 793687 71795 793743
rect 71881 793687 71937 793743
rect 72023 793687 72079 793743
rect 72165 793687 72221 793743
rect 72307 793687 72363 793743
rect 72449 793687 72505 793743
rect 72591 793687 72647 793743
rect 72733 793687 72789 793743
rect 72875 793687 72931 793743
rect 73017 793687 73073 793743
rect 73159 793687 73215 793743
rect 73301 793687 73357 793743
rect 71455 793545 71511 793601
rect 71597 793545 71653 793601
rect 71739 793545 71795 793601
rect 71881 793545 71937 793601
rect 72023 793545 72079 793601
rect 72165 793545 72221 793601
rect 72307 793545 72363 793601
rect 72449 793545 72505 793601
rect 72591 793545 72647 793601
rect 72733 793545 72789 793601
rect 72875 793545 72931 793601
rect 73017 793545 73073 793601
rect 73159 793545 73215 793601
rect 73301 793545 73357 793601
rect 71455 793403 71511 793459
rect 71597 793403 71653 793459
rect 71739 793403 71795 793459
rect 71881 793403 71937 793459
rect 72023 793403 72079 793459
rect 72165 793403 72221 793459
rect 72307 793403 72363 793459
rect 72449 793403 72505 793459
rect 72591 793403 72647 793459
rect 72733 793403 72789 793459
rect 72875 793403 72931 793459
rect 73017 793403 73073 793459
rect 73159 793403 73215 793459
rect 73301 793403 73357 793459
rect 71455 793261 71511 793317
rect 71597 793261 71653 793317
rect 71739 793261 71795 793317
rect 71881 793261 71937 793317
rect 72023 793261 72079 793317
rect 72165 793261 72221 793317
rect 72307 793261 72363 793317
rect 72449 793261 72505 793317
rect 72591 793261 72647 793317
rect 72733 793261 72789 793317
rect 72875 793261 72931 793317
rect 73017 793261 73073 793317
rect 73159 793261 73215 793317
rect 73301 793261 73357 793317
rect 71455 793119 71511 793175
rect 71597 793119 71653 793175
rect 71739 793119 71795 793175
rect 71881 793119 71937 793175
rect 72023 793119 72079 793175
rect 72165 793119 72221 793175
rect 72307 793119 72363 793175
rect 72449 793119 72505 793175
rect 72591 793119 72647 793175
rect 72733 793119 72789 793175
rect 72875 793119 72931 793175
rect 73017 793119 73073 793175
rect 73159 793119 73215 793175
rect 73301 793119 73357 793175
rect 71455 792977 71511 793033
rect 71597 792977 71653 793033
rect 71739 792977 71795 793033
rect 71881 792977 71937 793033
rect 72023 792977 72079 793033
rect 72165 792977 72221 793033
rect 72307 792977 72363 793033
rect 72449 792977 72505 793033
rect 72591 792977 72647 793033
rect 72733 792977 72789 793033
rect 72875 792977 72931 793033
rect 73017 792977 73073 793033
rect 73159 792977 73215 793033
rect 73301 792977 73357 793033
rect 71455 792835 71511 792891
rect 71597 792835 71653 792891
rect 71739 792835 71795 792891
rect 71881 792835 71937 792891
rect 72023 792835 72079 792891
rect 72165 792835 72221 792891
rect 72307 792835 72363 792891
rect 72449 792835 72505 792891
rect 72591 792835 72647 792891
rect 72733 792835 72789 792891
rect 72875 792835 72931 792891
rect 73017 792835 73073 792891
rect 73159 792835 73215 792891
rect 73301 792835 73357 792891
rect 71455 792693 71511 792749
rect 71597 792693 71653 792749
rect 71739 792693 71795 792749
rect 71881 792693 71937 792749
rect 72023 792693 72079 792749
rect 72165 792693 72221 792749
rect 72307 792693 72363 792749
rect 72449 792693 72505 792749
rect 72591 792693 72647 792749
rect 72733 792693 72789 792749
rect 72875 792693 72931 792749
rect 73017 792693 73073 792749
rect 73159 792693 73215 792749
rect 73301 792693 73357 792749
rect 71455 792551 71511 792607
rect 71597 792551 71653 792607
rect 71739 792551 71795 792607
rect 71881 792551 71937 792607
rect 72023 792551 72079 792607
rect 72165 792551 72221 792607
rect 72307 792551 72363 792607
rect 72449 792551 72505 792607
rect 72591 792551 72647 792607
rect 72733 792551 72789 792607
rect 72875 792551 72931 792607
rect 73017 792551 73073 792607
rect 73159 792551 73215 792607
rect 73301 792551 73357 792607
rect 71455 792409 71511 792465
rect 71597 792409 71653 792465
rect 71739 792409 71795 792465
rect 71881 792409 71937 792465
rect 72023 792409 72079 792465
rect 72165 792409 72221 792465
rect 72307 792409 72363 792465
rect 72449 792409 72505 792465
rect 72591 792409 72647 792465
rect 72733 792409 72789 792465
rect 72875 792409 72931 792465
rect 73017 792409 73073 792465
rect 73159 792409 73215 792465
rect 73301 792409 73357 792465
rect 71455 792267 71511 792323
rect 71597 792267 71653 792323
rect 71739 792267 71795 792323
rect 71881 792267 71937 792323
rect 72023 792267 72079 792323
rect 72165 792267 72221 792323
rect 72307 792267 72363 792323
rect 72449 792267 72505 792323
rect 72591 792267 72647 792323
rect 72733 792267 72789 792323
rect 72875 792267 72931 792323
rect 73017 792267 73073 792323
rect 73159 792267 73215 792323
rect 73301 792267 73357 792323
rect 71455 791743 71511 791799
rect 71597 791743 71653 791799
rect 71739 791743 71795 791799
rect 71881 791743 71937 791799
rect 72023 791743 72079 791799
rect 72165 791743 72221 791799
rect 72307 791743 72363 791799
rect 72449 791743 72505 791799
rect 72591 791743 72647 791799
rect 72733 791743 72789 791799
rect 72875 791743 72931 791799
rect 73017 791743 73073 791799
rect 73159 791743 73215 791799
rect 73301 791743 73357 791799
rect 71455 791601 71511 791657
rect 71597 791601 71653 791657
rect 71739 791601 71795 791657
rect 71881 791601 71937 791657
rect 72023 791601 72079 791657
rect 72165 791601 72221 791657
rect 72307 791601 72363 791657
rect 72449 791601 72505 791657
rect 72591 791601 72647 791657
rect 72733 791601 72789 791657
rect 72875 791601 72931 791657
rect 73017 791601 73073 791657
rect 73159 791601 73215 791657
rect 73301 791601 73357 791657
rect 71455 791459 71511 791515
rect 71597 791459 71653 791515
rect 71739 791459 71795 791515
rect 71881 791459 71937 791515
rect 72023 791459 72079 791515
rect 72165 791459 72221 791515
rect 72307 791459 72363 791515
rect 72449 791459 72505 791515
rect 72591 791459 72647 791515
rect 72733 791459 72789 791515
rect 72875 791459 72931 791515
rect 73017 791459 73073 791515
rect 73159 791459 73215 791515
rect 73301 791459 73357 791515
rect 71455 791317 71511 791373
rect 71597 791317 71653 791373
rect 71739 791317 71795 791373
rect 71881 791317 71937 791373
rect 72023 791317 72079 791373
rect 72165 791317 72221 791373
rect 72307 791317 72363 791373
rect 72449 791317 72505 791373
rect 72591 791317 72647 791373
rect 72733 791317 72789 791373
rect 72875 791317 72931 791373
rect 73017 791317 73073 791373
rect 73159 791317 73215 791373
rect 73301 791317 73357 791373
rect 71455 791175 71511 791231
rect 71597 791175 71653 791231
rect 71739 791175 71795 791231
rect 71881 791175 71937 791231
rect 72023 791175 72079 791231
rect 72165 791175 72221 791231
rect 72307 791175 72363 791231
rect 72449 791175 72505 791231
rect 72591 791175 72647 791231
rect 72733 791175 72789 791231
rect 72875 791175 72931 791231
rect 73017 791175 73073 791231
rect 73159 791175 73215 791231
rect 73301 791175 73357 791231
rect 71455 791033 71511 791089
rect 71597 791033 71653 791089
rect 71739 791033 71795 791089
rect 71881 791033 71937 791089
rect 72023 791033 72079 791089
rect 72165 791033 72221 791089
rect 72307 791033 72363 791089
rect 72449 791033 72505 791089
rect 72591 791033 72647 791089
rect 72733 791033 72789 791089
rect 72875 791033 72931 791089
rect 73017 791033 73073 791089
rect 73159 791033 73215 791089
rect 73301 791033 73357 791089
rect 71455 790891 71511 790947
rect 71597 790891 71653 790947
rect 71739 790891 71795 790947
rect 71881 790891 71937 790947
rect 72023 790891 72079 790947
rect 72165 790891 72221 790947
rect 72307 790891 72363 790947
rect 72449 790891 72505 790947
rect 72591 790891 72647 790947
rect 72733 790891 72789 790947
rect 72875 790891 72931 790947
rect 73017 790891 73073 790947
rect 73159 790891 73215 790947
rect 73301 790891 73357 790947
rect 71455 790749 71511 790805
rect 71597 790749 71653 790805
rect 71739 790749 71795 790805
rect 71881 790749 71937 790805
rect 72023 790749 72079 790805
rect 72165 790749 72221 790805
rect 72307 790749 72363 790805
rect 72449 790749 72505 790805
rect 72591 790749 72647 790805
rect 72733 790749 72789 790805
rect 72875 790749 72931 790805
rect 73017 790749 73073 790805
rect 73159 790749 73215 790805
rect 73301 790749 73357 790805
rect 71455 790607 71511 790663
rect 71597 790607 71653 790663
rect 71739 790607 71795 790663
rect 71881 790607 71937 790663
rect 72023 790607 72079 790663
rect 72165 790607 72221 790663
rect 72307 790607 72363 790663
rect 72449 790607 72505 790663
rect 72591 790607 72647 790663
rect 72733 790607 72789 790663
rect 72875 790607 72931 790663
rect 73017 790607 73073 790663
rect 73159 790607 73215 790663
rect 73301 790607 73357 790663
rect 71455 790465 71511 790521
rect 71597 790465 71653 790521
rect 71739 790465 71795 790521
rect 71881 790465 71937 790521
rect 72023 790465 72079 790521
rect 72165 790465 72221 790521
rect 72307 790465 72363 790521
rect 72449 790465 72505 790521
rect 72591 790465 72647 790521
rect 72733 790465 72789 790521
rect 72875 790465 72931 790521
rect 73017 790465 73073 790521
rect 73159 790465 73215 790521
rect 73301 790465 73357 790521
rect 71455 790323 71511 790379
rect 71597 790323 71653 790379
rect 71739 790323 71795 790379
rect 71881 790323 71937 790379
rect 72023 790323 72079 790379
rect 72165 790323 72221 790379
rect 72307 790323 72363 790379
rect 72449 790323 72505 790379
rect 72591 790323 72647 790379
rect 72733 790323 72789 790379
rect 72875 790323 72931 790379
rect 73017 790323 73073 790379
rect 73159 790323 73215 790379
rect 73301 790323 73357 790379
rect 71455 790181 71511 790237
rect 71597 790181 71653 790237
rect 71739 790181 71795 790237
rect 71881 790181 71937 790237
rect 72023 790181 72079 790237
rect 72165 790181 72221 790237
rect 72307 790181 72363 790237
rect 72449 790181 72505 790237
rect 72591 790181 72647 790237
rect 72733 790181 72789 790237
rect 72875 790181 72931 790237
rect 73017 790181 73073 790237
rect 73159 790181 73215 790237
rect 73301 790181 73357 790237
rect 71455 790039 71511 790095
rect 71597 790039 71653 790095
rect 71739 790039 71795 790095
rect 71881 790039 71937 790095
rect 72023 790039 72079 790095
rect 72165 790039 72221 790095
rect 72307 790039 72363 790095
rect 72449 790039 72505 790095
rect 72591 790039 72647 790095
rect 72733 790039 72789 790095
rect 72875 790039 72931 790095
rect 73017 790039 73073 790095
rect 73159 790039 73215 790095
rect 73301 790039 73357 790095
rect 71455 789897 71511 789953
rect 71597 789897 71653 789953
rect 71739 789897 71795 789953
rect 71881 789897 71937 789953
rect 72023 789897 72079 789953
rect 72165 789897 72221 789953
rect 72307 789897 72363 789953
rect 72449 789897 72505 789953
rect 72591 789897 72647 789953
rect 72733 789897 72789 789953
rect 72875 789897 72931 789953
rect 73017 789897 73073 789953
rect 73159 789897 73215 789953
rect 73301 789897 73357 789953
rect 700040 791610 700096 791666
rect 700182 791610 700238 791666
rect 700324 791610 700380 791666
rect 700466 791610 700522 791666
rect 700608 791610 700664 791666
rect 700750 791610 700806 791666
rect 700892 791610 700948 791666
rect 701034 791610 701090 791666
rect 701176 791610 701232 791666
rect 701318 791610 701374 791666
rect 701460 791610 701516 791666
rect 701602 791610 701658 791666
rect 701744 791610 701800 791666
rect 701886 791610 701942 791666
rect 700040 791468 700096 791524
rect 700182 791468 700238 791524
rect 700324 791468 700380 791524
rect 700466 791468 700522 791524
rect 700608 791468 700664 791524
rect 700750 791468 700806 791524
rect 700892 791468 700948 791524
rect 701034 791468 701090 791524
rect 701176 791468 701232 791524
rect 701318 791468 701374 791524
rect 701460 791468 701516 791524
rect 701602 791468 701658 791524
rect 701744 791468 701800 791524
rect 701886 791468 701942 791524
rect 700040 791326 700096 791382
rect 700182 791326 700238 791382
rect 700324 791326 700380 791382
rect 700466 791326 700522 791382
rect 700608 791326 700664 791382
rect 700750 791326 700806 791382
rect 700892 791326 700948 791382
rect 701034 791326 701090 791382
rect 701176 791326 701232 791382
rect 701318 791326 701374 791382
rect 701460 791326 701516 791382
rect 701602 791326 701658 791382
rect 701744 791326 701800 791382
rect 701886 791326 701942 791382
rect 700040 791184 700096 791240
rect 700182 791184 700238 791240
rect 700324 791184 700380 791240
rect 700466 791184 700522 791240
rect 700608 791184 700664 791240
rect 700750 791184 700806 791240
rect 700892 791184 700948 791240
rect 701034 791184 701090 791240
rect 701176 791184 701232 791240
rect 701318 791184 701374 791240
rect 701460 791184 701516 791240
rect 701602 791184 701658 791240
rect 701744 791184 701800 791240
rect 701886 791184 701942 791240
rect 700040 791042 700096 791098
rect 700182 791042 700238 791098
rect 700324 791042 700380 791098
rect 700466 791042 700522 791098
rect 700608 791042 700664 791098
rect 700750 791042 700806 791098
rect 700892 791042 700948 791098
rect 701034 791042 701090 791098
rect 701176 791042 701232 791098
rect 701318 791042 701374 791098
rect 701460 791042 701516 791098
rect 701602 791042 701658 791098
rect 701744 791042 701800 791098
rect 701886 791042 701942 791098
rect 700040 790900 700096 790956
rect 700182 790900 700238 790956
rect 700324 790900 700380 790956
rect 700466 790900 700522 790956
rect 700608 790900 700664 790956
rect 700750 790900 700806 790956
rect 700892 790900 700948 790956
rect 701034 790900 701090 790956
rect 701176 790900 701232 790956
rect 701318 790900 701374 790956
rect 701460 790900 701516 790956
rect 701602 790900 701658 790956
rect 701744 790900 701800 790956
rect 701886 790900 701942 790956
rect 700040 790758 700096 790814
rect 700182 790758 700238 790814
rect 700324 790758 700380 790814
rect 700466 790758 700522 790814
rect 700608 790758 700664 790814
rect 700750 790758 700806 790814
rect 700892 790758 700948 790814
rect 701034 790758 701090 790814
rect 701176 790758 701232 790814
rect 701318 790758 701374 790814
rect 701460 790758 701516 790814
rect 701602 790758 701658 790814
rect 701744 790758 701800 790814
rect 701886 790758 701942 790814
rect 700040 790616 700096 790672
rect 700182 790616 700238 790672
rect 700324 790616 700380 790672
rect 700466 790616 700522 790672
rect 700608 790616 700664 790672
rect 700750 790616 700806 790672
rect 700892 790616 700948 790672
rect 701034 790616 701090 790672
rect 701176 790616 701232 790672
rect 701318 790616 701374 790672
rect 701460 790616 701516 790672
rect 701602 790616 701658 790672
rect 701744 790616 701800 790672
rect 701886 790616 701942 790672
rect 700040 790474 700096 790530
rect 700182 790474 700238 790530
rect 700324 790474 700380 790530
rect 700466 790474 700522 790530
rect 700608 790474 700664 790530
rect 700750 790474 700806 790530
rect 700892 790474 700948 790530
rect 701034 790474 701090 790530
rect 701176 790474 701232 790530
rect 701318 790474 701374 790530
rect 701460 790474 701516 790530
rect 701602 790474 701658 790530
rect 701744 790474 701800 790530
rect 701886 790474 701942 790530
rect 700040 790332 700096 790388
rect 700182 790332 700238 790388
rect 700324 790332 700380 790388
rect 700466 790332 700522 790388
rect 700608 790332 700664 790388
rect 700750 790332 700806 790388
rect 700892 790332 700948 790388
rect 701034 790332 701090 790388
rect 701176 790332 701232 790388
rect 701318 790332 701374 790388
rect 701460 790332 701516 790388
rect 701602 790332 701658 790388
rect 701744 790332 701800 790388
rect 701886 790332 701942 790388
rect 700040 790190 700096 790246
rect 700182 790190 700238 790246
rect 700324 790190 700380 790246
rect 700466 790190 700522 790246
rect 700608 790190 700664 790246
rect 700750 790190 700806 790246
rect 700892 790190 700948 790246
rect 701034 790190 701090 790246
rect 701176 790190 701232 790246
rect 701318 790190 701374 790246
rect 701460 790190 701516 790246
rect 701602 790190 701658 790246
rect 701744 790190 701800 790246
rect 701886 790190 701942 790246
rect 700040 790048 700096 790104
rect 700182 790048 700238 790104
rect 700324 790048 700380 790104
rect 700466 790048 700522 790104
rect 700608 790048 700664 790104
rect 700750 790048 700806 790104
rect 700892 790048 700948 790104
rect 701034 790048 701090 790104
rect 701176 790048 701232 790104
rect 701318 790048 701374 790104
rect 701460 790048 701516 790104
rect 701602 790048 701658 790104
rect 701744 790048 701800 790104
rect 701886 790048 701942 790104
rect 700040 789906 700096 789962
rect 700182 789906 700238 789962
rect 700324 789906 700380 789962
rect 700466 789906 700522 789962
rect 700608 789906 700664 789962
rect 700750 789906 700806 789962
rect 700892 789906 700948 789962
rect 701034 789906 701090 789962
rect 701176 789906 701232 789962
rect 701318 789906 701374 789962
rect 701460 789906 701516 789962
rect 701602 789906 701658 789962
rect 701744 789906 701800 789962
rect 701886 789906 701942 789962
rect 71455 789037 71511 789093
rect 71597 789037 71653 789093
rect 71739 789037 71795 789093
rect 71881 789037 71937 789093
rect 72023 789037 72079 789093
rect 72165 789037 72221 789093
rect 72307 789037 72363 789093
rect 72449 789037 72505 789093
rect 72591 789037 72647 789093
rect 72733 789037 72789 789093
rect 72875 789037 72931 789093
rect 73017 789037 73073 789093
rect 73159 789037 73215 789093
rect 73301 789037 73357 789093
rect 71455 788895 71511 788951
rect 71597 788895 71653 788951
rect 71739 788895 71795 788951
rect 71881 788895 71937 788951
rect 72023 788895 72079 788951
rect 72165 788895 72221 788951
rect 72307 788895 72363 788951
rect 72449 788895 72505 788951
rect 72591 788895 72647 788951
rect 72733 788895 72789 788951
rect 72875 788895 72931 788951
rect 73017 788895 73073 788951
rect 73159 788895 73215 788951
rect 73301 788895 73357 788951
rect 71455 788753 71511 788809
rect 71597 788753 71653 788809
rect 71739 788753 71795 788809
rect 71881 788753 71937 788809
rect 72023 788753 72079 788809
rect 72165 788753 72221 788809
rect 72307 788753 72363 788809
rect 72449 788753 72505 788809
rect 72591 788753 72647 788809
rect 72733 788753 72789 788809
rect 72875 788753 72931 788809
rect 73017 788753 73073 788809
rect 73159 788753 73215 788809
rect 73301 788753 73357 788809
rect 71455 788611 71511 788667
rect 71597 788611 71653 788667
rect 71739 788611 71795 788667
rect 71881 788611 71937 788667
rect 72023 788611 72079 788667
rect 72165 788611 72221 788667
rect 72307 788611 72363 788667
rect 72449 788611 72505 788667
rect 72591 788611 72647 788667
rect 72733 788611 72789 788667
rect 72875 788611 72931 788667
rect 73017 788611 73073 788667
rect 73159 788611 73215 788667
rect 73301 788611 73357 788667
rect 71455 788469 71511 788525
rect 71597 788469 71653 788525
rect 71739 788469 71795 788525
rect 71881 788469 71937 788525
rect 72023 788469 72079 788525
rect 72165 788469 72221 788525
rect 72307 788469 72363 788525
rect 72449 788469 72505 788525
rect 72591 788469 72647 788525
rect 72733 788469 72789 788525
rect 72875 788469 72931 788525
rect 73017 788469 73073 788525
rect 73159 788469 73215 788525
rect 73301 788469 73357 788525
rect 71455 788327 71511 788383
rect 71597 788327 71653 788383
rect 71739 788327 71795 788383
rect 71881 788327 71937 788383
rect 72023 788327 72079 788383
rect 72165 788327 72221 788383
rect 72307 788327 72363 788383
rect 72449 788327 72505 788383
rect 72591 788327 72647 788383
rect 72733 788327 72789 788383
rect 72875 788327 72931 788383
rect 73017 788327 73073 788383
rect 73159 788327 73215 788383
rect 73301 788327 73357 788383
rect 71455 788185 71511 788241
rect 71597 788185 71653 788241
rect 71739 788185 71795 788241
rect 71881 788185 71937 788241
rect 72023 788185 72079 788241
rect 72165 788185 72221 788241
rect 72307 788185 72363 788241
rect 72449 788185 72505 788241
rect 72591 788185 72647 788241
rect 72733 788185 72789 788241
rect 72875 788185 72931 788241
rect 73017 788185 73073 788241
rect 73159 788185 73215 788241
rect 73301 788185 73357 788241
rect 71455 788043 71511 788099
rect 71597 788043 71653 788099
rect 71739 788043 71795 788099
rect 71881 788043 71937 788099
rect 72023 788043 72079 788099
rect 72165 788043 72221 788099
rect 72307 788043 72363 788099
rect 72449 788043 72505 788099
rect 72591 788043 72647 788099
rect 72733 788043 72789 788099
rect 72875 788043 72931 788099
rect 73017 788043 73073 788099
rect 73159 788043 73215 788099
rect 73301 788043 73357 788099
rect 71455 787901 71511 787957
rect 71597 787901 71653 787957
rect 71739 787901 71795 787957
rect 71881 787901 71937 787957
rect 72023 787901 72079 787957
rect 72165 787901 72221 787957
rect 72307 787901 72363 787957
rect 72449 787901 72505 787957
rect 72591 787901 72647 787957
rect 72733 787901 72789 787957
rect 72875 787901 72931 787957
rect 73017 787901 73073 787957
rect 73159 787901 73215 787957
rect 73301 787901 73357 787957
rect 71455 787759 71511 787815
rect 71597 787759 71653 787815
rect 71739 787759 71795 787815
rect 71881 787759 71937 787815
rect 72023 787759 72079 787815
rect 72165 787759 72221 787815
rect 72307 787759 72363 787815
rect 72449 787759 72505 787815
rect 72591 787759 72647 787815
rect 72733 787759 72789 787815
rect 72875 787759 72931 787815
rect 73017 787759 73073 787815
rect 73159 787759 73215 787815
rect 73301 787759 73357 787815
rect 71455 787617 71511 787673
rect 71597 787617 71653 787673
rect 71739 787617 71795 787673
rect 71881 787617 71937 787673
rect 72023 787617 72079 787673
rect 72165 787617 72221 787673
rect 72307 787617 72363 787673
rect 72449 787617 72505 787673
rect 72591 787617 72647 787673
rect 72733 787617 72789 787673
rect 72875 787617 72931 787673
rect 73017 787617 73073 787673
rect 73159 787617 73215 787673
rect 73301 787617 73357 787673
rect 71455 787475 71511 787531
rect 71597 787475 71653 787531
rect 71739 787475 71795 787531
rect 71881 787475 71937 787531
rect 72023 787475 72079 787531
rect 72165 787475 72221 787531
rect 72307 787475 72363 787531
rect 72449 787475 72505 787531
rect 72591 787475 72647 787531
rect 72733 787475 72789 787531
rect 72875 787475 72931 787531
rect 73017 787475 73073 787531
rect 73159 787475 73215 787531
rect 73301 787475 73357 787531
rect 71455 787333 71511 787389
rect 71597 787333 71653 787389
rect 71739 787333 71795 787389
rect 71881 787333 71937 787389
rect 72023 787333 72079 787389
rect 72165 787333 72221 787389
rect 72307 787333 72363 787389
rect 72449 787333 72505 787389
rect 72591 787333 72647 787389
rect 72733 787333 72789 787389
rect 72875 787333 72931 787389
rect 73017 787333 73073 787389
rect 73159 787333 73215 787389
rect 73301 787333 73357 787389
rect 71455 787191 71511 787247
rect 71597 787191 71653 787247
rect 71739 787191 71795 787247
rect 71881 787191 71937 787247
rect 72023 787191 72079 787247
rect 72165 787191 72221 787247
rect 72307 787191 72363 787247
rect 72449 787191 72505 787247
rect 72591 787191 72647 787247
rect 72733 787191 72789 787247
rect 72875 787191 72931 787247
rect 73017 787191 73073 787247
rect 73159 787191 73215 787247
rect 73301 787191 73357 787247
rect 700051 789123 700107 789179
rect 700193 789123 700249 789179
rect 700335 789123 700391 789179
rect 700477 789123 700533 789179
rect 700619 789123 700675 789179
rect 700761 789123 700817 789179
rect 700903 789123 700959 789179
rect 701045 789123 701101 789179
rect 701187 789123 701243 789179
rect 701329 789123 701385 789179
rect 701471 789123 701527 789179
rect 701613 789123 701669 789179
rect 701755 789123 701811 789179
rect 701897 789123 701953 789179
rect 700051 788981 700107 789037
rect 700193 788981 700249 789037
rect 700335 788981 700391 789037
rect 700477 788981 700533 789037
rect 700619 788981 700675 789037
rect 700761 788981 700817 789037
rect 700903 788981 700959 789037
rect 701045 788981 701101 789037
rect 701187 788981 701243 789037
rect 701329 788981 701385 789037
rect 701471 788981 701527 789037
rect 701613 788981 701669 789037
rect 701755 788981 701811 789037
rect 701897 788981 701953 789037
rect 700051 788839 700107 788895
rect 700193 788839 700249 788895
rect 700335 788839 700391 788895
rect 700477 788839 700533 788895
rect 700619 788839 700675 788895
rect 700761 788839 700817 788895
rect 700903 788839 700959 788895
rect 701045 788839 701101 788895
rect 701187 788839 701243 788895
rect 701329 788839 701385 788895
rect 701471 788839 701527 788895
rect 701613 788839 701669 788895
rect 701755 788839 701811 788895
rect 701897 788839 701953 788895
rect 700051 788697 700107 788753
rect 700193 788697 700249 788753
rect 700335 788697 700391 788753
rect 700477 788697 700533 788753
rect 700619 788697 700675 788753
rect 700761 788697 700817 788753
rect 700903 788697 700959 788753
rect 701045 788697 701101 788753
rect 701187 788697 701243 788753
rect 701329 788697 701385 788753
rect 701471 788697 701527 788753
rect 701613 788697 701669 788753
rect 701755 788697 701811 788753
rect 701897 788697 701953 788753
rect 700051 788555 700107 788611
rect 700193 788555 700249 788611
rect 700335 788555 700391 788611
rect 700477 788555 700533 788611
rect 700619 788555 700675 788611
rect 700761 788555 700817 788611
rect 700903 788555 700959 788611
rect 701045 788555 701101 788611
rect 701187 788555 701243 788611
rect 701329 788555 701385 788611
rect 701471 788555 701527 788611
rect 701613 788555 701669 788611
rect 701755 788555 701811 788611
rect 701897 788555 701953 788611
rect 700051 788413 700107 788469
rect 700193 788413 700249 788469
rect 700335 788413 700391 788469
rect 700477 788413 700533 788469
rect 700619 788413 700675 788469
rect 700761 788413 700817 788469
rect 700903 788413 700959 788469
rect 701045 788413 701101 788469
rect 701187 788413 701243 788469
rect 701329 788413 701385 788469
rect 701471 788413 701527 788469
rect 701613 788413 701669 788469
rect 701755 788413 701811 788469
rect 701897 788413 701953 788469
rect 700051 788271 700107 788327
rect 700193 788271 700249 788327
rect 700335 788271 700391 788327
rect 700477 788271 700533 788327
rect 700619 788271 700675 788327
rect 700761 788271 700817 788327
rect 700903 788271 700959 788327
rect 701045 788271 701101 788327
rect 701187 788271 701243 788327
rect 701329 788271 701385 788327
rect 701471 788271 701527 788327
rect 701613 788271 701669 788327
rect 701755 788271 701811 788327
rect 701897 788271 701953 788327
rect 700051 788129 700107 788185
rect 700193 788129 700249 788185
rect 700335 788129 700391 788185
rect 700477 788129 700533 788185
rect 700619 788129 700675 788185
rect 700761 788129 700817 788185
rect 700903 788129 700959 788185
rect 701045 788129 701101 788185
rect 701187 788129 701243 788185
rect 701329 788129 701385 788185
rect 701471 788129 701527 788185
rect 701613 788129 701669 788185
rect 701755 788129 701811 788185
rect 701897 788129 701953 788185
rect 700051 787987 700107 788043
rect 700193 787987 700249 788043
rect 700335 787987 700391 788043
rect 700477 787987 700533 788043
rect 700619 787987 700675 788043
rect 700761 787987 700817 788043
rect 700903 787987 700959 788043
rect 701045 787987 701101 788043
rect 701187 787987 701243 788043
rect 701329 787987 701385 788043
rect 701471 787987 701527 788043
rect 701613 787987 701669 788043
rect 701755 787987 701811 788043
rect 701897 787987 701953 788043
rect 700051 787845 700107 787901
rect 700193 787845 700249 787901
rect 700335 787845 700391 787901
rect 700477 787845 700533 787901
rect 700619 787845 700675 787901
rect 700761 787845 700817 787901
rect 700903 787845 700959 787901
rect 701045 787845 701101 787901
rect 701187 787845 701243 787901
rect 701329 787845 701385 787901
rect 701471 787845 701527 787901
rect 701613 787845 701669 787901
rect 701755 787845 701811 787901
rect 701897 787845 701953 787901
rect 700051 787703 700107 787759
rect 700193 787703 700249 787759
rect 700335 787703 700391 787759
rect 700477 787703 700533 787759
rect 700619 787703 700675 787759
rect 700761 787703 700817 787759
rect 700903 787703 700959 787759
rect 701045 787703 701101 787759
rect 701187 787703 701243 787759
rect 701329 787703 701385 787759
rect 701471 787703 701527 787759
rect 701613 787703 701669 787759
rect 701755 787703 701811 787759
rect 701897 787703 701953 787759
rect 700051 787561 700107 787617
rect 700193 787561 700249 787617
rect 700335 787561 700391 787617
rect 700477 787561 700533 787617
rect 700619 787561 700675 787617
rect 700761 787561 700817 787617
rect 700903 787561 700959 787617
rect 701045 787561 701101 787617
rect 701187 787561 701243 787617
rect 701329 787561 701385 787617
rect 701471 787561 701527 787617
rect 701613 787561 701669 787617
rect 701755 787561 701811 787617
rect 701897 787561 701953 787617
rect 700051 787419 700107 787475
rect 700193 787419 700249 787475
rect 700335 787419 700391 787475
rect 700477 787419 700533 787475
rect 700619 787419 700675 787475
rect 700761 787419 700817 787475
rect 700903 787419 700959 787475
rect 701045 787419 701101 787475
rect 701187 787419 701243 787475
rect 701329 787419 701385 787475
rect 701471 787419 701527 787475
rect 701613 787419 701669 787475
rect 701755 787419 701811 787475
rect 701897 787419 701953 787475
rect 700051 787277 700107 787333
rect 700193 787277 700249 787333
rect 700335 787277 700391 787333
rect 700477 787277 700533 787333
rect 700619 787277 700675 787333
rect 700761 787277 700817 787333
rect 700903 787277 700959 787333
rect 701045 787277 701101 787333
rect 701187 787277 701243 787333
rect 701329 787277 701385 787333
rect 701471 787277 701527 787333
rect 701613 787277 701669 787333
rect 701755 787277 701811 787333
rect 701897 787277 701953 787333
rect 71455 786667 71511 786723
rect 71597 786667 71653 786723
rect 71739 786667 71795 786723
rect 71881 786667 71937 786723
rect 72023 786667 72079 786723
rect 72165 786667 72221 786723
rect 72307 786667 72363 786723
rect 72449 786667 72505 786723
rect 72591 786667 72647 786723
rect 72733 786667 72789 786723
rect 72875 786667 72931 786723
rect 73017 786667 73073 786723
rect 73159 786667 73215 786723
rect 73301 786667 73357 786723
rect 71455 786525 71511 786581
rect 71597 786525 71653 786581
rect 71739 786525 71795 786581
rect 71881 786525 71937 786581
rect 72023 786525 72079 786581
rect 72165 786525 72221 786581
rect 72307 786525 72363 786581
rect 72449 786525 72505 786581
rect 72591 786525 72647 786581
rect 72733 786525 72789 786581
rect 72875 786525 72931 786581
rect 73017 786525 73073 786581
rect 73159 786525 73215 786581
rect 73301 786525 73357 786581
rect 71455 786383 71511 786439
rect 71597 786383 71653 786439
rect 71739 786383 71795 786439
rect 71881 786383 71937 786439
rect 72023 786383 72079 786439
rect 72165 786383 72221 786439
rect 72307 786383 72363 786439
rect 72449 786383 72505 786439
rect 72591 786383 72647 786439
rect 72733 786383 72789 786439
rect 72875 786383 72931 786439
rect 73017 786383 73073 786439
rect 73159 786383 73215 786439
rect 73301 786383 73357 786439
rect 71455 786241 71511 786297
rect 71597 786241 71653 786297
rect 71739 786241 71795 786297
rect 71881 786241 71937 786297
rect 72023 786241 72079 786297
rect 72165 786241 72221 786297
rect 72307 786241 72363 786297
rect 72449 786241 72505 786297
rect 72591 786241 72647 786297
rect 72733 786241 72789 786297
rect 72875 786241 72931 786297
rect 73017 786241 73073 786297
rect 73159 786241 73215 786297
rect 73301 786241 73357 786297
rect 71455 786099 71511 786155
rect 71597 786099 71653 786155
rect 71739 786099 71795 786155
rect 71881 786099 71937 786155
rect 72023 786099 72079 786155
rect 72165 786099 72221 786155
rect 72307 786099 72363 786155
rect 72449 786099 72505 786155
rect 72591 786099 72647 786155
rect 72733 786099 72789 786155
rect 72875 786099 72931 786155
rect 73017 786099 73073 786155
rect 73159 786099 73215 786155
rect 73301 786099 73357 786155
rect 71455 785957 71511 786013
rect 71597 785957 71653 786013
rect 71739 785957 71795 786013
rect 71881 785957 71937 786013
rect 72023 785957 72079 786013
rect 72165 785957 72221 786013
rect 72307 785957 72363 786013
rect 72449 785957 72505 786013
rect 72591 785957 72647 786013
rect 72733 785957 72789 786013
rect 72875 785957 72931 786013
rect 73017 785957 73073 786013
rect 73159 785957 73215 786013
rect 73301 785957 73357 786013
rect 71455 785815 71511 785871
rect 71597 785815 71653 785871
rect 71739 785815 71795 785871
rect 71881 785815 71937 785871
rect 72023 785815 72079 785871
rect 72165 785815 72221 785871
rect 72307 785815 72363 785871
rect 72449 785815 72505 785871
rect 72591 785815 72647 785871
rect 72733 785815 72789 785871
rect 72875 785815 72931 785871
rect 73017 785815 73073 785871
rect 73159 785815 73215 785871
rect 73301 785815 73357 785871
rect 71455 785673 71511 785729
rect 71597 785673 71653 785729
rect 71739 785673 71795 785729
rect 71881 785673 71937 785729
rect 72023 785673 72079 785729
rect 72165 785673 72221 785729
rect 72307 785673 72363 785729
rect 72449 785673 72505 785729
rect 72591 785673 72647 785729
rect 72733 785673 72789 785729
rect 72875 785673 72931 785729
rect 73017 785673 73073 785729
rect 73159 785673 73215 785729
rect 73301 785673 73357 785729
rect 71455 785531 71511 785587
rect 71597 785531 71653 785587
rect 71739 785531 71795 785587
rect 71881 785531 71937 785587
rect 72023 785531 72079 785587
rect 72165 785531 72221 785587
rect 72307 785531 72363 785587
rect 72449 785531 72505 785587
rect 72591 785531 72647 785587
rect 72733 785531 72789 785587
rect 72875 785531 72931 785587
rect 73017 785531 73073 785587
rect 73159 785531 73215 785587
rect 73301 785531 73357 785587
rect 71455 785389 71511 785445
rect 71597 785389 71653 785445
rect 71739 785389 71795 785445
rect 71881 785389 71937 785445
rect 72023 785389 72079 785445
rect 72165 785389 72221 785445
rect 72307 785389 72363 785445
rect 72449 785389 72505 785445
rect 72591 785389 72647 785445
rect 72733 785389 72789 785445
rect 72875 785389 72931 785445
rect 73017 785389 73073 785445
rect 73159 785389 73215 785445
rect 73301 785389 73357 785445
rect 71455 785247 71511 785303
rect 71597 785247 71653 785303
rect 71739 785247 71795 785303
rect 71881 785247 71937 785303
rect 72023 785247 72079 785303
rect 72165 785247 72221 785303
rect 72307 785247 72363 785303
rect 72449 785247 72505 785303
rect 72591 785247 72647 785303
rect 72733 785247 72789 785303
rect 72875 785247 72931 785303
rect 73017 785247 73073 785303
rect 73159 785247 73215 785303
rect 73301 785247 73357 785303
rect 71455 785105 71511 785161
rect 71597 785105 71653 785161
rect 71739 785105 71795 785161
rect 71881 785105 71937 785161
rect 72023 785105 72079 785161
rect 72165 785105 72221 785161
rect 72307 785105 72363 785161
rect 72449 785105 72505 785161
rect 72591 785105 72647 785161
rect 72733 785105 72789 785161
rect 72875 785105 72931 785161
rect 73017 785105 73073 785161
rect 73159 785105 73215 785161
rect 73301 785105 73357 785161
rect 71455 784963 71511 785019
rect 71597 784963 71653 785019
rect 71739 784963 71795 785019
rect 71881 784963 71937 785019
rect 72023 784963 72079 785019
rect 72165 784963 72221 785019
rect 72307 784963 72363 785019
rect 72449 784963 72505 785019
rect 72591 784963 72647 785019
rect 72733 784963 72789 785019
rect 72875 784963 72931 785019
rect 73017 784963 73073 785019
rect 73159 784963 73215 785019
rect 73301 784963 73357 785019
rect 71455 784821 71511 784877
rect 71597 784821 71653 784877
rect 71739 784821 71795 784877
rect 71881 784821 71937 784877
rect 72023 784821 72079 784877
rect 72165 784821 72221 784877
rect 72307 784821 72363 784877
rect 72449 784821 72505 784877
rect 72591 784821 72647 784877
rect 72733 784821 72789 784877
rect 72875 784821 72931 784877
rect 73017 784821 73073 784877
rect 73159 784821 73215 784877
rect 73301 784821 73357 784877
rect 700051 786753 700107 786809
rect 700193 786753 700249 786809
rect 700335 786753 700391 786809
rect 700477 786753 700533 786809
rect 700619 786753 700675 786809
rect 700761 786753 700817 786809
rect 700903 786753 700959 786809
rect 701045 786753 701101 786809
rect 701187 786753 701243 786809
rect 701329 786753 701385 786809
rect 701471 786753 701527 786809
rect 701613 786753 701669 786809
rect 701755 786753 701811 786809
rect 701897 786753 701953 786809
rect 700051 786611 700107 786667
rect 700193 786611 700249 786667
rect 700335 786611 700391 786667
rect 700477 786611 700533 786667
rect 700619 786611 700675 786667
rect 700761 786611 700817 786667
rect 700903 786611 700959 786667
rect 701045 786611 701101 786667
rect 701187 786611 701243 786667
rect 701329 786611 701385 786667
rect 701471 786611 701527 786667
rect 701613 786611 701669 786667
rect 701755 786611 701811 786667
rect 701897 786611 701953 786667
rect 700051 786469 700107 786525
rect 700193 786469 700249 786525
rect 700335 786469 700391 786525
rect 700477 786469 700533 786525
rect 700619 786469 700675 786525
rect 700761 786469 700817 786525
rect 700903 786469 700959 786525
rect 701045 786469 701101 786525
rect 701187 786469 701243 786525
rect 701329 786469 701385 786525
rect 701471 786469 701527 786525
rect 701613 786469 701669 786525
rect 701755 786469 701811 786525
rect 701897 786469 701953 786525
rect 700051 786327 700107 786383
rect 700193 786327 700249 786383
rect 700335 786327 700391 786383
rect 700477 786327 700533 786383
rect 700619 786327 700675 786383
rect 700761 786327 700817 786383
rect 700903 786327 700959 786383
rect 701045 786327 701101 786383
rect 701187 786327 701243 786383
rect 701329 786327 701385 786383
rect 701471 786327 701527 786383
rect 701613 786327 701669 786383
rect 701755 786327 701811 786383
rect 701897 786327 701953 786383
rect 700051 786185 700107 786241
rect 700193 786185 700249 786241
rect 700335 786185 700391 786241
rect 700477 786185 700533 786241
rect 700619 786185 700675 786241
rect 700761 786185 700817 786241
rect 700903 786185 700959 786241
rect 701045 786185 701101 786241
rect 701187 786185 701243 786241
rect 701329 786185 701385 786241
rect 701471 786185 701527 786241
rect 701613 786185 701669 786241
rect 701755 786185 701811 786241
rect 701897 786185 701953 786241
rect 700051 786043 700107 786099
rect 700193 786043 700249 786099
rect 700335 786043 700391 786099
rect 700477 786043 700533 786099
rect 700619 786043 700675 786099
rect 700761 786043 700817 786099
rect 700903 786043 700959 786099
rect 701045 786043 701101 786099
rect 701187 786043 701243 786099
rect 701329 786043 701385 786099
rect 701471 786043 701527 786099
rect 701613 786043 701669 786099
rect 701755 786043 701811 786099
rect 701897 786043 701953 786099
rect 700051 785901 700107 785957
rect 700193 785901 700249 785957
rect 700335 785901 700391 785957
rect 700477 785901 700533 785957
rect 700619 785901 700675 785957
rect 700761 785901 700817 785957
rect 700903 785901 700959 785957
rect 701045 785901 701101 785957
rect 701187 785901 701243 785957
rect 701329 785901 701385 785957
rect 701471 785901 701527 785957
rect 701613 785901 701669 785957
rect 701755 785901 701811 785957
rect 701897 785901 701953 785957
rect 700051 785759 700107 785815
rect 700193 785759 700249 785815
rect 700335 785759 700391 785815
rect 700477 785759 700533 785815
rect 700619 785759 700675 785815
rect 700761 785759 700817 785815
rect 700903 785759 700959 785815
rect 701045 785759 701101 785815
rect 701187 785759 701243 785815
rect 701329 785759 701385 785815
rect 701471 785759 701527 785815
rect 701613 785759 701669 785815
rect 701755 785759 701811 785815
rect 701897 785759 701953 785815
rect 700051 785617 700107 785673
rect 700193 785617 700249 785673
rect 700335 785617 700391 785673
rect 700477 785617 700533 785673
rect 700619 785617 700675 785673
rect 700761 785617 700817 785673
rect 700903 785617 700959 785673
rect 701045 785617 701101 785673
rect 701187 785617 701243 785673
rect 701329 785617 701385 785673
rect 701471 785617 701527 785673
rect 701613 785617 701669 785673
rect 701755 785617 701811 785673
rect 701897 785617 701953 785673
rect 700051 785475 700107 785531
rect 700193 785475 700249 785531
rect 700335 785475 700391 785531
rect 700477 785475 700533 785531
rect 700619 785475 700675 785531
rect 700761 785475 700817 785531
rect 700903 785475 700959 785531
rect 701045 785475 701101 785531
rect 701187 785475 701243 785531
rect 701329 785475 701385 785531
rect 701471 785475 701527 785531
rect 701613 785475 701669 785531
rect 701755 785475 701811 785531
rect 701897 785475 701953 785531
rect 700051 785333 700107 785389
rect 700193 785333 700249 785389
rect 700335 785333 700391 785389
rect 700477 785333 700533 785389
rect 700619 785333 700675 785389
rect 700761 785333 700817 785389
rect 700903 785333 700959 785389
rect 701045 785333 701101 785389
rect 701187 785333 701243 785389
rect 701329 785333 701385 785389
rect 701471 785333 701527 785389
rect 701613 785333 701669 785389
rect 701755 785333 701811 785389
rect 701897 785333 701953 785389
rect 700051 785191 700107 785247
rect 700193 785191 700249 785247
rect 700335 785191 700391 785247
rect 700477 785191 700533 785247
rect 700619 785191 700675 785247
rect 700761 785191 700817 785247
rect 700903 785191 700959 785247
rect 701045 785191 701101 785247
rect 701187 785191 701243 785247
rect 701329 785191 701385 785247
rect 701471 785191 701527 785247
rect 701613 785191 701669 785247
rect 701755 785191 701811 785247
rect 701897 785191 701953 785247
rect 700051 785049 700107 785105
rect 700193 785049 700249 785105
rect 700335 785049 700391 785105
rect 700477 785049 700533 785105
rect 700619 785049 700675 785105
rect 700761 785049 700817 785105
rect 700903 785049 700959 785105
rect 701045 785049 701101 785105
rect 701187 785049 701243 785105
rect 701329 785049 701385 785105
rect 701471 785049 701527 785105
rect 701613 785049 701669 785105
rect 701755 785049 701811 785105
rect 701897 785049 701953 785105
rect 700051 784907 700107 784963
rect 700193 784907 700249 784963
rect 700335 784907 700391 784963
rect 700477 784907 700533 784963
rect 700619 784907 700675 784963
rect 700761 784907 700817 784963
rect 700903 784907 700959 784963
rect 701045 784907 701101 784963
rect 701187 784907 701243 784963
rect 701329 784907 701385 784963
rect 701471 784907 701527 784963
rect 701613 784907 701669 784963
rect 701755 784907 701811 784963
rect 701897 784907 701953 784963
rect 71466 784038 71522 784094
rect 71608 784038 71664 784094
rect 71750 784038 71806 784094
rect 71892 784038 71948 784094
rect 72034 784038 72090 784094
rect 72176 784038 72232 784094
rect 72318 784038 72374 784094
rect 72460 784038 72516 784094
rect 72602 784038 72658 784094
rect 72744 784038 72800 784094
rect 72886 784038 72942 784094
rect 73028 784038 73084 784094
rect 73170 784038 73226 784094
rect 73312 784038 73368 784094
rect 71466 783896 71522 783952
rect 71608 783896 71664 783952
rect 71750 783896 71806 783952
rect 71892 783896 71948 783952
rect 72034 783896 72090 783952
rect 72176 783896 72232 783952
rect 72318 783896 72374 783952
rect 72460 783896 72516 783952
rect 72602 783896 72658 783952
rect 72744 783896 72800 783952
rect 72886 783896 72942 783952
rect 73028 783896 73084 783952
rect 73170 783896 73226 783952
rect 73312 783896 73368 783952
rect 71466 783754 71522 783810
rect 71608 783754 71664 783810
rect 71750 783754 71806 783810
rect 71892 783754 71948 783810
rect 72034 783754 72090 783810
rect 72176 783754 72232 783810
rect 72318 783754 72374 783810
rect 72460 783754 72516 783810
rect 72602 783754 72658 783810
rect 72744 783754 72800 783810
rect 72886 783754 72942 783810
rect 73028 783754 73084 783810
rect 73170 783754 73226 783810
rect 73312 783754 73368 783810
rect 71466 783612 71522 783668
rect 71608 783612 71664 783668
rect 71750 783612 71806 783668
rect 71892 783612 71948 783668
rect 72034 783612 72090 783668
rect 72176 783612 72232 783668
rect 72318 783612 72374 783668
rect 72460 783612 72516 783668
rect 72602 783612 72658 783668
rect 72744 783612 72800 783668
rect 72886 783612 72942 783668
rect 73028 783612 73084 783668
rect 73170 783612 73226 783668
rect 73312 783612 73368 783668
rect 71466 783470 71522 783526
rect 71608 783470 71664 783526
rect 71750 783470 71806 783526
rect 71892 783470 71948 783526
rect 72034 783470 72090 783526
rect 72176 783470 72232 783526
rect 72318 783470 72374 783526
rect 72460 783470 72516 783526
rect 72602 783470 72658 783526
rect 72744 783470 72800 783526
rect 72886 783470 72942 783526
rect 73028 783470 73084 783526
rect 73170 783470 73226 783526
rect 73312 783470 73368 783526
rect 71466 783328 71522 783384
rect 71608 783328 71664 783384
rect 71750 783328 71806 783384
rect 71892 783328 71948 783384
rect 72034 783328 72090 783384
rect 72176 783328 72232 783384
rect 72318 783328 72374 783384
rect 72460 783328 72516 783384
rect 72602 783328 72658 783384
rect 72744 783328 72800 783384
rect 72886 783328 72942 783384
rect 73028 783328 73084 783384
rect 73170 783328 73226 783384
rect 73312 783328 73368 783384
rect 71466 783186 71522 783242
rect 71608 783186 71664 783242
rect 71750 783186 71806 783242
rect 71892 783186 71948 783242
rect 72034 783186 72090 783242
rect 72176 783186 72232 783242
rect 72318 783186 72374 783242
rect 72460 783186 72516 783242
rect 72602 783186 72658 783242
rect 72744 783186 72800 783242
rect 72886 783186 72942 783242
rect 73028 783186 73084 783242
rect 73170 783186 73226 783242
rect 73312 783186 73368 783242
rect 71466 783044 71522 783100
rect 71608 783044 71664 783100
rect 71750 783044 71806 783100
rect 71892 783044 71948 783100
rect 72034 783044 72090 783100
rect 72176 783044 72232 783100
rect 72318 783044 72374 783100
rect 72460 783044 72516 783100
rect 72602 783044 72658 783100
rect 72744 783044 72800 783100
rect 72886 783044 72942 783100
rect 73028 783044 73084 783100
rect 73170 783044 73226 783100
rect 73312 783044 73368 783100
rect 71466 782902 71522 782958
rect 71608 782902 71664 782958
rect 71750 782902 71806 782958
rect 71892 782902 71948 782958
rect 72034 782902 72090 782958
rect 72176 782902 72232 782958
rect 72318 782902 72374 782958
rect 72460 782902 72516 782958
rect 72602 782902 72658 782958
rect 72744 782902 72800 782958
rect 72886 782902 72942 782958
rect 73028 782902 73084 782958
rect 73170 782902 73226 782958
rect 73312 782902 73368 782958
rect 71466 782760 71522 782816
rect 71608 782760 71664 782816
rect 71750 782760 71806 782816
rect 71892 782760 71948 782816
rect 72034 782760 72090 782816
rect 72176 782760 72232 782816
rect 72318 782760 72374 782816
rect 72460 782760 72516 782816
rect 72602 782760 72658 782816
rect 72744 782760 72800 782816
rect 72886 782760 72942 782816
rect 73028 782760 73084 782816
rect 73170 782760 73226 782816
rect 73312 782760 73368 782816
rect 71466 782618 71522 782674
rect 71608 782618 71664 782674
rect 71750 782618 71806 782674
rect 71892 782618 71948 782674
rect 72034 782618 72090 782674
rect 72176 782618 72232 782674
rect 72318 782618 72374 782674
rect 72460 782618 72516 782674
rect 72602 782618 72658 782674
rect 72744 782618 72800 782674
rect 72886 782618 72942 782674
rect 73028 782618 73084 782674
rect 73170 782618 73226 782674
rect 73312 782618 73368 782674
rect 71466 782476 71522 782532
rect 71608 782476 71664 782532
rect 71750 782476 71806 782532
rect 71892 782476 71948 782532
rect 72034 782476 72090 782532
rect 72176 782476 72232 782532
rect 72318 782476 72374 782532
rect 72460 782476 72516 782532
rect 72602 782476 72658 782532
rect 72744 782476 72800 782532
rect 72886 782476 72942 782532
rect 73028 782476 73084 782532
rect 73170 782476 73226 782532
rect 73312 782476 73368 782532
rect 71466 782334 71522 782390
rect 71608 782334 71664 782390
rect 71750 782334 71806 782390
rect 71892 782334 71948 782390
rect 72034 782334 72090 782390
rect 72176 782334 72232 782390
rect 72318 782334 72374 782390
rect 72460 782334 72516 782390
rect 72602 782334 72658 782390
rect 72744 782334 72800 782390
rect 72886 782334 72942 782390
rect 73028 782334 73084 782390
rect 73170 782334 73226 782390
rect 73312 782334 73368 782390
rect 700051 784047 700107 784103
rect 700193 784047 700249 784103
rect 700335 784047 700391 784103
rect 700477 784047 700533 784103
rect 700619 784047 700675 784103
rect 700761 784047 700817 784103
rect 700903 784047 700959 784103
rect 701045 784047 701101 784103
rect 701187 784047 701243 784103
rect 701329 784047 701385 784103
rect 701471 784047 701527 784103
rect 701613 784047 701669 784103
rect 701755 784047 701811 784103
rect 701897 784047 701953 784103
rect 700051 783905 700107 783961
rect 700193 783905 700249 783961
rect 700335 783905 700391 783961
rect 700477 783905 700533 783961
rect 700619 783905 700675 783961
rect 700761 783905 700817 783961
rect 700903 783905 700959 783961
rect 701045 783905 701101 783961
rect 701187 783905 701243 783961
rect 701329 783905 701385 783961
rect 701471 783905 701527 783961
rect 701613 783905 701669 783961
rect 701755 783905 701811 783961
rect 701897 783905 701953 783961
rect 700051 783763 700107 783819
rect 700193 783763 700249 783819
rect 700335 783763 700391 783819
rect 700477 783763 700533 783819
rect 700619 783763 700675 783819
rect 700761 783763 700817 783819
rect 700903 783763 700959 783819
rect 701045 783763 701101 783819
rect 701187 783763 701243 783819
rect 701329 783763 701385 783819
rect 701471 783763 701527 783819
rect 701613 783763 701669 783819
rect 701755 783763 701811 783819
rect 701897 783763 701953 783819
rect 700051 783621 700107 783677
rect 700193 783621 700249 783677
rect 700335 783621 700391 783677
rect 700477 783621 700533 783677
rect 700619 783621 700675 783677
rect 700761 783621 700817 783677
rect 700903 783621 700959 783677
rect 701045 783621 701101 783677
rect 701187 783621 701243 783677
rect 701329 783621 701385 783677
rect 701471 783621 701527 783677
rect 701613 783621 701669 783677
rect 701755 783621 701811 783677
rect 701897 783621 701953 783677
rect 700051 783479 700107 783535
rect 700193 783479 700249 783535
rect 700335 783479 700391 783535
rect 700477 783479 700533 783535
rect 700619 783479 700675 783535
rect 700761 783479 700817 783535
rect 700903 783479 700959 783535
rect 701045 783479 701101 783535
rect 701187 783479 701243 783535
rect 701329 783479 701385 783535
rect 701471 783479 701527 783535
rect 701613 783479 701669 783535
rect 701755 783479 701811 783535
rect 701897 783479 701953 783535
rect 700051 783337 700107 783393
rect 700193 783337 700249 783393
rect 700335 783337 700391 783393
rect 700477 783337 700533 783393
rect 700619 783337 700675 783393
rect 700761 783337 700817 783393
rect 700903 783337 700959 783393
rect 701045 783337 701101 783393
rect 701187 783337 701243 783393
rect 701329 783337 701385 783393
rect 701471 783337 701527 783393
rect 701613 783337 701669 783393
rect 701755 783337 701811 783393
rect 701897 783337 701953 783393
rect 700051 783195 700107 783251
rect 700193 783195 700249 783251
rect 700335 783195 700391 783251
rect 700477 783195 700533 783251
rect 700619 783195 700675 783251
rect 700761 783195 700817 783251
rect 700903 783195 700959 783251
rect 701045 783195 701101 783251
rect 701187 783195 701243 783251
rect 701329 783195 701385 783251
rect 701471 783195 701527 783251
rect 701613 783195 701669 783251
rect 701755 783195 701811 783251
rect 701897 783195 701953 783251
rect 700051 783053 700107 783109
rect 700193 783053 700249 783109
rect 700335 783053 700391 783109
rect 700477 783053 700533 783109
rect 700619 783053 700675 783109
rect 700761 783053 700817 783109
rect 700903 783053 700959 783109
rect 701045 783053 701101 783109
rect 701187 783053 701243 783109
rect 701329 783053 701385 783109
rect 701471 783053 701527 783109
rect 701613 783053 701669 783109
rect 701755 783053 701811 783109
rect 701897 783053 701953 783109
rect 700051 782911 700107 782967
rect 700193 782911 700249 782967
rect 700335 782911 700391 782967
rect 700477 782911 700533 782967
rect 700619 782911 700675 782967
rect 700761 782911 700817 782967
rect 700903 782911 700959 782967
rect 701045 782911 701101 782967
rect 701187 782911 701243 782967
rect 701329 782911 701385 782967
rect 701471 782911 701527 782967
rect 701613 782911 701669 782967
rect 701755 782911 701811 782967
rect 701897 782911 701953 782967
rect 700051 782769 700107 782825
rect 700193 782769 700249 782825
rect 700335 782769 700391 782825
rect 700477 782769 700533 782825
rect 700619 782769 700675 782825
rect 700761 782769 700817 782825
rect 700903 782769 700959 782825
rect 701045 782769 701101 782825
rect 701187 782769 701243 782825
rect 701329 782769 701385 782825
rect 701471 782769 701527 782825
rect 701613 782769 701669 782825
rect 701755 782769 701811 782825
rect 701897 782769 701953 782825
rect 700051 782627 700107 782683
rect 700193 782627 700249 782683
rect 700335 782627 700391 782683
rect 700477 782627 700533 782683
rect 700619 782627 700675 782683
rect 700761 782627 700817 782683
rect 700903 782627 700959 782683
rect 701045 782627 701101 782683
rect 701187 782627 701243 782683
rect 701329 782627 701385 782683
rect 701471 782627 701527 782683
rect 701613 782627 701669 782683
rect 701755 782627 701811 782683
rect 701897 782627 701953 782683
rect 700051 782485 700107 782541
rect 700193 782485 700249 782541
rect 700335 782485 700391 782541
rect 700477 782485 700533 782541
rect 700619 782485 700675 782541
rect 700761 782485 700817 782541
rect 700903 782485 700959 782541
rect 701045 782485 701101 782541
rect 701187 782485 701243 782541
rect 701329 782485 701385 782541
rect 701471 782485 701527 782541
rect 701613 782485 701669 782541
rect 701755 782485 701811 782541
rect 701897 782485 701953 782541
rect 700051 782343 700107 782399
rect 700193 782343 700249 782399
rect 700335 782343 700391 782399
rect 700477 782343 700533 782399
rect 700619 782343 700675 782399
rect 700761 782343 700817 782399
rect 700903 782343 700959 782399
rect 701045 782343 701101 782399
rect 701187 782343 701243 782399
rect 701329 782343 701385 782399
rect 701471 782343 701527 782399
rect 701613 782343 701669 782399
rect 701755 782343 701811 782399
rect 701897 782343 701953 782399
rect 700051 782201 700107 782257
rect 700193 782201 700249 782257
rect 700335 782201 700391 782257
rect 700477 782201 700533 782257
rect 700619 782201 700675 782257
rect 700761 782201 700817 782257
rect 700903 782201 700959 782257
rect 701045 782201 701101 782257
rect 701187 782201 701243 782257
rect 701329 782201 701385 782257
rect 701471 782201 701527 782257
rect 701613 782201 701669 782257
rect 701755 782201 701811 782257
rect 701897 782201 701953 782257
rect 700051 781677 700107 781733
rect 700193 781677 700249 781733
rect 700335 781677 700391 781733
rect 700477 781677 700533 781733
rect 700619 781677 700675 781733
rect 700761 781677 700817 781733
rect 700903 781677 700959 781733
rect 701045 781677 701101 781733
rect 701187 781677 701243 781733
rect 701329 781677 701385 781733
rect 701471 781677 701527 781733
rect 701613 781677 701669 781733
rect 701755 781677 701811 781733
rect 701897 781677 701953 781733
rect 700051 781535 700107 781591
rect 700193 781535 700249 781591
rect 700335 781535 700391 781591
rect 700477 781535 700533 781591
rect 700619 781535 700675 781591
rect 700761 781535 700817 781591
rect 700903 781535 700959 781591
rect 701045 781535 701101 781591
rect 701187 781535 701243 781591
rect 701329 781535 701385 781591
rect 701471 781535 701527 781591
rect 701613 781535 701669 781591
rect 701755 781535 701811 781591
rect 701897 781535 701953 781591
rect 700051 781393 700107 781449
rect 700193 781393 700249 781449
rect 700335 781393 700391 781449
rect 700477 781393 700533 781449
rect 700619 781393 700675 781449
rect 700761 781393 700817 781449
rect 700903 781393 700959 781449
rect 701045 781393 701101 781449
rect 701187 781393 701243 781449
rect 701329 781393 701385 781449
rect 701471 781393 701527 781449
rect 701613 781393 701669 781449
rect 701755 781393 701811 781449
rect 701897 781393 701953 781449
rect 700051 781251 700107 781307
rect 700193 781251 700249 781307
rect 700335 781251 700391 781307
rect 700477 781251 700533 781307
rect 700619 781251 700675 781307
rect 700761 781251 700817 781307
rect 700903 781251 700959 781307
rect 701045 781251 701101 781307
rect 701187 781251 701243 781307
rect 701329 781251 701385 781307
rect 701471 781251 701527 781307
rect 701613 781251 701669 781307
rect 701755 781251 701811 781307
rect 701897 781251 701953 781307
rect 700051 781109 700107 781165
rect 700193 781109 700249 781165
rect 700335 781109 700391 781165
rect 700477 781109 700533 781165
rect 700619 781109 700675 781165
rect 700761 781109 700817 781165
rect 700903 781109 700959 781165
rect 701045 781109 701101 781165
rect 701187 781109 701243 781165
rect 701329 781109 701385 781165
rect 701471 781109 701527 781165
rect 701613 781109 701669 781165
rect 701755 781109 701811 781165
rect 701897 781109 701953 781165
rect 700051 780967 700107 781023
rect 700193 780967 700249 781023
rect 700335 780967 700391 781023
rect 700477 780967 700533 781023
rect 700619 780967 700675 781023
rect 700761 780967 700817 781023
rect 700903 780967 700959 781023
rect 701045 780967 701101 781023
rect 701187 780967 701243 781023
rect 701329 780967 701385 781023
rect 701471 780967 701527 781023
rect 701613 780967 701669 781023
rect 701755 780967 701811 781023
rect 701897 780967 701953 781023
rect 700051 780825 700107 780881
rect 700193 780825 700249 780881
rect 700335 780825 700391 780881
rect 700477 780825 700533 780881
rect 700619 780825 700675 780881
rect 700761 780825 700817 780881
rect 700903 780825 700959 780881
rect 701045 780825 701101 780881
rect 701187 780825 701243 780881
rect 701329 780825 701385 780881
rect 701471 780825 701527 780881
rect 701613 780825 701669 780881
rect 701755 780825 701811 780881
rect 701897 780825 701953 780881
rect 700051 780683 700107 780739
rect 700193 780683 700249 780739
rect 700335 780683 700391 780739
rect 700477 780683 700533 780739
rect 700619 780683 700675 780739
rect 700761 780683 700817 780739
rect 700903 780683 700959 780739
rect 701045 780683 701101 780739
rect 701187 780683 701243 780739
rect 701329 780683 701385 780739
rect 701471 780683 701527 780739
rect 701613 780683 701669 780739
rect 701755 780683 701811 780739
rect 701897 780683 701953 780739
rect 700051 780541 700107 780597
rect 700193 780541 700249 780597
rect 700335 780541 700391 780597
rect 700477 780541 700533 780597
rect 700619 780541 700675 780597
rect 700761 780541 700817 780597
rect 700903 780541 700959 780597
rect 701045 780541 701101 780597
rect 701187 780541 701243 780597
rect 701329 780541 701385 780597
rect 701471 780541 701527 780597
rect 701613 780541 701669 780597
rect 701755 780541 701811 780597
rect 701897 780541 701953 780597
rect 700051 780399 700107 780455
rect 700193 780399 700249 780455
rect 700335 780399 700391 780455
rect 700477 780399 700533 780455
rect 700619 780399 700675 780455
rect 700761 780399 700817 780455
rect 700903 780399 700959 780455
rect 701045 780399 701101 780455
rect 701187 780399 701243 780455
rect 701329 780399 701385 780455
rect 701471 780399 701527 780455
rect 701613 780399 701669 780455
rect 701755 780399 701811 780455
rect 701897 780399 701953 780455
rect 700051 780257 700107 780313
rect 700193 780257 700249 780313
rect 700335 780257 700391 780313
rect 700477 780257 700533 780313
rect 700619 780257 700675 780313
rect 700761 780257 700817 780313
rect 700903 780257 700959 780313
rect 701045 780257 701101 780313
rect 701187 780257 701243 780313
rect 701329 780257 701385 780313
rect 701471 780257 701527 780313
rect 701613 780257 701669 780313
rect 701755 780257 701811 780313
rect 701897 780257 701953 780313
rect 700051 780115 700107 780171
rect 700193 780115 700249 780171
rect 700335 780115 700391 780171
rect 700477 780115 700533 780171
rect 700619 780115 700675 780171
rect 700761 780115 700817 780171
rect 700903 780115 700959 780171
rect 701045 780115 701101 780171
rect 701187 780115 701243 780171
rect 701329 780115 701385 780171
rect 701471 780115 701527 780171
rect 701613 780115 701669 780171
rect 701755 780115 701811 780171
rect 701897 780115 701953 780171
rect 700051 779973 700107 780029
rect 700193 779973 700249 780029
rect 700335 779973 700391 780029
rect 700477 779973 700533 780029
rect 700619 779973 700675 780029
rect 700761 779973 700817 780029
rect 700903 779973 700959 780029
rect 701045 779973 701101 780029
rect 701187 779973 701243 780029
rect 701329 779973 701385 780029
rect 701471 779973 701527 780029
rect 701613 779973 701669 780029
rect 701755 779973 701811 780029
rect 701897 779973 701953 780029
rect 700051 779831 700107 779887
rect 700193 779831 700249 779887
rect 700335 779831 700391 779887
rect 700477 779831 700533 779887
rect 700619 779831 700675 779887
rect 700761 779831 700817 779887
rect 700903 779831 700959 779887
rect 701045 779831 701101 779887
rect 701187 779831 701243 779887
rect 701329 779831 701385 779887
rect 701471 779831 701527 779887
rect 701613 779831 701669 779887
rect 701755 779831 701811 779887
rect 701897 779831 701953 779887
rect 700040 779054 700096 779110
rect 700182 779054 700238 779110
rect 700324 779054 700380 779110
rect 700466 779054 700522 779110
rect 700608 779054 700664 779110
rect 700750 779054 700806 779110
rect 700892 779054 700948 779110
rect 701034 779054 701090 779110
rect 701176 779054 701232 779110
rect 701318 779054 701374 779110
rect 701460 779054 701516 779110
rect 701602 779054 701658 779110
rect 701744 779054 701800 779110
rect 701886 779054 701942 779110
rect 700040 778912 700096 778968
rect 700182 778912 700238 778968
rect 700324 778912 700380 778968
rect 700466 778912 700522 778968
rect 700608 778912 700664 778968
rect 700750 778912 700806 778968
rect 700892 778912 700948 778968
rect 701034 778912 701090 778968
rect 701176 778912 701232 778968
rect 701318 778912 701374 778968
rect 701460 778912 701516 778968
rect 701602 778912 701658 778968
rect 701744 778912 701800 778968
rect 701886 778912 701942 778968
rect 700040 778770 700096 778826
rect 700182 778770 700238 778826
rect 700324 778770 700380 778826
rect 700466 778770 700522 778826
rect 700608 778770 700664 778826
rect 700750 778770 700806 778826
rect 700892 778770 700948 778826
rect 701034 778770 701090 778826
rect 701176 778770 701232 778826
rect 701318 778770 701374 778826
rect 701460 778770 701516 778826
rect 701602 778770 701658 778826
rect 701744 778770 701800 778826
rect 701886 778770 701942 778826
rect 700040 778628 700096 778684
rect 700182 778628 700238 778684
rect 700324 778628 700380 778684
rect 700466 778628 700522 778684
rect 700608 778628 700664 778684
rect 700750 778628 700806 778684
rect 700892 778628 700948 778684
rect 701034 778628 701090 778684
rect 701176 778628 701232 778684
rect 701318 778628 701374 778684
rect 701460 778628 701516 778684
rect 701602 778628 701658 778684
rect 701744 778628 701800 778684
rect 701886 778628 701942 778684
rect 700040 778486 700096 778542
rect 700182 778486 700238 778542
rect 700324 778486 700380 778542
rect 700466 778486 700522 778542
rect 700608 778486 700664 778542
rect 700750 778486 700806 778542
rect 700892 778486 700948 778542
rect 701034 778486 701090 778542
rect 701176 778486 701232 778542
rect 701318 778486 701374 778542
rect 701460 778486 701516 778542
rect 701602 778486 701658 778542
rect 701744 778486 701800 778542
rect 701886 778486 701942 778542
rect 700040 778344 700096 778400
rect 700182 778344 700238 778400
rect 700324 778344 700380 778400
rect 700466 778344 700522 778400
rect 700608 778344 700664 778400
rect 700750 778344 700806 778400
rect 700892 778344 700948 778400
rect 701034 778344 701090 778400
rect 701176 778344 701232 778400
rect 701318 778344 701374 778400
rect 701460 778344 701516 778400
rect 701602 778344 701658 778400
rect 701744 778344 701800 778400
rect 701886 778344 701942 778400
rect 700040 778202 700096 778258
rect 700182 778202 700238 778258
rect 700324 778202 700380 778258
rect 700466 778202 700522 778258
rect 700608 778202 700664 778258
rect 700750 778202 700806 778258
rect 700892 778202 700948 778258
rect 701034 778202 701090 778258
rect 701176 778202 701232 778258
rect 701318 778202 701374 778258
rect 701460 778202 701516 778258
rect 701602 778202 701658 778258
rect 701744 778202 701800 778258
rect 701886 778202 701942 778258
rect 700040 778060 700096 778116
rect 700182 778060 700238 778116
rect 700324 778060 700380 778116
rect 700466 778060 700522 778116
rect 700608 778060 700664 778116
rect 700750 778060 700806 778116
rect 700892 778060 700948 778116
rect 701034 778060 701090 778116
rect 701176 778060 701232 778116
rect 701318 778060 701374 778116
rect 701460 778060 701516 778116
rect 701602 778060 701658 778116
rect 701744 778060 701800 778116
rect 701886 778060 701942 778116
rect 700040 777918 700096 777974
rect 700182 777918 700238 777974
rect 700324 777918 700380 777974
rect 700466 777918 700522 777974
rect 700608 777918 700664 777974
rect 700750 777918 700806 777974
rect 700892 777918 700948 777974
rect 701034 777918 701090 777974
rect 701176 777918 701232 777974
rect 701318 777918 701374 777974
rect 701460 777918 701516 777974
rect 701602 777918 701658 777974
rect 701744 777918 701800 777974
rect 701886 777918 701942 777974
rect 700040 777776 700096 777832
rect 700182 777776 700238 777832
rect 700324 777776 700380 777832
rect 700466 777776 700522 777832
rect 700608 777776 700664 777832
rect 700750 777776 700806 777832
rect 700892 777776 700948 777832
rect 701034 777776 701090 777832
rect 701176 777776 701232 777832
rect 701318 777776 701374 777832
rect 701460 777776 701516 777832
rect 701602 777776 701658 777832
rect 701744 777776 701800 777832
rect 701886 777776 701942 777832
rect 700040 777634 700096 777690
rect 700182 777634 700238 777690
rect 700324 777634 700380 777690
rect 700466 777634 700522 777690
rect 700608 777634 700664 777690
rect 700750 777634 700806 777690
rect 700892 777634 700948 777690
rect 701034 777634 701090 777690
rect 701176 777634 701232 777690
rect 701318 777634 701374 777690
rect 701460 777634 701516 777690
rect 701602 777634 701658 777690
rect 701744 777634 701800 777690
rect 701886 777634 701942 777690
rect 700040 777492 700096 777548
rect 700182 777492 700238 777548
rect 700324 777492 700380 777548
rect 700466 777492 700522 777548
rect 700608 777492 700664 777548
rect 700750 777492 700806 777548
rect 700892 777492 700948 777548
rect 701034 777492 701090 777548
rect 701176 777492 701232 777548
rect 701318 777492 701374 777548
rect 701460 777492 701516 777548
rect 701602 777492 701658 777548
rect 701744 777492 701800 777548
rect 701886 777492 701942 777548
rect 700040 777350 700096 777406
rect 700182 777350 700238 777406
rect 700324 777350 700380 777406
rect 700466 777350 700522 777406
rect 700608 777350 700664 777406
rect 700750 777350 700806 777406
rect 700892 777350 700948 777406
rect 701034 777350 701090 777406
rect 701176 777350 701232 777406
rect 701318 777350 701374 777406
rect 701460 777350 701516 777406
rect 701602 777350 701658 777406
rect 701744 777350 701800 777406
rect 701886 777350 701942 777406
rect 700040 490610 700096 490666
rect 700182 490610 700238 490666
rect 700324 490610 700380 490666
rect 700466 490610 700522 490666
rect 700608 490610 700664 490666
rect 700750 490610 700806 490666
rect 700892 490610 700948 490666
rect 701034 490610 701090 490666
rect 701176 490610 701232 490666
rect 701318 490610 701374 490666
rect 701460 490610 701516 490666
rect 701602 490610 701658 490666
rect 701744 490610 701800 490666
rect 701886 490610 701942 490666
rect 700040 490468 700096 490524
rect 700182 490468 700238 490524
rect 700324 490468 700380 490524
rect 700466 490468 700522 490524
rect 700608 490468 700664 490524
rect 700750 490468 700806 490524
rect 700892 490468 700948 490524
rect 701034 490468 701090 490524
rect 701176 490468 701232 490524
rect 701318 490468 701374 490524
rect 701460 490468 701516 490524
rect 701602 490468 701658 490524
rect 701744 490468 701800 490524
rect 701886 490468 701942 490524
rect 700040 490326 700096 490382
rect 700182 490326 700238 490382
rect 700324 490326 700380 490382
rect 700466 490326 700522 490382
rect 700608 490326 700664 490382
rect 700750 490326 700806 490382
rect 700892 490326 700948 490382
rect 701034 490326 701090 490382
rect 701176 490326 701232 490382
rect 701318 490326 701374 490382
rect 701460 490326 701516 490382
rect 701602 490326 701658 490382
rect 701744 490326 701800 490382
rect 701886 490326 701942 490382
rect 700040 490184 700096 490240
rect 700182 490184 700238 490240
rect 700324 490184 700380 490240
rect 700466 490184 700522 490240
rect 700608 490184 700664 490240
rect 700750 490184 700806 490240
rect 700892 490184 700948 490240
rect 701034 490184 701090 490240
rect 701176 490184 701232 490240
rect 701318 490184 701374 490240
rect 701460 490184 701516 490240
rect 701602 490184 701658 490240
rect 701744 490184 701800 490240
rect 701886 490184 701942 490240
rect 700040 490042 700096 490098
rect 700182 490042 700238 490098
rect 700324 490042 700380 490098
rect 700466 490042 700522 490098
rect 700608 490042 700664 490098
rect 700750 490042 700806 490098
rect 700892 490042 700948 490098
rect 701034 490042 701090 490098
rect 701176 490042 701232 490098
rect 701318 490042 701374 490098
rect 701460 490042 701516 490098
rect 701602 490042 701658 490098
rect 701744 490042 701800 490098
rect 701886 490042 701942 490098
rect 700040 489900 700096 489956
rect 700182 489900 700238 489956
rect 700324 489900 700380 489956
rect 700466 489900 700522 489956
rect 700608 489900 700664 489956
rect 700750 489900 700806 489956
rect 700892 489900 700948 489956
rect 701034 489900 701090 489956
rect 701176 489900 701232 489956
rect 701318 489900 701374 489956
rect 701460 489900 701516 489956
rect 701602 489900 701658 489956
rect 701744 489900 701800 489956
rect 701886 489900 701942 489956
rect 700040 489758 700096 489814
rect 700182 489758 700238 489814
rect 700324 489758 700380 489814
rect 700466 489758 700522 489814
rect 700608 489758 700664 489814
rect 700750 489758 700806 489814
rect 700892 489758 700948 489814
rect 701034 489758 701090 489814
rect 701176 489758 701232 489814
rect 701318 489758 701374 489814
rect 701460 489758 701516 489814
rect 701602 489758 701658 489814
rect 701744 489758 701800 489814
rect 701886 489758 701942 489814
rect 700040 489616 700096 489672
rect 700182 489616 700238 489672
rect 700324 489616 700380 489672
rect 700466 489616 700522 489672
rect 700608 489616 700664 489672
rect 700750 489616 700806 489672
rect 700892 489616 700948 489672
rect 701034 489616 701090 489672
rect 701176 489616 701232 489672
rect 701318 489616 701374 489672
rect 701460 489616 701516 489672
rect 701602 489616 701658 489672
rect 701744 489616 701800 489672
rect 701886 489616 701942 489672
rect 700040 489474 700096 489530
rect 700182 489474 700238 489530
rect 700324 489474 700380 489530
rect 700466 489474 700522 489530
rect 700608 489474 700664 489530
rect 700750 489474 700806 489530
rect 700892 489474 700948 489530
rect 701034 489474 701090 489530
rect 701176 489474 701232 489530
rect 701318 489474 701374 489530
rect 701460 489474 701516 489530
rect 701602 489474 701658 489530
rect 701744 489474 701800 489530
rect 701886 489474 701942 489530
rect 700040 489332 700096 489388
rect 700182 489332 700238 489388
rect 700324 489332 700380 489388
rect 700466 489332 700522 489388
rect 700608 489332 700664 489388
rect 700750 489332 700806 489388
rect 700892 489332 700948 489388
rect 701034 489332 701090 489388
rect 701176 489332 701232 489388
rect 701318 489332 701374 489388
rect 701460 489332 701516 489388
rect 701602 489332 701658 489388
rect 701744 489332 701800 489388
rect 701886 489332 701942 489388
rect 700040 489190 700096 489246
rect 700182 489190 700238 489246
rect 700324 489190 700380 489246
rect 700466 489190 700522 489246
rect 700608 489190 700664 489246
rect 700750 489190 700806 489246
rect 700892 489190 700948 489246
rect 701034 489190 701090 489246
rect 701176 489190 701232 489246
rect 701318 489190 701374 489246
rect 701460 489190 701516 489246
rect 701602 489190 701658 489246
rect 701744 489190 701800 489246
rect 701886 489190 701942 489246
rect 700040 489048 700096 489104
rect 700182 489048 700238 489104
rect 700324 489048 700380 489104
rect 700466 489048 700522 489104
rect 700608 489048 700664 489104
rect 700750 489048 700806 489104
rect 700892 489048 700948 489104
rect 701034 489048 701090 489104
rect 701176 489048 701232 489104
rect 701318 489048 701374 489104
rect 701460 489048 701516 489104
rect 701602 489048 701658 489104
rect 701744 489048 701800 489104
rect 701886 489048 701942 489104
rect 700040 488906 700096 488962
rect 700182 488906 700238 488962
rect 700324 488906 700380 488962
rect 700466 488906 700522 488962
rect 700608 488906 700664 488962
rect 700750 488906 700806 488962
rect 700892 488906 700948 488962
rect 701034 488906 701090 488962
rect 701176 488906 701232 488962
rect 701318 488906 701374 488962
rect 701460 488906 701516 488962
rect 701602 488906 701658 488962
rect 701744 488906 701800 488962
rect 701886 488906 701942 488962
rect 700051 488123 700107 488179
rect 700193 488123 700249 488179
rect 700335 488123 700391 488179
rect 700477 488123 700533 488179
rect 700619 488123 700675 488179
rect 700761 488123 700817 488179
rect 700903 488123 700959 488179
rect 701045 488123 701101 488179
rect 701187 488123 701243 488179
rect 701329 488123 701385 488179
rect 701471 488123 701527 488179
rect 701613 488123 701669 488179
rect 701755 488123 701811 488179
rect 701897 488123 701953 488179
rect 700051 487981 700107 488037
rect 700193 487981 700249 488037
rect 700335 487981 700391 488037
rect 700477 487981 700533 488037
rect 700619 487981 700675 488037
rect 700761 487981 700817 488037
rect 700903 487981 700959 488037
rect 701045 487981 701101 488037
rect 701187 487981 701243 488037
rect 701329 487981 701385 488037
rect 701471 487981 701527 488037
rect 701613 487981 701669 488037
rect 701755 487981 701811 488037
rect 701897 487981 701953 488037
rect 700051 487839 700107 487895
rect 700193 487839 700249 487895
rect 700335 487839 700391 487895
rect 700477 487839 700533 487895
rect 700619 487839 700675 487895
rect 700761 487839 700817 487895
rect 700903 487839 700959 487895
rect 701045 487839 701101 487895
rect 701187 487839 701243 487895
rect 701329 487839 701385 487895
rect 701471 487839 701527 487895
rect 701613 487839 701669 487895
rect 701755 487839 701811 487895
rect 701897 487839 701953 487895
rect 700051 487697 700107 487753
rect 700193 487697 700249 487753
rect 700335 487697 700391 487753
rect 700477 487697 700533 487753
rect 700619 487697 700675 487753
rect 700761 487697 700817 487753
rect 700903 487697 700959 487753
rect 701045 487697 701101 487753
rect 701187 487697 701243 487753
rect 701329 487697 701385 487753
rect 701471 487697 701527 487753
rect 701613 487697 701669 487753
rect 701755 487697 701811 487753
rect 701897 487697 701953 487753
rect 700051 487555 700107 487611
rect 700193 487555 700249 487611
rect 700335 487555 700391 487611
rect 700477 487555 700533 487611
rect 700619 487555 700675 487611
rect 700761 487555 700817 487611
rect 700903 487555 700959 487611
rect 701045 487555 701101 487611
rect 701187 487555 701243 487611
rect 701329 487555 701385 487611
rect 701471 487555 701527 487611
rect 701613 487555 701669 487611
rect 701755 487555 701811 487611
rect 701897 487555 701953 487611
rect 700051 487413 700107 487469
rect 700193 487413 700249 487469
rect 700335 487413 700391 487469
rect 700477 487413 700533 487469
rect 700619 487413 700675 487469
rect 700761 487413 700817 487469
rect 700903 487413 700959 487469
rect 701045 487413 701101 487469
rect 701187 487413 701243 487469
rect 701329 487413 701385 487469
rect 701471 487413 701527 487469
rect 701613 487413 701669 487469
rect 701755 487413 701811 487469
rect 701897 487413 701953 487469
rect 700051 487271 700107 487327
rect 700193 487271 700249 487327
rect 700335 487271 700391 487327
rect 700477 487271 700533 487327
rect 700619 487271 700675 487327
rect 700761 487271 700817 487327
rect 700903 487271 700959 487327
rect 701045 487271 701101 487327
rect 701187 487271 701243 487327
rect 701329 487271 701385 487327
rect 701471 487271 701527 487327
rect 701613 487271 701669 487327
rect 701755 487271 701811 487327
rect 701897 487271 701953 487327
rect 700051 487129 700107 487185
rect 700193 487129 700249 487185
rect 700335 487129 700391 487185
rect 700477 487129 700533 487185
rect 700619 487129 700675 487185
rect 700761 487129 700817 487185
rect 700903 487129 700959 487185
rect 701045 487129 701101 487185
rect 701187 487129 701243 487185
rect 701329 487129 701385 487185
rect 701471 487129 701527 487185
rect 701613 487129 701669 487185
rect 701755 487129 701811 487185
rect 701897 487129 701953 487185
rect 700051 486987 700107 487043
rect 700193 486987 700249 487043
rect 700335 486987 700391 487043
rect 700477 486987 700533 487043
rect 700619 486987 700675 487043
rect 700761 486987 700817 487043
rect 700903 486987 700959 487043
rect 701045 486987 701101 487043
rect 701187 486987 701243 487043
rect 701329 486987 701385 487043
rect 701471 486987 701527 487043
rect 701613 486987 701669 487043
rect 701755 486987 701811 487043
rect 701897 486987 701953 487043
rect 700051 486845 700107 486901
rect 700193 486845 700249 486901
rect 700335 486845 700391 486901
rect 700477 486845 700533 486901
rect 700619 486845 700675 486901
rect 700761 486845 700817 486901
rect 700903 486845 700959 486901
rect 701045 486845 701101 486901
rect 701187 486845 701243 486901
rect 701329 486845 701385 486901
rect 701471 486845 701527 486901
rect 701613 486845 701669 486901
rect 701755 486845 701811 486901
rect 701897 486845 701953 486901
rect 700051 486703 700107 486759
rect 700193 486703 700249 486759
rect 700335 486703 700391 486759
rect 700477 486703 700533 486759
rect 700619 486703 700675 486759
rect 700761 486703 700817 486759
rect 700903 486703 700959 486759
rect 701045 486703 701101 486759
rect 701187 486703 701243 486759
rect 701329 486703 701385 486759
rect 701471 486703 701527 486759
rect 701613 486703 701669 486759
rect 701755 486703 701811 486759
rect 701897 486703 701953 486759
rect 700051 486561 700107 486617
rect 700193 486561 700249 486617
rect 700335 486561 700391 486617
rect 700477 486561 700533 486617
rect 700619 486561 700675 486617
rect 700761 486561 700817 486617
rect 700903 486561 700959 486617
rect 701045 486561 701101 486617
rect 701187 486561 701243 486617
rect 701329 486561 701385 486617
rect 701471 486561 701527 486617
rect 701613 486561 701669 486617
rect 701755 486561 701811 486617
rect 701897 486561 701953 486617
rect 700051 486419 700107 486475
rect 700193 486419 700249 486475
rect 700335 486419 700391 486475
rect 700477 486419 700533 486475
rect 700619 486419 700675 486475
rect 700761 486419 700817 486475
rect 700903 486419 700959 486475
rect 701045 486419 701101 486475
rect 701187 486419 701243 486475
rect 701329 486419 701385 486475
rect 701471 486419 701527 486475
rect 701613 486419 701669 486475
rect 701755 486419 701811 486475
rect 701897 486419 701953 486475
rect 700051 486277 700107 486333
rect 700193 486277 700249 486333
rect 700335 486277 700391 486333
rect 700477 486277 700533 486333
rect 700619 486277 700675 486333
rect 700761 486277 700817 486333
rect 700903 486277 700959 486333
rect 701045 486277 701101 486333
rect 701187 486277 701243 486333
rect 701329 486277 701385 486333
rect 701471 486277 701527 486333
rect 701613 486277 701669 486333
rect 701755 486277 701811 486333
rect 701897 486277 701953 486333
rect 700051 485753 700107 485809
rect 700193 485753 700249 485809
rect 700335 485753 700391 485809
rect 700477 485753 700533 485809
rect 700619 485753 700675 485809
rect 700761 485753 700817 485809
rect 700903 485753 700959 485809
rect 701045 485753 701101 485809
rect 701187 485753 701243 485809
rect 701329 485753 701385 485809
rect 701471 485753 701527 485809
rect 701613 485753 701669 485809
rect 701755 485753 701811 485809
rect 701897 485753 701953 485809
rect 700051 485611 700107 485667
rect 700193 485611 700249 485667
rect 700335 485611 700391 485667
rect 700477 485611 700533 485667
rect 700619 485611 700675 485667
rect 700761 485611 700817 485667
rect 700903 485611 700959 485667
rect 701045 485611 701101 485667
rect 701187 485611 701243 485667
rect 701329 485611 701385 485667
rect 701471 485611 701527 485667
rect 701613 485611 701669 485667
rect 701755 485611 701811 485667
rect 701897 485611 701953 485667
rect 700051 485469 700107 485525
rect 700193 485469 700249 485525
rect 700335 485469 700391 485525
rect 700477 485469 700533 485525
rect 700619 485469 700675 485525
rect 700761 485469 700817 485525
rect 700903 485469 700959 485525
rect 701045 485469 701101 485525
rect 701187 485469 701243 485525
rect 701329 485469 701385 485525
rect 701471 485469 701527 485525
rect 701613 485469 701669 485525
rect 701755 485469 701811 485525
rect 701897 485469 701953 485525
rect 700051 485327 700107 485383
rect 700193 485327 700249 485383
rect 700335 485327 700391 485383
rect 700477 485327 700533 485383
rect 700619 485327 700675 485383
rect 700761 485327 700817 485383
rect 700903 485327 700959 485383
rect 701045 485327 701101 485383
rect 701187 485327 701243 485383
rect 701329 485327 701385 485383
rect 701471 485327 701527 485383
rect 701613 485327 701669 485383
rect 701755 485327 701811 485383
rect 701897 485327 701953 485383
rect 700051 485185 700107 485241
rect 700193 485185 700249 485241
rect 700335 485185 700391 485241
rect 700477 485185 700533 485241
rect 700619 485185 700675 485241
rect 700761 485185 700817 485241
rect 700903 485185 700959 485241
rect 701045 485185 701101 485241
rect 701187 485185 701243 485241
rect 701329 485185 701385 485241
rect 701471 485185 701527 485241
rect 701613 485185 701669 485241
rect 701755 485185 701811 485241
rect 701897 485185 701953 485241
rect 700051 485043 700107 485099
rect 700193 485043 700249 485099
rect 700335 485043 700391 485099
rect 700477 485043 700533 485099
rect 700619 485043 700675 485099
rect 700761 485043 700817 485099
rect 700903 485043 700959 485099
rect 701045 485043 701101 485099
rect 701187 485043 701243 485099
rect 701329 485043 701385 485099
rect 701471 485043 701527 485099
rect 701613 485043 701669 485099
rect 701755 485043 701811 485099
rect 701897 485043 701953 485099
rect 700051 484901 700107 484957
rect 700193 484901 700249 484957
rect 700335 484901 700391 484957
rect 700477 484901 700533 484957
rect 700619 484901 700675 484957
rect 700761 484901 700817 484957
rect 700903 484901 700959 484957
rect 701045 484901 701101 484957
rect 701187 484901 701243 484957
rect 701329 484901 701385 484957
rect 701471 484901 701527 484957
rect 701613 484901 701669 484957
rect 701755 484901 701811 484957
rect 701897 484901 701953 484957
rect 700051 484759 700107 484815
rect 700193 484759 700249 484815
rect 700335 484759 700391 484815
rect 700477 484759 700533 484815
rect 700619 484759 700675 484815
rect 700761 484759 700817 484815
rect 700903 484759 700959 484815
rect 701045 484759 701101 484815
rect 701187 484759 701243 484815
rect 701329 484759 701385 484815
rect 701471 484759 701527 484815
rect 701613 484759 701669 484815
rect 701755 484759 701811 484815
rect 701897 484759 701953 484815
rect 700051 484617 700107 484673
rect 700193 484617 700249 484673
rect 700335 484617 700391 484673
rect 700477 484617 700533 484673
rect 700619 484617 700675 484673
rect 700761 484617 700817 484673
rect 700903 484617 700959 484673
rect 701045 484617 701101 484673
rect 701187 484617 701243 484673
rect 701329 484617 701385 484673
rect 701471 484617 701527 484673
rect 701613 484617 701669 484673
rect 701755 484617 701811 484673
rect 701897 484617 701953 484673
rect 700051 484475 700107 484531
rect 700193 484475 700249 484531
rect 700335 484475 700391 484531
rect 700477 484475 700533 484531
rect 700619 484475 700675 484531
rect 700761 484475 700817 484531
rect 700903 484475 700959 484531
rect 701045 484475 701101 484531
rect 701187 484475 701243 484531
rect 701329 484475 701385 484531
rect 701471 484475 701527 484531
rect 701613 484475 701669 484531
rect 701755 484475 701811 484531
rect 701897 484475 701953 484531
rect 700051 484333 700107 484389
rect 700193 484333 700249 484389
rect 700335 484333 700391 484389
rect 700477 484333 700533 484389
rect 700619 484333 700675 484389
rect 700761 484333 700817 484389
rect 700903 484333 700959 484389
rect 701045 484333 701101 484389
rect 701187 484333 701243 484389
rect 701329 484333 701385 484389
rect 701471 484333 701527 484389
rect 701613 484333 701669 484389
rect 701755 484333 701811 484389
rect 701897 484333 701953 484389
rect 700051 484191 700107 484247
rect 700193 484191 700249 484247
rect 700335 484191 700391 484247
rect 700477 484191 700533 484247
rect 700619 484191 700675 484247
rect 700761 484191 700817 484247
rect 700903 484191 700959 484247
rect 701045 484191 701101 484247
rect 701187 484191 701243 484247
rect 701329 484191 701385 484247
rect 701471 484191 701527 484247
rect 701613 484191 701669 484247
rect 701755 484191 701811 484247
rect 701897 484191 701953 484247
rect 700051 484049 700107 484105
rect 700193 484049 700249 484105
rect 700335 484049 700391 484105
rect 700477 484049 700533 484105
rect 700619 484049 700675 484105
rect 700761 484049 700817 484105
rect 700903 484049 700959 484105
rect 701045 484049 701101 484105
rect 701187 484049 701243 484105
rect 701329 484049 701385 484105
rect 701471 484049 701527 484105
rect 701613 484049 701669 484105
rect 701755 484049 701811 484105
rect 701897 484049 701953 484105
rect 700051 483907 700107 483963
rect 700193 483907 700249 483963
rect 700335 483907 700391 483963
rect 700477 483907 700533 483963
rect 700619 483907 700675 483963
rect 700761 483907 700817 483963
rect 700903 483907 700959 483963
rect 701045 483907 701101 483963
rect 701187 483907 701243 483963
rect 701329 483907 701385 483963
rect 701471 483907 701527 483963
rect 701613 483907 701669 483963
rect 701755 483907 701811 483963
rect 701897 483907 701953 483963
rect 700051 483047 700107 483103
rect 700193 483047 700249 483103
rect 700335 483047 700391 483103
rect 700477 483047 700533 483103
rect 700619 483047 700675 483103
rect 700761 483047 700817 483103
rect 700903 483047 700959 483103
rect 701045 483047 701101 483103
rect 701187 483047 701243 483103
rect 701329 483047 701385 483103
rect 701471 483047 701527 483103
rect 701613 483047 701669 483103
rect 701755 483047 701811 483103
rect 701897 483047 701953 483103
rect 700051 482905 700107 482961
rect 700193 482905 700249 482961
rect 700335 482905 700391 482961
rect 700477 482905 700533 482961
rect 700619 482905 700675 482961
rect 700761 482905 700817 482961
rect 700903 482905 700959 482961
rect 701045 482905 701101 482961
rect 701187 482905 701243 482961
rect 701329 482905 701385 482961
rect 701471 482905 701527 482961
rect 701613 482905 701669 482961
rect 701755 482905 701811 482961
rect 701897 482905 701953 482961
rect 700051 482763 700107 482819
rect 700193 482763 700249 482819
rect 700335 482763 700391 482819
rect 700477 482763 700533 482819
rect 700619 482763 700675 482819
rect 700761 482763 700817 482819
rect 700903 482763 700959 482819
rect 701045 482763 701101 482819
rect 701187 482763 701243 482819
rect 701329 482763 701385 482819
rect 701471 482763 701527 482819
rect 701613 482763 701669 482819
rect 701755 482763 701811 482819
rect 701897 482763 701953 482819
rect 700051 482621 700107 482677
rect 700193 482621 700249 482677
rect 700335 482621 700391 482677
rect 700477 482621 700533 482677
rect 700619 482621 700675 482677
rect 700761 482621 700817 482677
rect 700903 482621 700959 482677
rect 701045 482621 701101 482677
rect 701187 482621 701243 482677
rect 701329 482621 701385 482677
rect 701471 482621 701527 482677
rect 701613 482621 701669 482677
rect 701755 482621 701811 482677
rect 701897 482621 701953 482677
rect 700051 482479 700107 482535
rect 700193 482479 700249 482535
rect 700335 482479 700391 482535
rect 700477 482479 700533 482535
rect 700619 482479 700675 482535
rect 700761 482479 700817 482535
rect 700903 482479 700959 482535
rect 701045 482479 701101 482535
rect 701187 482479 701243 482535
rect 701329 482479 701385 482535
rect 701471 482479 701527 482535
rect 701613 482479 701669 482535
rect 701755 482479 701811 482535
rect 701897 482479 701953 482535
rect 700051 482337 700107 482393
rect 700193 482337 700249 482393
rect 700335 482337 700391 482393
rect 700477 482337 700533 482393
rect 700619 482337 700675 482393
rect 700761 482337 700817 482393
rect 700903 482337 700959 482393
rect 701045 482337 701101 482393
rect 701187 482337 701243 482393
rect 701329 482337 701385 482393
rect 701471 482337 701527 482393
rect 701613 482337 701669 482393
rect 701755 482337 701811 482393
rect 701897 482337 701953 482393
rect 700051 482195 700107 482251
rect 700193 482195 700249 482251
rect 700335 482195 700391 482251
rect 700477 482195 700533 482251
rect 700619 482195 700675 482251
rect 700761 482195 700817 482251
rect 700903 482195 700959 482251
rect 701045 482195 701101 482251
rect 701187 482195 701243 482251
rect 701329 482195 701385 482251
rect 701471 482195 701527 482251
rect 701613 482195 701669 482251
rect 701755 482195 701811 482251
rect 701897 482195 701953 482251
rect 700051 482053 700107 482109
rect 700193 482053 700249 482109
rect 700335 482053 700391 482109
rect 700477 482053 700533 482109
rect 700619 482053 700675 482109
rect 700761 482053 700817 482109
rect 700903 482053 700959 482109
rect 701045 482053 701101 482109
rect 701187 482053 701243 482109
rect 701329 482053 701385 482109
rect 701471 482053 701527 482109
rect 701613 482053 701669 482109
rect 701755 482053 701811 482109
rect 701897 482053 701953 482109
rect 700051 481911 700107 481967
rect 700193 481911 700249 481967
rect 700335 481911 700391 481967
rect 700477 481911 700533 481967
rect 700619 481911 700675 481967
rect 700761 481911 700817 481967
rect 700903 481911 700959 481967
rect 701045 481911 701101 481967
rect 701187 481911 701243 481967
rect 701329 481911 701385 481967
rect 701471 481911 701527 481967
rect 701613 481911 701669 481967
rect 701755 481911 701811 481967
rect 701897 481911 701953 481967
rect 700051 481769 700107 481825
rect 700193 481769 700249 481825
rect 700335 481769 700391 481825
rect 700477 481769 700533 481825
rect 700619 481769 700675 481825
rect 700761 481769 700817 481825
rect 700903 481769 700959 481825
rect 701045 481769 701101 481825
rect 701187 481769 701243 481825
rect 701329 481769 701385 481825
rect 701471 481769 701527 481825
rect 701613 481769 701669 481825
rect 701755 481769 701811 481825
rect 701897 481769 701953 481825
rect 700051 481627 700107 481683
rect 700193 481627 700249 481683
rect 700335 481627 700391 481683
rect 700477 481627 700533 481683
rect 700619 481627 700675 481683
rect 700761 481627 700817 481683
rect 700903 481627 700959 481683
rect 701045 481627 701101 481683
rect 701187 481627 701243 481683
rect 701329 481627 701385 481683
rect 701471 481627 701527 481683
rect 701613 481627 701669 481683
rect 701755 481627 701811 481683
rect 701897 481627 701953 481683
rect 700051 481485 700107 481541
rect 700193 481485 700249 481541
rect 700335 481485 700391 481541
rect 700477 481485 700533 481541
rect 700619 481485 700675 481541
rect 700761 481485 700817 481541
rect 700903 481485 700959 481541
rect 701045 481485 701101 481541
rect 701187 481485 701243 481541
rect 701329 481485 701385 481541
rect 701471 481485 701527 481541
rect 701613 481485 701669 481541
rect 701755 481485 701811 481541
rect 701897 481485 701953 481541
rect 700051 481343 700107 481399
rect 700193 481343 700249 481399
rect 700335 481343 700391 481399
rect 700477 481343 700533 481399
rect 700619 481343 700675 481399
rect 700761 481343 700817 481399
rect 700903 481343 700959 481399
rect 701045 481343 701101 481399
rect 701187 481343 701243 481399
rect 701329 481343 701385 481399
rect 701471 481343 701527 481399
rect 701613 481343 701669 481399
rect 701755 481343 701811 481399
rect 701897 481343 701953 481399
rect 700051 481201 700107 481257
rect 700193 481201 700249 481257
rect 700335 481201 700391 481257
rect 700477 481201 700533 481257
rect 700619 481201 700675 481257
rect 700761 481201 700817 481257
rect 700903 481201 700959 481257
rect 701045 481201 701101 481257
rect 701187 481201 701243 481257
rect 701329 481201 701385 481257
rect 701471 481201 701527 481257
rect 701613 481201 701669 481257
rect 701755 481201 701811 481257
rect 701897 481201 701953 481257
rect 700051 480677 700107 480733
rect 700193 480677 700249 480733
rect 700335 480677 700391 480733
rect 700477 480677 700533 480733
rect 700619 480677 700675 480733
rect 700761 480677 700817 480733
rect 700903 480677 700959 480733
rect 701045 480677 701101 480733
rect 701187 480677 701243 480733
rect 701329 480677 701385 480733
rect 701471 480677 701527 480733
rect 701613 480677 701669 480733
rect 701755 480677 701811 480733
rect 701897 480677 701953 480733
rect 700051 480535 700107 480591
rect 700193 480535 700249 480591
rect 700335 480535 700391 480591
rect 700477 480535 700533 480591
rect 700619 480535 700675 480591
rect 700761 480535 700817 480591
rect 700903 480535 700959 480591
rect 701045 480535 701101 480591
rect 701187 480535 701243 480591
rect 701329 480535 701385 480591
rect 701471 480535 701527 480591
rect 701613 480535 701669 480591
rect 701755 480535 701811 480591
rect 701897 480535 701953 480591
rect 700051 480393 700107 480449
rect 700193 480393 700249 480449
rect 700335 480393 700391 480449
rect 700477 480393 700533 480449
rect 700619 480393 700675 480449
rect 700761 480393 700817 480449
rect 700903 480393 700959 480449
rect 701045 480393 701101 480449
rect 701187 480393 701243 480449
rect 701329 480393 701385 480449
rect 701471 480393 701527 480449
rect 701613 480393 701669 480449
rect 701755 480393 701811 480449
rect 701897 480393 701953 480449
rect 700051 480251 700107 480307
rect 700193 480251 700249 480307
rect 700335 480251 700391 480307
rect 700477 480251 700533 480307
rect 700619 480251 700675 480307
rect 700761 480251 700817 480307
rect 700903 480251 700959 480307
rect 701045 480251 701101 480307
rect 701187 480251 701243 480307
rect 701329 480251 701385 480307
rect 701471 480251 701527 480307
rect 701613 480251 701669 480307
rect 701755 480251 701811 480307
rect 701897 480251 701953 480307
rect 700051 480109 700107 480165
rect 700193 480109 700249 480165
rect 700335 480109 700391 480165
rect 700477 480109 700533 480165
rect 700619 480109 700675 480165
rect 700761 480109 700817 480165
rect 700903 480109 700959 480165
rect 701045 480109 701101 480165
rect 701187 480109 701243 480165
rect 701329 480109 701385 480165
rect 701471 480109 701527 480165
rect 701613 480109 701669 480165
rect 701755 480109 701811 480165
rect 701897 480109 701953 480165
rect 700051 479967 700107 480023
rect 700193 479967 700249 480023
rect 700335 479967 700391 480023
rect 700477 479967 700533 480023
rect 700619 479967 700675 480023
rect 700761 479967 700817 480023
rect 700903 479967 700959 480023
rect 701045 479967 701101 480023
rect 701187 479967 701243 480023
rect 701329 479967 701385 480023
rect 701471 479967 701527 480023
rect 701613 479967 701669 480023
rect 701755 479967 701811 480023
rect 701897 479967 701953 480023
rect 700051 479825 700107 479881
rect 700193 479825 700249 479881
rect 700335 479825 700391 479881
rect 700477 479825 700533 479881
rect 700619 479825 700675 479881
rect 700761 479825 700817 479881
rect 700903 479825 700959 479881
rect 701045 479825 701101 479881
rect 701187 479825 701243 479881
rect 701329 479825 701385 479881
rect 701471 479825 701527 479881
rect 701613 479825 701669 479881
rect 701755 479825 701811 479881
rect 701897 479825 701953 479881
rect 700051 479683 700107 479739
rect 700193 479683 700249 479739
rect 700335 479683 700391 479739
rect 700477 479683 700533 479739
rect 700619 479683 700675 479739
rect 700761 479683 700817 479739
rect 700903 479683 700959 479739
rect 701045 479683 701101 479739
rect 701187 479683 701243 479739
rect 701329 479683 701385 479739
rect 701471 479683 701527 479739
rect 701613 479683 701669 479739
rect 701755 479683 701811 479739
rect 701897 479683 701953 479739
rect 700051 479541 700107 479597
rect 700193 479541 700249 479597
rect 700335 479541 700391 479597
rect 700477 479541 700533 479597
rect 700619 479541 700675 479597
rect 700761 479541 700817 479597
rect 700903 479541 700959 479597
rect 701045 479541 701101 479597
rect 701187 479541 701243 479597
rect 701329 479541 701385 479597
rect 701471 479541 701527 479597
rect 701613 479541 701669 479597
rect 701755 479541 701811 479597
rect 701897 479541 701953 479597
rect 700051 479399 700107 479455
rect 700193 479399 700249 479455
rect 700335 479399 700391 479455
rect 700477 479399 700533 479455
rect 700619 479399 700675 479455
rect 700761 479399 700817 479455
rect 700903 479399 700959 479455
rect 701045 479399 701101 479455
rect 701187 479399 701243 479455
rect 701329 479399 701385 479455
rect 701471 479399 701527 479455
rect 701613 479399 701669 479455
rect 701755 479399 701811 479455
rect 701897 479399 701953 479455
rect 700051 479257 700107 479313
rect 700193 479257 700249 479313
rect 700335 479257 700391 479313
rect 700477 479257 700533 479313
rect 700619 479257 700675 479313
rect 700761 479257 700817 479313
rect 700903 479257 700959 479313
rect 701045 479257 701101 479313
rect 701187 479257 701243 479313
rect 701329 479257 701385 479313
rect 701471 479257 701527 479313
rect 701613 479257 701669 479313
rect 701755 479257 701811 479313
rect 701897 479257 701953 479313
rect 700051 479115 700107 479171
rect 700193 479115 700249 479171
rect 700335 479115 700391 479171
rect 700477 479115 700533 479171
rect 700619 479115 700675 479171
rect 700761 479115 700817 479171
rect 700903 479115 700959 479171
rect 701045 479115 701101 479171
rect 701187 479115 701243 479171
rect 701329 479115 701385 479171
rect 701471 479115 701527 479171
rect 701613 479115 701669 479171
rect 701755 479115 701811 479171
rect 701897 479115 701953 479171
rect 700051 478973 700107 479029
rect 700193 478973 700249 479029
rect 700335 478973 700391 479029
rect 700477 478973 700533 479029
rect 700619 478973 700675 479029
rect 700761 478973 700817 479029
rect 700903 478973 700959 479029
rect 701045 478973 701101 479029
rect 701187 478973 701243 479029
rect 701329 478973 701385 479029
rect 701471 478973 701527 479029
rect 701613 478973 701669 479029
rect 701755 478973 701811 479029
rect 701897 478973 701953 479029
rect 700051 478831 700107 478887
rect 700193 478831 700249 478887
rect 700335 478831 700391 478887
rect 700477 478831 700533 478887
rect 700619 478831 700675 478887
rect 700761 478831 700817 478887
rect 700903 478831 700959 478887
rect 701045 478831 701101 478887
rect 701187 478831 701243 478887
rect 701329 478831 701385 478887
rect 701471 478831 701527 478887
rect 701613 478831 701669 478887
rect 701755 478831 701811 478887
rect 701897 478831 701953 478887
rect 700040 478054 700096 478110
rect 700182 478054 700238 478110
rect 700324 478054 700380 478110
rect 700466 478054 700522 478110
rect 700608 478054 700664 478110
rect 700750 478054 700806 478110
rect 700892 478054 700948 478110
rect 701034 478054 701090 478110
rect 701176 478054 701232 478110
rect 701318 478054 701374 478110
rect 701460 478054 701516 478110
rect 701602 478054 701658 478110
rect 701744 478054 701800 478110
rect 701886 478054 701942 478110
rect 700040 477912 700096 477968
rect 700182 477912 700238 477968
rect 700324 477912 700380 477968
rect 700466 477912 700522 477968
rect 700608 477912 700664 477968
rect 700750 477912 700806 477968
rect 700892 477912 700948 477968
rect 701034 477912 701090 477968
rect 701176 477912 701232 477968
rect 701318 477912 701374 477968
rect 701460 477912 701516 477968
rect 701602 477912 701658 477968
rect 701744 477912 701800 477968
rect 701886 477912 701942 477968
rect 700040 477770 700096 477826
rect 700182 477770 700238 477826
rect 700324 477770 700380 477826
rect 700466 477770 700522 477826
rect 700608 477770 700664 477826
rect 700750 477770 700806 477826
rect 700892 477770 700948 477826
rect 701034 477770 701090 477826
rect 701176 477770 701232 477826
rect 701318 477770 701374 477826
rect 701460 477770 701516 477826
rect 701602 477770 701658 477826
rect 701744 477770 701800 477826
rect 701886 477770 701942 477826
rect 700040 477628 700096 477684
rect 700182 477628 700238 477684
rect 700324 477628 700380 477684
rect 700466 477628 700522 477684
rect 700608 477628 700664 477684
rect 700750 477628 700806 477684
rect 700892 477628 700948 477684
rect 701034 477628 701090 477684
rect 701176 477628 701232 477684
rect 701318 477628 701374 477684
rect 701460 477628 701516 477684
rect 701602 477628 701658 477684
rect 701744 477628 701800 477684
rect 701886 477628 701942 477684
rect 700040 477486 700096 477542
rect 700182 477486 700238 477542
rect 700324 477486 700380 477542
rect 700466 477486 700522 477542
rect 700608 477486 700664 477542
rect 700750 477486 700806 477542
rect 700892 477486 700948 477542
rect 701034 477486 701090 477542
rect 701176 477486 701232 477542
rect 701318 477486 701374 477542
rect 701460 477486 701516 477542
rect 701602 477486 701658 477542
rect 701744 477486 701800 477542
rect 701886 477486 701942 477542
rect 700040 477344 700096 477400
rect 700182 477344 700238 477400
rect 700324 477344 700380 477400
rect 700466 477344 700522 477400
rect 700608 477344 700664 477400
rect 700750 477344 700806 477400
rect 700892 477344 700948 477400
rect 701034 477344 701090 477400
rect 701176 477344 701232 477400
rect 701318 477344 701374 477400
rect 701460 477344 701516 477400
rect 701602 477344 701658 477400
rect 701744 477344 701800 477400
rect 701886 477344 701942 477400
rect 700040 477202 700096 477258
rect 700182 477202 700238 477258
rect 700324 477202 700380 477258
rect 700466 477202 700522 477258
rect 700608 477202 700664 477258
rect 700750 477202 700806 477258
rect 700892 477202 700948 477258
rect 701034 477202 701090 477258
rect 701176 477202 701232 477258
rect 701318 477202 701374 477258
rect 701460 477202 701516 477258
rect 701602 477202 701658 477258
rect 701744 477202 701800 477258
rect 701886 477202 701942 477258
rect 700040 477060 700096 477116
rect 700182 477060 700238 477116
rect 700324 477060 700380 477116
rect 700466 477060 700522 477116
rect 700608 477060 700664 477116
rect 700750 477060 700806 477116
rect 700892 477060 700948 477116
rect 701034 477060 701090 477116
rect 701176 477060 701232 477116
rect 701318 477060 701374 477116
rect 701460 477060 701516 477116
rect 701602 477060 701658 477116
rect 701744 477060 701800 477116
rect 701886 477060 701942 477116
rect 700040 476918 700096 476974
rect 700182 476918 700238 476974
rect 700324 476918 700380 476974
rect 700466 476918 700522 476974
rect 700608 476918 700664 476974
rect 700750 476918 700806 476974
rect 700892 476918 700948 476974
rect 701034 476918 701090 476974
rect 701176 476918 701232 476974
rect 701318 476918 701374 476974
rect 701460 476918 701516 476974
rect 701602 476918 701658 476974
rect 701744 476918 701800 476974
rect 701886 476918 701942 476974
rect 700040 476776 700096 476832
rect 700182 476776 700238 476832
rect 700324 476776 700380 476832
rect 700466 476776 700522 476832
rect 700608 476776 700664 476832
rect 700750 476776 700806 476832
rect 700892 476776 700948 476832
rect 701034 476776 701090 476832
rect 701176 476776 701232 476832
rect 701318 476776 701374 476832
rect 701460 476776 701516 476832
rect 701602 476776 701658 476832
rect 701744 476776 701800 476832
rect 701886 476776 701942 476832
rect 700040 476634 700096 476690
rect 700182 476634 700238 476690
rect 700324 476634 700380 476690
rect 700466 476634 700522 476690
rect 700608 476634 700664 476690
rect 700750 476634 700806 476690
rect 700892 476634 700948 476690
rect 701034 476634 701090 476690
rect 701176 476634 701232 476690
rect 701318 476634 701374 476690
rect 701460 476634 701516 476690
rect 701602 476634 701658 476690
rect 701744 476634 701800 476690
rect 701886 476634 701942 476690
rect 700040 476492 700096 476548
rect 700182 476492 700238 476548
rect 700324 476492 700380 476548
rect 700466 476492 700522 476548
rect 700608 476492 700664 476548
rect 700750 476492 700806 476548
rect 700892 476492 700948 476548
rect 701034 476492 701090 476548
rect 701176 476492 701232 476548
rect 701318 476492 701374 476548
rect 701460 476492 701516 476548
rect 701602 476492 701658 476548
rect 701744 476492 701800 476548
rect 701886 476492 701942 476548
rect 700040 476350 700096 476406
rect 700182 476350 700238 476406
rect 700324 476350 700380 476406
rect 700466 476350 700522 476406
rect 700608 476350 700664 476406
rect 700750 476350 700806 476406
rect 700892 476350 700948 476406
rect 701034 476350 701090 476406
rect 701176 476350 701232 476406
rect 701318 476350 701374 476406
rect 701460 476350 701516 476406
rect 701602 476350 701658 476406
rect 701744 476350 701800 476406
rect 701886 476350 701942 476406
rect 73866 468594 73922 468650
rect 74008 468594 74064 468650
rect 74150 468594 74206 468650
rect 74292 468594 74348 468650
rect 74434 468594 74490 468650
rect 74576 468594 74632 468650
rect 74718 468594 74774 468650
rect 74860 468594 74916 468650
rect 75002 468594 75058 468650
rect 75144 468594 75200 468650
rect 75286 468594 75342 468650
rect 73866 468452 73922 468508
rect 74008 468452 74064 468508
rect 74150 468452 74206 468508
rect 74292 468452 74348 468508
rect 74434 468452 74490 468508
rect 74576 468452 74632 468508
rect 74718 468452 74774 468508
rect 74860 468452 74916 468508
rect 75002 468452 75058 468508
rect 75144 468452 75200 468508
rect 75286 468452 75342 468508
rect 73866 468310 73922 468366
rect 74008 468310 74064 468366
rect 74150 468310 74206 468366
rect 74292 468310 74348 468366
rect 74434 468310 74490 468366
rect 74576 468310 74632 468366
rect 74718 468310 74774 468366
rect 74860 468310 74916 468366
rect 75002 468310 75058 468366
rect 75144 468310 75200 468366
rect 75286 468310 75342 468366
rect 73866 468168 73922 468224
rect 74008 468168 74064 468224
rect 74150 468168 74206 468224
rect 74292 468168 74348 468224
rect 74434 468168 74490 468224
rect 74576 468168 74632 468224
rect 74718 468168 74774 468224
rect 74860 468168 74916 468224
rect 75002 468168 75058 468224
rect 75144 468168 75200 468224
rect 75286 468168 75342 468224
rect 73866 468026 73922 468082
rect 74008 468026 74064 468082
rect 74150 468026 74206 468082
rect 74292 468026 74348 468082
rect 74434 468026 74490 468082
rect 74576 468026 74632 468082
rect 74718 468026 74774 468082
rect 74860 468026 74916 468082
rect 75002 468026 75058 468082
rect 75144 468026 75200 468082
rect 75286 468026 75342 468082
rect 73866 467884 73922 467940
rect 74008 467884 74064 467940
rect 74150 467884 74206 467940
rect 74292 467884 74348 467940
rect 74434 467884 74490 467940
rect 74576 467884 74632 467940
rect 74718 467884 74774 467940
rect 74860 467884 74916 467940
rect 75002 467884 75058 467940
rect 75144 467884 75200 467940
rect 75286 467884 75342 467940
rect 73866 467742 73922 467798
rect 74008 467742 74064 467798
rect 74150 467742 74206 467798
rect 74292 467742 74348 467798
rect 74434 467742 74490 467798
rect 74576 467742 74632 467798
rect 74718 467742 74774 467798
rect 74860 467742 74916 467798
rect 75002 467742 75058 467798
rect 75144 467742 75200 467798
rect 75286 467742 75342 467798
rect 73866 467600 73922 467656
rect 74008 467600 74064 467656
rect 74150 467600 74206 467656
rect 74292 467600 74348 467656
rect 74434 467600 74490 467656
rect 74576 467600 74632 467656
rect 74718 467600 74774 467656
rect 74860 467600 74916 467656
rect 75002 467600 75058 467656
rect 75144 467600 75200 467656
rect 75286 467600 75342 467656
rect 73866 467458 73922 467514
rect 74008 467458 74064 467514
rect 74150 467458 74206 467514
rect 74292 467458 74348 467514
rect 74434 467458 74490 467514
rect 74576 467458 74632 467514
rect 74718 467458 74774 467514
rect 74860 467458 74916 467514
rect 75002 467458 75058 467514
rect 75144 467458 75200 467514
rect 75286 467458 75342 467514
rect 73866 467316 73922 467372
rect 74008 467316 74064 467372
rect 74150 467316 74206 467372
rect 74292 467316 74348 467372
rect 74434 467316 74490 467372
rect 74576 467316 74632 467372
rect 74718 467316 74774 467372
rect 74860 467316 74916 467372
rect 75002 467316 75058 467372
rect 75144 467316 75200 467372
rect 75286 467316 75342 467372
rect 73866 467174 73922 467230
rect 74008 467174 74064 467230
rect 74150 467174 74206 467230
rect 74292 467174 74348 467230
rect 74434 467174 74490 467230
rect 74576 467174 74632 467230
rect 74718 467174 74774 467230
rect 74860 467174 74916 467230
rect 75002 467174 75058 467230
rect 75144 467174 75200 467230
rect 75286 467174 75342 467230
rect 73866 467032 73922 467088
rect 74008 467032 74064 467088
rect 74150 467032 74206 467088
rect 74292 467032 74348 467088
rect 74434 467032 74490 467088
rect 74576 467032 74632 467088
rect 74718 467032 74774 467088
rect 74860 467032 74916 467088
rect 75002 467032 75058 467088
rect 75144 467032 75200 467088
rect 75286 467032 75342 467088
rect 73866 466890 73922 466946
rect 74008 466890 74064 466946
rect 74150 466890 74206 466946
rect 74292 466890 74348 466946
rect 74434 466890 74490 466946
rect 74576 466890 74632 466946
rect 74718 466890 74774 466946
rect 74860 466890 74916 466946
rect 75002 466890 75058 466946
rect 75144 466890 75200 466946
rect 75286 466890 75342 466946
rect 73855 466113 73911 466169
rect 73997 466113 74053 466169
rect 74139 466113 74195 466169
rect 74281 466113 74337 466169
rect 74423 466113 74479 466169
rect 74565 466113 74621 466169
rect 74707 466113 74763 466169
rect 74849 466113 74905 466169
rect 74991 466113 75047 466169
rect 75133 466113 75189 466169
rect 75275 466113 75331 466169
rect 73855 465971 73911 466027
rect 73997 465971 74053 466027
rect 74139 465971 74195 466027
rect 74281 465971 74337 466027
rect 74423 465971 74479 466027
rect 74565 465971 74621 466027
rect 74707 465971 74763 466027
rect 74849 465971 74905 466027
rect 74991 465971 75047 466027
rect 75133 465971 75189 466027
rect 75275 465971 75331 466027
rect 73855 465829 73911 465885
rect 73997 465829 74053 465885
rect 74139 465829 74195 465885
rect 74281 465829 74337 465885
rect 74423 465829 74479 465885
rect 74565 465829 74621 465885
rect 74707 465829 74763 465885
rect 74849 465829 74905 465885
rect 74991 465829 75047 465885
rect 75133 465829 75189 465885
rect 75275 465829 75331 465885
rect 73855 465687 73911 465743
rect 73997 465687 74053 465743
rect 74139 465687 74195 465743
rect 74281 465687 74337 465743
rect 74423 465687 74479 465743
rect 74565 465687 74621 465743
rect 74707 465687 74763 465743
rect 74849 465687 74905 465743
rect 74991 465687 75047 465743
rect 75133 465687 75189 465743
rect 75275 465687 75331 465743
rect 73855 465545 73911 465601
rect 73997 465545 74053 465601
rect 74139 465545 74195 465601
rect 74281 465545 74337 465601
rect 74423 465545 74479 465601
rect 74565 465545 74621 465601
rect 74707 465545 74763 465601
rect 74849 465545 74905 465601
rect 74991 465545 75047 465601
rect 75133 465545 75189 465601
rect 75275 465545 75331 465601
rect 73855 465403 73911 465459
rect 73997 465403 74053 465459
rect 74139 465403 74195 465459
rect 74281 465403 74337 465459
rect 74423 465403 74479 465459
rect 74565 465403 74621 465459
rect 74707 465403 74763 465459
rect 74849 465403 74905 465459
rect 74991 465403 75047 465459
rect 75133 465403 75189 465459
rect 75275 465403 75331 465459
rect 73855 465261 73911 465317
rect 73997 465261 74053 465317
rect 74139 465261 74195 465317
rect 74281 465261 74337 465317
rect 74423 465261 74479 465317
rect 74565 465261 74621 465317
rect 74707 465261 74763 465317
rect 74849 465261 74905 465317
rect 74991 465261 75047 465317
rect 75133 465261 75189 465317
rect 75275 465261 75331 465317
rect 73855 465119 73911 465175
rect 73997 465119 74053 465175
rect 74139 465119 74195 465175
rect 74281 465119 74337 465175
rect 74423 465119 74479 465175
rect 74565 465119 74621 465175
rect 74707 465119 74763 465175
rect 74849 465119 74905 465175
rect 74991 465119 75047 465175
rect 75133 465119 75189 465175
rect 75275 465119 75331 465175
rect 73855 464977 73911 465033
rect 73997 464977 74053 465033
rect 74139 464977 74195 465033
rect 74281 464977 74337 465033
rect 74423 464977 74479 465033
rect 74565 464977 74621 465033
rect 74707 464977 74763 465033
rect 74849 464977 74905 465033
rect 74991 464977 75047 465033
rect 75133 464977 75189 465033
rect 75275 464977 75331 465033
rect 73855 464835 73911 464891
rect 73997 464835 74053 464891
rect 74139 464835 74195 464891
rect 74281 464835 74337 464891
rect 74423 464835 74479 464891
rect 74565 464835 74621 464891
rect 74707 464835 74763 464891
rect 74849 464835 74905 464891
rect 74991 464835 75047 464891
rect 75133 464835 75189 464891
rect 75275 464835 75331 464891
rect 73855 464693 73911 464749
rect 73997 464693 74053 464749
rect 74139 464693 74195 464749
rect 74281 464693 74337 464749
rect 74423 464693 74479 464749
rect 74565 464693 74621 464749
rect 74707 464693 74763 464749
rect 74849 464693 74905 464749
rect 74991 464693 75047 464749
rect 75133 464693 75189 464749
rect 75275 464693 75331 464749
rect 73855 464551 73911 464607
rect 73997 464551 74053 464607
rect 74139 464551 74195 464607
rect 74281 464551 74337 464607
rect 74423 464551 74479 464607
rect 74565 464551 74621 464607
rect 74707 464551 74763 464607
rect 74849 464551 74905 464607
rect 74991 464551 75047 464607
rect 75133 464551 75189 464607
rect 75275 464551 75331 464607
rect 73855 464409 73911 464465
rect 73997 464409 74053 464465
rect 74139 464409 74195 464465
rect 74281 464409 74337 464465
rect 74423 464409 74479 464465
rect 74565 464409 74621 464465
rect 74707 464409 74763 464465
rect 74849 464409 74905 464465
rect 74991 464409 75047 464465
rect 75133 464409 75189 464465
rect 75275 464409 75331 464465
rect 73855 464267 73911 464323
rect 73997 464267 74053 464323
rect 74139 464267 74195 464323
rect 74281 464267 74337 464323
rect 74423 464267 74479 464323
rect 74565 464267 74621 464323
rect 74707 464267 74763 464323
rect 74849 464267 74905 464323
rect 74991 464267 75047 464323
rect 75133 464267 75189 464323
rect 75275 464267 75331 464323
rect 73855 463743 73911 463799
rect 73997 463743 74053 463799
rect 74139 463743 74195 463799
rect 74281 463743 74337 463799
rect 74423 463743 74479 463799
rect 74565 463743 74621 463799
rect 74707 463743 74763 463799
rect 74849 463743 74905 463799
rect 74991 463743 75047 463799
rect 75133 463743 75189 463799
rect 75275 463743 75331 463799
rect 73855 463601 73911 463657
rect 73997 463601 74053 463657
rect 74139 463601 74195 463657
rect 74281 463601 74337 463657
rect 74423 463601 74479 463657
rect 74565 463601 74621 463657
rect 74707 463601 74763 463657
rect 74849 463601 74905 463657
rect 74991 463601 75047 463657
rect 75133 463601 75189 463657
rect 75275 463601 75331 463657
rect 73855 463459 73911 463515
rect 73997 463459 74053 463515
rect 74139 463459 74195 463515
rect 74281 463459 74337 463515
rect 74423 463459 74479 463515
rect 74565 463459 74621 463515
rect 74707 463459 74763 463515
rect 74849 463459 74905 463515
rect 74991 463459 75047 463515
rect 75133 463459 75189 463515
rect 75275 463459 75331 463515
rect 73855 463317 73911 463373
rect 73997 463317 74053 463373
rect 74139 463317 74195 463373
rect 74281 463317 74337 463373
rect 74423 463317 74479 463373
rect 74565 463317 74621 463373
rect 74707 463317 74763 463373
rect 74849 463317 74905 463373
rect 74991 463317 75047 463373
rect 75133 463317 75189 463373
rect 75275 463317 75331 463373
rect 73855 463175 73911 463231
rect 73997 463175 74053 463231
rect 74139 463175 74195 463231
rect 74281 463175 74337 463231
rect 74423 463175 74479 463231
rect 74565 463175 74621 463231
rect 74707 463175 74763 463231
rect 74849 463175 74905 463231
rect 74991 463175 75047 463231
rect 75133 463175 75189 463231
rect 75275 463175 75331 463231
rect 73855 463033 73911 463089
rect 73997 463033 74053 463089
rect 74139 463033 74195 463089
rect 74281 463033 74337 463089
rect 74423 463033 74479 463089
rect 74565 463033 74621 463089
rect 74707 463033 74763 463089
rect 74849 463033 74905 463089
rect 74991 463033 75047 463089
rect 75133 463033 75189 463089
rect 75275 463033 75331 463089
rect 73855 462891 73911 462947
rect 73997 462891 74053 462947
rect 74139 462891 74195 462947
rect 74281 462891 74337 462947
rect 74423 462891 74479 462947
rect 74565 462891 74621 462947
rect 74707 462891 74763 462947
rect 74849 462891 74905 462947
rect 74991 462891 75047 462947
rect 75133 462891 75189 462947
rect 75275 462891 75331 462947
rect 73855 462749 73911 462805
rect 73997 462749 74053 462805
rect 74139 462749 74195 462805
rect 74281 462749 74337 462805
rect 74423 462749 74479 462805
rect 74565 462749 74621 462805
rect 74707 462749 74763 462805
rect 74849 462749 74905 462805
rect 74991 462749 75047 462805
rect 75133 462749 75189 462805
rect 75275 462749 75331 462805
rect 73855 462607 73911 462663
rect 73997 462607 74053 462663
rect 74139 462607 74195 462663
rect 74281 462607 74337 462663
rect 74423 462607 74479 462663
rect 74565 462607 74621 462663
rect 74707 462607 74763 462663
rect 74849 462607 74905 462663
rect 74991 462607 75047 462663
rect 75133 462607 75189 462663
rect 75275 462607 75331 462663
rect 73855 462465 73911 462521
rect 73997 462465 74053 462521
rect 74139 462465 74195 462521
rect 74281 462465 74337 462521
rect 74423 462465 74479 462521
rect 74565 462465 74621 462521
rect 74707 462465 74763 462521
rect 74849 462465 74905 462521
rect 74991 462465 75047 462521
rect 75133 462465 75189 462521
rect 75275 462465 75331 462521
rect 73855 462323 73911 462379
rect 73997 462323 74053 462379
rect 74139 462323 74195 462379
rect 74281 462323 74337 462379
rect 74423 462323 74479 462379
rect 74565 462323 74621 462379
rect 74707 462323 74763 462379
rect 74849 462323 74905 462379
rect 74991 462323 75047 462379
rect 75133 462323 75189 462379
rect 75275 462323 75331 462379
rect 73855 462181 73911 462237
rect 73997 462181 74053 462237
rect 74139 462181 74195 462237
rect 74281 462181 74337 462237
rect 74423 462181 74479 462237
rect 74565 462181 74621 462237
rect 74707 462181 74763 462237
rect 74849 462181 74905 462237
rect 74991 462181 75047 462237
rect 75133 462181 75189 462237
rect 75275 462181 75331 462237
rect 73855 462039 73911 462095
rect 73997 462039 74053 462095
rect 74139 462039 74195 462095
rect 74281 462039 74337 462095
rect 74423 462039 74479 462095
rect 74565 462039 74621 462095
rect 74707 462039 74763 462095
rect 74849 462039 74905 462095
rect 74991 462039 75047 462095
rect 75133 462039 75189 462095
rect 75275 462039 75331 462095
rect 73855 461897 73911 461953
rect 73997 461897 74053 461953
rect 74139 461897 74195 461953
rect 74281 461897 74337 461953
rect 74423 461897 74479 461953
rect 74565 461897 74621 461953
rect 74707 461897 74763 461953
rect 74849 461897 74905 461953
rect 74991 461897 75047 461953
rect 75133 461897 75189 461953
rect 75275 461897 75331 461953
rect 73855 461037 73911 461093
rect 73997 461037 74053 461093
rect 74139 461037 74195 461093
rect 74281 461037 74337 461093
rect 74423 461037 74479 461093
rect 74565 461037 74621 461093
rect 74707 461037 74763 461093
rect 74849 461037 74905 461093
rect 74991 461037 75047 461093
rect 75133 461037 75189 461093
rect 75275 461037 75331 461093
rect 73855 460895 73911 460951
rect 73997 460895 74053 460951
rect 74139 460895 74195 460951
rect 74281 460895 74337 460951
rect 74423 460895 74479 460951
rect 74565 460895 74621 460951
rect 74707 460895 74763 460951
rect 74849 460895 74905 460951
rect 74991 460895 75047 460951
rect 75133 460895 75189 460951
rect 75275 460895 75331 460951
rect 73855 460753 73911 460809
rect 73997 460753 74053 460809
rect 74139 460753 74195 460809
rect 74281 460753 74337 460809
rect 74423 460753 74479 460809
rect 74565 460753 74621 460809
rect 74707 460753 74763 460809
rect 74849 460753 74905 460809
rect 74991 460753 75047 460809
rect 75133 460753 75189 460809
rect 75275 460753 75331 460809
rect 73855 460611 73911 460667
rect 73997 460611 74053 460667
rect 74139 460611 74195 460667
rect 74281 460611 74337 460667
rect 74423 460611 74479 460667
rect 74565 460611 74621 460667
rect 74707 460611 74763 460667
rect 74849 460611 74905 460667
rect 74991 460611 75047 460667
rect 75133 460611 75189 460667
rect 75275 460611 75331 460667
rect 73855 460469 73911 460525
rect 73997 460469 74053 460525
rect 74139 460469 74195 460525
rect 74281 460469 74337 460525
rect 74423 460469 74479 460525
rect 74565 460469 74621 460525
rect 74707 460469 74763 460525
rect 74849 460469 74905 460525
rect 74991 460469 75047 460525
rect 75133 460469 75189 460525
rect 75275 460469 75331 460525
rect 73855 460327 73911 460383
rect 73997 460327 74053 460383
rect 74139 460327 74195 460383
rect 74281 460327 74337 460383
rect 74423 460327 74479 460383
rect 74565 460327 74621 460383
rect 74707 460327 74763 460383
rect 74849 460327 74905 460383
rect 74991 460327 75047 460383
rect 75133 460327 75189 460383
rect 75275 460327 75331 460383
rect 73855 460185 73911 460241
rect 73997 460185 74053 460241
rect 74139 460185 74195 460241
rect 74281 460185 74337 460241
rect 74423 460185 74479 460241
rect 74565 460185 74621 460241
rect 74707 460185 74763 460241
rect 74849 460185 74905 460241
rect 74991 460185 75047 460241
rect 75133 460185 75189 460241
rect 75275 460185 75331 460241
rect 73855 460043 73911 460099
rect 73997 460043 74053 460099
rect 74139 460043 74195 460099
rect 74281 460043 74337 460099
rect 74423 460043 74479 460099
rect 74565 460043 74621 460099
rect 74707 460043 74763 460099
rect 74849 460043 74905 460099
rect 74991 460043 75047 460099
rect 75133 460043 75189 460099
rect 75275 460043 75331 460099
rect 73855 459901 73911 459957
rect 73997 459901 74053 459957
rect 74139 459901 74195 459957
rect 74281 459901 74337 459957
rect 74423 459901 74479 459957
rect 74565 459901 74621 459957
rect 74707 459901 74763 459957
rect 74849 459901 74905 459957
rect 74991 459901 75047 459957
rect 75133 459901 75189 459957
rect 75275 459901 75331 459957
rect 73855 459759 73911 459815
rect 73997 459759 74053 459815
rect 74139 459759 74195 459815
rect 74281 459759 74337 459815
rect 74423 459759 74479 459815
rect 74565 459759 74621 459815
rect 74707 459759 74763 459815
rect 74849 459759 74905 459815
rect 74991 459759 75047 459815
rect 75133 459759 75189 459815
rect 75275 459759 75331 459815
rect 73855 459617 73911 459673
rect 73997 459617 74053 459673
rect 74139 459617 74195 459673
rect 74281 459617 74337 459673
rect 74423 459617 74479 459673
rect 74565 459617 74621 459673
rect 74707 459617 74763 459673
rect 74849 459617 74905 459673
rect 74991 459617 75047 459673
rect 75133 459617 75189 459673
rect 75275 459617 75331 459673
rect 73855 459475 73911 459531
rect 73997 459475 74053 459531
rect 74139 459475 74195 459531
rect 74281 459475 74337 459531
rect 74423 459475 74479 459531
rect 74565 459475 74621 459531
rect 74707 459475 74763 459531
rect 74849 459475 74905 459531
rect 74991 459475 75047 459531
rect 75133 459475 75189 459531
rect 75275 459475 75331 459531
rect 73855 459333 73911 459389
rect 73997 459333 74053 459389
rect 74139 459333 74195 459389
rect 74281 459333 74337 459389
rect 74423 459333 74479 459389
rect 74565 459333 74621 459389
rect 74707 459333 74763 459389
rect 74849 459333 74905 459389
rect 74991 459333 75047 459389
rect 75133 459333 75189 459389
rect 75275 459333 75331 459389
rect 73855 459191 73911 459247
rect 73997 459191 74053 459247
rect 74139 459191 74195 459247
rect 74281 459191 74337 459247
rect 74423 459191 74479 459247
rect 74565 459191 74621 459247
rect 74707 459191 74763 459247
rect 74849 459191 74905 459247
rect 74991 459191 75047 459247
rect 75133 459191 75189 459247
rect 75275 459191 75331 459247
rect 73855 458667 73911 458723
rect 73997 458667 74053 458723
rect 74139 458667 74195 458723
rect 74281 458667 74337 458723
rect 74423 458667 74479 458723
rect 74565 458667 74621 458723
rect 74707 458667 74763 458723
rect 74849 458667 74905 458723
rect 74991 458667 75047 458723
rect 75133 458667 75189 458723
rect 75275 458667 75331 458723
rect 73855 458525 73911 458581
rect 73997 458525 74053 458581
rect 74139 458525 74195 458581
rect 74281 458525 74337 458581
rect 74423 458525 74479 458581
rect 74565 458525 74621 458581
rect 74707 458525 74763 458581
rect 74849 458525 74905 458581
rect 74991 458525 75047 458581
rect 75133 458525 75189 458581
rect 75275 458525 75331 458581
rect 73855 458383 73911 458439
rect 73997 458383 74053 458439
rect 74139 458383 74195 458439
rect 74281 458383 74337 458439
rect 74423 458383 74479 458439
rect 74565 458383 74621 458439
rect 74707 458383 74763 458439
rect 74849 458383 74905 458439
rect 74991 458383 75047 458439
rect 75133 458383 75189 458439
rect 75275 458383 75331 458439
rect 73855 458241 73911 458297
rect 73997 458241 74053 458297
rect 74139 458241 74195 458297
rect 74281 458241 74337 458297
rect 74423 458241 74479 458297
rect 74565 458241 74621 458297
rect 74707 458241 74763 458297
rect 74849 458241 74905 458297
rect 74991 458241 75047 458297
rect 75133 458241 75189 458297
rect 75275 458241 75331 458297
rect 73855 458099 73911 458155
rect 73997 458099 74053 458155
rect 74139 458099 74195 458155
rect 74281 458099 74337 458155
rect 74423 458099 74479 458155
rect 74565 458099 74621 458155
rect 74707 458099 74763 458155
rect 74849 458099 74905 458155
rect 74991 458099 75047 458155
rect 75133 458099 75189 458155
rect 75275 458099 75331 458155
rect 73855 457957 73911 458013
rect 73997 457957 74053 458013
rect 74139 457957 74195 458013
rect 74281 457957 74337 458013
rect 74423 457957 74479 458013
rect 74565 457957 74621 458013
rect 74707 457957 74763 458013
rect 74849 457957 74905 458013
rect 74991 457957 75047 458013
rect 75133 457957 75189 458013
rect 75275 457957 75331 458013
rect 73855 457815 73911 457871
rect 73997 457815 74053 457871
rect 74139 457815 74195 457871
rect 74281 457815 74337 457871
rect 74423 457815 74479 457871
rect 74565 457815 74621 457871
rect 74707 457815 74763 457871
rect 74849 457815 74905 457871
rect 74991 457815 75047 457871
rect 75133 457815 75189 457871
rect 75275 457815 75331 457871
rect 73855 457673 73911 457729
rect 73997 457673 74053 457729
rect 74139 457673 74195 457729
rect 74281 457673 74337 457729
rect 74423 457673 74479 457729
rect 74565 457673 74621 457729
rect 74707 457673 74763 457729
rect 74849 457673 74905 457729
rect 74991 457673 75047 457729
rect 75133 457673 75189 457729
rect 75275 457673 75331 457729
rect 73855 457531 73911 457587
rect 73997 457531 74053 457587
rect 74139 457531 74195 457587
rect 74281 457531 74337 457587
rect 74423 457531 74479 457587
rect 74565 457531 74621 457587
rect 74707 457531 74763 457587
rect 74849 457531 74905 457587
rect 74991 457531 75047 457587
rect 75133 457531 75189 457587
rect 75275 457531 75331 457587
rect 73855 457389 73911 457445
rect 73997 457389 74053 457445
rect 74139 457389 74195 457445
rect 74281 457389 74337 457445
rect 74423 457389 74479 457445
rect 74565 457389 74621 457445
rect 74707 457389 74763 457445
rect 74849 457389 74905 457445
rect 74991 457389 75047 457445
rect 75133 457389 75189 457445
rect 75275 457389 75331 457445
rect 73855 457247 73911 457303
rect 73997 457247 74053 457303
rect 74139 457247 74195 457303
rect 74281 457247 74337 457303
rect 74423 457247 74479 457303
rect 74565 457247 74621 457303
rect 74707 457247 74763 457303
rect 74849 457247 74905 457303
rect 74991 457247 75047 457303
rect 75133 457247 75189 457303
rect 75275 457247 75331 457303
rect 73855 457105 73911 457161
rect 73997 457105 74053 457161
rect 74139 457105 74195 457161
rect 74281 457105 74337 457161
rect 74423 457105 74479 457161
rect 74565 457105 74621 457161
rect 74707 457105 74763 457161
rect 74849 457105 74905 457161
rect 74991 457105 75047 457161
rect 75133 457105 75189 457161
rect 75275 457105 75331 457161
rect 73855 456963 73911 457019
rect 73997 456963 74053 457019
rect 74139 456963 74195 457019
rect 74281 456963 74337 457019
rect 74423 456963 74479 457019
rect 74565 456963 74621 457019
rect 74707 456963 74763 457019
rect 74849 456963 74905 457019
rect 74991 456963 75047 457019
rect 75133 456963 75189 457019
rect 75275 456963 75331 457019
rect 73855 456821 73911 456877
rect 73997 456821 74053 456877
rect 74139 456821 74195 456877
rect 74281 456821 74337 456877
rect 74423 456821 74479 456877
rect 74565 456821 74621 456877
rect 74707 456821 74763 456877
rect 74849 456821 74905 456877
rect 74991 456821 75047 456877
rect 75133 456821 75189 456877
rect 75275 456821 75331 456877
rect 73866 456038 73922 456094
rect 74008 456038 74064 456094
rect 74150 456038 74206 456094
rect 74292 456038 74348 456094
rect 74434 456038 74490 456094
rect 74576 456038 74632 456094
rect 74718 456038 74774 456094
rect 74860 456038 74916 456094
rect 75002 456038 75058 456094
rect 75144 456038 75200 456094
rect 75286 456038 75342 456094
rect 73866 455896 73922 455952
rect 74008 455896 74064 455952
rect 74150 455896 74206 455952
rect 74292 455896 74348 455952
rect 74434 455896 74490 455952
rect 74576 455896 74632 455952
rect 74718 455896 74774 455952
rect 74860 455896 74916 455952
rect 75002 455896 75058 455952
rect 75144 455896 75200 455952
rect 75286 455896 75342 455952
rect 73866 455754 73922 455810
rect 74008 455754 74064 455810
rect 74150 455754 74206 455810
rect 74292 455754 74348 455810
rect 74434 455754 74490 455810
rect 74576 455754 74632 455810
rect 74718 455754 74774 455810
rect 74860 455754 74916 455810
rect 75002 455754 75058 455810
rect 75144 455754 75200 455810
rect 75286 455754 75342 455810
rect 73866 455612 73922 455668
rect 74008 455612 74064 455668
rect 74150 455612 74206 455668
rect 74292 455612 74348 455668
rect 74434 455612 74490 455668
rect 74576 455612 74632 455668
rect 74718 455612 74774 455668
rect 74860 455612 74916 455668
rect 75002 455612 75058 455668
rect 75144 455612 75200 455668
rect 75286 455612 75342 455668
rect 73866 455470 73922 455526
rect 74008 455470 74064 455526
rect 74150 455470 74206 455526
rect 74292 455470 74348 455526
rect 74434 455470 74490 455526
rect 74576 455470 74632 455526
rect 74718 455470 74774 455526
rect 74860 455470 74916 455526
rect 75002 455470 75058 455526
rect 75144 455470 75200 455526
rect 75286 455470 75342 455526
rect 73866 455328 73922 455384
rect 74008 455328 74064 455384
rect 74150 455328 74206 455384
rect 74292 455328 74348 455384
rect 74434 455328 74490 455384
rect 74576 455328 74632 455384
rect 74718 455328 74774 455384
rect 74860 455328 74916 455384
rect 75002 455328 75058 455384
rect 75144 455328 75200 455384
rect 75286 455328 75342 455384
rect 73866 455186 73922 455242
rect 74008 455186 74064 455242
rect 74150 455186 74206 455242
rect 74292 455186 74348 455242
rect 74434 455186 74490 455242
rect 74576 455186 74632 455242
rect 74718 455186 74774 455242
rect 74860 455186 74916 455242
rect 75002 455186 75058 455242
rect 75144 455186 75200 455242
rect 75286 455186 75342 455242
rect 73866 455044 73922 455100
rect 74008 455044 74064 455100
rect 74150 455044 74206 455100
rect 74292 455044 74348 455100
rect 74434 455044 74490 455100
rect 74576 455044 74632 455100
rect 74718 455044 74774 455100
rect 74860 455044 74916 455100
rect 75002 455044 75058 455100
rect 75144 455044 75200 455100
rect 75286 455044 75342 455100
rect 73866 454902 73922 454958
rect 74008 454902 74064 454958
rect 74150 454902 74206 454958
rect 74292 454902 74348 454958
rect 74434 454902 74490 454958
rect 74576 454902 74632 454958
rect 74718 454902 74774 454958
rect 74860 454902 74916 454958
rect 75002 454902 75058 454958
rect 75144 454902 75200 454958
rect 75286 454902 75342 454958
rect 73866 454760 73922 454816
rect 74008 454760 74064 454816
rect 74150 454760 74206 454816
rect 74292 454760 74348 454816
rect 74434 454760 74490 454816
rect 74576 454760 74632 454816
rect 74718 454760 74774 454816
rect 74860 454760 74916 454816
rect 75002 454760 75058 454816
rect 75144 454760 75200 454816
rect 75286 454760 75342 454816
rect 73866 454618 73922 454674
rect 74008 454618 74064 454674
rect 74150 454618 74206 454674
rect 74292 454618 74348 454674
rect 74434 454618 74490 454674
rect 74576 454618 74632 454674
rect 74718 454618 74774 454674
rect 74860 454618 74916 454674
rect 75002 454618 75058 454674
rect 75144 454618 75200 454674
rect 75286 454618 75342 454674
rect 73866 454476 73922 454532
rect 74008 454476 74064 454532
rect 74150 454476 74206 454532
rect 74292 454476 74348 454532
rect 74434 454476 74490 454532
rect 74576 454476 74632 454532
rect 74718 454476 74774 454532
rect 74860 454476 74916 454532
rect 75002 454476 75058 454532
rect 75144 454476 75200 454532
rect 75286 454476 75342 454532
rect 73866 454334 73922 454390
rect 74008 454334 74064 454390
rect 74150 454334 74206 454390
rect 74292 454334 74348 454390
rect 74434 454334 74490 454390
rect 74576 454334 74632 454390
rect 74718 454334 74774 454390
rect 74860 454334 74916 454390
rect 75002 454334 75058 454390
rect 75144 454334 75200 454390
rect 75286 454334 75342 454390
rect 702440 447610 702496 447666
rect 702582 447610 702638 447666
rect 702724 447610 702780 447666
rect 702866 447610 702922 447666
rect 703008 447610 703064 447666
rect 703150 447610 703206 447666
rect 703292 447610 703348 447666
rect 703434 447610 703490 447666
rect 703576 447610 703632 447666
rect 703718 447610 703774 447666
rect 703860 447610 703916 447666
rect 704002 447610 704058 447666
rect 704144 447610 704200 447666
rect 704286 447610 704342 447666
rect 702440 447468 702496 447524
rect 702582 447468 702638 447524
rect 702724 447468 702780 447524
rect 702866 447468 702922 447524
rect 703008 447468 703064 447524
rect 703150 447468 703206 447524
rect 703292 447468 703348 447524
rect 703434 447468 703490 447524
rect 703576 447468 703632 447524
rect 703718 447468 703774 447524
rect 703860 447468 703916 447524
rect 704002 447468 704058 447524
rect 704144 447468 704200 447524
rect 704286 447468 704342 447524
rect 702440 447326 702496 447382
rect 702582 447326 702638 447382
rect 702724 447326 702780 447382
rect 702866 447326 702922 447382
rect 703008 447326 703064 447382
rect 703150 447326 703206 447382
rect 703292 447326 703348 447382
rect 703434 447326 703490 447382
rect 703576 447326 703632 447382
rect 703718 447326 703774 447382
rect 703860 447326 703916 447382
rect 704002 447326 704058 447382
rect 704144 447326 704200 447382
rect 704286 447326 704342 447382
rect 702440 447184 702496 447240
rect 702582 447184 702638 447240
rect 702724 447184 702780 447240
rect 702866 447184 702922 447240
rect 703008 447184 703064 447240
rect 703150 447184 703206 447240
rect 703292 447184 703348 447240
rect 703434 447184 703490 447240
rect 703576 447184 703632 447240
rect 703718 447184 703774 447240
rect 703860 447184 703916 447240
rect 704002 447184 704058 447240
rect 704144 447184 704200 447240
rect 704286 447184 704342 447240
rect 702440 447042 702496 447098
rect 702582 447042 702638 447098
rect 702724 447042 702780 447098
rect 702866 447042 702922 447098
rect 703008 447042 703064 447098
rect 703150 447042 703206 447098
rect 703292 447042 703348 447098
rect 703434 447042 703490 447098
rect 703576 447042 703632 447098
rect 703718 447042 703774 447098
rect 703860 447042 703916 447098
rect 704002 447042 704058 447098
rect 704144 447042 704200 447098
rect 704286 447042 704342 447098
rect 702440 446900 702496 446956
rect 702582 446900 702638 446956
rect 702724 446900 702780 446956
rect 702866 446900 702922 446956
rect 703008 446900 703064 446956
rect 703150 446900 703206 446956
rect 703292 446900 703348 446956
rect 703434 446900 703490 446956
rect 703576 446900 703632 446956
rect 703718 446900 703774 446956
rect 703860 446900 703916 446956
rect 704002 446900 704058 446956
rect 704144 446900 704200 446956
rect 704286 446900 704342 446956
rect 702440 446758 702496 446814
rect 702582 446758 702638 446814
rect 702724 446758 702780 446814
rect 702866 446758 702922 446814
rect 703008 446758 703064 446814
rect 703150 446758 703206 446814
rect 703292 446758 703348 446814
rect 703434 446758 703490 446814
rect 703576 446758 703632 446814
rect 703718 446758 703774 446814
rect 703860 446758 703916 446814
rect 704002 446758 704058 446814
rect 704144 446758 704200 446814
rect 704286 446758 704342 446814
rect 702440 446616 702496 446672
rect 702582 446616 702638 446672
rect 702724 446616 702780 446672
rect 702866 446616 702922 446672
rect 703008 446616 703064 446672
rect 703150 446616 703206 446672
rect 703292 446616 703348 446672
rect 703434 446616 703490 446672
rect 703576 446616 703632 446672
rect 703718 446616 703774 446672
rect 703860 446616 703916 446672
rect 704002 446616 704058 446672
rect 704144 446616 704200 446672
rect 704286 446616 704342 446672
rect 702440 446474 702496 446530
rect 702582 446474 702638 446530
rect 702724 446474 702780 446530
rect 702866 446474 702922 446530
rect 703008 446474 703064 446530
rect 703150 446474 703206 446530
rect 703292 446474 703348 446530
rect 703434 446474 703490 446530
rect 703576 446474 703632 446530
rect 703718 446474 703774 446530
rect 703860 446474 703916 446530
rect 704002 446474 704058 446530
rect 704144 446474 704200 446530
rect 704286 446474 704342 446530
rect 702440 446332 702496 446388
rect 702582 446332 702638 446388
rect 702724 446332 702780 446388
rect 702866 446332 702922 446388
rect 703008 446332 703064 446388
rect 703150 446332 703206 446388
rect 703292 446332 703348 446388
rect 703434 446332 703490 446388
rect 703576 446332 703632 446388
rect 703718 446332 703774 446388
rect 703860 446332 703916 446388
rect 704002 446332 704058 446388
rect 704144 446332 704200 446388
rect 704286 446332 704342 446388
rect 702440 446190 702496 446246
rect 702582 446190 702638 446246
rect 702724 446190 702780 446246
rect 702866 446190 702922 446246
rect 703008 446190 703064 446246
rect 703150 446190 703206 446246
rect 703292 446190 703348 446246
rect 703434 446190 703490 446246
rect 703576 446190 703632 446246
rect 703718 446190 703774 446246
rect 703860 446190 703916 446246
rect 704002 446190 704058 446246
rect 704144 446190 704200 446246
rect 704286 446190 704342 446246
rect 702440 446048 702496 446104
rect 702582 446048 702638 446104
rect 702724 446048 702780 446104
rect 702866 446048 702922 446104
rect 703008 446048 703064 446104
rect 703150 446048 703206 446104
rect 703292 446048 703348 446104
rect 703434 446048 703490 446104
rect 703576 446048 703632 446104
rect 703718 446048 703774 446104
rect 703860 446048 703916 446104
rect 704002 446048 704058 446104
rect 704144 446048 704200 446104
rect 704286 446048 704342 446104
rect 702440 445906 702496 445962
rect 702582 445906 702638 445962
rect 702724 445906 702780 445962
rect 702866 445906 702922 445962
rect 703008 445906 703064 445962
rect 703150 445906 703206 445962
rect 703292 445906 703348 445962
rect 703434 445906 703490 445962
rect 703576 445906 703632 445962
rect 703718 445906 703774 445962
rect 703860 445906 703916 445962
rect 704002 445906 704058 445962
rect 704144 445906 704200 445962
rect 704286 445906 704342 445962
rect 702451 445123 702507 445179
rect 702593 445123 702649 445179
rect 702735 445123 702791 445179
rect 702877 445123 702933 445179
rect 703019 445123 703075 445179
rect 703161 445123 703217 445179
rect 703303 445123 703359 445179
rect 703445 445123 703501 445179
rect 703587 445123 703643 445179
rect 703729 445123 703785 445179
rect 703871 445123 703927 445179
rect 704013 445123 704069 445179
rect 704155 445123 704211 445179
rect 704297 445123 704353 445179
rect 702451 444981 702507 445037
rect 702593 444981 702649 445037
rect 702735 444981 702791 445037
rect 702877 444981 702933 445037
rect 703019 444981 703075 445037
rect 703161 444981 703217 445037
rect 703303 444981 703359 445037
rect 703445 444981 703501 445037
rect 703587 444981 703643 445037
rect 703729 444981 703785 445037
rect 703871 444981 703927 445037
rect 704013 444981 704069 445037
rect 704155 444981 704211 445037
rect 704297 444981 704353 445037
rect 702451 444839 702507 444895
rect 702593 444839 702649 444895
rect 702735 444839 702791 444895
rect 702877 444839 702933 444895
rect 703019 444839 703075 444895
rect 703161 444839 703217 444895
rect 703303 444839 703359 444895
rect 703445 444839 703501 444895
rect 703587 444839 703643 444895
rect 703729 444839 703785 444895
rect 703871 444839 703927 444895
rect 704013 444839 704069 444895
rect 704155 444839 704211 444895
rect 704297 444839 704353 444895
rect 702451 444697 702507 444753
rect 702593 444697 702649 444753
rect 702735 444697 702791 444753
rect 702877 444697 702933 444753
rect 703019 444697 703075 444753
rect 703161 444697 703217 444753
rect 703303 444697 703359 444753
rect 703445 444697 703501 444753
rect 703587 444697 703643 444753
rect 703729 444697 703785 444753
rect 703871 444697 703927 444753
rect 704013 444697 704069 444753
rect 704155 444697 704211 444753
rect 704297 444697 704353 444753
rect 702451 444555 702507 444611
rect 702593 444555 702649 444611
rect 702735 444555 702791 444611
rect 702877 444555 702933 444611
rect 703019 444555 703075 444611
rect 703161 444555 703217 444611
rect 703303 444555 703359 444611
rect 703445 444555 703501 444611
rect 703587 444555 703643 444611
rect 703729 444555 703785 444611
rect 703871 444555 703927 444611
rect 704013 444555 704069 444611
rect 704155 444555 704211 444611
rect 704297 444555 704353 444611
rect 702451 444413 702507 444469
rect 702593 444413 702649 444469
rect 702735 444413 702791 444469
rect 702877 444413 702933 444469
rect 703019 444413 703075 444469
rect 703161 444413 703217 444469
rect 703303 444413 703359 444469
rect 703445 444413 703501 444469
rect 703587 444413 703643 444469
rect 703729 444413 703785 444469
rect 703871 444413 703927 444469
rect 704013 444413 704069 444469
rect 704155 444413 704211 444469
rect 704297 444413 704353 444469
rect 702451 444271 702507 444327
rect 702593 444271 702649 444327
rect 702735 444271 702791 444327
rect 702877 444271 702933 444327
rect 703019 444271 703075 444327
rect 703161 444271 703217 444327
rect 703303 444271 703359 444327
rect 703445 444271 703501 444327
rect 703587 444271 703643 444327
rect 703729 444271 703785 444327
rect 703871 444271 703927 444327
rect 704013 444271 704069 444327
rect 704155 444271 704211 444327
rect 704297 444271 704353 444327
rect 702451 444129 702507 444185
rect 702593 444129 702649 444185
rect 702735 444129 702791 444185
rect 702877 444129 702933 444185
rect 703019 444129 703075 444185
rect 703161 444129 703217 444185
rect 703303 444129 703359 444185
rect 703445 444129 703501 444185
rect 703587 444129 703643 444185
rect 703729 444129 703785 444185
rect 703871 444129 703927 444185
rect 704013 444129 704069 444185
rect 704155 444129 704211 444185
rect 704297 444129 704353 444185
rect 702451 443987 702507 444043
rect 702593 443987 702649 444043
rect 702735 443987 702791 444043
rect 702877 443987 702933 444043
rect 703019 443987 703075 444043
rect 703161 443987 703217 444043
rect 703303 443987 703359 444043
rect 703445 443987 703501 444043
rect 703587 443987 703643 444043
rect 703729 443987 703785 444043
rect 703871 443987 703927 444043
rect 704013 443987 704069 444043
rect 704155 443987 704211 444043
rect 704297 443987 704353 444043
rect 702451 443845 702507 443901
rect 702593 443845 702649 443901
rect 702735 443845 702791 443901
rect 702877 443845 702933 443901
rect 703019 443845 703075 443901
rect 703161 443845 703217 443901
rect 703303 443845 703359 443901
rect 703445 443845 703501 443901
rect 703587 443845 703643 443901
rect 703729 443845 703785 443901
rect 703871 443845 703927 443901
rect 704013 443845 704069 443901
rect 704155 443845 704211 443901
rect 704297 443845 704353 443901
rect 702451 443703 702507 443759
rect 702593 443703 702649 443759
rect 702735 443703 702791 443759
rect 702877 443703 702933 443759
rect 703019 443703 703075 443759
rect 703161 443703 703217 443759
rect 703303 443703 703359 443759
rect 703445 443703 703501 443759
rect 703587 443703 703643 443759
rect 703729 443703 703785 443759
rect 703871 443703 703927 443759
rect 704013 443703 704069 443759
rect 704155 443703 704211 443759
rect 704297 443703 704353 443759
rect 702451 443561 702507 443617
rect 702593 443561 702649 443617
rect 702735 443561 702791 443617
rect 702877 443561 702933 443617
rect 703019 443561 703075 443617
rect 703161 443561 703217 443617
rect 703303 443561 703359 443617
rect 703445 443561 703501 443617
rect 703587 443561 703643 443617
rect 703729 443561 703785 443617
rect 703871 443561 703927 443617
rect 704013 443561 704069 443617
rect 704155 443561 704211 443617
rect 704297 443561 704353 443617
rect 702451 443419 702507 443475
rect 702593 443419 702649 443475
rect 702735 443419 702791 443475
rect 702877 443419 702933 443475
rect 703019 443419 703075 443475
rect 703161 443419 703217 443475
rect 703303 443419 703359 443475
rect 703445 443419 703501 443475
rect 703587 443419 703643 443475
rect 703729 443419 703785 443475
rect 703871 443419 703927 443475
rect 704013 443419 704069 443475
rect 704155 443419 704211 443475
rect 704297 443419 704353 443475
rect 702451 443277 702507 443333
rect 702593 443277 702649 443333
rect 702735 443277 702791 443333
rect 702877 443277 702933 443333
rect 703019 443277 703075 443333
rect 703161 443277 703217 443333
rect 703303 443277 703359 443333
rect 703445 443277 703501 443333
rect 703587 443277 703643 443333
rect 703729 443277 703785 443333
rect 703871 443277 703927 443333
rect 704013 443277 704069 443333
rect 704155 443277 704211 443333
rect 704297 443277 704353 443333
rect 702451 442753 702507 442809
rect 702593 442753 702649 442809
rect 702735 442753 702791 442809
rect 702877 442753 702933 442809
rect 703019 442753 703075 442809
rect 703161 442753 703217 442809
rect 703303 442753 703359 442809
rect 703445 442753 703501 442809
rect 703587 442753 703643 442809
rect 703729 442753 703785 442809
rect 703871 442753 703927 442809
rect 704013 442753 704069 442809
rect 704155 442753 704211 442809
rect 704297 442753 704353 442809
rect 702451 442611 702507 442667
rect 702593 442611 702649 442667
rect 702735 442611 702791 442667
rect 702877 442611 702933 442667
rect 703019 442611 703075 442667
rect 703161 442611 703217 442667
rect 703303 442611 703359 442667
rect 703445 442611 703501 442667
rect 703587 442611 703643 442667
rect 703729 442611 703785 442667
rect 703871 442611 703927 442667
rect 704013 442611 704069 442667
rect 704155 442611 704211 442667
rect 704297 442611 704353 442667
rect 702451 442469 702507 442525
rect 702593 442469 702649 442525
rect 702735 442469 702791 442525
rect 702877 442469 702933 442525
rect 703019 442469 703075 442525
rect 703161 442469 703217 442525
rect 703303 442469 703359 442525
rect 703445 442469 703501 442525
rect 703587 442469 703643 442525
rect 703729 442469 703785 442525
rect 703871 442469 703927 442525
rect 704013 442469 704069 442525
rect 704155 442469 704211 442525
rect 704297 442469 704353 442525
rect 702451 442327 702507 442383
rect 702593 442327 702649 442383
rect 702735 442327 702791 442383
rect 702877 442327 702933 442383
rect 703019 442327 703075 442383
rect 703161 442327 703217 442383
rect 703303 442327 703359 442383
rect 703445 442327 703501 442383
rect 703587 442327 703643 442383
rect 703729 442327 703785 442383
rect 703871 442327 703927 442383
rect 704013 442327 704069 442383
rect 704155 442327 704211 442383
rect 704297 442327 704353 442383
rect 702451 442185 702507 442241
rect 702593 442185 702649 442241
rect 702735 442185 702791 442241
rect 702877 442185 702933 442241
rect 703019 442185 703075 442241
rect 703161 442185 703217 442241
rect 703303 442185 703359 442241
rect 703445 442185 703501 442241
rect 703587 442185 703643 442241
rect 703729 442185 703785 442241
rect 703871 442185 703927 442241
rect 704013 442185 704069 442241
rect 704155 442185 704211 442241
rect 704297 442185 704353 442241
rect 702451 442043 702507 442099
rect 702593 442043 702649 442099
rect 702735 442043 702791 442099
rect 702877 442043 702933 442099
rect 703019 442043 703075 442099
rect 703161 442043 703217 442099
rect 703303 442043 703359 442099
rect 703445 442043 703501 442099
rect 703587 442043 703643 442099
rect 703729 442043 703785 442099
rect 703871 442043 703927 442099
rect 704013 442043 704069 442099
rect 704155 442043 704211 442099
rect 704297 442043 704353 442099
rect 702451 441901 702507 441957
rect 702593 441901 702649 441957
rect 702735 441901 702791 441957
rect 702877 441901 702933 441957
rect 703019 441901 703075 441957
rect 703161 441901 703217 441957
rect 703303 441901 703359 441957
rect 703445 441901 703501 441957
rect 703587 441901 703643 441957
rect 703729 441901 703785 441957
rect 703871 441901 703927 441957
rect 704013 441901 704069 441957
rect 704155 441901 704211 441957
rect 704297 441901 704353 441957
rect 702451 441759 702507 441815
rect 702593 441759 702649 441815
rect 702735 441759 702791 441815
rect 702877 441759 702933 441815
rect 703019 441759 703075 441815
rect 703161 441759 703217 441815
rect 703303 441759 703359 441815
rect 703445 441759 703501 441815
rect 703587 441759 703643 441815
rect 703729 441759 703785 441815
rect 703871 441759 703927 441815
rect 704013 441759 704069 441815
rect 704155 441759 704211 441815
rect 704297 441759 704353 441815
rect 702451 441617 702507 441673
rect 702593 441617 702649 441673
rect 702735 441617 702791 441673
rect 702877 441617 702933 441673
rect 703019 441617 703075 441673
rect 703161 441617 703217 441673
rect 703303 441617 703359 441673
rect 703445 441617 703501 441673
rect 703587 441617 703643 441673
rect 703729 441617 703785 441673
rect 703871 441617 703927 441673
rect 704013 441617 704069 441673
rect 704155 441617 704211 441673
rect 704297 441617 704353 441673
rect 702451 441475 702507 441531
rect 702593 441475 702649 441531
rect 702735 441475 702791 441531
rect 702877 441475 702933 441531
rect 703019 441475 703075 441531
rect 703161 441475 703217 441531
rect 703303 441475 703359 441531
rect 703445 441475 703501 441531
rect 703587 441475 703643 441531
rect 703729 441475 703785 441531
rect 703871 441475 703927 441531
rect 704013 441475 704069 441531
rect 704155 441475 704211 441531
rect 704297 441475 704353 441531
rect 702451 441333 702507 441389
rect 702593 441333 702649 441389
rect 702735 441333 702791 441389
rect 702877 441333 702933 441389
rect 703019 441333 703075 441389
rect 703161 441333 703217 441389
rect 703303 441333 703359 441389
rect 703445 441333 703501 441389
rect 703587 441333 703643 441389
rect 703729 441333 703785 441389
rect 703871 441333 703927 441389
rect 704013 441333 704069 441389
rect 704155 441333 704211 441389
rect 704297 441333 704353 441389
rect 702451 441191 702507 441247
rect 702593 441191 702649 441247
rect 702735 441191 702791 441247
rect 702877 441191 702933 441247
rect 703019 441191 703075 441247
rect 703161 441191 703217 441247
rect 703303 441191 703359 441247
rect 703445 441191 703501 441247
rect 703587 441191 703643 441247
rect 703729 441191 703785 441247
rect 703871 441191 703927 441247
rect 704013 441191 704069 441247
rect 704155 441191 704211 441247
rect 704297 441191 704353 441247
rect 702451 441049 702507 441105
rect 702593 441049 702649 441105
rect 702735 441049 702791 441105
rect 702877 441049 702933 441105
rect 703019 441049 703075 441105
rect 703161 441049 703217 441105
rect 703303 441049 703359 441105
rect 703445 441049 703501 441105
rect 703587 441049 703643 441105
rect 703729 441049 703785 441105
rect 703871 441049 703927 441105
rect 704013 441049 704069 441105
rect 704155 441049 704211 441105
rect 704297 441049 704353 441105
rect 702451 440907 702507 440963
rect 702593 440907 702649 440963
rect 702735 440907 702791 440963
rect 702877 440907 702933 440963
rect 703019 440907 703075 440963
rect 703161 440907 703217 440963
rect 703303 440907 703359 440963
rect 703445 440907 703501 440963
rect 703587 440907 703643 440963
rect 703729 440907 703785 440963
rect 703871 440907 703927 440963
rect 704013 440907 704069 440963
rect 704155 440907 704211 440963
rect 704297 440907 704353 440963
rect 702451 440047 702507 440103
rect 702593 440047 702649 440103
rect 702735 440047 702791 440103
rect 702877 440047 702933 440103
rect 703019 440047 703075 440103
rect 703161 440047 703217 440103
rect 703303 440047 703359 440103
rect 703445 440047 703501 440103
rect 703587 440047 703643 440103
rect 703729 440047 703785 440103
rect 703871 440047 703927 440103
rect 704013 440047 704069 440103
rect 704155 440047 704211 440103
rect 704297 440047 704353 440103
rect 702451 439905 702507 439961
rect 702593 439905 702649 439961
rect 702735 439905 702791 439961
rect 702877 439905 702933 439961
rect 703019 439905 703075 439961
rect 703161 439905 703217 439961
rect 703303 439905 703359 439961
rect 703445 439905 703501 439961
rect 703587 439905 703643 439961
rect 703729 439905 703785 439961
rect 703871 439905 703927 439961
rect 704013 439905 704069 439961
rect 704155 439905 704211 439961
rect 704297 439905 704353 439961
rect 702451 439763 702507 439819
rect 702593 439763 702649 439819
rect 702735 439763 702791 439819
rect 702877 439763 702933 439819
rect 703019 439763 703075 439819
rect 703161 439763 703217 439819
rect 703303 439763 703359 439819
rect 703445 439763 703501 439819
rect 703587 439763 703643 439819
rect 703729 439763 703785 439819
rect 703871 439763 703927 439819
rect 704013 439763 704069 439819
rect 704155 439763 704211 439819
rect 704297 439763 704353 439819
rect 702451 439621 702507 439677
rect 702593 439621 702649 439677
rect 702735 439621 702791 439677
rect 702877 439621 702933 439677
rect 703019 439621 703075 439677
rect 703161 439621 703217 439677
rect 703303 439621 703359 439677
rect 703445 439621 703501 439677
rect 703587 439621 703643 439677
rect 703729 439621 703785 439677
rect 703871 439621 703927 439677
rect 704013 439621 704069 439677
rect 704155 439621 704211 439677
rect 704297 439621 704353 439677
rect 702451 439479 702507 439535
rect 702593 439479 702649 439535
rect 702735 439479 702791 439535
rect 702877 439479 702933 439535
rect 703019 439479 703075 439535
rect 703161 439479 703217 439535
rect 703303 439479 703359 439535
rect 703445 439479 703501 439535
rect 703587 439479 703643 439535
rect 703729 439479 703785 439535
rect 703871 439479 703927 439535
rect 704013 439479 704069 439535
rect 704155 439479 704211 439535
rect 704297 439479 704353 439535
rect 702451 439337 702507 439393
rect 702593 439337 702649 439393
rect 702735 439337 702791 439393
rect 702877 439337 702933 439393
rect 703019 439337 703075 439393
rect 703161 439337 703217 439393
rect 703303 439337 703359 439393
rect 703445 439337 703501 439393
rect 703587 439337 703643 439393
rect 703729 439337 703785 439393
rect 703871 439337 703927 439393
rect 704013 439337 704069 439393
rect 704155 439337 704211 439393
rect 704297 439337 704353 439393
rect 702451 439195 702507 439251
rect 702593 439195 702649 439251
rect 702735 439195 702791 439251
rect 702877 439195 702933 439251
rect 703019 439195 703075 439251
rect 703161 439195 703217 439251
rect 703303 439195 703359 439251
rect 703445 439195 703501 439251
rect 703587 439195 703643 439251
rect 703729 439195 703785 439251
rect 703871 439195 703927 439251
rect 704013 439195 704069 439251
rect 704155 439195 704211 439251
rect 704297 439195 704353 439251
rect 702451 439053 702507 439109
rect 702593 439053 702649 439109
rect 702735 439053 702791 439109
rect 702877 439053 702933 439109
rect 703019 439053 703075 439109
rect 703161 439053 703217 439109
rect 703303 439053 703359 439109
rect 703445 439053 703501 439109
rect 703587 439053 703643 439109
rect 703729 439053 703785 439109
rect 703871 439053 703927 439109
rect 704013 439053 704069 439109
rect 704155 439053 704211 439109
rect 704297 439053 704353 439109
rect 702451 438911 702507 438967
rect 702593 438911 702649 438967
rect 702735 438911 702791 438967
rect 702877 438911 702933 438967
rect 703019 438911 703075 438967
rect 703161 438911 703217 438967
rect 703303 438911 703359 438967
rect 703445 438911 703501 438967
rect 703587 438911 703643 438967
rect 703729 438911 703785 438967
rect 703871 438911 703927 438967
rect 704013 438911 704069 438967
rect 704155 438911 704211 438967
rect 704297 438911 704353 438967
rect 702451 438769 702507 438825
rect 702593 438769 702649 438825
rect 702735 438769 702791 438825
rect 702877 438769 702933 438825
rect 703019 438769 703075 438825
rect 703161 438769 703217 438825
rect 703303 438769 703359 438825
rect 703445 438769 703501 438825
rect 703587 438769 703643 438825
rect 703729 438769 703785 438825
rect 703871 438769 703927 438825
rect 704013 438769 704069 438825
rect 704155 438769 704211 438825
rect 704297 438769 704353 438825
rect 702451 438627 702507 438683
rect 702593 438627 702649 438683
rect 702735 438627 702791 438683
rect 702877 438627 702933 438683
rect 703019 438627 703075 438683
rect 703161 438627 703217 438683
rect 703303 438627 703359 438683
rect 703445 438627 703501 438683
rect 703587 438627 703643 438683
rect 703729 438627 703785 438683
rect 703871 438627 703927 438683
rect 704013 438627 704069 438683
rect 704155 438627 704211 438683
rect 704297 438627 704353 438683
rect 702451 438485 702507 438541
rect 702593 438485 702649 438541
rect 702735 438485 702791 438541
rect 702877 438485 702933 438541
rect 703019 438485 703075 438541
rect 703161 438485 703217 438541
rect 703303 438485 703359 438541
rect 703445 438485 703501 438541
rect 703587 438485 703643 438541
rect 703729 438485 703785 438541
rect 703871 438485 703927 438541
rect 704013 438485 704069 438541
rect 704155 438485 704211 438541
rect 704297 438485 704353 438541
rect 702451 438343 702507 438399
rect 702593 438343 702649 438399
rect 702735 438343 702791 438399
rect 702877 438343 702933 438399
rect 703019 438343 703075 438399
rect 703161 438343 703217 438399
rect 703303 438343 703359 438399
rect 703445 438343 703501 438399
rect 703587 438343 703643 438399
rect 703729 438343 703785 438399
rect 703871 438343 703927 438399
rect 704013 438343 704069 438399
rect 704155 438343 704211 438399
rect 704297 438343 704353 438399
rect 702451 438201 702507 438257
rect 702593 438201 702649 438257
rect 702735 438201 702791 438257
rect 702877 438201 702933 438257
rect 703019 438201 703075 438257
rect 703161 438201 703217 438257
rect 703303 438201 703359 438257
rect 703445 438201 703501 438257
rect 703587 438201 703643 438257
rect 703729 438201 703785 438257
rect 703871 438201 703927 438257
rect 704013 438201 704069 438257
rect 704155 438201 704211 438257
rect 704297 438201 704353 438257
rect 702451 437677 702507 437733
rect 702593 437677 702649 437733
rect 702735 437677 702791 437733
rect 702877 437677 702933 437733
rect 703019 437677 703075 437733
rect 703161 437677 703217 437733
rect 703303 437677 703359 437733
rect 703445 437677 703501 437733
rect 703587 437677 703643 437733
rect 703729 437677 703785 437733
rect 703871 437677 703927 437733
rect 704013 437677 704069 437733
rect 704155 437677 704211 437733
rect 704297 437677 704353 437733
rect 702451 437535 702507 437591
rect 702593 437535 702649 437591
rect 702735 437535 702791 437591
rect 702877 437535 702933 437591
rect 703019 437535 703075 437591
rect 703161 437535 703217 437591
rect 703303 437535 703359 437591
rect 703445 437535 703501 437591
rect 703587 437535 703643 437591
rect 703729 437535 703785 437591
rect 703871 437535 703927 437591
rect 704013 437535 704069 437591
rect 704155 437535 704211 437591
rect 704297 437535 704353 437591
rect 702451 437393 702507 437449
rect 702593 437393 702649 437449
rect 702735 437393 702791 437449
rect 702877 437393 702933 437449
rect 703019 437393 703075 437449
rect 703161 437393 703217 437449
rect 703303 437393 703359 437449
rect 703445 437393 703501 437449
rect 703587 437393 703643 437449
rect 703729 437393 703785 437449
rect 703871 437393 703927 437449
rect 704013 437393 704069 437449
rect 704155 437393 704211 437449
rect 704297 437393 704353 437449
rect 702451 437251 702507 437307
rect 702593 437251 702649 437307
rect 702735 437251 702791 437307
rect 702877 437251 702933 437307
rect 703019 437251 703075 437307
rect 703161 437251 703217 437307
rect 703303 437251 703359 437307
rect 703445 437251 703501 437307
rect 703587 437251 703643 437307
rect 703729 437251 703785 437307
rect 703871 437251 703927 437307
rect 704013 437251 704069 437307
rect 704155 437251 704211 437307
rect 704297 437251 704353 437307
rect 702451 437109 702507 437165
rect 702593 437109 702649 437165
rect 702735 437109 702791 437165
rect 702877 437109 702933 437165
rect 703019 437109 703075 437165
rect 703161 437109 703217 437165
rect 703303 437109 703359 437165
rect 703445 437109 703501 437165
rect 703587 437109 703643 437165
rect 703729 437109 703785 437165
rect 703871 437109 703927 437165
rect 704013 437109 704069 437165
rect 704155 437109 704211 437165
rect 704297 437109 704353 437165
rect 702451 436967 702507 437023
rect 702593 436967 702649 437023
rect 702735 436967 702791 437023
rect 702877 436967 702933 437023
rect 703019 436967 703075 437023
rect 703161 436967 703217 437023
rect 703303 436967 703359 437023
rect 703445 436967 703501 437023
rect 703587 436967 703643 437023
rect 703729 436967 703785 437023
rect 703871 436967 703927 437023
rect 704013 436967 704069 437023
rect 704155 436967 704211 437023
rect 704297 436967 704353 437023
rect 702451 436825 702507 436881
rect 702593 436825 702649 436881
rect 702735 436825 702791 436881
rect 702877 436825 702933 436881
rect 703019 436825 703075 436881
rect 703161 436825 703217 436881
rect 703303 436825 703359 436881
rect 703445 436825 703501 436881
rect 703587 436825 703643 436881
rect 703729 436825 703785 436881
rect 703871 436825 703927 436881
rect 704013 436825 704069 436881
rect 704155 436825 704211 436881
rect 704297 436825 704353 436881
rect 702451 436683 702507 436739
rect 702593 436683 702649 436739
rect 702735 436683 702791 436739
rect 702877 436683 702933 436739
rect 703019 436683 703075 436739
rect 703161 436683 703217 436739
rect 703303 436683 703359 436739
rect 703445 436683 703501 436739
rect 703587 436683 703643 436739
rect 703729 436683 703785 436739
rect 703871 436683 703927 436739
rect 704013 436683 704069 436739
rect 704155 436683 704211 436739
rect 704297 436683 704353 436739
rect 702451 436541 702507 436597
rect 702593 436541 702649 436597
rect 702735 436541 702791 436597
rect 702877 436541 702933 436597
rect 703019 436541 703075 436597
rect 703161 436541 703217 436597
rect 703303 436541 703359 436597
rect 703445 436541 703501 436597
rect 703587 436541 703643 436597
rect 703729 436541 703785 436597
rect 703871 436541 703927 436597
rect 704013 436541 704069 436597
rect 704155 436541 704211 436597
rect 704297 436541 704353 436597
rect 702451 436399 702507 436455
rect 702593 436399 702649 436455
rect 702735 436399 702791 436455
rect 702877 436399 702933 436455
rect 703019 436399 703075 436455
rect 703161 436399 703217 436455
rect 703303 436399 703359 436455
rect 703445 436399 703501 436455
rect 703587 436399 703643 436455
rect 703729 436399 703785 436455
rect 703871 436399 703927 436455
rect 704013 436399 704069 436455
rect 704155 436399 704211 436455
rect 704297 436399 704353 436455
rect 702451 436257 702507 436313
rect 702593 436257 702649 436313
rect 702735 436257 702791 436313
rect 702877 436257 702933 436313
rect 703019 436257 703075 436313
rect 703161 436257 703217 436313
rect 703303 436257 703359 436313
rect 703445 436257 703501 436313
rect 703587 436257 703643 436313
rect 703729 436257 703785 436313
rect 703871 436257 703927 436313
rect 704013 436257 704069 436313
rect 704155 436257 704211 436313
rect 704297 436257 704353 436313
rect 702451 436115 702507 436171
rect 702593 436115 702649 436171
rect 702735 436115 702791 436171
rect 702877 436115 702933 436171
rect 703019 436115 703075 436171
rect 703161 436115 703217 436171
rect 703303 436115 703359 436171
rect 703445 436115 703501 436171
rect 703587 436115 703643 436171
rect 703729 436115 703785 436171
rect 703871 436115 703927 436171
rect 704013 436115 704069 436171
rect 704155 436115 704211 436171
rect 704297 436115 704353 436171
rect 702440 435054 702496 435110
rect 702582 435054 702638 435110
rect 702724 435054 702780 435110
rect 702866 435054 702922 435110
rect 703008 435054 703064 435110
rect 703150 435054 703206 435110
rect 703292 435054 703348 435110
rect 703434 435054 703490 435110
rect 703576 435054 703632 435110
rect 703718 435054 703774 435110
rect 703860 435054 703916 435110
rect 704002 435054 704058 435110
rect 704144 435054 704200 435110
rect 704286 435054 704342 435110
rect 702440 434912 702496 434968
rect 702582 434912 702638 434968
rect 702724 434912 702780 434968
rect 702866 434912 702922 434968
rect 703008 434912 703064 434968
rect 703150 434912 703206 434968
rect 703292 434912 703348 434968
rect 703434 434912 703490 434968
rect 703576 434912 703632 434968
rect 703718 434912 703774 434968
rect 703860 434912 703916 434968
rect 704002 434912 704058 434968
rect 704144 434912 704200 434968
rect 704286 434912 704342 434968
rect 702440 434770 702496 434826
rect 702582 434770 702638 434826
rect 702724 434770 702780 434826
rect 702866 434770 702922 434826
rect 703008 434770 703064 434826
rect 703150 434770 703206 434826
rect 703292 434770 703348 434826
rect 703434 434770 703490 434826
rect 703576 434770 703632 434826
rect 703718 434770 703774 434826
rect 703860 434770 703916 434826
rect 704002 434770 704058 434826
rect 704144 434770 704200 434826
rect 704286 434770 704342 434826
rect 702440 434628 702496 434684
rect 702582 434628 702638 434684
rect 702724 434628 702780 434684
rect 702866 434628 702922 434684
rect 703008 434628 703064 434684
rect 703150 434628 703206 434684
rect 703292 434628 703348 434684
rect 703434 434628 703490 434684
rect 703576 434628 703632 434684
rect 703718 434628 703774 434684
rect 703860 434628 703916 434684
rect 704002 434628 704058 434684
rect 704144 434628 704200 434684
rect 704286 434628 704342 434684
rect 702440 434486 702496 434542
rect 702582 434486 702638 434542
rect 702724 434486 702780 434542
rect 702866 434486 702922 434542
rect 703008 434486 703064 434542
rect 703150 434486 703206 434542
rect 703292 434486 703348 434542
rect 703434 434486 703490 434542
rect 703576 434486 703632 434542
rect 703718 434486 703774 434542
rect 703860 434486 703916 434542
rect 704002 434486 704058 434542
rect 704144 434486 704200 434542
rect 704286 434486 704342 434542
rect 702440 434344 702496 434400
rect 702582 434344 702638 434400
rect 702724 434344 702780 434400
rect 702866 434344 702922 434400
rect 703008 434344 703064 434400
rect 703150 434344 703206 434400
rect 703292 434344 703348 434400
rect 703434 434344 703490 434400
rect 703576 434344 703632 434400
rect 703718 434344 703774 434400
rect 703860 434344 703916 434400
rect 704002 434344 704058 434400
rect 704144 434344 704200 434400
rect 704286 434344 704342 434400
rect 702440 434202 702496 434258
rect 702582 434202 702638 434258
rect 702724 434202 702780 434258
rect 702866 434202 702922 434258
rect 703008 434202 703064 434258
rect 703150 434202 703206 434258
rect 703292 434202 703348 434258
rect 703434 434202 703490 434258
rect 703576 434202 703632 434258
rect 703718 434202 703774 434258
rect 703860 434202 703916 434258
rect 704002 434202 704058 434258
rect 704144 434202 704200 434258
rect 704286 434202 704342 434258
rect 702440 434060 702496 434116
rect 702582 434060 702638 434116
rect 702724 434060 702780 434116
rect 702866 434060 702922 434116
rect 703008 434060 703064 434116
rect 703150 434060 703206 434116
rect 703292 434060 703348 434116
rect 703434 434060 703490 434116
rect 703576 434060 703632 434116
rect 703718 434060 703774 434116
rect 703860 434060 703916 434116
rect 704002 434060 704058 434116
rect 704144 434060 704200 434116
rect 704286 434060 704342 434116
rect 702440 433918 702496 433974
rect 702582 433918 702638 433974
rect 702724 433918 702780 433974
rect 702866 433918 702922 433974
rect 703008 433918 703064 433974
rect 703150 433918 703206 433974
rect 703292 433918 703348 433974
rect 703434 433918 703490 433974
rect 703576 433918 703632 433974
rect 703718 433918 703774 433974
rect 703860 433918 703916 433974
rect 704002 433918 704058 433974
rect 704144 433918 704200 433974
rect 704286 433918 704342 433974
rect 702440 433776 702496 433832
rect 702582 433776 702638 433832
rect 702724 433776 702780 433832
rect 702866 433776 702922 433832
rect 703008 433776 703064 433832
rect 703150 433776 703206 433832
rect 703292 433776 703348 433832
rect 703434 433776 703490 433832
rect 703576 433776 703632 433832
rect 703718 433776 703774 433832
rect 703860 433776 703916 433832
rect 704002 433776 704058 433832
rect 704144 433776 704200 433832
rect 704286 433776 704342 433832
rect 702440 433634 702496 433690
rect 702582 433634 702638 433690
rect 702724 433634 702780 433690
rect 702866 433634 702922 433690
rect 703008 433634 703064 433690
rect 703150 433634 703206 433690
rect 703292 433634 703348 433690
rect 703434 433634 703490 433690
rect 703576 433634 703632 433690
rect 703718 433634 703774 433690
rect 703860 433634 703916 433690
rect 704002 433634 704058 433690
rect 704144 433634 704200 433690
rect 704286 433634 704342 433690
rect 702440 433492 702496 433548
rect 702582 433492 702638 433548
rect 702724 433492 702780 433548
rect 702866 433492 702922 433548
rect 703008 433492 703064 433548
rect 703150 433492 703206 433548
rect 703292 433492 703348 433548
rect 703434 433492 703490 433548
rect 703576 433492 703632 433548
rect 703718 433492 703774 433548
rect 703860 433492 703916 433548
rect 704002 433492 704058 433548
rect 704144 433492 704200 433548
rect 704286 433492 704342 433548
rect 702440 433350 702496 433406
rect 702582 433350 702638 433406
rect 702724 433350 702780 433406
rect 702866 433350 702922 433406
rect 703008 433350 703064 433406
rect 703150 433350 703206 433406
rect 703292 433350 703348 433406
rect 703434 433350 703490 433406
rect 703576 433350 703632 433406
rect 703718 433350 703774 433406
rect 703860 433350 703916 433406
rect 704002 433350 704058 433406
rect 704144 433350 704200 433406
rect 704286 433350 704342 433406
rect 71466 427594 71522 427650
rect 71608 427594 71664 427650
rect 71750 427594 71806 427650
rect 71892 427594 71948 427650
rect 72034 427594 72090 427650
rect 72176 427594 72232 427650
rect 72318 427594 72374 427650
rect 72460 427594 72516 427650
rect 72602 427594 72658 427650
rect 72744 427594 72800 427650
rect 72886 427594 72942 427650
rect 73028 427594 73084 427650
rect 73170 427594 73226 427650
rect 73312 427594 73368 427650
rect 71466 427452 71522 427508
rect 71608 427452 71664 427508
rect 71750 427452 71806 427508
rect 71892 427452 71948 427508
rect 72034 427452 72090 427508
rect 72176 427452 72232 427508
rect 72318 427452 72374 427508
rect 72460 427452 72516 427508
rect 72602 427452 72658 427508
rect 72744 427452 72800 427508
rect 72886 427452 72942 427508
rect 73028 427452 73084 427508
rect 73170 427452 73226 427508
rect 73312 427452 73368 427508
rect 71466 427310 71522 427366
rect 71608 427310 71664 427366
rect 71750 427310 71806 427366
rect 71892 427310 71948 427366
rect 72034 427310 72090 427366
rect 72176 427310 72232 427366
rect 72318 427310 72374 427366
rect 72460 427310 72516 427366
rect 72602 427310 72658 427366
rect 72744 427310 72800 427366
rect 72886 427310 72942 427366
rect 73028 427310 73084 427366
rect 73170 427310 73226 427366
rect 73312 427310 73368 427366
rect 71466 427168 71522 427224
rect 71608 427168 71664 427224
rect 71750 427168 71806 427224
rect 71892 427168 71948 427224
rect 72034 427168 72090 427224
rect 72176 427168 72232 427224
rect 72318 427168 72374 427224
rect 72460 427168 72516 427224
rect 72602 427168 72658 427224
rect 72744 427168 72800 427224
rect 72886 427168 72942 427224
rect 73028 427168 73084 427224
rect 73170 427168 73226 427224
rect 73312 427168 73368 427224
rect 71466 427026 71522 427082
rect 71608 427026 71664 427082
rect 71750 427026 71806 427082
rect 71892 427026 71948 427082
rect 72034 427026 72090 427082
rect 72176 427026 72232 427082
rect 72318 427026 72374 427082
rect 72460 427026 72516 427082
rect 72602 427026 72658 427082
rect 72744 427026 72800 427082
rect 72886 427026 72942 427082
rect 73028 427026 73084 427082
rect 73170 427026 73226 427082
rect 73312 427026 73368 427082
rect 71466 426884 71522 426940
rect 71608 426884 71664 426940
rect 71750 426884 71806 426940
rect 71892 426884 71948 426940
rect 72034 426884 72090 426940
rect 72176 426884 72232 426940
rect 72318 426884 72374 426940
rect 72460 426884 72516 426940
rect 72602 426884 72658 426940
rect 72744 426884 72800 426940
rect 72886 426884 72942 426940
rect 73028 426884 73084 426940
rect 73170 426884 73226 426940
rect 73312 426884 73368 426940
rect 71466 426742 71522 426798
rect 71608 426742 71664 426798
rect 71750 426742 71806 426798
rect 71892 426742 71948 426798
rect 72034 426742 72090 426798
rect 72176 426742 72232 426798
rect 72318 426742 72374 426798
rect 72460 426742 72516 426798
rect 72602 426742 72658 426798
rect 72744 426742 72800 426798
rect 72886 426742 72942 426798
rect 73028 426742 73084 426798
rect 73170 426742 73226 426798
rect 73312 426742 73368 426798
rect 71466 426600 71522 426656
rect 71608 426600 71664 426656
rect 71750 426600 71806 426656
rect 71892 426600 71948 426656
rect 72034 426600 72090 426656
rect 72176 426600 72232 426656
rect 72318 426600 72374 426656
rect 72460 426600 72516 426656
rect 72602 426600 72658 426656
rect 72744 426600 72800 426656
rect 72886 426600 72942 426656
rect 73028 426600 73084 426656
rect 73170 426600 73226 426656
rect 73312 426600 73368 426656
rect 71466 426458 71522 426514
rect 71608 426458 71664 426514
rect 71750 426458 71806 426514
rect 71892 426458 71948 426514
rect 72034 426458 72090 426514
rect 72176 426458 72232 426514
rect 72318 426458 72374 426514
rect 72460 426458 72516 426514
rect 72602 426458 72658 426514
rect 72744 426458 72800 426514
rect 72886 426458 72942 426514
rect 73028 426458 73084 426514
rect 73170 426458 73226 426514
rect 73312 426458 73368 426514
rect 71466 426316 71522 426372
rect 71608 426316 71664 426372
rect 71750 426316 71806 426372
rect 71892 426316 71948 426372
rect 72034 426316 72090 426372
rect 72176 426316 72232 426372
rect 72318 426316 72374 426372
rect 72460 426316 72516 426372
rect 72602 426316 72658 426372
rect 72744 426316 72800 426372
rect 72886 426316 72942 426372
rect 73028 426316 73084 426372
rect 73170 426316 73226 426372
rect 73312 426316 73368 426372
rect 71466 426174 71522 426230
rect 71608 426174 71664 426230
rect 71750 426174 71806 426230
rect 71892 426174 71948 426230
rect 72034 426174 72090 426230
rect 72176 426174 72232 426230
rect 72318 426174 72374 426230
rect 72460 426174 72516 426230
rect 72602 426174 72658 426230
rect 72744 426174 72800 426230
rect 72886 426174 72942 426230
rect 73028 426174 73084 426230
rect 73170 426174 73226 426230
rect 73312 426174 73368 426230
rect 71466 426032 71522 426088
rect 71608 426032 71664 426088
rect 71750 426032 71806 426088
rect 71892 426032 71948 426088
rect 72034 426032 72090 426088
rect 72176 426032 72232 426088
rect 72318 426032 72374 426088
rect 72460 426032 72516 426088
rect 72602 426032 72658 426088
rect 72744 426032 72800 426088
rect 72886 426032 72942 426088
rect 73028 426032 73084 426088
rect 73170 426032 73226 426088
rect 73312 426032 73368 426088
rect 71466 425890 71522 425946
rect 71608 425890 71664 425946
rect 71750 425890 71806 425946
rect 71892 425890 71948 425946
rect 72034 425890 72090 425946
rect 72176 425890 72232 425946
rect 72318 425890 72374 425946
rect 72460 425890 72516 425946
rect 72602 425890 72658 425946
rect 72744 425890 72800 425946
rect 72886 425890 72942 425946
rect 73028 425890 73084 425946
rect 73170 425890 73226 425946
rect 73312 425890 73368 425946
rect 71455 425113 71511 425169
rect 71597 425113 71653 425169
rect 71739 425113 71795 425169
rect 71881 425113 71937 425169
rect 72023 425113 72079 425169
rect 72165 425113 72221 425169
rect 72307 425113 72363 425169
rect 72449 425113 72505 425169
rect 72591 425113 72647 425169
rect 72733 425113 72789 425169
rect 72875 425113 72931 425169
rect 73017 425113 73073 425169
rect 73159 425113 73215 425169
rect 73301 425113 73357 425169
rect 71455 424971 71511 425027
rect 71597 424971 71653 425027
rect 71739 424971 71795 425027
rect 71881 424971 71937 425027
rect 72023 424971 72079 425027
rect 72165 424971 72221 425027
rect 72307 424971 72363 425027
rect 72449 424971 72505 425027
rect 72591 424971 72647 425027
rect 72733 424971 72789 425027
rect 72875 424971 72931 425027
rect 73017 424971 73073 425027
rect 73159 424971 73215 425027
rect 73301 424971 73357 425027
rect 71455 424829 71511 424885
rect 71597 424829 71653 424885
rect 71739 424829 71795 424885
rect 71881 424829 71937 424885
rect 72023 424829 72079 424885
rect 72165 424829 72221 424885
rect 72307 424829 72363 424885
rect 72449 424829 72505 424885
rect 72591 424829 72647 424885
rect 72733 424829 72789 424885
rect 72875 424829 72931 424885
rect 73017 424829 73073 424885
rect 73159 424829 73215 424885
rect 73301 424829 73357 424885
rect 71455 424687 71511 424743
rect 71597 424687 71653 424743
rect 71739 424687 71795 424743
rect 71881 424687 71937 424743
rect 72023 424687 72079 424743
rect 72165 424687 72221 424743
rect 72307 424687 72363 424743
rect 72449 424687 72505 424743
rect 72591 424687 72647 424743
rect 72733 424687 72789 424743
rect 72875 424687 72931 424743
rect 73017 424687 73073 424743
rect 73159 424687 73215 424743
rect 73301 424687 73357 424743
rect 71455 424545 71511 424601
rect 71597 424545 71653 424601
rect 71739 424545 71795 424601
rect 71881 424545 71937 424601
rect 72023 424545 72079 424601
rect 72165 424545 72221 424601
rect 72307 424545 72363 424601
rect 72449 424545 72505 424601
rect 72591 424545 72647 424601
rect 72733 424545 72789 424601
rect 72875 424545 72931 424601
rect 73017 424545 73073 424601
rect 73159 424545 73215 424601
rect 73301 424545 73357 424601
rect 71455 424403 71511 424459
rect 71597 424403 71653 424459
rect 71739 424403 71795 424459
rect 71881 424403 71937 424459
rect 72023 424403 72079 424459
rect 72165 424403 72221 424459
rect 72307 424403 72363 424459
rect 72449 424403 72505 424459
rect 72591 424403 72647 424459
rect 72733 424403 72789 424459
rect 72875 424403 72931 424459
rect 73017 424403 73073 424459
rect 73159 424403 73215 424459
rect 73301 424403 73357 424459
rect 71455 424261 71511 424317
rect 71597 424261 71653 424317
rect 71739 424261 71795 424317
rect 71881 424261 71937 424317
rect 72023 424261 72079 424317
rect 72165 424261 72221 424317
rect 72307 424261 72363 424317
rect 72449 424261 72505 424317
rect 72591 424261 72647 424317
rect 72733 424261 72789 424317
rect 72875 424261 72931 424317
rect 73017 424261 73073 424317
rect 73159 424261 73215 424317
rect 73301 424261 73357 424317
rect 71455 424119 71511 424175
rect 71597 424119 71653 424175
rect 71739 424119 71795 424175
rect 71881 424119 71937 424175
rect 72023 424119 72079 424175
rect 72165 424119 72221 424175
rect 72307 424119 72363 424175
rect 72449 424119 72505 424175
rect 72591 424119 72647 424175
rect 72733 424119 72789 424175
rect 72875 424119 72931 424175
rect 73017 424119 73073 424175
rect 73159 424119 73215 424175
rect 73301 424119 73357 424175
rect 71455 423977 71511 424033
rect 71597 423977 71653 424033
rect 71739 423977 71795 424033
rect 71881 423977 71937 424033
rect 72023 423977 72079 424033
rect 72165 423977 72221 424033
rect 72307 423977 72363 424033
rect 72449 423977 72505 424033
rect 72591 423977 72647 424033
rect 72733 423977 72789 424033
rect 72875 423977 72931 424033
rect 73017 423977 73073 424033
rect 73159 423977 73215 424033
rect 73301 423977 73357 424033
rect 71455 423835 71511 423891
rect 71597 423835 71653 423891
rect 71739 423835 71795 423891
rect 71881 423835 71937 423891
rect 72023 423835 72079 423891
rect 72165 423835 72221 423891
rect 72307 423835 72363 423891
rect 72449 423835 72505 423891
rect 72591 423835 72647 423891
rect 72733 423835 72789 423891
rect 72875 423835 72931 423891
rect 73017 423835 73073 423891
rect 73159 423835 73215 423891
rect 73301 423835 73357 423891
rect 71455 423693 71511 423749
rect 71597 423693 71653 423749
rect 71739 423693 71795 423749
rect 71881 423693 71937 423749
rect 72023 423693 72079 423749
rect 72165 423693 72221 423749
rect 72307 423693 72363 423749
rect 72449 423693 72505 423749
rect 72591 423693 72647 423749
rect 72733 423693 72789 423749
rect 72875 423693 72931 423749
rect 73017 423693 73073 423749
rect 73159 423693 73215 423749
rect 73301 423693 73357 423749
rect 71455 423551 71511 423607
rect 71597 423551 71653 423607
rect 71739 423551 71795 423607
rect 71881 423551 71937 423607
rect 72023 423551 72079 423607
rect 72165 423551 72221 423607
rect 72307 423551 72363 423607
rect 72449 423551 72505 423607
rect 72591 423551 72647 423607
rect 72733 423551 72789 423607
rect 72875 423551 72931 423607
rect 73017 423551 73073 423607
rect 73159 423551 73215 423607
rect 73301 423551 73357 423607
rect 71455 423409 71511 423465
rect 71597 423409 71653 423465
rect 71739 423409 71795 423465
rect 71881 423409 71937 423465
rect 72023 423409 72079 423465
rect 72165 423409 72221 423465
rect 72307 423409 72363 423465
rect 72449 423409 72505 423465
rect 72591 423409 72647 423465
rect 72733 423409 72789 423465
rect 72875 423409 72931 423465
rect 73017 423409 73073 423465
rect 73159 423409 73215 423465
rect 73301 423409 73357 423465
rect 71455 423267 71511 423323
rect 71597 423267 71653 423323
rect 71739 423267 71795 423323
rect 71881 423267 71937 423323
rect 72023 423267 72079 423323
rect 72165 423267 72221 423323
rect 72307 423267 72363 423323
rect 72449 423267 72505 423323
rect 72591 423267 72647 423323
rect 72733 423267 72789 423323
rect 72875 423267 72931 423323
rect 73017 423267 73073 423323
rect 73159 423267 73215 423323
rect 73301 423267 73357 423323
rect 71455 422743 71511 422799
rect 71597 422743 71653 422799
rect 71739 422743 71795 422799
rect 71881 422743 71937 422799
rect 72023 422743 72079 422799
rect 72165 422743 72221 422799
rect 72307 422743 72363 422799
rect 72449 422743 72505 422799
rect 72591 422743 72647 422799
rect 72733 422743 72789 422799
rect 72875 422743 72931 422799
rect 73017 422743 73073 422799
rect 73159 422743 73215 422799
rect 73301 422743 73357 422799
rect 71455 422601 71511 422657
rect 71597 422601 71653 422657
rect 71739 422601 71795 422657
rect 71881 422601 71937 422657
rect 72023 422601 72079 422657
rect 72165 422601 72221 422657
rect 72307 422601 72363 422657
rect 72449 422601 72505 422657
rect 72591 422601 72647 422657
rect 72733 422601 72789 422657
rect 72875 422601 72931 422657
rect 73017 422601 73073 422657
rect 73159 422601 73215 422657
rect 73301 422601 73357 422657
rect 71455 422459 71511 422515
rect 71597 422459 71653 422515
rect 71739 422459 71795 422515
rect 71881 422459 71937 422515
rect 72023 422459 72079 422515
rect 72165 422459 72221 422515
rect 72307 422459 72363 422515
rect 72449 422459 72505 422515
rect 72591 422459 72647 422515
rect 72733 422459 72789 422515
rect 72875 422459 72931 422515
rect 73017 422459 73073 422515
rect 73159 422459 73215 422515
rect 73301 422459 73357 422515
rect 71455 422317 71511 422373
rect 71597 422317 71653 422373
rect 71739 422317 71795 422373
rect 71881 422317 71937 422373
rect 72023 422317 72079 422373
rect 72165 422317 72221 422373
rect 72307 422317 72363 422373
rect 72449 422317 72505 422373
rect 72591 422317 72647 422373
rect 72733 422317 72789 422373
rect 72875 422317 72931 422373
rect 73017 422317 73073 422373
rect 73159 422317 73215 422373
rect 73301 422317 73357 422373
rect 71455 422175 71511 422231
rect 71597 422175 71653 422231
rect 71739 422175 71795 422231
rect 71881 422175 71937 422231
rect 72023 422175 72079 422231
rect 72165 422175 72221 422231
rect 72307 422175 72363 422231
rect 72449 422175 72505 422231
rect 72591 422175 72647 422231
rect 72733 422175 72789 422231
rect 72875 422175 72931 422231
rect 73017 422175 73073 422231
rect 73159 422175 73215 422231
rect 73301 422175 73357 422231
rect 71455 422033 71511 422089
rect 71597 422033 71653 422089
rect 71739 422033 71795 422089
rect 71881 422033 71937 422089
rect 72023 422033 72079 422089
rect 72165 422033 72221 422089
rect 72307 422033 72363 422089
rect 72449 422033 72505 422089
rect 72591 422033 72647 422089
rect 72733 422033 72789 422089
rect 72875 422033 72931 422089
rect 73017 422033 73073 422089
rect 73159 422033 73215 422089
rect 73301 422033 73357 422089
rect 71455 421891 71511 421947
rect 71597 421891 71653 421947
rect 71739 421891 71795 421947
rect 71881 421891 71937 421947
rect 72023 421891 72079 421947
rect 72165 421891 72221 421947
rect 72307 421891 72363 421947
rect 72449 421891 72505 421947
rect 72591 421891 72647 421947
rect 72733 421891 72789 421947
rect 72875 421891 72931 421947
rect 73017 421891 73073 421947
rect 73159 421891 73215 421947
rect 73301 421891 73357 421947
rect 71455 421749 71511 421805
rect 71597 421749 71653 421805
rect 71739 421749 71795 421805
rect 71881 421749 71937 421805
rect 72023 421749 72079 421805
rect 72165 421749 72221 421805
rect 72307 421749 72363 421805
rect 72449 421749 72505 421805
rect 72591 421749 72647 421805
rect 72733 421749 72789 421805
rect 72875 421749 72931 421805
rect 73017 421749 73073 421805
rect 73159 421749 73215 421805
rect 73301 421749 73357 421805
rect 71455 421607 71511 421663
rect 71597 421607 71653 421663
rect 71739 421607 71795 421663
rect 71881 421607 71937 421663
rect 72023 421607 72079 421663
rect 72165 421607 72221 421663
rect 72307 421607 72363 421663
rect 72449 421607 72505 421663
rect 72591 421607 72647 421663
rect 72733 421607 72789 421663
rect 72875 421607 72931 421663
rect 73017 421607 73073 421663
rect 73159 421607 73215 421663
rect 73301 421607 73357 421663
rect 71455 421465 71511 421521
rect 71597 421465 71653 421521
rect 71739 421465 71795 421521
rect 71881 421465 71937 421521
rect 72023 421465 72079 421521
rect 72165 421465 72221 421521
rect 72307 421465 72363 421521
rect 72449 421465 72505 421521
rect 72591 421465 72647 421521
rect 72733 421465 72789 421521
rect 72875 421465 72931 421521
rect 73017 421465 73073 421521
rect 73159 421465 73215 421521
rect 73301 421465 73357 421521
rect 71455 421323 71511 421379
rect 71597 421323 71653 421379
rect 71739 421323 71795 421379
rect 71881 421323 71937 421379
rect 72023 421323 72079 421379
rect 72165 421323 72221 421379
rect 72307 421323 72363 421379
rect 72449 421323 72505 421379
rect 72591 421323 72647 421379
rect 72733 421323 72789 421379
rect 72875 421323 72931 421379
rect 73017 421323 73073 421379
rect 73159 421323 73215 421379
rect 73301 421323 73357 421379
rect 71455 421181 71511 421237
rect 71597 421181 71653 421237
rect 71739 421181 71795 421237
rect 71881 421181 71937 421237
rect 72023 421181 72079 421237
rect 72165 421181 72221 421237
rect 72307 421181 72363 421237
rect 72449 421181 72505 421237
rect 72591 421181 72647 421237
rect 72733 421181 72789 421237
rect 72875 421181 72931 421237
rect 73017 421181 73073 421237
rect 73159 421181 73215 421237
rect 73301 421181 73357 421237
rect 71455 421039 71511 421095
rect 71597 421039 71653 421095
rect 71739 421039 71795 421095
rect 71881 421039 71937 421095
rect 72023 421039 72079 421095
rect 72165 421039 72221 421095
rect 72307 421039 72363 421095
rect 72449 421039 72505 421095
rect 72591 421039 72647 421095
rect 72733 421039 72789 421095
rect 72875 421039 72931 421095
rect 73017 421039 73073 421095
rect 73159 421039 73215 421095
rect 73301 421039 73357 421095
rect 71455 420897 71511 420953
rect 71597 420897 71653 420953
rect 71739 420897 71795 420953
rect 71881 420897 71937 420953
rect 72023 420897 72079 420953
rect 72165 420897 72221 420953
rect 72307 420897 72363 420953
rect 72449 420897 72505 420953
rect 72591 420897 72647 420953
rect 72733 420897 72789 420953
rect 72875 420897 72931 420953
rect 73017 420897 73073 420953
rect 73159 420897 73215 420953
rect 73301 420897 73357 420953
rect 71455 420037 71511 420093
rect 71597 420037 71653 420093
rect 71739 420037 71795 420093
rect 71881 420037 71937 420093
rect 72023 420037 72079 420093
rect 72165 420037 72221 420093
rect 72307 420037 72363 420093
rect 72449 420037 72505 420093
rect 72591 420037 72647 420093
rect 72733 420037 72789 420093
rect 72875 420037 72931 420093
rect 73017 420037 73073 420093
rect 73159 420037 73215 420093
rect 73301 420037 73357 420093
rect 71455 419895 71511 419951
rect 71597 419895 71653 419951
rect 71739 419895 71795 419951
rect 71881 419895 71937 419951
rect 72023 419895 72079 419951
rect 72165 419895 72221 419951
rect 72307 419895 72363 419951
rect 72449 419895 72505 419951
rect 72591 419895 72647 419951
rect 72733 419895 72789 419951
rect 72875 419895 72931 419951
rect 73017 419895 73073 419951
rect 73159 419895 73215 419951
rect 73301 419895 73357 419951
rect 71455 419753 71511 419809
rect 71597 419753 71653 419809
rect 71739 419753 71795 419809
rect 71881 419753 71937 419809
rect 72023 419753 72079 419809
rect 72165 419753 72221 419809
rect 72307 419753 72363 419809
rect 72449 419753 72505 419809
rect 72591 419753 72647 419809
rect 72733 419753 72789 419809
rect 72875 419753 72931 419809
rect 73017 419753 73073 419809
rect 73159 419753 73215 419809
rect 73301 419753 73357 419809
rect 71455 419611 71511 419667
rect 71597 419611 71653 419667
rect 71739 419611 71795 419667
rect 71881 419611 71937 419667
rect 72023 419611 72079 419667
rect 72165 419611 72221 419667
rect 72307 419611 72363 419667
rect 72449 419611 72505 419667
rect 72591 419611 72647 419667
rect 72733 419611 72789 419667
rect 72875 419611 72931 419667
rect 73017 419611 73073 419667
rect 73159 419611 73215 419667
rect 73301 419611 73357 419667
rect 71455 419469 71511 419525
rect 71597 419469 71653 419525
rect 71739 419469 71795 419525
rect 71881 419469 71937 419525
rect 72023 419469 72079 419525
rect 72165 419469 72221 419525
rect 72307 419469 72363 419525
rect 72449 419469 72505 419525
rect 72591 419469 72647 419525
rect 72733 419469 72789 419525
rect 72875 419469 72931 419525
rect 73017 419469 73073 419525
rect 73159 419469 73215 419525
rect 73301 419469 73357 419525
rect 71455 419327 71511 419383
rect 71597 419327 71653 419383
rect 71739 419327 71795 419383
rect 71881 419327 71937 419383
rect 72023 419327 72079 419383
rect 72165 419327 72221 419383
rect 72307 419327 72363 419383
rect 72449 419327 72505 419383
rect 72591 419327 72647 419383
rect 72733 419327 72789 419383
rect 72875 419327 72931 419383
rect 73017 419327 73073 419383
rect 73159 419327 73215 419383
rect 73301 419327 73357 419383
rect 71455 419185 71511 419241
rect 71597 419185 71653 419241
rect 71739 419185 71795 419241
rect 71881 419185 71937 419241
rect 72023 419185 72079 419241
rect 72165 419185 72221 419241
rect 72307 419185 72363 419241
rect 72449 419185 72505 419241
rect 72591 419185 72647 419241
rect 72733 419185 72789 419241
rect 72875 419185 72931 419241
rect 73017 419185 73073 419241
rect 73159 419185 73215 419241
rect 73301 419185 73357 419241
rect 71455 419043 71511 419099
rect 71597 419043 71653 419099
rect 71739 419043 71795 419099
rect 71881 419043 71937 419099
rect 72023 419043 72079 419099
rect 72165 419043 72221 419099
rect 72307 419043 72363 419099
rect 72449 419043 72505 419099
rect 72591 419043 72647 419099
rect 72733 419043 72789 419099
rect 72875 419043 72931 419099
rect 73017 419043 73073 419099
rect 73159 419043 73215 419099
rect 73301 419043 73357 419099
rect 71455 418901 71511 418957
rect 71597 418901 71653 418957
rect 71739 418901 71795 418957
rect 71881 418901 71937 418957
rect 72023 418901 72079 418957
rect 72165 418901 72221 418957
rect 72307 418901 72363 418957
rect 72449 418901 72505 418957
rect 72591 418901 72647 418957
rect 72733 418901 72789 418957
rect 72875 418901 72931 418957
rect 73017 418901 73073 418957
rect 73159 418901 73215 418957
rect 73301 418901 73357 418957
rect 71455 418759 71511 418815
rect 71597 418759 71653 418815
rect 71739 418759 71795 418815
rect 71881 418759 71937 418815
rect 72023 418759 72079 418815
rect 72165 418759 72221 418815
rect 72307 418759 72363 418815
rect 72449 418759 72505 418815
rect 72591 418759 72647 418815
rect 72733 418759 72789 418815
rect 72875 418759 72931 418815
rect 73017 418759 73073 418815
rect 73159 418759 73215 418815
rect 73301 418759 73357 418815
rect 71455 418617 71511 418673
rect 71597 418617 71653 418673
rect 71739 418617 71795 418673
rect 71881 418617 71937 418673
rect 72023 418617 72079 418673
rect 72165 418617 72221 418673
rect 72307 418617 72363 418673
rect 72449 418617 72505 418673
rect 72591 418617 72647 418673
rect 72733 418617 72789 418673
rect 72875 418617 72931 418673
rect 73017 418617 73073 418673
rect 73159 418617 73215 418673
rect 73301 418617 73357 418673
rect 71455 418475 71511 418531
rect 71597 418475 71653 418531
rect 71739 418475 71795 418531
rect 71881 418475 71937 418531
rect 72023 418475 72079 418531
rect 72165 418475 72221 418531
rect 72307 418475 72363 418531
rect 72449 418475 72505 418531
rect 72591 418475 72647 418531
rect 72733 418475 72789 418531
rect 72875 418475 72931 418531
rect 73017 418475 73073 418531
rect 73159 418475 73215 418531
rect 73301 418475 73357 418531
rect 71455 418333 71511 418389
rect 71597 418333 71653 418389
rect 71739 418333 71795 418389
rect 71881 418333 71937 418389
rect 72023 418333 72079 418389
rect 72165 418333 72221 418389
rect 72307 418333 72363 418389
rect 72449 418333 72505 418389
rect 72591 418333 72647 418389
rect 72733 418333 72789 418389
rect 72875 418333 72931 418389
rect 73017 418333 73073 418389
rect 73159 418333 73215 418389
rect 73301 418333 73357 418389
rect 71455 418191 71511 418247
rect 71597 418191 71653 418247
rect 71739 418191 71795 418247
rect 71881 418191 71937 418247
rect 72023 418191 72079 418247
rect 72165 418191 72221 418247
rect 72307 418191 72363 418247
rect 72449 418191 72505 418247
rect 72591 418191 72647 418247
rect 72733 418191 72789 418247
rect 72875 418191 72931 418247
rect 73017 418191 73073 418247
rect 73159 418191 73215 418247
rect 73301 418191 73357 418247
rect 71455 417667 71511 417723
rect 71597 417667 71653 417723
rect 71739 417667 71795 417723
rect 71881 417667 71937 417723
rect 72023 417667 72079 417723
rect 72165 417667 72221 417723
rect 72307 417667 72363 417723
rect 72449 417667 72505 417723
rect 72591 417667 72647 417723
rect 72733 417667 72789 417723
rect 72875 417667 72931 417723
rect 73017 417667 73073 417723
rect 73159 417667 73215 417723
rect 73301 417667 73357 417723
rect 71455 417525 71511 417581
rect 71597 417525 71653 417581
rect 71739 417525 71795 417581
rect 71881 417525 71937 417581
rect 72023 417525 72079 417581
rect 72165 417525 72221 417581
rect 72307 417525 72363 417581
rect 72449 417525 72505 417581
rect 72591 417525 72647 417581
rect 72733 417525 72789 417581
rect 72875 417525 72931 417581
rect 73017 417525 73073 417581
rect 73159 417525 73215 417581
rect 73301 417525 73357 417581
rect 71455 417383 71511 417439
rect 71597 417383 71653 417439
rect 71739 417383 71795 417439
rect 71881 417383 71937 417439
rect 72023 417383 72079 417439
rect 72165 417383 72221 417439
rect 72307 417383 72363 417439
rect 72449 417383 72505 417439
rect 72591 417383 72647 417439
rect 72733 417383 72789 417439
rect 72875 417383 72931 417439
rect 73017 417383 73073 417439
rect 73159 417383 73215 417439
rect 73301 417383 73357 417439
rect 71455 417241 71511 417297
rect 71597 417241 71653 417297
rect 71739 417241 71795 417297
rect 71881 417241 71937 417297
rect 72023 417241 72079 417297
rect 72165 417241 72221 417297
rect 72307 417241 72363 417297
rect 72449 417241 72505 417297
rect 72591 417241 72647 417297
rect 72733 417241 72789 417297
rect 72875 417241 72931 417297
rect 73017 417241 73073 417297
rect 73159 417241 73215 417297
rect 73301 417241 73357 417297
rect 71455 417099 71511 417155
rect 71597 417099 71653 417155
rect 71739 417099 71795 417155
rect 71881 417099 71937 417155
rect 72023 417099 72079 417155
rect 72165 417099 72221 417155
rect 72307 417099 72363 417155
rect 72449 417099 72505 417155
rect 72591 417099 72647 417155
rect 72733 417099 72789 417155
rect 72875 417099 72931 417155
rect 73017 417099 73073 417155
rect 73159 417099 73215 417155
rect 73301 417099 73357 417155
rect 71455 416957 71511 417013
rect 71597 416957 71653 417013
rect 71739 416957 71795 417013
rect 71881 416957 71937 417013
rect 72023 416957 72079 417013
rect 72165 416957 72221 417013
rect 72307 416957 72363 417013
rect 72449 416957 72505 417013
rect 72591 416957 72647 417013
rect 72733 416957 72789 417013
rect 72875 416957 72931 417013
rect 73017 416957 73073 417013
rect 73159 416957 73215 417013
rect 73301 416957 73357 417013
rect 71455 416815 71511 416871
rect 71597 416815 71653 416871
rect 71739 416815 71795 416871
rect 71881 416815 71937 416871
rect 72023 416815 72079 416871
rect 72165 416815 72221 416871
rect 72307 416815 72363 416871
rect 72449 416815 72505 416871
rect 72591 416815 72647 416871
rect 72733 416815 72789 416871
rect 72875 416815 72931 416871
rect 73017 416815 73073 416871
rect 73159 416815 73215 416871
rect 73301 416815 73357 416871
rect 71455 416673 71511 416729
rect 71597 416673 71653 416729
rect 71739 416673 71795 416729
rect 71881 416673 71937 416729
rect 72023 416673 72079 416729
rect 72165 416673 72221 416729
rect 72307 416673 72363 416729
rect 72449 416673 72505 416729
rect 72591 416673 72647 416729
rect 72733 416673 72789 416729
rect 72875 416673 72931 416729
rect 73017 416673 73073 416729
rect 73159 416673 73215 416729
rect 73301 416673 73357 416729
rect 71455 416531 71511 416587
rect 71597 416531 71653 416587
rect 71739 416531 71795 416587
rect 71881 416531 71937 416587
rect 72023 416531 72079 416587
rect 72165 416531 72221 416587
rect 72307 416531 72363 416587
rect 72449 416531 72505 416587
rect 72591 416531 72647 416587
rect 72733 416531 72789 416587
rect 72875 416531 72931 416587
rect 73017 416531 73073 416587
rect 73159 416531 73215 416587
rect 73301 416531 73357 416587
rect 71455 416389 71511 416445
rect 71597 416389 71653 416445
rect 71739 416389 71795 416445
rect 71881 416389 71937 416445
rect 72023 416389 72079 416445
rect 72165 416389 72221 416445
rect 72307 416389 72363 416445
rect 72449 416389 72505 416445
rect 72591 416389 72647 416445
rect 72733 416389 72789 416445
rect 72875 416389 72931 416445
rect 73017 416389 73073 416445
rect 73159 416389 73215 416445
rect 73301 416389 73357 416445
rect 71455 416247 71511 416303
rect 71597 416247 71653 416303
rect 71739 416247 71795 416303
rect 71881 416247 71937 416303
rect 72023 416247 72079 416303
rect 72165 416247 72221 416303
rect 72307 416247 72363 416303
rect 72449 416247 72505 416303
rect 72591 416247 72647 416303
rect 72733 416247 72789 416303
rect 72875 416247 72931 416303
rect 73017 416247 73073 416303
rect 73159 416247 73215 416303
rect 73301 416247 73357 416303
rect 71455 416105 71511 416161
rect 71597 416105 71653 416161
rect 71739 416105 71795 416161
rect 71881 416105 71937 416161
rect 72023 416105 72079 416161
rect 72165 416105 72221 416161
rect 72307 416105 72363 416161
rect 72449 416105 72505 416161
rect 72591 416105 72647 416161
rect 72733 416105 72789 416161
rect 72875 416105 72931 416161
rect 73017 416105 73073 416161
rect 73159 416105 73215 416161
rect 73301 416105 73357 416161
rect 71455 415963 71511 416019
rect 71597 415963 71653 416019
rect 71739 415963 71795 416019
rect 71881 415963 71937 416019
rect 72023 415963 72079 416019
rect 72165 415963 72221 416019
rect 72307 415963 72363 416019
rect 72449 415963 72505 416019
rect 72591 415963 72647 416019
rect 72733 415963 72789 416019
rect 72875 415963 72931 416019
rect 73017 415963 73073 416019
rect 73159 415963 73215 416019
rect 73301 415963 73357 416019
rect 71455 415821 71511 415877
rect 71597 415821 71653 415877
rect 71739 415821 71795 415877
rect 71881 415821 71937 415877
rect 72023 415821 72079 415877
rect 72165 415821 72221 415877
rect 72307 415821 72363 415877
rect 72449 415821 72505 415877
rect 72591 415821 72647 415877
rect 72733 415821 72789 415877
rect 72875 415821 72931 415877
rect 73017 415821 73073 415877
rect 73159 415821 73215 415877
rect 73301 415821 73357 415877
rect 71466 415038 71522 415094
rect 71608 415038 71664 415094
rect 71750 415038 71806 415094
rect 71892 415038 71948 415094
rect 72034 415038 72090 415094
rect 72176 415038 72232 415094
rect 72318 415038 72374 415094
rect 72460 415038 72516 415094
rect 72602 415038 72658 415094
rect 72744 415038 72800 415094
rect 72886 415038 72942 415094
rect 73028 415038 73084 415094
rect 73170 415038 73226 415094
rect 73312 415038 73368 415094
rect 71466 414896 71522 414952
rect 71608 414896 71664 414952
rect 71750 414896 71806 414952
rect 71892 414896 71948 414952
rect 72034 414896 72090 414952
rect 72176 414896 72232 414952
rect 72318 414896 72374 414952
rect 72460 414896 72516 414952
rect 72602 414896 72658 414952
rect 72744 414896 72800 414952
rect 72886 414896 72942 414952
rect 73028 414896 73084 414952
rect 73170 414896 73226 414952
rect 73312 414896 73368 414952
rect 71466 414754 71522 414810
rect 71608 414754 71664 414810
rect 71750 414754 71806 414810
rect 71892 414754 71948 414810
rect 72034 414754 72090 414810
rect 72176 414754 72232 414810
rect 72318 414754 72374 414810
rect 72460 414754 72516 414810
rect 72602 414754 72658 414810
rect 72744 414754 72800 414810
rect 72886 414754 72942 414810
rect 73028 414754 73084 414810
rect 73170 414754 73226 414810
rect 73312 414754 73368 414810
rect 71466 414612 71522 414668
rect 71608 414612 71664 414668
rect 71750 414612 71806 414668
rect 71892 414612 71948 414668
rect 72034 414612 72090 414668
rect 72176 414612 72232 414668
rect 72318 414612 72374 414668
rect 72460 414612 72516 414668
rect 72602 414612 72658 414668
rect 72744 414612 72800 414668
rect 72886 414612 72942 414668
rect 73028 414612 73084 414668
rect 73170 414612 73226 414668
rect 73312 414612 73368 414668
rect 71466 414470 71522 414526
rect 71608 414470 71664 414526
rect 71750 414470 71806 414526
rect 71892 414470 71948 414526
rect 72034 414470 72090 414526
rect 72176 414470 72232 414526
rect 72318 414470 72374 414526
rect 72460 414470 72516 414526
rect 72602 414470 72658 414526
rect 72744 414470 72800 414526
rect 72886 414470 72942 414526
rect 73028 414470 73084 414526
rect 73170 414470 73226 414526
rect 73312 414470 73368 414526
rect 71466 414328 71522 414384
rect 71608 414328 71664 414384
rect 71750 414328 71806 414384
rect 71892 414328 71948 414384
rect 72034 414328 72090 414384
rect 72176 414328 72232 414384
rect 72318 414328 72374 414384
rect 72460 414328 72516 414384
rect 72602 414328 72658 414384
rect 72744 414328 72800 414384
rect 72886 414328 72942 414384
rect 73028 414328 73084 414384
rect 73170 414328 73226 414384
rect 73312 414328 73368 414384
rect 71466 414186 71522 414242
rect 71608 414186 71664 414242
rect 71750 414186 71806 414242
rect 71892 414186 71948 414242
rect 72034 414186 72090 414242
rect 72176 414186 72232 414242
rect 72318 414186 72374 414242
rect 72460 414186 72516 414242
rect 72602 414186 72658 414242
rect 72744 414186 72800 414242
rect 72886 414186 72942 414242
rect 73028 414186 73084 414242
rect 73170 414186 73226 414242
rect 73312 414186 73368 414242
rect 71466 414044 71522 414100
rect 71608 414044 71664 414100
rect 71750 414044 71806 414100
rect 71892 414044 71948 414100
rect 72034 414044 72090 414100
rect 72176 414044 72232 414100
rect 72318 414044 72374 414100
rect 72460 414044 72516 414100
rect 72602 414044 72658 414100
rect 72744 414044 72800 414100
rect 72886 414044 72942 414100
rect 73028 414044 73084 414100
rect 73170 414044 73226 414100
rect 73312 414044 73368 414100
rect 71466 413902 71522 413958
rect 71608 413902 71664 413958
rect 71750 413902 71806 413958
rect 71892 413902 71948 413958
rect 72034 413902 72090 413958
rect 72176 413902 72232 413958
rect 72318 413902 72374 413958
rect 72460 413902 72516 413958
rect 72602 413902 72658 413958
rect 72744 413902 72800 413958
rect 72886 413902 72942 413958
rect 73028 413902 73084 413958
rect 73170 413902 73226 413958
rect 73312 413902 73368 413958
rect 71466 413760 71522 413816
rect 71608 413760 71664 413816
rect 71750 413760 71806 413816
rect 71892 413760 71948 413816
rect 72034 413760 72090 413816
rect 72176 413760 72232 413816
rect 72318 413760 72374 413816
rect 72460 413760 72516 413816
rect 72602 413760 72658 413816
rect 72744 413760 72800 413816
rect 72886 413760 72942 413816
rect 73028 413760 73084 413816
rect 73170 413760 73226 413816
rect 73312 413760 73368 413816
rect 71466 413618 71522 413674
rect 71608 413618 71664 413674
rect 71750 413618 71806 413674
rect 71892 413618 71948 413674
rect 72034 413618 72090 413674
rect 72176 413618 72232 413674
rect 72318 413618 72374 413674
rect 72460 413618 72516 413674
rect 72602 413618 72658 413674
rect 72744 413618 72800 413674
rect 72886 413618 72942 413674
rect 73028 413618 73084 413674
rect 73170 413618 73226 413674
rect 73312 413618 73368 413674
rect 71466 413476 71522 413532
rect 71608 413476 71664 413532
rect 71750 413476 71806 413532
rect 71892 413476 71948 413532
rect 72034 413476 72090 413532
rect 72176 413476 72232 413532
rect 72318 413476 72374 413532
rect 72460 413476 72516 413532
rect 72602 413476 72658 413532
rect 72744 413476 72800 413532
rect 72886 413476 72942 413532
rect 73028 413476 73084 413532
rect 73170 413476 73226 413532
rect 73312 413476 73368 413532
rect 71466 413334 71522 413390
rect 71608 413334 71664 413390
rect 71750 413334 71806 413390
rect 71892 413334 71948 413390
rect 72034 413334 72090 413390
rect 72176 413334 72232 413390
rect 72318 413334 72374 413390
rect 72460 413334 72516 413390
rect 72602 413334 72658 413390
rect 72744 413334 72800 413390
rect 72886 413334 72942 413390
rect 73028 413334 73084 413390
rect 73170 413334 73226 413390
rect 73312 413334 73368 413390
rect 702440 404610 702496 404666
rect 702582 404610 702638 404666
rect 702724 404610 702780 404666
rect 702866 404610 702922 404666
rect 703008 404610 703064 404666
rect 703150 404610 703206 404666
rect 703292 404610 703348 404666
rect 703434 404610 703490 404666
rect 703576 404610 703632 404666
rect 703718 404610 703774 404666
rect 703860 404610 703916 404666
rect 704002 404610 704058 404666
rect 704144 404610 704200 404666
rect 704286 404610 704342 404666
rect 702440 404468 702496 404524
rect 702582 404468 702638 404524
rect 702724 404468 702780 404524
rect 702866 404468 702922 404524
rect 703008 404468 703064 404524
rect 703150 404468 703206 404524
rect 703292 404468 703348 404524
rect 703434 404468 703490 404524
rect 703576 404468 703632 404524
rect 703718 404468 703774 404524
rect 703860 404468 703916 404524
rect 704002 404468 704058 404524
rect 704144 404468 704200 404524
rect 704286 404468 704342 404524
rect 702440 404326 702496 404382
rect 702582 404326 702638 404382
rect 702724 404326 702780 404382
rect 702866 404326 702922 404382
rect 703008 404326 703064 404382
rect 703150 404326 703206 404382
rect 703292 404326 703348 404382
rect 703434 404326 703490 404382
rect 703576 404326 703632 404382
rect 703718 404326 703774 404382
rect 703860 404326 703916 404382
rect 704002 404326 704058 404382
rect 704144 404326 704200 404382
rect 704286 404326 704342 404382
rect 702440 404184 702496 404240
rect 702582 404184 702638 404240
rect 702724 404184 702780 404240
rect 702866 404184 702922 404240
rect 703008 404184 703064 404240
rect 703150 404184 703206 404240
rect 703292 404184 703348 404240
rect 703434 404184 703490 404240
rect 703576 404184 703632 404240
rect 703718 404184 703774 404240
rect 703860 404184 703916 404240
rect 704002 404184 704058 404240
rect 704144 404184 704200 404240
rect 704286 404184 704342 404240
rect 702440 404042 702496 404098
rect 702582 404042 702638 404098
rect 702724 404042 702780 404098
rect 702866 404042 702922 404098
rect 703008 404042 703064 404098
rect 703150 404042 703206 404098
rect 703292 404042 703348 404098
rect 703434 404042 703490 404098
rect 703576 404042 703632 404098
rect 703718 404042 703774 404098
rect 703860 404042 703916 404098
rect 704002 404042 704058 404098
rect 704144 404042 704200 404098
rect 704286 404042 704342 404098
rect 702440 403900 702496 403956
rect 702582 403900 702638 403956
rect 702724 403900 702780 403956
rect 702866 403900 702922 403956
rect 703008 403900 703064 403956
rect 703150 403900 703206 403956
rect 703292 403900 703348 403956
rect 703434 403900 703490 403956
rect 703576 403900 703632 403956
rect 703718 403900 703774 403956
rect 703860 403900 703916 403956
rect 704002 403900 704058 403956
rect 704144 403900 704200 403956
rect 704286 403900 704342 403956
rect 702440 403758 702496 403814
rect 702582 403758 702638 403814
rect 702724 403758 702780 403814
rect 702866 403758 702922 403814
rect 703008 403758 703064 403814
rect 703150 403758 703206 403814
rect 703292 403758 703348 403814
rect 703434 403758 703490 403814
rect 703576 403758 703632 403814
rect 703718 403758 703774 403814
rect 703860 403758 703916 403814
rect 704002 403758 704058 403814
rect 704144 403758 704200 403814
rect 704286 403758 704342 403814
rect 702440 403616 702496 403672
rect 702582 403616 702638 403672
rect 702724 403616 702780 403672
rect 702866 403616 702922 403672
rect 703008 403616 703064 403672
rect 703150 403616 703206 403672
rect 703292 403616 703348 403672
rect 703434 403616 703490 403672
rect 703576 403616 703632 403672
rect 703718 403616 703774 403672
rect 703860 403616 703916 403672
rect 704002 403616 704058 403672
rect 704144 403616 704200 403672
rect 704286 403616 704342 403672
rect 702440 403474 702496 403530
rect 702582 403474 702638 403530
rect 702724 403474 702780 403530
rect 702866 403474 702922 403530
rect 703008 403474 703064 403530
rect 703150 403474 703206 403530
rect 703292 403474 703348 403530
rect 703434 403474 703490 403530
rect 703576 403474 703632 403530
rect 703718 403474 703774 403530
rect 703860 403474 703916 403530
rect 704002 403474 704058 403530
rect 704144 403474 704200 403530
rect 704286 403474 704342 403530
rect 702440 403332 702496 403388
rect 702582 403332 702638 403388
rect 702724 403332 702780 403388
rect 702866 403332 702922 403388
rect 703008 403332 703064 403388
rect 703150 403332 703206 403388
rect 703292 403332 703348 403388
rect 703434 403332 703490 403388
rect 703576 403332 703632 403388
rect 703718 403332 703774 403388
rect 703860 403332 703916 403388
rect 704002 403332 704058 403388
rect 704144 403332 704200 403388
rect 704286 403332 704342 403388
rect 702440 403190 702496 403246
rect 702582 403190 702638 403246
rect 702724 403190 702780 403246
rect 702866 403190 702922 403246
rect 703008 403190 703064 403246
rect 703150 403190 703206 403246
rect 703292 403190 703348 403246
rect 703434 403190 703490 403246
rect 703576 403190 703632 403246
rect 703718 403190 703774 403246
rect 703860 403190 703916 403246
rect 704002 403190 704058 403246
rect 704144 403190 704200 403246
rect 704286 403190 704342 403246
rect 702440 403048 702496 403104
rect 702582 403048 702638 403104
rect 702724 403048 702780 403104
rect 702866 403048 702922 403104
rect 703008 403048 703064 403104
rect 703150 403048 703206 403104
rect 703292 403048 703348 403104
rect 703434 403048 703490 403104
rect 703576 403048 703632 403104
rect 703718 403048 703774 403104
rect 703860 403048 703916 403104
rect 704002 403048 704058 403104
rect 704144 403048 704200 403104
rect 704286 403048 704342 403104
rect 702440 402906 702496 402962
rect 702582 402906 702638 402962
rect 702724 402906 702780 402962
rect 702866 402906 702922 402962
rect 703008 402906 703064 402962
rect 703150 402906 703206 402962
rect 703292 402906 703348 402962
rect 703434 402906 703490 402962
rect 703576 402906 703632 402962
rect 703718 402906 703774 402962
rect 703860 402906 703916 402962
rect 704002 402906 704058 402962
rect 704144 402906 704200 402962
rect 704286 402906 704342 402962
rect 702451 402123 702507 402179
rect 702593 402123 702649 402179
rect 702735 402123 702791 402179
rect 702877 402123 702933 402179
rect 703019 402123 703075 402179
rect 703161 402123 703217 402179
rect 703303 402123 703359 402179
rect 703445 402123 703501 402179
rect 703587 402123 703643 402179
rect 703729 402123 703785 402179
rect 703871 402123 703927 402179
rect 704013 402123 704069 402179
rect 704155 402123 704211 402179
rect 704297 402123 704353 402179
rect 702451 401981 702507 402037
rect 702593 401981 702649 402037
rect 702735 401981 702791 402037
rect 702877 401981 702933 402037
rect 703019 401981 703075 402037
rect 703161 401981 703217 402037
rect 703303 401981 703359 402037
rect 703445 401981 703501 402037
rect 703587 401981 703643 402037
rect 703729 401981 703785 402037
rect 703871 401981 703927 402037
rect 704013 401981 704069 402037
rect 704155 401981 704211 402037
rect 704297 401981 704353 402037
rect 702451 401839 702507 401895
rect 702593 401839 702649 401895
rect 702735 401839 702791 401895
rect 702877 401839 702933 401895
rect 703019 401839 703075 401895
rect 703161 401839 703217 401895
rect 703303 401839 703359 401895
rect 703445 401839 703501 401895
rect 703587 401839 703643 401895
rect 703729 401839 703785 401895
rect 703871 401839 703927 401895
rect 704013 401839 704069 401895
rect 704155 401839 704211 401895
rect 704297 401839 704353 401895
rect 702451 401697 702507 401753
rect 702593 401697 702649 401753
rect 702735 401697 702791 401753
rect 702877 401697 702933 401753
rect 703019 401697 703075 401753
rect 703161 401697 703217 401753
rect 703303 401697 703359 401753
rect 703445 401697 703501 401753
rect 703587 401697 703643 401753
rect 703729 401697 703785 401753
rect 703871 401697 703927 401753
rect 704013 401697 704069 401753
rect 704155 401697 704211 401753
rect 704297 401697 704353 401753
rect 702451 401555 702507 401611
rect 702593 401555 702649 401611
rect 702735 401555 702791 401611
rect 702877 401555 702933 401611
rect 703019 401555 703075 401611
rect 703161 401555 703217 401611
rect 703303 401555 703359 401611
rect 703445 401555 703501 401611
rect 703587 401555 703643 401611
rect 703729 401555 703785 401611
rect 703871 401555 703927 401611
rect 704013 401555 704069 401611
rect 704155 401555 704211 401611
rect 704297 401555 704353 401611
rect 702451 401413 702507 401469
rect 702593 401413 702649 401469
rect 702735 401413 702791 401469
rect 702877 401413 702933 401469
rect 703019 401413 703075 401469
rect 703161 401413 703217 401469
rect 703303 401413 703359 401469
rect 703445 401413 703501 401469
rect 703587 401413 703643 401469
rect 703729 401413 703785 401469
rect 703871 401413 703927 401469
rect 704013 401413 704069 401469
rect 704155 401413 704211 401469
rect 704297 401413 704353 401469
rect 702451 401271 702507 401327
rect 702593 401271 702649 401327
rect 702735 401271 702791 401327
rect 702877 401271 702933 401327
rect 703019 401271 703075 401327
rect 703161 401271 703217 401327
rect 703303 401271 703359 401327
rect 703445 401271 703501 401327
rect 703587 401271 703643 401327
rect 703729 401271 703785 401327
rect 703871 401271 703927 401327
rect 704013 401271 704069 401327
rect 704155 401271 704211 401327
rect 704297 401271 704353 401327
rect 702451 401129 702507 401185
rect 702593 401129 702649 401185
rect 702735 401129 702791 401185
rect 702877 401129 702933 401185
rect 703019 401129 703075 401185
rect 703161 401129 703217 401185
rect 703303 401129 703359 401185
rect 703445 401129 703501 401185
rect 703587 401129 703643 401185
rect 703729 401129 703785 401185
rect 703871 401129 703927 401185
rect 704013 401129 704069 401185
rect 704155 401129 704211 401185
rect 704297 401129 704353 401185
rect 702451 400987 702507 401043
rect 702593 400987 702649 401043
rect 702735 400987 702791 401043
rect 702877 400987 702933 401043
rect 703019 400987 703075 401043
rect 703161 400987 703217 401043
rect 703303 400987 703359 401043
rect 703445 400987 703501 401043
rect 703587 400987 703643 401043
rect 703729 400987 703785 401043
rect 703871 400987 703927 401043
rect 704013 400987 704069 401043
rect 704155 400987 704211 401043
rect 704297 400987 704353 401043
rect 702451 400845 702507 400901
rect 702593 400845 702649 400901
rect 702735 400845 702791 400901
rect 702877 400845 702933 400901
rect 703019 400845 703075 400901
rect 703161 400845 703217 400901
rect 703303 400845 703359 400901
rect 703445 400845 703501 400901
rect 703587 400845 703643 400901
rect 703729 400845 703785 400901
rect 703871 400845 703927 400901
rect 704013 400845 704069 400901
rect 704155 400845 704211 400901
rect 704297 400845 704353 400901
rect 702451 400703 702507 400759
rect 702593 400703 702649 400759
rect 702735 400703 702791 400759
rect 702877 400703 702933 400759
rect 703019 400703 703075 400759
rect 703161 400703 703217 400759
rect 703303 400703 703359 400759
rect 703445 400703 703501 400759
rect 703587 400703 703643 400759
rect 703729 400703 703785 400759
rect 703871 400703 703927 400759
rect 704013 400703 704069 400759
rect 704155 400703 704211 400759
rect 704297 400703 704353 400759
rect 702451 400561 702507 400617
rect 702593 400561 702649 400617
rect 702735 400561 702791 400617
rect 702877 400561 702933 400617
rect 703019 400561 703075 400617
rect 703161 400561 703217 400617
rect 703303 400561 703359 400617
rect 703445 400561 703501 400617
rect 703587 400561 703643 400617
rect 703729 400561 703785 400617
rect 703871 400561 703927 400617
rect 704013 400561 704069 400617
rect 704155 400561 704211 400617
rect 704297 400561 704353 400617
rect 702451 400419 702507 400475
rect 702593 400419 702649 400475
rect 702735 400419 702791 400475
rect 702877 400419 702933 400475
rect 703019 400419 703075 400475
rect 703161 400419 703217 400475
rect 703303 400419 703359 400475
rect 703445 400419 703501 400475
rect 703587 400419 703643 400475
rect 703729 400419 703785 400475
rect 703871 400419 703927 400475
rect 704013 400419 704069 400475
rect 704155 400419 704211 400475
rect 704297 400419 704353 400475
rect 702451 400277 702507 400333
rect 702593 400277 702649 400333
rect 702735 400277 702791 400333
rect 702877 400277 702933 400333
rect 703019 400277 703075 400333
rect 703161 400277 703217 400333
rect 703303 400277 703359 400333
rect 703445 400277 703501 400333
rect 703587 400277 703643 400333
rect 703729 400277 703785 400333
rect 703871 400277 703927 400333
rect 704013 400277 704069 400333
rect 704155 400277 704211 400333
rect 704297 400277 704353 400333
rect 702451 399753 702507 399809
rect 702593 399753 702649 399809
rect 702735 399753 702791 399809
rect 702877 399753 702933 399809
rect 703019 399753 703075 399809
rect 703161 399753 703217 399809
rect 703303 399753 703359 399809
rect 703445 399753 703501 399809
rect 703587 399753 703643 399809
rect 703729 399753 703785 399809
rect 703871 399753 703927 399809
rect 704013 399753 704069 399809
rect 704155 399753 704211 399809
rect 704297 399753 704353 399809
rect 702451 399611 702507 399667
rect 702593 399611 702649 399667
rect 702735 399611 702791 399667
rect 702877 399611 702933 399667
rect 703019 399611 703075 399667
rect 703161 399611 703217 399667
rect 703303 399611 703359 399667
rect 703445 399611 703501 399667
rect 703587 399611 703643 399667
rect 703729 399611 703785 399667
rect 703871 399611 703927 399667
rect 704013 399611 704069 399667
rect 704155 399611 704211 399667
rect 704297 399611 704353 399667
rect 702451 399469 702507 399525
rect 702593 399469 702649 399525
rect 702735 399469 702791 399525
rect 702877 399469 702933 399525
rect 703019 399469 703075 399525
rect 703161 399469 703217 399525
rect 703303 399469 703359 399525
rect 703445 399469 703501 399525
rect 703587 399469 703643 399525
rect 703729 399469 703785 399525
rect 703871 399469 703927 399525
rect 704013 399469 704069 399525
rect 704155 399469 704211 399525
rect 704297 399469 704353 399525
rect 702451 399327 702507 399383
rect 702593 399327 702649 399383
rect 702735 399327 702791 399383
rect 702877 399327 702933 399383
rect 703019 399327 703075 399383
rect 703161 399327 703217 399383
rect 703303 399327 703359 399383
rect 703445 399327 703501 399383
rect 703587 399327 703643 399383
rect 703729 399327 703785 399383
rect 703871 399327 703927 399383
rect 704013 399327 704069 399383
rect 704155 399327 704211 399383
rect 704297 399327 704353 399383
rect 702451 399185 702507 399241
rect 702593 399185 702649 399241
rect 702735 399185 702791 399241
rect 702877 399185 702933 399241
rect 703019 399185 703075 399241
rect 703161 399185 703217 399241
rect 703303 399185 703359 399241
rect 703445 399185 703501 399241
rect 703587 399185 703643 399241
rect 703729 399185 703785 399241
rect 703871 399185 703927 399241
rect 704013 399185 704069 399241
rect 704155 399185 704211 399241
rect 704297 399185 704353 399241
rect 702451 399043 702507 399099
rect 702593 399043 702649 399099
rect 702735 399043 702791 399099
rect 702877 399043 702933 399099
rect 703019 399043 703075 399099
rect 703161 399043 703217 399099
rect 703303 399043 703359 399099
rect 703445 399043 703501 399099
rect 703587 399043 703643 399099
rect 703729 399043 703785 399099
rect 703871 399043 703927 399099
rect 704013 399043 704069 399099
rect 704155 399043 704211 399099
rect 704297 399043 704353 399099
rect 702451 398901 702507 398957
rect 702593 398901 702649 398957
rect 702735 398901 702791 398957
rect 702877 398901 702933 398957
rect 703019 398901 703075 398957
rect 703161 398901 703217 398957
rect 703303 398901 703359 398957
rect 703445 398901 703501 398957
rect 703587 398901 703643 398957
rect 703729 398901 703785 398957
rect 703871 398901 703927 398957
rect 704013 398901 704069 398957
rect 704155 398901 704211 398957
rect 704297 398901 704353 398957
rect 702451 398759 702507 398815
rect 702593 398759 702649 398815
rect 702735 398759 702791 398815
rect 702877 398759 702933 398815
rect 703019 398759 703075 398815
rect 703161 398759 703217 398815
rect 703303 398759 703359 398815
rect 703445 398759 703501 398815
rect 703587 398759 703643 398815
rect 703729 398759 703785 398815
rect 703871 398759 703927 398815
rect 704013 398759 704069 398815
rect 704155 398759 704211 398815
rect 704297 398759 704353 398815
rect 702451 398617 702507 398673
rect 702593 398617 702649 398673
rect 702735 398617 702791 398673
rect 702877 398617 702933 398673
rect 703019 398617 703075 398673
rect 703161 398617 703217 398673
rect 703303 398617 703359 398673
rect 703445 398617 703501 398673
rect 703587 398617 703643 398673
rect 703729 398617 703785 398673
rect 703871 398617 703927 398673
rect 704013 398617 704069 398673
rect 704155 398617 704211 398673
rect 704297 398617 704353 398673
rect 702451 398475 702507 398531
rect 702593 398475 702649 398531
rect 702735 398475 702791 398531
rect 702877 398475 702933 398531
rect 703019 398475 703075 398531
rect 703161 398475 703217 398531
rect 703303 398475 703359 398531
rect 703445 398475 703501 398531
rect 703587 398475 703643 398531
rect 703729 398475 703785 398531
rect 703871 398475 703927 398531
rect 704013 398475 704069 398531
rect 704155 398475 704211 398531
rect 704297 398475 704353 398531
rect 702451 398333 702507 398389
rect 702593 398333 702649 398389
rect 702735 398333 702791 398389
rect 702877 398333 702933 398389
rect 703019 398333 703075 398389
rect 703161 398333 703217 398389
rect 703303 398333 703359 398389
rect 703445 398333 703501 398389
rect 703587 398333 703643 398389
rect 703729 398333 703785 398389
rect 703871 398333 703927 398389
rect 704013 398333 704069 398389
rect 704155 398333 704211 398389
rect 704297 398333 704353 398389
rect 702451 398191 702507 398247
rect 702593 398191 702649 398247
rect 702735 398191 702791 398247
rect 702877 398191 702933 398247
rect 703019 398191 703075 398247
rect 703161 398191 703217 398247
rect 703303 398191 703359 398247
rect 703445 398191 703501 398247
rect 703587 398191 703643 398247
rect 703729 398191 703785 398247
rect 703871 398191 703927 398247
rect 704013 398191 704069 398247
rect 704155 398191 704211 398247
rect 704297 398191 704353 398247
rect 702451 398049 702507 398105
rect 702593 398049 702649 398105
rect 702735 398049 702791 398105
rect 702877 398049 702933 398105
rect 703019 398049 703075 398105
rect 703161 398049 703217 398105
rect 703303 398049 703359 398105
rect 703445 398049 703501 398105
rect 703587 398049 703643 398105
rect 703729 398049 703785 398105
rect 703871 398049 703927 398105
rect 704013 398049 704069 398105
rect 704155 398049 704211 398105
rect 704297 398049 704353 398105
rect 702451 397907 702507 397963
rect 702593 397907 702649 397963
rect 702735 397907 702791 397963
rect 702877 397907 702933 397963
rect 703019 397907 703075 397963
rect 703161 397907 703217 397963
rect 703303 397907 703359 397963
rect 703445 397907 703501 397963
rect 703587 397907 703643 397963
rect 703729 397907 703785 397963
rect 703871 397907 703927 397963
rect 704013 397907 704069 397963
rect 704155 397907 704211 397963
rect 704297 397907 704353 397963
rect 702451 397047 702507 397103
rect 702593 397047 702649 397103
rect 702735 397047 702791 397103
rect 702877 397047 702933 397103
rect 703019 397047 703075 397103
rect 703161 397047 703217 397103
rect 703303 397047 703359 397103
rect 703445 397047 703501 397103
rect 703587 397047 703643 397103
rect 703729 397047 703785 397103
rect 703871 397047 703927 397103
rect 704013 397047 704069 397103
rect 704155 397047 704211 397103
rect 704297 397047 704353 397103
rect 702451 396905 702507 396961
rect 702593 396905 702649 396961
rect 702735 396905 702791 396961
rect 702877 396905 702933 396961
rect 703019 396905 703075 396961
rect 703161 396905 703217 396961
rect 703303 396905 703359 396961
rect 703445 396905 703501 396961
rect 703587 396905 703643 396961
rect 703729 396905 703785 396961
rect 703871 396905 703927 396961
rect 704013 396905 704069 396961
rect 704155 396905 704211 396961
rect 704297 396905 704353 396961
rect 702451 396763 702507 396819
rect 702593 396763 702649 396819
rect 702735 396763 702791 396819
rect 702877 396763 702933 396819
rect 703019 396763 703075 396819
rect 703161 396763 703217 396819
rect 703303 396763 703359 396819
rect 703445 396763 703501 396819
rect 703587 396763 703643 396819
rect 703729 396763 703785 396819
rect 703871 396763 703927 396819
rect 704013 396763 704069 396819
rect 704155 396763 704211 396819
rect 704297 396763 704353 396819
rect 702451 396621 702507 396677
rect 702593 396621 702649 396677
rect 702735 396621 702791 396677
rect 702877 396621 702933 396677
rect 703019 396621 703075 396677
rect 703161 396621 703217 396677
rect 703303 396621 703359 396677
rect 703445 396621 703501 396677
rect 703587 396621 703643 396677
rect 703729 396621 703785 396677
rect 703871 396621 703927 396677
rect 704013 396621 704069 396677
rect 704155 396621 704211 396677
rect 704297 396621 704353 396677
rect 702451 396479 702507 396535
rect 702593 396479 702649 396535
rect 702735 396479 702791 396535
rect 702877 396479 702933 396535
rect 703019 396479 703075 396535
rect 703161 396479 703217 396535
rect 703303 396479 703359 396535
rect 703445 396479 703501 396535
rect 703587 396479 703643 396535
rect 703729 396479 703785 396535
rect 703871 396479 703927 396535
rect 704013 396479 704069 396535
rect 704155 396479 704211 396535
rect 704297 396479 704353 396535
rect 702451 396337 702507 396393
rect 702593 396337 702649 396393
rect 702735 396337 702791 396393
rect 702877 396337 702933 396393
rect 703019 396337 703075 396393
rect 703161 396337 703217 396393
rect 703303 396337 703359 396393
rect 703445 396337 703501 396393
rect 703587 396337 703643 396393
rect 703729 396337 703785 396393
rect 703871 396337 703927 396393
rect 704013 396337 704069 396393
rect 704155 396337 704211 396393
rect 704297 396337 704353 396393
rect 702451 396195 702507 396251
rect 702593 396195 702649 396251
rect 702735 396195 702791 396251
rect 702877 396195 702933 396251
rect 703019 396195 703075 396251
rect 703161 396195 703217 396251
rect 703303 396195 703359 396251
rect 703445 396195 703501 396251
rect 703587 396195 703643 396251
rect 703729 396195 703785 396251
rect 703871 396195 703927 396251
rect 704013 396195 704069 396251
rect 704155 396195 704211 396251
rect 704297 396195 704353 396251
rect 702451 396053 702507 396109
rect 702593 396053 702649 396109
rect 702735 396053 702791 396109
rect 702877 396053 702933 396109
rect 703019 396053 703075 396109
rect 703161 396053 703217 396109
rect 703303 396053 703359 396109
rect 703445 396053 703501 396109
rect 703587 396053 703643 396109
rect 703729 396053 703785 396109
rect 703871 396053 703927 396109
rect 704013 396053 704069 396109
rect 704155 396053 704211 396109
rect 704297 396053 704353 396109
rect 702451 395911 702507 395967
rect 702593 395911 702649 395967
rect 702735 395911 702791 395967
rect 702877 395911 702933 395967
rect 703019 395911 703075 395967
rect 703161 395911 703217 395967
rect 703303 395911 703359 395967
rect 703445 395911 703501 395967
rect 703587 395911 703643 395967
rect 703729 395911 703785 395967
rect 703871 395911 703927 395967
rect 704013 395911 704069 395967
rect 704155 395911 704211 395967
rect 704297 395911 704353 395967
rect 702451 395769 702507 395825
rect 702593 395769 702649 395825
rect 702735 395769 702791 395825
rect 702877 395769 702933 395825
rect 703019 395769 703075 395825
rect 703161 395769 703217 395825
rect 703303 395769 703359 395825
rect 703445 395769 703501 395825
rect 703587 395769 703643 395825
rect 703729 395769 703785 395825
rect 703871 395769 703927 395825
rect 704013 395769 704069 395825
rect 704155 395769 704211 395825
rect 704297 395769 704353 395825
rect 702451 395627 702507 395683
rect 702593 395627 702649 395683
rect 702735 395627 702791 395683
rect 702877 395627 702933 395683
rect 703019 395627 703075 395683
rect 703161 395627 703217 395683
rect 703303 395627 703359 395683
rect 703445 395627 703501 395683
rect 703587 395627 703643 395683
rect 703729 395627 703785 395683
rect 703871 395627 703927 395683
rect 704013 395627 704069 395683
rect 704155 395627 704211 395683
rect 704297 395627 704353 395683
rect 702451 395485 702507 395541
rect 702593 395485 702649 395541
rect 702735 395485 702791 395541
rect 702877 395485 702933 395541
rect 703019 395485 703075 395541
rect 703161 395485 703217 395541
rect 703303 395485 703359 395541
rect 703445 395485 703501 395541
rect 703587 395485 703643 395541
rect 703729 395485 703785 395541
rect 703871 395485 703927 395541
rect 704013 395485 704069 395541
rect 704155 395485 704211 395541
rect 704297 395485 704353 395541
rect 702451 395343 702507 395399
rect 702593 395343 702649 395399
rect 702735 395343 702791 395399
rect 702877 395343 702933 395399
rect 703019 395343 703075 395399
rect 703161 395343 703217 395399
rect 703303 395343 703359 395399
rect 703445 395343 703501 395399
rect 703587 395343 703643 395399
rect 703729 395343 703785 395399
rect 703871 395343 703927 395399
rect 704013 395343 704069 395399
rect 704155 395343 704211 395399
rect 704297 395343 704353 395399
rect 702451 395201 702507 395257
rect 702593 395201 702649 395257
rect 702735 395201 702791 395257
rect 702877 395201 702933 395257
rect 703019 395201 703075 395257
rect 703161 395201 703217 395257
rect 703303 395201 703359 395257
rect 703445 395201 703501 395257
rect 703587 395201 703643 395257
rect 703729 395201 703785 395257
rect 703871 395201 703927 395257
rect 704013 395201 704069 395257
rect 704155 395201 704211 395257
rect 704297 395201 704353 395257
rect 702451 394677 702507 394733
rect 702593 394677 702649 394733
rect 702735 394677 702791 394733
rect 702877 394677 702933 394733
rect 703019 394677 703075 394733
rect 703161 394677 703217 394733
rect 703303 394677 703359 394733
rect 703445 394677 703501 394733
rect 703587 394677 703643 394733
rect 703729 394677 703785 394733
rect 703871 394677 703927 394733
rect 704013 394677 704069 394733
rect 704155 394677 704211 394733
rect 704297 394677 704353 394733
rect 702451 394535 702507 394591
rect 702593 394535 702649 394591
rect 702735 394535 702791 394591
rect 702877 394535 702933 394591
rect 703019 394535 703075 394591
rect 703161 394535 703217 394591
rect 703303 394535 703359 394591
rect 703445 394535 703501 394591
rect 703587 394535 703643 394591
rect 703729 394535 703785 394591
rect 703871 394535 703927 394591
rect 704013 394535 704069 394591
rect 704155 394535 704211 394591
rect 704297 394535 704353 394591
rect 702451 394393 702507 394449
rect 702593 394393 702649 394449
rect 702735 394393 702791 394449
rect 702877 394393 702933 394449
rect 703019 394393 703075 394449
rect 703161 394393 703217 394449
rect 703303 394393 703359 394449
rect 703445 394393 703501 394449
rect 703587 394393 703643 394449
rect 703729 394393 703785 394449
rect 703871 394393 703927 394449
rect 704013 394393 704069 394449
rect 704155 394393 704211 394449
rect 704297 394393 704353 394449
rect 702451 394251 702507 394307
rect 702593 394251 702649 394307
rect 702735 394251 702791 394307
rect 702877 394251 702933 394307
rect 703019 394251 703075 394307
rect 703161 394251 703217 394307
rect 703303 394251 703359 394307
rect 703445 394251 703501 394307
rect 703587 394251 703643 394307
rect 703729 394251 703785 394307
rect 703871 394251 703927 394307
rect 704013 394251 704069 394307
rect 704155 394251 704211 394307
rect 704297 394251 704353 394307
rect 702451 394109 702507 394165
rect 702593 394109 702649 394165
rect 702735 394109 702791 394165
rect 702877 394109 702933 394165
rect 703019 394109 703075 394165
rect 703161 394109 703217 394165
rect 703303 394109 703359 394165
rect 703445 394109 703501 394165
rect 703587 394109 703643 394165
rect 703729 394109 703785 394165
rect 703871 394109 703927 394165
rect 704013 394109 704069 394165
rect 704155 394109 704211 394165
rect 704297 394109 704353 394165
rect 702451 393967 702507 394023
rect 702593 393967 702649 394023
rect 702735 393967 702791 394023
rect 702877 393967 702933 394023
rect 703019 393967 703075 394023
rect 703161 393967 703217 394023
rect 703303 393967 703359 394023
rect 703445 393967 703501 394023
rect 703587 393967 703643 394023
rect 703729 393967 703785 394023
rect 703871 393967 703927 394023
rect 704013 393967 704069 394023
rect 704155 393967 704211 394023
rect 704297 393967 704353 394023
rect 702451 393825 702507 393881
rect 702593 393825 702649 393881
rect 702735 393825 702791 393881
rect 702877 393825 702933 393881
rect 703019 393825 703075 393881
rect 703161 393825 703217 393881
rect 703303 393825 703359 393881
rect 703445 393825 703501 393881
rect 703587 393825 703643 393881
rect 703729 393825 703785 393881
rect 703871 393825 703927 393881
rect 704013 393825 704069 393881
rect 704155 393825 704211 393881
rect 704297 393825 704353 393881
rect 702451 393683 702507 393739
rect 702593 393683 702649 393739
rect 702735 393683 702791 393739
rect 702877 393683 702933 393739
rect 703019 393683 703075 393739
rect 703161 393683 703217 393739
rect 703303 393683 703359 393739
rect 703445 393683 703501 393739
rect 703587 393683 703643 393739
rect 703729 393683 703785 393739
rect 703871 393683 703927 393739
rect 704013 393683 704069 393739
rect 704155 393683 704211 393739
rect 704297 393683 704353 393739
rect 702451 393541 702507 393597
rect 702593 393541 702649 393597
rect 702735 393541 702791 393597
rect 702877 393541 702933 393597
rect 703019 393541 703075 393597
rect 703161 393541 703217 393597
rect 703303 393541 703359 393597
rect 703445 393541 703501 393597
rect 703587 393541 703643 393597
rect 703729 393541 703785 393597
rect 703871 393541 703927 393597
rect 704013 393541 704069 393597
rect 704155 393541 704211 393597
rect 704297 393541 704353 393597
rect 702451 393399 702507 393455
rect 702593 393399 702649 393455
rect 702735 393399 702791 393455
rect 702877 393399 702933 393455
rect 703019 393399 703075 393455
rect 703161 393399 703217 393455
rect 703303 393399 703359 393455
rect 703445 393399 703501 393455
rect 703587 393399 703643 393455
rect 703729 393399 703785 393455
rect 703871 393399 703927 393455
rect 704013 393399 704069 393455
rect 704155 393399 704211 393455
rect 704297 393399 704353 393455
rect 702451 393257 702507 393313
rect 702593 393257 702649 393313
rect 702735 393257 702791 393313
rect 702877 393257 702933 393313
rect 703019 393257 703075 393313
rect 703161 393257 703217 393313
rect 703303 393257 703359 393313
rect 703445 393257 703501 393313
rect 703587 393257 703643 393313
rect 703729 393257 703785 393313
rect 703871 393257 703927 393313
rect 704013 393257 704069 393313
rect 704155 393257 704211 393313
rect 704297 393257 704353 393313
rect 702451 393115 702507 393171
rect 702593 393115 702649 393171
rect 702735 393115 702791 393171
rect 702877 393115 702933 393171
rect 703019 393115 703075 393171
rect 703161 393115 703217 393171
rect 703303 393115 703359 393171
rect 703445 393115 703501 393171
rect 703587 393115 703643 393171
rect 703729 393115 703785 393171
rect 703871 393115 703927 393171
rect 704013 393115 704069 393171
rect 704155 393115 704211 393171
rect 704297 393115 704353 393171
rect 702451 392973 702507 393029
rect 702593 392973 702649 393029
rect 702735 392973 702791 393029
rect 702877 392973 702933 393029
rect 703019 392973 703075 393029
rect 703161 392973 703217 393029
rect 703303 392973 703359 393029
rect 703445 392973 703501 393029
rect 703587 392973 703643 393029
rect 703729 392973 703785 393029
rect 703871 392973 703927 393029
rect 704013 392973 704069 393029
rect 704155 392973 704211 393029
rect 704297 392973 704353 393029
rect 702451 392831 702507 392887
rect 702593 392831 702649 392887
rect 702735 392831 702791 392887
rect 702877 392831 702933 392887
rect 703019 392831 703075 392887
rect 703161 392831 703217 392887
rect 703303 392831 703359 392887
rect 703445 392831 703501 392887
rect 703587 392831 703643 392887
rect 703729 392831 703785 392887
rect 703871 392831 703927 392887
rect 704013 392831 704069 392887
rect 704155 392831 704211 392887
rect 704297 392831 704353 392887
rect 702440 392054 702496 392110
rect 702582 392054 702638 392110
rect 702724 392054 702780 392110
rect 702866 392054 702922 392110
rect 703008 392054 703064 392110
rect 703150 392054 703206 392110
rect 703292 392054 703348 392110
rect 703434 392054 703490 392110
rect 703576 392054 703632 392110
rect 703718 392054 703774 392110
rect 703860 392054 703916 392110
rect 704002 392054 704058 392110
rect 704144 392054 704200 392110
rect 704286 392054 704342 392110
rect 702440 391912 702496 391968
rect 702582 391912 702638 391968
rect 702724 391912 702780 391968
rect 702866 391912 702922 391968
rect 703008 391912 703064 391968
rect 703150 391912 703206 391968
rect 703292 391912 703348 391968
rect 703434 391912 703490 391968
rect 703576 391912 703632 391968
rect 703718 391912 703774 391968
rect 703860 391912 703916 391968
rect 704002 391912 704058 391968
rect 704144 391912 704200 391968
rect 704286 391912 704342 391968
rect 702440 391770 702496 391826
rect 702582 391770 702638 391826
rect 702724 391770 702780 391826
rect 702866 391770 702922 391826
rect 703008 391770 703064 391826
rect 703150 391770 703206 391826
rect 703292 391770 703348 391826
rect 703434 391770 703490 391826
rect 703576 391770 703632 391826
rect 703718 391770 703774 391826
rect 703860 391770 703916 391826
rect 704002 391770 704058 391826
rect 704144 391770 704200 391826
rect 704286 391770 704342 391826
rect 702440 391628 702496 391684
rect 702582 391628 702638 391684
rect 702724 391628 702780 391684
rect 702866 391628 702922 391684
rect 703008 391628 703064 391684
rect 703150 391628 703206 391684
rect 703292 391628 703348 391684
rect 703434 391628 703490 391684
rect 703576 391628 703632 391684
rect 703718 391628 703774 391684
rect 703860 391628 703916 391684
rect 704002 391628 704058 391684
rect 704144 391628 704200 391684
rect 704286 391628 704342 391684
rect 702440 391486 702496 391542
rect 702582 391486 702638 391542
rect 702724 391486 702780 391542
rect 702866 391486 702922 391542
rect 703008 391486 703064 391542
rect 703150 391486 703206 391542
rect 703292 391486 703348 391542
rect 703434 391486 703490 391542
rect 703576 391486 703632 391542
rect 703718 391486 703774 391542
rect 703860 391486 703916 391542
rect 704002 391486 704058 391542
rect 704144 391486 704200 391542
rect 704286 391486 704342 391542
rect 702440 391344 702496 391400
rect 702582 391344 702638 391400
rect 702724 391344 702780 391400
rect 702866 391344 702922 391400
rect 703008 391344 703064 391400
rect 703150 391344 703206 391400
rect 703292 391344 703348 391400
rect 703434 391344 703490 391400
rect 703576 391344 703632 391400
rect 703718 391344 703774 391400
rect 703860 391344 703916 391400
rect 704002 391344 704058 391400
rect 704144 391344 704200 391400
rect 704286 391344 704342 391400
rect 702440 391202 702496 391258
rect 702582 391202 702638 391258
rect 702724 391202 702780 391258
rect 702866 391202 702922 391258
rect 703008 391202 703064 391258
rect 703150 391202 703206 391258
rect 703292 391202 703348 391258
rect 703434 391202 703490 391258
rect 703576 391202 703632 391258
rect 703718 391202 703774 391258
rect 703860 391202 703916 391258
rect 704002 391202 704058 391258
rect 704144 391202 704200 391258
rect 704286 391202 704342 391258
rect 702440 391060 702496 391116
rect 702582 391060 702638 391116
rect 702724 391060 702780 391116
rect 702866 391060 702922 391116
rect 703008 391060 703064 391116
rect 703150 391060 703206 391116
rect 703292 391060 703348 391116
rect 703434 391060 703490 391116
rect 703576 391060 703632 391116
rect 703718 391060 703774 391116
rect 703860 391060 703916 391116
rect 704002 391060 704058 391116
rect 704144 391060 704200 391116
rect 704286 391060 704342 391116
rect 702440 390918 702496 390974
rect 702582 390918 702638 390974
rect 702724 390918 702780 390974
rect 702866 390918 702922 390974
rect 703008 390918 703064 390974
rect 703150 390918 703206 390974
rect 703292 390918 703348 390974
rect 703434 390918 703490 390974
rect 703576 390918 703632 390974
rect 703718 390918 703774 390974
rect 703860 390918 703916 390974
rect 704002 390918 704058 390974
rect 704144 390918 704200 390974
rect 704286 390918 704342 390974
rect 702440 390776 702496 390832
rect 702582 390776 702638 390832
rect 702724 390776 702780 390832
rect 702866 390776 702922 390832
rect 703008 390776 703064 390832
rect 703150 390776 703206 390832
rect 703292 390776 703348 390832
rect 703434 390776 703490 390832
rect 703576 390776 703632 390832
rect 703718 390776 703774 390832
rect 703860 390776 703916 390832
rect 704002 390776 704058 390832
rect 704144 390776 704200 390832
rect 704286 390776 704342 390832
rect 702440 390634 702496 390690
rect 702582 390634 702638 390690
rect 702724 390634 702780 390690
rect 702866 390634 702922 390690
rect 703008 390634 703064 390690
rect 703150 390634 703206 390690
rect 703292 390634 703348 390690
rect 703434 390634 703490 390690
rect 703576 390634 703632 390690
rect 703718 390634 703774 390690
rect 703860 390634 703916 390690
rect 704002 390634 704058 390690
rect 704144 390634 704200 390690
rect 704286 390634 704342 390690
rect 702440 390492 702496 390548
rect 702582 390492 702638 390548
rect 702724 390492 702780 390548
rect 702866 390492 702922 390548
rect 703008 390492 703064 390548
rect 703150 390492 703206 390548
rect 703292 390492 703348 390548
rect 703434 390492 703490 390548
rect 703576 390492 703632 390548
rect 703718 390492 703774 390548
rect 703860 390492 703916 390548
rect 704002 390492 704058 390548
rect 704144 390492 704200 390548
rect 704286 390492 704342 390548
rect 702440 390350 702496 390406
rect 702582 390350 702638 390406
rect 702724 390350 702780 390406
rect 702866 390350 702922 390406
rect 703008 390350 703064 390406
rect 703150 390350 703206 390406
rect 703292 390350 703348 390406
rect 703434 390350 703490 390406
rect 703576 390350 703632 390406
rect 703718 390350 703774 390406
rect 703860 390350 703916 390406
rect 704002 390350 704058 390406
rect 704144 390350 704200 390406
rect 704286 390350 704342 390406
rect 73866 140594 73922 140650
rect 74008 140594 74064 140650
rect 74150 140594 74206 140650
rect 74292 140594 74348 140650
rect 74434 140594 74490 140650
rect 74576 140594 74632 140650
rect 74718 140594 74774 140650
rect 74860 140594 74916 140650
rect 75002 140594 75058 140650
rect 75144 140594 75200 140650
rect 75286 140594 75342 140650
rect 73866 140452 73922 140508
rect 74008 140452 74064 140508
rect 74150 140452 74206 140508
rect 74292 140452 74348 140508
rect 74434 140452 74490 140508
rect 74576 140452 74632 140508
rect 74718 140452 74774 140508
rect 74860 140452 74916 140508
rect 75002 140452 75058 140508
rect 75144 140452 75200 140508
rect 75286 140452 75342 140508
rect 73866 140310 73922 140366
rect 74008 140310 74064 140366
rect 74150 140310 74206 140366
rect 74292 140310 74348 140366
rect 74434 140310 74490 140366
rect 74576 140310 74632 140366
rect 74718 140310 74774 140366
rect 74860 140310 74916 140366
rect 75002 140310 75058 140366
rect 75144 140310 75200 140366
rect 75286 140310 75342 140366
rect 73866 140168 73922 140224
rect 74008 140168 74064 140224
rect 74150 140168 74206 140224
rect 74292 140168 74348 140224
rect 74434 140168 74490 140224
rect 74576 140168 74632 140224
rect 74718 140168 74774 140224
rect 74860 140168 74916 140224
rect 75002 140168 75058 140224
rect 75144 140168 75200 140224
rect 75286 140168 75342 140224
rect 73866 140026 73922 140082
rect 74008 140026 74064 140082
rect 74150 140026 74206 140082
rect 74292 140026 74348 140082
rect 74434 140026 74490 140082
rect 74576 140026 74632 140082
rect 74718 140026 74774 140082
rect 74860 140026 74916 140082
rect 75002 140026 75058 140082
rect 75144 140026 75200 140082
rect 75286 140026 75342 140082
rect 73866 139884 73922 139940
rect 74008 139884 74064 139940
rect 74150 139884 74206 139940
rect 74292 139884 74348 139940
rect 74434 139884 74490 139940
rect 74576 139884 74632 139940
rect 74718 139884 74774 139940
rect 74860 139884 74916 139940
rect 75002 139884 75058 139940
rect 75144 139884 75200 139940
rect 75286 139884 75342 139940
rect 73866 139742 73922 139798
rect 74008 139742 74064 139798
rect 74150 139742 74206 139798
rect 74292 139742 74348 139798
rect 74434 139742 74490 139798
rect 74576 139742 74632 139798
rect 74718 139742 74774 139798
rect 74860 139742 74916 139798
rect 75002 139742 75058 139798
rect 75144 139742 75200 139798
rect 75286 139742 75342 139798
rect 73866 139600 73922 139656
rect 74008 139600 74064 139656
rect 74150 139600 74206 139656
rect 74292 139600 74348 139656
rect 74434 139600 74490 139656
rect 74576 139600 74632 139656
rect 74718 139600 74774 139656
rect 74860 139600 74916 139656
rect 75002 139600 75058 139656
rect 75144 139600 75200 139656
rect 75286 139600 75342 139656
rect 73866 139458 73922 139514
rect 74008 139458 74064 139514
rect 74150 139458 74206 139514
rect 74292 139458 74348 139514
rect 74434 139458 74490 139514
rect 74576 139458 74632 139514
rect 74718 139458 74774 139514
rect 74860 139458 74916 139514
rect 75002 139458 75058 139514
rect 75144 139458 75200 139514
rect 75286 139458 75342 139514
rect 73866 139316 73922 139372
rect 74008 139316 74064 139372
rect 74150 139316 74206 139372
rect 74292 139316 74348 139372
rect 74434 139316 74490 139372
rect 74576 139316 74632 139372
rect 74718 139316 74774 139372
rect 74860 139316 74916 139372
rect 75002 139316 75058 139372
rect 75144 139316 75200 139372
rect 75286 139316 75342 139372
rect 73866 139174 73922 139230
rect 74008 139174 74064 139230
rect 74150 139174 74206 139230
rect 74292 139174 74348 139230
rect 74434 139174 74490 139230
rect 74576 139174 74632 139230
rect 74718 139174 74774 139230
rect 74860 139174 74916 139230
rect 75002 139174 75058 139230
rect 75144 139174 75200 139230
rect 75286 139174 75342 139230
rect 73866 139032 73922 139088
rect 74008 139032 74064 139088
rect 74150 139032 74206 139088
rect 74292 139032 74348 139088
rect 74434 139032 74490 139088
rect 74576 139032 74632 139088
rect 74718 139032 74774 139088
rect 74860 139032 74916 139088
rect 75002 139032 75058 139088
rect 75144 139032 75200 139088
rect 75286 139032 75342 139088
rect 73866 138890 73922 138946
rect 74008 138890 74064 138946
rect 74150 138890 74206 138946
rect 74292 138890 74348 138946
rect 74434 138890 74490 138946
rect 74576 138890 74632 138946
rect 74718 138890 74774 138946
rect 74860 138890 74916 138946
rect 75002 138890 75058 138946
rect 75144 138890 75200 138946
rect 75286 138890 75342 138946
rect 73855 138113 73911 138169
rect 73997 138113 74053 138169
rect 74139 138113 74195 138169
rect 74281 138113 74337 138169
rect 74423 138113 74479 138169
rect 74565 138113 74621 138169
rect 74707 138113 74763 138169
rect 74849 138113 74905 138169
rect 74991 138113 75047 138169
rect 75133 138113 75189 138169
rect 75275 138113 75331 138169
rect 73855 137971 73911 138027
rect 73997 137971 74053 138027
rect 74139 137971 74195 138027
rect 74281 137971 74337 138027
rect 74423 137971 74479 138027
rect 74565 137971 74621 138027
rect 74707 137971 74763 138027
rect 74849 137971 74905 138027
rect 74991 137971 75047 138027
rect 75133 137971 75189 138027
rect 75275 137971 75331 138027
rect 73855 137829 73911 137885
rect 73997 137829 74053 137885
rect 74139 137829 74195 137885
rect 74281 137829 74337 137885
rect 74423 137829 74479 137885
rect 74565 137829 74621 137885
rect 74707 137829 74763 137885
rect 74849 137829 74905 137885
rect 74991 137829 75047 137885
rect 75133 137829 75189 137885
rect 75275 137829 75331 137885
rect 73855 137687 73911 137743
rect 73997 137687 74053 137743
rect 74139 137687 74195 137743
rect 74281 137687 74337 137743
rect 74423 137687 74479 137743
rect 74565 137687 74621 137743
rect 74707 137687 74763 137743
rect 74849 137687 74905 137743
rect 74991 137687 75047 137743
rect 75133 137687 75189 137743
rect 75275 137687 75331 137743
rect 73855 137545 73911 137601
rect 73997 137545 74053 137601
rect 74139 137545 74195 137601
rect 74281 137545 74337 137601
rect 74423 137545 74479 137601
rect 74565 137545 74621 137601
rect 74707 137545 74763 137601
rect 74849 137545 74905 137601
rect 74991 137545 75047 137601
rect 75133 137545 75189 137601
rect 75275 137545 75331 137601
rect 73855 137403 73911 137459
rect 73997 137403 74053 137459
rect 74139 137403 74195 137459
rect 74281 137403 74337 137459
rect 74423 137403 74479 137459
rect 74565 137403 74621 137459
rect 74707 137403 74763 137459
rect 74849 137403 74905 137459
rect 74991 137403 75047 137459
rect 75133 137403 75189 137459
rect 75275 137403 75331 137459
rect 73855 137261 73911 137317
rect 73997 137261 74053 137317
rect 74139 137261 74195 137317
rect 74281 137261 74337 137317
rect 74423 137261 74479 137317
rect 74565 137261 74621 137317
rect 74707 137261 74763 137317
rect 74849 137261 74905 137317
rect 74991 137261 75047 137317
rect 75133 137261 75189 137317
rect 75275 137261 75331 137317
rect 73855 137119 73911 137175
rect 73997 137119 74053 137175
rect 74139 137119 74195 137175
rect 74281 137119 74337 137175
rect 74423 137119 74479 137175
rect 74565 137119 74621 137175
rect 74707 137119 74763 137175
rect 74849 137119 74905 137175
rect 74991 137119 75047 137175
rect 75133 137119 75189 137175
rect 75275 137119 75331 137175
rect 73855 136977 73911 137033
rect 73997 136977 74053 137033
rect 74139 136977 74195 137033
rect 74281 136977 74337 137033
rect 74423 136977 74479 137033
rect 74565 136977 74621 137033
rect 74707 136977 74763 137033
rect 74849 136977 74905 137033
rect 74991 136977 75047 137033
rect 75133 136977 75189 137033
rect 75275 136977 75331 137033
rect 73855 136835 73911 136891
rect 73997 136835 74053 136891
rect 74139 136835 74195 136891
rect 74281 136835 74337 136891
rect 74423 136835 74479 136891
rect 74565 136835 74621 136891
rect 74707 136835 74763 136891
rect 74849 136835 74905 136891
rect 74991 136835 75047 136891
rect 75133 136835 75189 136891
rect 75275 136835 75331 136891
rect 73855 136693 73911 136749
rect 73997 136693 74053 136749
rect 74139 136693 74195 136749
rect 74281 136693 74337 136749
rect 74423 136693 74479 136749
rect 74565 136693 74621 136749
rect 74707 136693 74763 136749
rect 74849 136693 74905 136749
rect 74991 136693 75047 136749
rect 75133 136693 75189 136749
rect 75275 136693 75331 136749
rect 73855 136551 73911 136607
rect 73997 136551 74053 136607
rect 74139 136551 74195 136607
rect 74281 136551 74337 136607
rect 74423 136551 74479 136607
rect 74565 136551 74621 136607
rect 74707 136551 74763 136607
rect 74849 136551 74905 136607
rect 74991 136551 75047 136607
rect 75133 136551 75189 136607
rect 75275 136551 75331 136607
rect 73855 136409 73911 136465
rect 73997 136409 74053 136465
rect 74139 136409 74195 136465
rect 74281 136409 74337 136465
rect 74423 136409 74479 136465
rect 74565 136409 74621 136465
rect 74707 136409 74763 136465
rect 74849 136409 74905 136465
rect 74991 136409 75047 136465
rect 75133 136409 75189 136465
rect 75275 136409 75331 136465
rect 73855 136267 73911 136323
rect 73997 136267 74053 136323
rect 74139 136267 74195 136323
rect 74281 136267 74337 136323
rect 74423 136267 74479 136323
rect 74565 136267 74621 136323
rect 74707 136267 74763 136323
rect 74849 136267 74905 136323
rect 74991 136267 75047 136323
rect 75133 136267 75189 136323
rect 75275 136267 75331 136323
rect 73855 135743 73911 135799
rect 73997 135743 74053 135799
rect 74139 135743 74195 135799
rect 74281 135743 74337 135799
rect 74423 135743 74479 135799
rect 74565 135743 74621 135799
rect 74707 135743 74763 135799
rect 74849 135743 74905 135799
rect 74991 135743 75047 135799
rect 75133 135743 75189 135799
rect 75275 135743 75331 135799
rect 73855 135601 73911 135657
rect 73997 135601 74053 135657
rect 74139 135601 74195 135657
rect 74281 135601 74337 135657
rect 74423 135601 74479 135657
rect 74565 135601 74621 135657
rect 74707 135601 74763 135657
rect 74849 135601 74905 135657
rect 74991 135601 75047 135657
rect 75133 135601 75189 135657
rect 75275 135601 75331 135657
rect 73855 135459 73911 135515
rect 73997 135459 74053 135515
rect 74139 135459 74195 135515
rect 74281 135459 74337 135515
rect 74423 135459 74479 135515
rect 74565 135459 74621 135515
rect 74707 135459 74763 135515
rect 74849 135459 74905 135515
rect 74991 135459 75047 135515
rect 75133 135459 75189 135515
rect 75275 135459 75331 135515
rect 73855 135317 73911 135373
rect 73997 135317 74053 135373
rect 74139 135317 74195 135373
rect 74281 135317 74337 135373
rect 74423 135317 74479 135373
rect 74565 135317 74621 135373
rect 74707 135317 74763 135373
rect 74849 135317 74905 135373
rect 74991 135317 75047 135373
rect 75133 135317 75189 135373
rect 75275 135317 75331 135373
rect 73855 135175 73911 135231
rect 73997 135175 74053 135231
rect 74139 135175 74195 135231
rect 74281 135175 74337 135231
rect 74423 135175 74479 135231
rect 74565 135175 74621 135231
rect 74707 135175 74763 135231
rect 74849 135175 74905 135231
rect 74991 135175 75047 135231
rect 75133 135175 75189 135231
rect 75275 135175 75331 135231
rect 73855 135033 73911 135089
rect 73997 135033 74053 135089
rect 74139 135033 74195 135089
rect 74281 135033 74337 135089
rect 74423 135033 74479 135089
rect 74565 135033 74621 135089
rect 74707 135033 74763 135089
rect 74849 135033 74905 135089
rect 74991 135033 75047 135089
rect 75133 135033 75189 135089
rect 75275 135033 75331 135089
rect 73855 134891 73911 134947
rect 73997 134891 74053 134947
rect 74139 134891 74195 134947
rect 74281 134891 74337 134947
rect 74423 134891 74479 134947
rect 74565 134891 74621 134947
rect 74707 134891 74763 134947
rect 74849 134891 74905 134947
rect 74991 134891 75047 134947
rect 75133 134891 75189 134947
rect 75275 134891 75331 134947
rect 73855 134749 73911 134805
rect 73997 134749 74053 134805
rect 74139 134749 74195 134805
rect 74281 134749 74337 134805
rect 74423 134749 74479 134805
rect 74565 134749 74621 134805
rect 74707 134749 74763 134805
rect 74849 134749 74905 134805
rect 74991 134749 75047 134805
rect 75133 134749 75189 134805
rect 75275 134749 75331 134805
rect 73855 134607 73911 134663
rect 73997 134607 74053 134663
rect 74139 134607 74195 134663
rect 74281 134607 74337 134663
rect 74423 134607 74479 134663
rect 74565 134607 74621 134663
rect 74707 134607 74763 134663
rect 74849 134607 74905 134663
rect 74991 134607 75047 134663
rect 75133 134607 75189 134663
rect 75275 134607 75331 134663
rect 73855 134465 73911 134521
rect 73997 134465 74053 134521
rect 74139 134465 74195 134521
rect 74281 134465 74337 134521
rect 74423 134465 74479 134521
rect 74565 134465 74621 134521
rect 74707 134465 74763 134521
rect 74849 134465 74905 134521
rect 74991 134465 75047 134521
rect 75133 134465 75189 134521
rect 75275 134465 75331 134521
rect 73855 134323 73911 134379
rect 73997 134323 74053 134379
rect 74139 134323 74195 134379
rect 74281 134323 74337 134379
rect 74423 134323 74479 134379
rect 74565 134323 74621 134379
rect 74707 134323 74763 134379
rect 74849 134323 74905 134379
rect 74991 134323 75047 134379
rect 75133 134323 75189 134379
rect 75275 134323 75331 134379
rect 73855 134181 73911 134237
rect 73997 134181 74053 134237
rect 74139 134181 74195 134237
rect 74281 134181 74337 134237
rect 74423 134181 74479 134237
rect 74565 134181 74621 134237
rect 74707 134181 74763 134237
rect 74849 134181 74905 134237
rect 74991 134181 75047 134237
rect 75133 134181 75189 134237
rect 75275 134181 75331 134237
rect 73855 134039 73911 134095
rect 73997 134039 74053 134095
rect 74139 134039 74195 134095
rect 74281 134039 74337 134095
rect 74423 134039 74479 134095
rect 74565 134039 74621 134095
rect 74707 134039 74763 134095
rect 74849 134039 74905 134095
rect 74991 134039 75047 134095
rect 75133 134039 75189 134095
rect 75275 134039 75331 134095
rect 73855 133897 73911 133953
rect 73997 133897 74053 133953
rect 74139 133897 74195 133953
rect 74281 133897 74337 133953
rect 74423 133897 74479 133953
rect 74565 133897 74621 133953
rect 74707 133897 74763 133953
rect 74849 133897 74905 133953
rect 74991 133897 75047 133953
rect 75133 133897 75189 133953
rect 75275 133897 75331 133953
rect 73855 133037 73911 133093
rect 73997 133037 74053 133093
rect 74139 133037 74195 133093
rect 74281 133037 74337 133093
rect 74423 133037 74479 133093
rect 74565 133037 74621 133093
rect 74707 133037 74763 133093
rect 74849 133037 74905 133093
rect 74991 133037 75047 133093
rect 75133 133037 75189 133093
rect 75275 133037 75331 133093
rect 73855 132895 73911 132951
rect 73997 132895 74053 132951
rect 74139 132895 74195 132951
rect 74281 132895 74337 132951
rect 74423 132895 74479 132951
rect 74565 132895 74621 132951
rect 74707 132895 74763 132951
rect 74849 132895 74905 132951
rect 74991 132895 75047 132951
rect 75133 132895 75189 132951
rect 75275 132895 75331 132951
rect 73855 132753 73911 132809
rect 73997 132753 74053 132809
rect 74139 132753 74195 132809
rect 74281 132753 74337 132809
rect 74423 132753 74479 132809
rect 74565 132753 74621 132809
rect 74707 132753 74763 132809
rect 74849 132753 74905 132809
rect 74991 132753 75047 132809
rect 75133 132753 75189 132809
rect 75275 132753 75331 132809
rect 73855 132611 73911 132667
rect 73997 132611 74053 132667
rect 74139 132611 74195 132667
rect 74281 132611 74337 132667
rect 74423 132611 74479 132667
rect 74565 132611 74621 132667
rect 74707 132611 74763 132667
rect 74849 132611 74905 132667
rect 74991 132611 75047 132667
rect 75133 132611 75189 132667
rect 75275 132611 75331 132667
rect 73855 132469 73911 132525
rect 73997 132469 74053 132525
rect 74139 132469 74195 132525
rect 74281 132469 74337 132525
rect 74423 132469 74479 132525
rect 74565 132469 74621 132525
rect 74707 132469 74763 132525
rect 74849 132469 74905 132525
rect 74991 132469 75047 132525
rect 75133 132469 75189 132525
rect 75275 132469 75331 132525
rect 73855 132327 73911 132383
rect 73997 132327 74053 132383
rect 74139 132327 74195 132383
rect 74281 132327 74337 132383
rect 74423 132327 74479 132383
rect 74565 132327 74621 132383
rect 74707 132327 74763 132383
rect 74849 132327 74905 132383
rect 74991 132327 75047 132383
rect 75133 132327 75189 132383
rect 75275 132327 75331 132383
rect 73855 132185 73911 132241
rect 73997 132185 74053 132241
rect 74139 132185 74195 132241
rect 74281 132185 74337 132241
rect 74423 132185 74479 132241
rect 74565 132185 74621 132241
rect 74707 132185 74763 132241
rect 74849 132185 74905 132241
rect 74991 132185 75047 132241
rect 75133 132185 75189 132241
rect 75275 132185 75331 132241
rect 73855 132043 73911 132099
rect 73997 132043 74053 132099
rect 74139 132043 74195 132099
rect 74281 132043 74337 132099
rect 74423 132043 74479 132099
rect 74565 132043 74621 132099
rect 74707 132043 74763 132099
rect 74849 132043 74905 132099
rect 74991 132043 75047 132099
rect 75133 132043 75189 132099
rect 75275 132043 75331 132099
rect 73855 131901 73911 131957
rect 73997 131901 74053 131957
rect 74139 131901 74195 131957
rect 74281 131901 74337 131957
rect 74423 131901 74479 131957
rect 74565 131901 74621 131957
rect 74707 131901 74763 131957
rect 74849 131901 74905 131957
rect 74991 131901 75047 131957
rect 75133 131901 75189 131957
rect 75275 131901 75331 131957
rect 73855 131759 73911 131815
rect 73997 131759 74053 131815
rect 74139 131759 74195 131815
rect 74281 131759 74337 131815
rect 74423 131759 74479 131815
rect 74565 131759 74621 131815
rect 74707 131759 74763 131815
rect 74849 131759 74905 131815
rect 74991 131759 75047 131815
rect 75133 131759 75189 131815
rect 75275 131759 75331 131815
rect 73855 131617 73911 131673
rect 73997 131617 74053 131673
rect 74139 131617 74195 131673
rect 74281 131617 74337 131673
rect 74423 131617 74479 131673
rect 74565 131617 74621 131673
rect 74707 131617 74763 131673
rect 74849 131617 74905 131673
rect 74991 131617 75047 131673
rect 75133 131617 75189 131673
rect 75275 131617 75331 131673
rect 73855 131475 73911 131531
rect 73997 131475 74053 131531
rect 74139 131475 74195 131531
rect 74281 131475 74337 131531
rect 74423 131475 74479 131531
rect 74565 131475 74621 131531
rect 74707 131475 74763 131531
rect 74849 131475 74905 131531
rect 74991 131475 75047 131531
rect 75133 131475 75189 131531
rect 75275 131475 75331 131531
rect 73855 131333 73911 131389
rect 73997 131333 74053 131389
rect 74139 131333 74195 131389
rect 74281 131333 74337 131389
rect 74423 131333 74479 131389
rect 74565 131333 74621 131389
rect 74707 131333 74763 131389
rect 74849 131333 74905 131389
rect 74991 131333 75047 131389
rect 75133 131333 75189 131389
rect 75275 131333 75331 131389
rect 73855 131191 73911 131247
rect 73997 131191 74053 131247
rect 74139 131191 74195 131247
rect 74281 131191 74337 131247
rect 74423 131191 74479 131247
rect 74565 131191 74621 131247
rect 74707 131191 74763 131247
rect 74849 131191 74905 131247
rect 74991 131191 75047 131247
rect 75133 131191 75189 131247
rect 75275 131191 75331 131247
rect 73855 130667 73911 130723
rect 73997 130667 74053 130723
rect 74139 130667 74195 130723
rect 74281 130667 74337 130723
rect 74423 130667 74479 130723
rect 74565 130667 74621 130723
rect 74707 130667 74763 130723
rect 74849 130667 74905 130723
rect 74991 130667 75047 130723
rect 75133 130667 75189 130723
rect 75275 130667 75331 130723
rect 73855 130525 73911 130581
rect 73997 130525 74053 130581
rect 74139 130525 74195 130581
rect 74281 130525 74337 130581
rect 74423 130525 74479 130581
rect 74565 130525 74621 130581
rect 74707 130525 74763 130581
rect 74849 130525 74905 130581
rect 74991 130525 75047 130581
rect 75133 130525 75189 130581
rect 75275 130525 75331 130581
rect 73855 130383 73911 130439
rect 73997 130383 74053 130439
rect 74139 130383 74195 130439
rect 74281 130383 74337 130439
rect 74423 130383 74479 130439
rect 74565 130383 74621 130439
rect 74707 130383 74763 130439
rect 74849 130383 74905 130439
rect 74991 130383 75047 130439
rect 75133 130383 75189 130439
rect 75275 130383 75331 130439
rect 73855 130241 73911 130297
rect 73997 130241 74053 130297
rect 74139 130241 74195 130297
rect 74281 130241 74337 130297
rect 74423 130241 74479 130297
rect 74565 130241 74621 130297
rect 74707 130241 74763 130297
rect 74849 130241 74905 130297
rect 74991 130241 75047 130297
rect 75133 130241 75189 130297
rect 75275 130241 75331 130297
rect 73855 130099 73911 130155
rect 73997 130099 74053 130155
rect 74139 130099 74195 130155
rect 74281 130099 74337 130155
rect 74423 130099 74479 130155
rect 74565 130099 74621 130155
rect 74707 130099 74763 130155
rect 74849 130099 74905 130155
rect 74991 130099 75047 130155
rect 75133 130099 75189 130155
rect 75275 130099 75331 130155
rect 73855 129957 73911 130013
rect 73997 129957 74053 130013
rect 74139 129957 74195 130013
rect 74281 129957 74337 130013
rect 74423 129957 74479 130013
rect 74565 129957 74621 130013
rect 74707 129957 74763 130013
rect 74849 129957 74905 130013
rect 74991 129957 75047 130013
rect 75133 129957 75189 130013
rect 75275 129957 75331 130013
rect 73855 129815 73911 129871
rect 73997 129815 74053 129871
rect 74139 129815 74195 129871
rect 74281 129815 74337 129871
rect 74423 129815 74479 129871
rect 74565 129815 74621 129871
rect 74707 129815 74763 129871
rect 74849 129815 74905 129871
rect 74991 129815 75047 129871
rect 75133 129815 75189 129871
rect 75275 129815 75331 129871
rect 73855 129673 73911 129729
rect 73997 129673 74053 129729
rect 74139 129673 74195 129729
rect 74281 129673 74337 129729
rect 74423 129673 74479 129729
rect 74565 129673 74621 129729
rect 74707 129673 74763 129729
rect 74849 129673 74905 129729
rect 74991 129673 75047 129729
rect 75133 129673 75189 129729
rect 75275 129673 75331 129729
rect 73855 129531 73911 129587
rect 73997 129531 74053 129587
rect 74139 129531 74195 129587
rect 74281 129531 74337 129587
rect 74423 129531 74479 129587
rect 74565 129531 74621 129587
rect 74707 129531 74763 129587
rect 74849 129531 74905 129587
rect 74991 129531 75047 129587
rect 75133 129531 75189 129587
rect 75275 129531 75331 129587
rect 73855 129389 73911 129445
rect 73997 129389 74053 129445
rect 74139 129389 74195 129445
rect 74281 129389 74337 129445
rect 74423 129389 74479 129445
rect 74565 129389 74621 129445
rect 74707 129389 74763 129445
rect 74849 129389 74905 129445
rect 74991 129389 75047 129445
rect 75133 129389 75189 129445
rect 75275 129389 75331 129445
rect 73855 129247 73911 129303
rect 73997 129247 74053 129303
rect 74139 129247 74195 129303
rect 74281 129247 74337 129303
rect 74423 129247 74479 129303
rect 74565 129247 74621 129303
rect 74707 129247 74763 129303
rect 74849 129247 74905 129303
rect 74991 129247 75047 129303
rect 75133 129247 75189 129303
rect 75275 129247 75331 129303
rect 73855 129105 73911 129161
rect 73997 129105 74053 129161
rect 74139 129105 74195 129161
rect 74281 129105 74337 129161
rect 74423 129105 74479 129161
rect 74565 129105 74621 129161
rect 74707 129105 74763 129161
rect 74849 129105 74905 129161
rect 74991 129105 75047 129161
rect 75133 129105 75189 129161
rect 75275 129105 75331 129161
rect 73855 128963 73911 129019
rect 73997 128963 74053 129019
rect 74139 128963 74195 129019
rect 74281 128963 74337 129019
rect 74423 128963 74479 129019
rect 74565 128963 74621 129019
rect 74707 128963 74763 129019
rect 74849 128963 74905 129019
rect 74991 128963 75047 129019
rect 75133 128963 75189 129019
rect 75275 128963 75331 129019
rect 73855 128821 73911 128877
rect 73997 128821 74053 128877
rect 74139 128821 74195 128877
rect 74281 128821 74337 128877
rect 74423 128821 74479 128877
rect 74565 128821 74621 128877
rect 74707 128821 74763 128877
rect 74849 128821 74905 128877
rect 74991 128821 75047 128877
rect 75133 128821 75189 128877
rect 75275 128821 75331 128877
rect 73866 128038 73922 128094
rect 74008 128038 74064 128094
rect 74150 128038 74206 128094
rect 74292 128038 74348 128094
rect 74434 128038 74490 128094
rect 74576 128038 74632 128094
rect 74718 128038 74774 128094
rect 74860 128038 74916 128094
rect 75002 128038 75058 128094
rect 75144 128038 75200 128094
rect 75286 128038 75342 128094
rect 73866 127896 73922 127952
rect 74008 127896 74064 127952
rect 74150 127896 74206 127952
rect 74292 127896 74348 127952
rect 74434 127896 74490 127952
rect 74576 127896 74632 127952
rect 74718 127896 74774 127952
rect 74860 127896 74916 127952
rect 75002 127896 75058 127952
rect 75144 127896 75200 127952
rect 75286 127896 75342 127952
rect 73866 127754 73922 127810
rect 74008 127754 74064 127810
rect 74150 127754 74206 127810
rect 74292 127754 74348 127810
rect 74434 127754 74490 127810
rect 74576 127754 74632 127810
rect 74718 127754 74774 127810
rect 74860 127754 74916 127810
rect 75002 127754 75058 127810
rect 75144 127754 75200 127810
rect 75286 127754 75342 127810
rect 73866 127612 73922 127668
rect 74008 127612 74064 127668
rect 74150 127612 74206 127668
rect 74292 127612 74348 127668
rect 74434 127612 74490 127668
rect 74576 127612 74632 127668
rect 74718 127612 74774 127668
rect 74860 127612 74916 127668
rect 75002 127612 75058 127668
rect 75144 127612 75200 127668
rect 75286 127612 75342 127668
rect 73866 127470 73922 127526
rect 74008 127470 74064 127526
rect 74150 127470 74206 127526
rect 74292 127470 74348 127526
rect 74434 127470 74490 127526
rect 74576 127470 74632 127526
rect 74718 127470 74774 127526
rect 74860 127470 74916 127526
rect 75002 127470 75058 127526
rect 75144 127470 75200 127526
rect 75286 127470 75342 127526
rect 73866 127328 73922 127384
rect 74008 127328 74064 127384
rect 74150 127328 74206 127384
rect 74292 127328 74348 127384
rect 74434 127328 74490 127384
rect 74576 127328 74632 127384
rect 74718 127328 74774 127384
rect 74860 127328 74916 127384
rect 75002 127328 75058 127384
rect 75144 127328 75200 127384
rect 75286 127328 75342 127384
rect 73866 127186 73922 127242
rect 74008 127186 74064 127242
rect 74150 127186 74206 127242
rect 74292 127186 74348 127242
rect 74434 127186 74490 127242
rect 74576 127186 74632 127242
rect 74718 127186 74774 127242
rect 74860 127186 74916 127242
rect 75002 127186 75058 127242
rect 75144 127186 75200 127242
rect 75286 127186 75342 127242
rect 73866 127044 73922 127100
rect 74008 127044 74064 127100
rect 74150 127044 74206 127100
rect 74292 127044 74348 127100
rect 74434 127044 74490 127100
rect 74576 127044 74632 127100
rect 74718 127044 74774 127100
rect 74860 127044 74916 127100
rect 75002 127044 75058 127100
rect 75144 127044 75200 127100
rect 75286 127044 75342 127100
rect 73866 126902 73922 126958
rect 74008 126902 74064 126958
rect 74150 126902 74206 126958
rect 74292 126902 74348 126958
rect 74434 126902 74490 126958
rect 74576 126902 74632 126958
rect 74718 126902 74774 126958
rect 74860 126902 74916 126958
rect 75002 126902 75058 126958
rect 75144 126902 75200 126958
rect 75286 126902 75342 126958
rect 73866 126760 73922 126816
rect 74008 126760 74064 126816
rect 74150 126760 74206 126816
rect 74292 126760 74348 126816
rect 74434 126760 74490 126816
rect 74576 126760 74632 126816
rect 74718 126760 74774 126816
rect 74860 126760 74916 126816
rect 75002 126760 75058 126816
rect 75144 126760 75200 126816
rect 75286 126760 75342 126816
rect 73866 126618 73922 126674
rect 74008 126618 74064 126674
rect 74150 126618 74206 126674
rect 74292 126618 74348 126674
rect 74434 126618 74490 126674
rect 74576 126618 74632 126674
rect 74718 126618 74774 126674
rect 74860 126618 74916 126674
rect 75002 126618 75058 126674
rect 75144 126618 75200 126674
rect 75286 126618 75342 126674
rect 73866 126476 73922 126532
rect 74008 126476 74064 126532
rect 74150 126476 74206 126532
rect 74292 126476 74348 126532
rect 74434 126476 74490 126532
rect 74576 126476 74632 126532
rect 74718 126476 74774 126532
rect 74860 126476 74916 126532
rect 75002 126476 75058 126532
rect 75144 126476 75200 126532
rect 75286 126476 75342 126532
rect 73866 126334 73922 126390
rect 74008 126334 74064 126390
rect 74150 126334 74206 126390
rect 74292 126334 74348 126390
rect 74434 126334 74490 126390
rect 74576 126334 74632 126390
rect 74718 126334 74774 126390
rect 74860 126334 74916 126390
rect 75002 126334 75058 126390
rect 75144 126334 75200 126390
rect 75286 126334 75342 126390
rect 73866 99594 73922 99650
rect 74008 99594 74064 99650
rect 74150 99594 74206 99650
rect 74292 99594 74348 99650
rect 74434 99594 74490 99650
rect 74576 99594 74632 99650
rect 74718 99594 74774 99650
rect 74860 99594 74916 99650
rect 75002 99594 75058 99650
rect 75144 99594 75200 99650
rect 75286 99594 75342 99650
rect 73866 99452 73922 99508
rect 74008 99452 74064 99508
rect 74150 99452 74206 99508
rect 74292 99452 74348 99508
rect 74434 99452 74490 99508
rect 74576 99452 74632 99508
rect 74718 99452 74774 99508
rect 74860 99452 74916 99508
rect 75002 99452 75058 99508
rect 75144 99452 75200 99508
rect 75286 99452 75342 99508
rect 73866 99310 73922 99366
rect 74008 99310 74064 99366
rect 74150 99310 74206 99366
rect 74292 99310 74348 99366
rect 74434 99310 74490 99366
rect 74576 99310 74632 99366
rect 74718 99310 74774 99366
rect 74860 99310 74916 99366
rect 75002 99310 75058 99366
rect 75144 99310 75200 99366
rect 75286 99310 75342 99366
rect 73866 99168 73922 99224
rect 74008 99168 74064 99224
rect 74150 99168 74206 99224
rect 74292 99168 74348 99224
rect 74434 99168 74490 99224
rect 74576 99168 74632 99224
rect 74718 99168 74774 99224
rect 74860 99168 74916 99224
rect 75002 99168 75058 99224
rect 75144 99168 75200 99224
rect 75286 99168 75342 99224
rect 73866 99026 73922 99082
rect 74008 99026 74064 99082
rect 74150 99026 74206 99082
rect 74292 99026 74348 99082
rect 74434 99026 74490 99082
rect 74576 99026 74632 99082
rect 74718 99026 74774 99082
rect 74860 99026 74916 99082
rect 75002 99026 75058 99082
rect 75144 99026 75200 99082
rect 75286 99026 75342 99082
rect 73866 98884 73922 98940
rect 74008 98884 74064 98940
rect 74150 98884 74206 98940
rect 74292 98884 74348 98940
rect 74434 98884 74490 98940
rect 74576 98884 74632 98940
rect 74718 98884 74774 98940
rect 74860 98884 74916 98940
rect 75002 98884 75058 98940
rect 75144 98884 75200 98940
rect 75286 98884 75342 98940
rect 73866 98742 73922 98798
rect 74008 98742 74064 98798
rect 74150 98742 74206 98798
rect 74292 98742 74348 98798
rect 74434 98742 74490 98798
rect 74576 98742 74632 98798
rect 74718 98742 74774 98798
rect 74860 98742 74916 98798
rect 75002 98742 75058 98798
rect 75144 98742 75200 98798
rect 75286 98742 75342 98798
rect 73866 98600 73922 98656
rect 74008 98600 74064 98656
rect 74150 98600 74206 98656
rect 74292 98600 74348 98656
rect 74434 98600 74490 98656
rect 74576 98600 74632 98656
rect 74718 98600 74774 98656
rect 74860 98600 74916 98656
rect 75002 98600 75058 98656
rect 75144 98600 75200 98656
rect 75286 98600 75342 98656
rect 73866 98458 73922 98514
rect 74008 98458 74064 98514
rect 74150 98458 74206 98514
rect 74292 98458 74348 98514
rect 74434 98458 74490 98514
rect 74576 98458 74632 98514
rect 74718 98458 74774 98514
rect 74860 98458 74916 98514
rect 75002 98458 75058 98514
rect 75144 98458 75200 98514
rect 75286 98458 75342 98514
rect 73866 98316 73922 98372
rect 74008 98316 74064 98372
rect 74150 98316 74206 98372
rect 74292 98316 74348 98372
rect 74434 98316 74490 98372
rect 74576 98316 74632 98372
rect 74718 98316 74774 98372
rect 74860 98316 74916 98372
rect 75002 98316 75058 98372
rect 75144 98316 75200 98372
rect 75286 98316 75342 98372
rect 73866 98174 73922 98230
rect 74008 98174 74064 98230
rect 74150 98174 74206 98230
rect 74292 98174 74348 98230
rect 74434 98174 74490 98230
rect 74576 98174 74632 98230
rect 74718 98174 74774 98230
rect 74860 98174 74916 98230
rect 75002 98174 75058 98230
rect 75144 98174 75200 98230
rect 75286 98174 75342 98230
rect 73866 98032 73922 98088
rect 74008 98032 74064 98088
rect 74150 98032 74206 98088
rect 74292 98032 74348 98088
rect 74434 98032 74490 98088
rect 74576 98032 74632 98088
rect 74718 98032 74774 98088
rect 74860 98032 74916 98088
rect 75002 98032 75058 98088
rect 75144 98032 75200 98088
rect 75286 98032 75342 98088
rect 73866 97890 73922 97946
rect 74008 97890 74064 97946
rect 74150 97890 74206 97946
rect 74292 97890 74348 97946
rect 74434 97890 74490 97946
rect 74576 97890 74632 97946
rect 74718 97890 74774 97946
rect 74860 97890 74916 97946
rect 75002 97890 75058 97946
rect 75144 97890 75200 97946
rect 75286 97890 75342 97946
rect 73855 97113 73911 97169
rect 73997 97113 74053 97169
rect 74139 97113 74195 97169
rect 74281 97113 74337 97169
rect 74423 97113 74479 97169
rect 74565 97113 74621 97169
rect 74707 97113 74763 97169
rect 74849 97113 74905 97169
rect 74991 97113 75047 97169
rect 75133 97113 75189 97169
rect 75275 97113 75331 97169
rect 73855 96971 73911 97027
rect 73997 96971 74053 97027
rect 74139 96971 74195 97027
rect 74281 96971 74337 97027
rect 74423 96971 74479 97027
rect 74565 96971 74621 97027
rect 74707 96971 74763 97027
rect 74849 96971 74905 97027
rect 74991 96971 75047 97027
rect 75133 96971 75189 97027
rect 75275 96971 75331 97027
rect 73855 96829 73911 96885
rect 73997 96829 74053 96885
rect 74139 96829 74195 96885
rect 74281 96829 74337 96885
rect 74423 96829 74479 96885
rect 74565 96829 74621 96885
rect 74707 96829 74763 96885
rect 74849 96829 74905 96885
rect 74991 96829 75047 96885
rect 75133 96829 75189 96885
rect 75275 96829 75331 96885
rect 73855 96687 73911 96743
rect 73997 96687 74053 96743
rect 74139 96687 74195 96743
rect 74281 96687 74337 96743
rect 74423 96687 74479 96743
rect 74565 96687 74621 96743
rect 74707 96687 74763 96743
rect 74849 96687 74905 96743
rect 74991 96687 75047 96743
rect 75133 96687 75189 96743
rect 75275 96687 75331 96743
rect 73855 96545 73911 96601
rect 73997 96545 74053 96601
rect 74139 96545 74195 96601
rect 74281 96545 74337 96601
rect 74423 96545 74479 96601
rect 74565 96545 74621 96601
rect 74707 96545 74763 96601
rect 74849 96545 74905 96601
rect 74991 96545 75047 96601
rect 75133 96545 75189 96601
rect 75275 96545 75331 96601
rect 73855 96403 73911 96459
rect 73997 96403 74053 96459
rect 74139 96403 74195 96459
rect 74281 96403 74337 96459
rect 74423 96403 74479 96459
rect 74565 96403 74621 96459
rect 74707 96403 74763 96459
rect 74849 96403 74905 96459
rect 74991 96403 75047 96459
rect 75133 96403 75189 96459
rect 75275 96403 75331 96459
rect 73855 96261 73911 96317
rect 73997 96261 74053 96317
rect 74139 96261 74195 96317
rect 74281 96261 74337 96317
rect 74423 96261 74479 96317
rect 74565 96261 74621 96317
rect 74707 96261 74763 96317
rect 74849 96261 74905 96317
rect 74991 96261 75047 96317
rect 75133 96261 75189 96317
rect 75275 96261 75331 96317
rect 73855 96119 73911 96175
rect 73997 96119 74053 96175
rect 74139 96119 74195 96175
rect 74281 96119 74337 96175
rect 74423 96119 74479 96175
rect 74565 96119 74621 96175
rect 74707 96119 74763 96175
rect 74849 96119 74905 96175
rect 74991 96119 75047 96175
rect 75133 96119 75189 96175
rect 75275 96119 75331 96175
rect 73855 95977 73911 96033
rect 73997 95977 74053 96033
rect 74139 95977 74195 96033
rect 74281 95977 74337 96033
rect 74423 95977 74479 96033
rect 74565 95977 74621 96033
rect 74707 95977 74763 96033
rect 74849 95977 74905 96033
rect 74991 95977 75047 96033
rect 75133 95977 75189 96033
rect 75275 95977 75331 96033
rect 73855 95835 73911 95891
rect 73997 95835 74053 95891
rect 74139 95835 74195 95891
rect 74281 95835 74337 95891
rect 74423 95835 74479 95891
rect 74565 95835 74621 95891
rect 74707 95835 74763 95891
rect 74849 95835 74905 95891
rect 74991 95835 75047 95891
rect 75133 95835 75189 95891
rect 75275 95835 75331 95891
rect 73855 95693 73911 95749
rect 73997 95693 74053 95749
rect 74139 95693 74195 95749
rect 74281 95693 74337 95749
rect 74423 95693 74479 95749
rect 74565 95693 74621 95749
rect 74707 95693 74763 95749
rect 74849 95693 74905 95749
rect 74991 95693 75047 95749
rect 75133 95693 75189 95749
rect 75275 95693 75331 95749
rect 73855 95551 73911 95607
rect 73997 95551 74053 95607
rect 74139 95551 74195 95607
rect 74281 95551 74337 95607
rect 74423 95551 74479 95607
rect 74565 95551 74621 95607
rect 74707 95551 74763 95607
rect 74849 95551 74905 95607
rect 74991 95551 75047 95607
rect 75133 95551 75189 95607
rect 75275 95551 75331 95607
rect 73855 95409 73911 95465
rect 73997 95409 74053 95465
rect 74139 95409 74195 95465
rect 74281 95409 74337 95465
rect 74423 95409 74479 95465
rect 74565 95409 74621 95465
rect 74707 95409 74763 95465
rect 74849 95409 74905 95465
rect 74991 95409 75047 95465
rect 75133 95409 75189 95465
rect 75275 95409 75331 95465
rect 73855 95267 73911 95323
rect 73997 95267 74053 95323
rect 74139 95267 74195 95323
rect 74281 95267 74337 95323
rect 74423 95267 74479 95323
rect 74565 95267 74621 95323
rect 74707 95267 74763 95323
rect 74849 95267 74905 95323
rect 74991 95267 75047 95323
rect 75133 95267 75189 95323
rect 75275 95267 75331 95323
rect 73855 94743 73911 94799
rect 73997 94743 74053 94799
rect 74139 94743 74195 94799
rect 74281 94743 74337 94799
rect 74423 94743 74479 94799
rect 74565 94743 74621 94799
rect 74707 94743 74763 94799
rect 74849 94743 74905 94799
rect 74991 94743 75047 94799
rect 75133 94743 75189 94799
rect 75275 94743 75331 94799
rect 73855 94601 73911 94657
rect 73997 94601 74053 94657
rect 74139 94601 74195 94657
rect 74281 94601 74337 94657
rect 74423 94601 74479 94657
rect 74565 94601 74621 94657
rect 74707 94601 74763 94657
rect 74849 94601 74905 94657
rect 74991 94601 75047 94657
rect 75133 94601 75189 94657
rect 75275 94601 75331 94657
rect 73855 94459 73911 94515
rect 73997 94459 74053 94515
rect 74139 94459 74195 94515
rect 74281 94459 74337 94515
rect 74423 94459 74479 94515
rect 74565 94459 74621 94515
rect 74707 94459 74763 94515
rect 74849 94459 74905 94515
rect 74991 94459 75047 94515
rect 75133 94459 75189 94515
rect 75275 94459 75331 94515
rect 73855 94317 73911 94373
rect 73997 94317 74053 94373
rect 74139 94317 74195 94373
rect 74281 94317 74337 94373
rect 74423 94317 74479 94373
rect 74565 94317 74621 94373
rect 74707 94317 74763 94373
rect 74849 94317 74905 94373
rect 74991 94317 75047 94373
rect 75133 94317 75189 94373
rect 75275 94317 75331 94373
rect 73855 94175 73911 94231
rect 73997 94175 74053 94231
rect 74139 94175 74195 94231
rect 74281 94175 74337 94231
rect 74423 94175 74479 94231
rect 74565 94175 74621 94231
rect 74707 94175 74763 94231
rect 74849 94175 74905 94231
rect 74991 94175 75047 94231
rect 75133 94175 75189 94231
rect 75275 94175 75331 94231
rect 73855 94033 73911 94089
rect 73997 94033 74053 94089
rect 74139 94033 74195 94089
rect 74281 94033 74337 94089
rect 74423 94033 74479 94089
rect 74565 94033 74621 94089
rect 74707 94033 74763 94089
rect 74849 94033 74905 94089
rect 74991 94033 75047 94089
rect 75133 94033 75189 94089
rect 75275 94033 75331 94089
rect 73855 93891 73911 93947
rect 73997 93891 74053 93947
rect 74139 93891 74195 93947
rect 74281 93891 74337 93947
rect 74423 93891 74479 93947
rect 74565 93891 74621 93947
rect 74707 93891 74763 93947
rect 74849 93891 74905 93947
rect 74991 93891 75047 93947
rect 75133 93891 75189 93947
rect 75275 93891 75331 93947
rect 73855 93749 73911 93805
rect 73997 93749 74053 93805
rect 74139 93749 74195 93805
rect 74281 93749 74337 93805
rect 74423 93749 74479 93805
rect 74565 93749 74621 93805
rect 74707 93749 74763 93805
rect 74849 93749 74905 93805
rect 74991 93749 75047 93805
rect 75133 93749 75189 93805
rect 75275 93749 75331 93805
rect 73855 93607 73911 93663
rect 73997 93607 74053 93663
rect 74139 93607 74195 93663
rect 74281 93607 74337 93663
rect 74423 93607 74479 93663
rect 74565 93607 74621 93663
rect 74707 93607 74763 93663
rect 74849 93607 74905 93663
rect 74991 93607 75047 93663
rect 75133 93607 75189 93663
rect 75275 93607 75331 93663
rect 73855 93465 73911 93521
rect 73997 93465 74053 93521
rect 74139 93465 74195 93521
rect 74281 93465 74337 93521
rect 74423 93465 74479 93521
rect 74565 93465 74621 93521
rect 74707 93465 74763 93521
rect 74849 93465 74905 93521
rect 74991 93465 75047 93521
rect 75133 93465 75189 93521
rect 75275 93465 75331 93521
rect 73855 93323 73911 93379
rect 73997 93323 74053 93379
rect 74139 93323 74195 93379
rect 74281 93323 74337 93379
rect 74423 93323 74479 93379
rect 74565 93323 74621 93379
rect 74707 93323 74763 93379
rect 74849 93323 74905 93379
rect 74991 93323 75047 93379
rect 75133 93323 75189 93379
rect 75275 93323 75331 93379
rect 73855 93181 73911 93237
rect 73997 93181 74053 93237
rect 74139 93181 74195 93237
rect 74281 93181 74337 93237
rect 74423 93181 74479 93237
rect 74565 93181 74621 93237
rect 74707 93181 74763 93237
rect 74849 93181 74905 93237
rect 74991 93181 75047 93237
rect 75133 93181 75189 93237
rect 75275 93181 75331 93237
rect 73855 93039 73911 93095
rect 73997 93039 74053 93095
rect 74139 93039 74195 93095
rect 74281 93039 74337 93095
rect 74423 93039 74479 93095
rect 74565 93039 74621 93095
rect 74707 93039 74763 93095
rect 74849 93039 74905 93095
rect 74991 93039 75047 93095
rect 75133 93039 75189 93095
rect 75275 93039 75331 93095
rect 73855 92897 73911 92953
rect 73997 92897 74053 92953
rect 74139 92897 74195 92953
rect 74281 92897 74337 92953
rect 74423 92897 74479 92953
rect 74565 92897 74621 92953
rect 74707 92897 74763 92953
rect 74849 92897 74905 92953
rect 74991 92897 75047 92953
rect 75133 92897 75189 92953
rect 75275 92897 75331 92953
rect 73855 92037 73911 92093
rect 73997 92037 74053 92093
rect 74139 92037 74195 92093
rect 74281 92037 74337 92093
rect 74423 92037 74479 92093
rect 74565 92037 74621 92093
rect 74707 92037 74763 92093
rect 74849 92037 74905 92093
rect 74991 92037 75047 92093
rect 75133 92037 75189 92093
rect 75275 92037 75331 92093
rect 73855 91895 73911 91951
rect 73997 91895 74053 91951
rect 74139 91895 74195 91951
rect 74281 91895 74337 91951
rect 74423 91895 74479 91951
rect 74565 91895 74621 91951
rect 74707 91895 74763 91951
rect 74849 91895 74905 91951
rect 74991 91895 75047 91951
rect 75133 91895 75189 91951
rect 75275 91895 75331 91951
rect 73855 91753 73911 91809
rect 73997 91753 74053 91809
rect 74139 91753 74195 91809
rect 74281 91753 74337 91809
rect 74423 91753 74479 91809
rect 74565 91753 74621 91809
rect 74707 91753 74763 91809
rect 74849 91753 74905 91809
rect 74991 91753 75047 91809
rect 75133 91753 75189 91809
rect 75275 91753 75331 91809
rect 73855 91611 73911 91667
rect 73997 91611 74053 91667
rect 74139 91611 74195 91667
rect 74281 91611 74337 91667
rect 74423 91611 74479 91667
rect 74565 91611 74621 91667
rect 74707 91611 74763 91667
rect 74849 91611 74905 91667
rect 74991 91611 75047 91667
rect 75133 91611 75189 91667
rect 75275 91611 75331 91667
rect 73855 91469 73911 91525
rect 73997 91469 74053 91525
rect 74139 91469 74195 91525
rect 74281 91469 74337 91525
rect 74423 91469 74479 91525
rect 74565 91469 74621 91525
rect 74707 91469 74763 91525
rect 74849 91469 74905 91525
rect 74991 91469 75047 91525
rect 75133 91469 75189 91525
rect 75275 91469 75331 91525
rect 73855 91327 73911 91383
rect 73997 91327 74053 91383
rect 74139 91327 74195 91383
rect 74281 91327 74337 91383
rect 74423 91327 74479 91383
rect 74565 91327 74621 91383
rect 74707 91327 74763 91383
rect 74849 91327 74905 91383
rect 74991 91327 75047 91383
rect 75133 91327 75189 91383
rect 75275 91327 75331 91383
rect 73855 91185 73911 91241
rect 73997 91185 74053 91241
rect 74139 91185 74195 91241
rect 74281 91185 74337 91241
rect 74423 91185 74479 91241
rect 74565 91185 74621 91241
rect 74707 91185 74763 91241
rect 74849 91185 74905 91241
rect 74991 91185 75047 91241
rect 75133 91185 75189 91241
rect 75275 91185 75331 91241
rect 73855 91043 73911 91099
rect 73997 91043 74053 91099
rect 74139 91043 74195 91099
rect 74281 91043 74337 91099
rect 74423 91043 74479 91099
rect 74565 91043 74621 91099
rect 74707 91043 74763 91099
rect 74849 91043 74905 91099
rect 74991 91043 75047 91099
rect 75133 91043 75189 91099
rect 75275 91043 75331 91099
rect 73855 90901 73911 90957
rect 73997 90901 74053 90957
rect 74139 90901 74195 90957
rect 74281 90901 74337 90957
rect 74423 90901 74479 90957
rect 74565 90901 74621 90957
rect 74707 90901 74763 90957
rect 74849 90901 74905 90957
rect 74991 90901 75047 90957
rect 75133 90901 75189 90957
rect 75275 90901 75331 90957
rect 73855 90759 73911 90815
rect 73997 90759 74053 90815
rect 74139 90759 74195 90815
rect 74281 90759 74337 90815
rect 74423 90759 74479 90815
rect 74565 90759 74621 90815
rect 74707 90759 74763 90815
rect 74849 90759 74905 90815
rect 74991 90759 75047 90815
rect 75133 90759 75189 90815
rect 75275 90759 75331 90815
rect 73855 90617 73911 90673
rect 73997 90617 74053 90673
rect 74139 90617 74195 90673
rect 74281 90617 74337 90673
rect 74423 90617 74479 90673
rect 74565 90617 74621 90673
rect 74707 90617 74763 90673
rect 74849 90617 74905 90673
rect 74991 90617 75047 90673
rect 75133 90617 75189 90673
rect 75275 90617 75331 90673
rect 73855 90475 73911 90531
rect 73997 90475 74053 90531
rect 74139 90475 74195 90531
rect 74281 90475 74337 90531
rect 74423 90475 74479 90531
rect 74565 90475 74621 90531
rect 74707 90475 74763 90531
rect 74849 90475 74905 90531
rect 74991 90475 75047 90531
rect 75133 90475 75189 90531
rect 75275 90475 75331 90531
rect 73855 90333 73911 90389
rect 73997 90333 74053 90389
rect 74139 90333 74195 90389
rect 74281 90333 74337 90389
rect 74423 90333 74479 90389
rect 74565 90333 74621 90389
rect 74707 90333 74763 90389
rect 74849 90333 74905 90389
rect 74991 90333 75047 90389
rect 75133 90333 75189 90389
rect 75275 90333 75331 90389
rect 73855 90191 73911 90247
rect 73997 90191 74053 90247
rect 74139 90191 74195 90247
rect 74281 90191 74337 90247
rect 74423 90191 74479 90247
rect 74565 90191 74621 90247
rect 74707 90191 74763 90247
rect 74849 90191 74905 90247
rect 74991 90191 75047 90247
rect 75133 90191 75189 90247
rect 75275 90191 75331 90247
rect 73855 89667 73911 89723
rect 73997 89667 74053 89723
rect 74139 89667 74195 89723
rect 74281 89667 74337 89723
rect 74423 89667 74479 89723
rect 74565 89667 74621 89723
rect 74707 89667 74763 89723
rect 74849 89667 74905 89723
rect 74991 89667 75047 89723
rect 75133 89667 75189 89723
rect 75275 89667 75331 89723
rect 73855 89525 73911 89581
rect 73997 89525 74053 89581
rect 74139 89525 74195 89581
rect 74281 89525 74337 89581
rect 74423 89525 74479 89581
rect 74565 89525 74621 89581
rect 74707 89525 74763 89581
rect 74849 89525 74905 89581
rect 74991 89525 75047 89581
rect 75133 89525 75189 89581
rect 75275 89525 75331 89581
rect 73855 89383 73911 89439
rect 73997 89383 74053 89439
rect 74139 89383 74195 89439
rect 74281 89383 74337 89439
rect 74423 89383 74479 89439
rect 74565 89383 74621 89439
rect 74707 89383 74763 89439
rect 74849 89383 74905 89439
rect 74991 89383 75047 89439
rect 75133 89383 75189 89439
rect 75275 89383 75331 89439
rect 73855 89241 73911 89297
rect 73997 89241 74053 89297
rect 74139 89241 74195 89297
rect 74281 89241 74337 89297
rect 74423 89241 74479 89297
rect 74565 89241 74621 89297
rect 74707 89241 74763 89297
rect 74849 89241 74905 89297
rect 74991 89241 75047 89297
rect 75133 89241 75189 89297
rect 75275 89241 75331 89297
rect 73855 89099 73911 89155
rect 73997 89099 74053 89155
rect 74139 89099 74195 89155
rect 74281 89099 74337 89155
rect 74423 89099 74479 89155
rect 74565 89099 74621 89155
rect 74707 89099 74763 89155
rect 74849 89099 74905 89155
rect 74991 89099 75047 89155
rect 75133 89099 75189 89155
rect 75275 89099 75331 89155
rect 73855 88957 73911 89013
rect 73997 88957 74053 89013
rect 74139 88957 74195 89013
rect 74281 88957 74337 89013
rect 74423 88957 74479 89013
rect 74565 88957 74621 89013
rect 74707 88957 74763 89013
rect 74849 88957 74905 89013
rect 74991 88957 75047 89013
rect 75133 88957 75189 89013
rect 75275 88957 75331 89013
rect 73855 88815 73911 88871
rect 73997 88815 74053 88871
rect 74139 88815 74195 88871
rect 74281 88815 74337 88871
rect 74423 88815 74479 88871
rect 74565 88815 74621 88871
rect 74707 88815 74763 88871
rect 74849 88815 74905 88871
rect 74991 88815 75047 88871
rect 75133 88815 75189 88871
rect 75275 88815 75331 88871
rect 73855 88673 73911 88729
rect 73997 88673 74053 88729
rect 74139 88673 74195 88729
rect 74281 88673 74337 88729
rect 74423 88673 74479 88729
rect 74565 88673 74621 88729
rect 74707 88673 74763 88729
rect 74849 88673 74905 88729
rect 74991 88673 75047 88729
rect 75133 88673 75189 88729
rect 75275 88673 75331 88729
rect 73855 88531 73911 88587
rect 73997 88531 74053 88587
rect 74139 88531 74195 88587
rect 74281 88531 74337 88587
rect 74423 88531 74479 88587
rect 74565 88531 74621 88587
rect 74707 88531 74763 88587
rect 74849 88531 74905 88587
rect 74991 88531 75047 88587
rect 75133 88531 75189 88587
rect 75275 88531 75331 88587
rect 73855 88389 73911 88445
rect 73997 88389 74053 88445
rect 74139 88389 74195 88445
rect 74281 88389 74337 88445
rect 74423 88389 74479 88445
rect 74565 88389 74621 88445
rect 74707 88389 74763 88445
rect 74849 88389 74905 88445
rect 74991 88389 75047 88445
rect 75133 88389 75189 88445
rect 75275 88389 75331 88445
rect 73855 88247 73911 88303
rect 73997 88247 74053 88303
rect 74139 88247 74195 88303
rect 74281 88247 74337 88303
rect 74423 88247 74479 88303
rect 74565 88247 74621 88303
rect 74707 88247 74763 88303
rect 74849 88247 74905 88303
rect 74991 88247 75047 88303
rect 75133 88247 75189 88303
rect 75275 88247 75331 88303
rect 73855 88105 73911 88161
rect 73997 88105 74053 88161
rect 74139 88105 74195 88161
rect 74281 88105 74337 88161
rect 74423 88105 74479 88161
rect 74565 88105 74621 88161
rect 74707 88105 74763 88161
rect 74849 88105 74905 88161
rect 74991 88105 75047 88161
rect 75133 88105 75189 88161
rect 75275 88105 75331 88161
rect 73855 87963 73911 88019
rect 73997 87963 74053 88019
rect 74139 87963 74195 88019
rect 74281 87963 74337 88019
rect 74423 87963 74479 88019
rect 74565 87963 74621 88019
rect 74707 87963 74763 88019
rect 74849 87963 74905 88019
rect 74991 87963 75047 88019
rect 75133 87963 75189 88019
rect 75275 87963 75331 88019
rect 73855 87821 73911 87877
rect 73997 87821 74053 87877
rect 74139 87821 74195 87877
rect 74281 87821 74337 87877
rect 74423 87821 74479 87877
rect 74565 87821 74621 87877
rect 74707 87821 74763 87877
rect 74849 87821 74905 87877
rect 74991 87821 75047 87877
rect 75133 87821 75189 87877
rect 75275 87821 75331 87877
rect 73866 87038 73922 87094
rect 74008 87038 74064 87094
rect 74150 87038 74206 87094
rect 74292 87038 74348 87094
rect 74434 87038 74490 87094
rect 74576 87038 74632 87094
rect 74718 87038 74774 87094
rect 74860 87038 74916 87094
rect 75002 87038 75058 87094
rect 75144 87038 75200 87094
rect 75286 87038 75342 87094
rect 73866 86896 73922 86952
rect 74008 86896 74064 86952
rect 74150 86896 74206 86952
rect 74292 86896 74348 86952
rect 74434 86896 74490 86952
rect 74576 86896 74632 86952
rect 74718 86896 74774 86952
rect 74860 86896 74916 86952
rect 75002 86896 75058 86952
rect 75144 86896 75200 86952
rect 75286 86896 75342 86952
rect 73866 86754 73922 86810
rect 74008 86754 74064 86810
rect 74150 86754 74206 86810
rect 74292 86754 74348 86810
rect 74434 86754 74490 86810
rect 74576 86754 74632 86810
rect 74718 86754 74774 86810
rect 74860 86754 74916 86810
rect 75002 86754 75058 86810
rect 75144 86754 75200 86810
rect 75286 86754 75342 86810
rect 73866 86612 73922 86668
rect 74008 86612 74064 86668
rect 74150 86612 74206 86668
rect 74292 86612 74348 86668
rect 74434 86612 74490 86668
rect 74576 86612 74632 86668
rect 74718 86612 74774 86668
rect 74860 86612 74916 86668
rect 75002 86612 75058 86668
rect 75144 86612 75200 86668
rect 75286 86612 75342 86668
rect 73866 86470 73922 86526
rect 74008 86470 74064 86526
rect 74150 86470 74206 86526
rect 74292 86470 74348 86526
rect 74434 86470 74490 86526
rect 74576 86470 74632 86526
rect 74718 86470 74774 86526
rect 74860 86470 74916 86526
rect 75002 86470 75058 86526
rect 75144 86470 75200 86526
rect 75286 86470 75342 86526
rect 73866 86328 73922 86384
rect 74008 86328 74064 86384
rect 74150 86328 74206 86384
rect 74292 86328 74348 86384
rect 74434 86328 74490 86384
rect 74576 86328 74632 86384
rect 74718 86328 74774 86384
rect 74860 86328 74916 86384
rect 75002 86328 75058 86384
rect 75144 86328 75200 86384
rect 75286 86328 75342 86384
rect 73866 86186 73922 86242
rect 74008 86186 74064 86242
rect 74150 86186 74206 86242
rect 74292 86186 74348 86242
rect 74434 86186 74490 86242
rect 74576 86186 74632 86242
rect 74718 86186 74774 86242
rect 74860 86186 74916 86242
rect 75002 86186 75058 86242
rect 75144 86186 75200 86242
rect 75286 86186 75342 86242
rect 73866 86044 73922 86100
rect 74008 86044 74064 86100
rect 74150 86044 74206 86100
rect 74292 86044 74348 86100
rect 74434 86044 74490 86100
rect 74576 86044 74632 86100
rect 74718 86044 74774 86100
rect 74860 86044 74916 86100
rect 75002 86044 75058 86100
rect 75144 86044 75200 86100
rect 75286 86044 75342 86100
rect 73866 85902 73922 85958
rect 74008 85902 74064 85958
rect 74150 85902 74206 85958
rect 74292 85902 74348 85958
rect 74434 85902 74490 85958
rect 74576 85902 74632 85958
rect 74718 85902 74774 85958
rect 74860 85902 74916 85958
rect 75002 85902 75058 85958
rect 75144 85902 75200 85958
rect 75286 85902 75342 85958
rect 73866 85760 73922 85816
rect 74008 85760 74064 85816
rect 74150 85760 74206 85816
rect 74292 85760 74348 85816
rect 74434 85760 74490 85816
rect 74576 85760 74632 85816
rect 74718 85760 74774 85816
rect 74860 85760 74916 85816
rect 75002 85760 75058 85816
rect 75144 85760 75200 85816
rect 75286 85760 75342 85816
rect 73866 85618 73922 85674
rect 74008 85618 74064 85674
rect 74150 85618 74206 85674
rect 74292 85618 74348 85674
rect 74434 85618 74490 85674
rect 74576 85618 74632 85674
rect 74718 85618 74774 85674
rect 74860 85618 74916 85674
rect 75002 85618 75058 85674
rect 75144 85618 75200 85674
rect 75286 85618 75342 85674
rect 73866 85476 73922 85532
rect 74008 85476 74064 85532
rect 74150 85476 74206 85532
rect 74292 85476 74348 85532
rect 74434 85476 74490 85532
rect 74576 85476 74632 85532
rect 74718 85476 74774 85532
rect 74860 85476 74916 85532
rect 75002 85476 75058 85532
rect 75144 85476 75200 85532
rect 75286 85476 75342 85532
rect 73866 85334 73922 85390
rect 74008 85334 74064 85390
rect 74150 85334 74206 85390
rect 74292 85334 74348 85390
rect 74434 85334 74490 85390
rect 74576 85334 74632 85390
rect 74718 85334 74774 85390
rect 74860 85334 74916 85390
rect 75002 85334 75058 85390
rect 75144 85334 75200 85390
rect 75286 85334 75342 85390
rect 655343 75979 655399 76035
rect 655485 75979 655541 76035
rect 655627 75979 655683 76035
rect 655769 75979 655825 76035
rect 655911 75979 655967 76035
rect 656053 75979 656109 76035
rect 656195 75979 656251 76035
rect 656337 75979 656393 76035
rect 655343 75889 655382 75893
rect 655382 75889 655399 75893
rect 655485 75889 655506 75893
rect 655506 75889 655541 75893
rect 655627 75889 655630 75893
rect 655630 75889 655683 75893
rect 655769 75889 655822 75893
rect 655822 75889 655825 75893
rect 655911 75889 655946 75893
rect 655946 75889 655967 75893
rect 656053 75889 656070 75893
rect 656070 75889 656109 75893
rect 656195 75889 656250 75893
rect 656250 75889 656251 75893
rect 656337 75889 656374 75893
rect 656374 75889 656393 75893
rect 655343 75837 655399 75889
rect 655485 75837 655541 75889
rect 655627 75837 655683 75889
rect 655769 75837 655825 75889
rect 655911 75837 655967 75889
rect 656053 75837 656109 75889
rect 656195 75837 656251 75889
rect 656337 75837 656393 75889
rect 655343 75697 655399 75751
rect 655485 75697 655541 75751
rect 655627 75697 655683 75751
rect 655769 75697 655825 75751
rect 655911 75697 655967 75751
rect 656053 75697 656109 75751
rect 656195 75697 656251 75751
rect 656337 75697 656393 75751
rect 655343 75695 655382 75697
rect 655382 75695 655399 75697
rect 655485 75695 655506 75697
rect 655506 75695 655541 75697
rect 655627 75695 655630 75697
rect 655630 75695 655683 75697
rect 655769 75695 655822 75697
rect 655822 75695 655825 75697
rect 655911 75695 655946 75697
rect 655946 75695 655967 75697
rect 656053 75695 656070 75697
rect 656070 75695 656109 75697
rect 656195 75695 656250 75697
rect 656250 75695 656251 75697
rect 656337 75695 656374 75697
rect 656374 75695 656393 75697
rect 655343 75573 655399 75609
rect 655485 75573 655541 75609
rect 655627 75573 655683 75609
rect 655769 75573 655825 75609
rect 655911 75573 655967 75609
rect 656053 75573 656109 75609
rect 656195 75573 656251 75609
rect 656337 75573 656393 75609
rect 655343 75553 655382 75573
rect 655382 75553 655399 75573
rect 655485 75553 655506 75573
rect 655506 75553 655541 75573
rect 655627 75553 655630 75573
rect 655630 75553 655683 75573
rect 655769 75553 655822 75573
rect 655822 75553 655825 75573
rect 655911 75553 655946 75573
rect 655946 75553 655967 75573
rect 656053 75553 656070 75573
rect 656070 75553 656109 75573
rect 656195 75553 656250 75573
rect 656250 75553 656251 75573
rect 656337 75553 656374 75573
rect 656374 75553 656393 75573
rect 655343 75449 655399 75467
rect 655485 75449 655541 75467
rect 655627 75449 655683 75467
rect 655769 75449 655825 75467
rect 655911 75449 655967 75467
rect 656053 75449 656109 75467
rect 656195 75449 656251 75467
rect 656337 75449 656393 75467
rect 655343 75411 655382 75449
rect 655382 75411 655399 75449
rect 655485 75411 655506 75449
rect 655506 75411 655541 75449
rect 655627 75411 655630 75449
rect 655630 75411 655683 75449
rect 655769 75411 655822 75449
rect 655822 75411 655825 75449
rect 655911 75411 655946 75449
rect 655946 75411 655967 75449
rect 656053 75411 656070 75449
rect 656070 75411 656109 75449
rect 656195 75411 656250 75449
rect 656250 75411 656251 75449
rect 656337 75411 656374 75449
rect 656374 75411 656393 75449
rect 655343 75269 655382 75325
rect 655382 75269 655399 75325
rect 655485 75269 655506 75325
rect 655506 75269 655541 75325
rect 655627 75269 655630 75325
rect 655630 75269 655683 75325
rect 655769 75269 655822 75325
rect 655822 75269 655825 75325
rect 655911 75269 655946 75325
rect 655946 75269 655967 75325
rect 656053 75269 656070 75325
rect 656070 75269 656109 75325
rect 656195 75269 656250 75325
rect 656250 75269 656251 75325
rect 656337 75269 656374 75325
rect 656374 75269 656393 75325
rect 655343 75145 655382 75183
rect 655382 75145 655399 75183
rect 655485 75145 655506 75183
rect 655506 75145 655541 75183
rect 655627 75145 655630 75183
rect 655630 75145 655683 75183
rect 655769 75145 655822 75183
rect 655822 75145 655825 75183
rect 655911 75145 655946 75183
rect 655946 75145 655967 75183
rect 656053 75145 656070 75183
rect 656070 75145 656109 75183
rect 656195 75145 656250 75183
rect 656250 75145 656251 75183
rect 656337 75145 656374 75183
rect 656374 75145 656393 75183
rect 655343 75127 655399 75145
rect 655485 75127 655541 75145
rect 655627 75127 655683 75145
rect 655769 75127 655825 75145
rect 655911 75127 655967 75145
rect 656053 75127 656109 75145
rect 656195 75127 656251 75145
rect 656337 75127 656393 75145
rect 655343 75021 655382 75041
rect 655382 75021 655399 75041
rect 655485 75021 655506 75041
rect 655506 75021 655541 75041
rect 655627 75021 655630 75041
rect 655630 75021 655683 75041
rect 655769 75021 655822 75041
rect 655822 75021 655825 75041
rect 655911 75021 655946 75041
rect 655946 75021 655967 75041
rect 656053 75021 656070 75041
rect 656070 75021 656109 75041
rect 656195 75021 656250 75041
rect 656250 75021 656251 75041
rect 656337 75021 656374 75041
rect 656374 75021 656393 75041
rect 655343 74985 655399 75021
rect 655485 74985 655541 75021
rect 655627 74985 655683 75021
rect 655769 74985 655825 75021
rect 655911 74985 655967 75021
rect 656053 74985 656109 75021
rect 656195 74985 656251 75021
rect 656337 74985 656393 75021
rect 655343 74897 655382 74899
rect 655382 74897 655399 74899
rect 655485 74897 655506 74899
rect 655506 74897 655541 74899
rect 655627 74897 655630 74899
rect 655630 74897 655683 74899
rect 655769 74897 655822 74899
rect 655822 74897 655825 74899
rect 655911 74897 655946 74899
rect 655946 74897 655967 74899
rect 656053 74897 656070 74899
rect 656070 74897 656109 74899
rect 656195 74897 656250 74899
rect 656250 74897 656251 74899
rect 656337 74897 656374 74899
rect 656374 74897 656393 74899
rect 655343 74843 655399 74897
rect 655485 74843 655541 74897
rect 655627 74843 655683 74897
rect 655769 74843 655825 74897
rect 655911 74843 655967 74897
rect 656053 74843 656109 74897
rect 656195 74843 656251 74897
rect 656337 74843 656393 74897
rect 655343 74705 655399 74757
rect 655485 74705 655541 74757
rect 655627 74705 655683 74757
rect 655769 74705 655825 74757
rect 655911 74705 655967 74757
rect 656053 74705 656109 74757
rect 656195 74705 656251 74757
rect 656337 74705 656393 74757
rect 655343 74701 655382 74705
rect 655382 74701 655399 74705
rect 655485 74701 655506 74705
rect 655506 74701 655541 74705
rect 655627 74701 655630 74705
rect 655630 74701 655683 74705
rect 655769 74701 655822 74705
rect 655822 74701 655825 74705
rect 655911 74701 655946 74705
rect 655946 74701 655967 74705
rect 656053 74701 656070 74705
rect 656070 74701 656109 74705
rect 656195 74701 656250 74705
rect 656250 74701 656251 74705
rect 656337 74701 656374 74705
rect 656374 74701 656393 74705
rect 655343 74581 655399 74615
rect 655485 74581 655541 74615
rect 655627 74581 655683 74615
rect 655769 74581 655825 74615
rect 655911 74581 655967 74615
rect 656053 74581 656109 74615
rect 656195 74581 656251 74615
rect 656337 74581 656393 74615
rect 655343 74559 655382 74581
rect 655382 74559 655399 74581
rect 655485 74559 655506 74581
rect 655506 74559 655541 74581
rect 655627 74559 655630 74581
rect 655630 74559 655683 74581
rect 655769 74559 655822 74581
rect 655822 74559 655825 74581
rect 655911 74559 655946 74581
rect 655946 74559 655967 74581
rect 656053 74559 656070 74581
rect 656070 74559 656109 74581
rect 656195 74559 656250 74581
rect 656250 74559 656251 74581
rect 656337 74559 656374 74581
rect 656374 74559 656393 74581
rect 657823 75979 657879 76035
rect 657965 75979 658021 76035
rect 658107 75979 658163 76035
rect 658249 75979 658305 76035
rect 658391 75979 658447 76035
rect 658533 75979 658589 76035
rect 658675 75979 658731 76035
rect 658817 75979 658873 76035
rect 658959 75979 659015 76035
rect 659101 75979 659157 76035
rect 659243 75979 659299 76035
rect 659385 75979 659441 76035
rect 659527 75979 659583 76035
rect 659669 75979 659725 76035
rect 657823 75889 657862 75893
rect 657862 75889 657879 75893
rect 657965 75889 657986 75893
rect 657986 75889 658021 75893
rect 658107 75889 658110 75893
rect 658110 75889 658163 75893
rect 658249 75889 658302 75893
rect 658302 75889 658305 75893
rect 658391 75889 658426 75893
rect 658426 75889 658447 75893
rect 658533 75889 658550 75893
rect 658550 75889 658589 75893
rect 658675 75889 658730 75893
rect 658730 75889 658731 75893
rect 658817 75889 658854 75893
rect 658854 75889 658873 75893
rect 658959 75889 658978 75893
rect 658978 75889 659015 75893
rect 659101 75889 659102 75893
rect 659102 75889 659157 75893
rect 659243 75889 659294 75893
rect 659294 75889 659299 75893
rect 659385 75889 659418 75893
rect 659418 75889 659441 75893
rect 659527 75889 659542 75893
rect 659542 75889 659583 75893
rect 659669 75889 659722 75893
rect 659722 75889 659725 75893
rect 657823 75837 657879 75889
rect 657965 75837 658021 75889
rect 658107 75837 658163 75889
rect 658249 75837 658305 75889
rect 658391 75837 658447 75889
rect 658533 75837 658589 75889
rect 658675 75837 658731 75889
rect 658817 75837 658873 75889
rect 658959 75837 659015 75889
rect 659101 75837 659157 75889
rect 659243 75837 659299 75889
rect 659385 75837 659441 75889
rect 659527 75837 659583 75889
rect 659669 75837 659725 75889
rect 657823 75697 657879 75751
rect 657965 75697 658021 75751
rect 658107 75697 658163 75751
rect 658249 75697 658305 75751
rect 658391 75697 658447 75751
rect 658533 75697 658589 75751
rect 658675 75697 658731 75751
rect 658817 75697 658873 75751
rect 658959 75697 659015 75751
rect 659101 75697 659157 75751
rect 659243 75697 659299 75751
rect 659385 75697 659441 75751
rect 659527 75697 659583 75751
rect 659669 75697 659725 75751
rect 657823 75695 657862 75697
rect 657862 75695 657879 75697
rect 657965 75695 657986 75697
rect 657986 75695 658021 75697
rect 658107 75695 658110 75697
rect 658110 75695 658163 75697
rect 658249 75695 658302 75697
rect 658302 75695 658305 75697
rect 658391 75695 658426 75697
rect 658426 75695 658447 75697
rect 658533 75695 658550 75697
rect 658550 75695 658589 75697
rect 658675 75695 658730 75697
rect 658730 75695 658731 75697
rect 658817 75695 658854 75697
rect 658854 75695 658873 75697
rect 658959 75695 658978 75697
rect 658978 75695 659015 75697
rect 659101 75695 659102 75697
rect 659102 75695 659157 75697
rect 659243 75695 659294 75697
rect 659294 75695 659299 75697
rect 659385 75695 659418 75697
rect 659418 75695 659441 75697
rect 659527 75695 659542 75697
rect 659542 75695 659583 75697
rect 659669 75695 659722 75697
rect 659722 75695 659725 75697
rect 657823 75573 657879 75609
rect 657965 75573 658021 75609
rect 658107 75573 658163 75609
rect 658249 75573 658305 75609
rect 658391 75573 658447 75609
rect 658533 75573 658589 75609
rect 658675 75573 658731 75609
rect 658817 75573 658873 75609
rect 658959 75573 659015 75609
rect 659101 75573 659157 75609
rect 659243 75573 659299 75609
rect 659385 75573 659441 75609
rect 659527 75573 659583 75609
rect 659669 75573 659725 75609
rect 657823 75553 657862 75573
rect 657862 75553 657879 75573
rect 657965 75553 657986 75573
rect 657986 75553 658021 75573
rect 658107 75553 658110 75573
rect 658110 75553 658163 75573
rect 658249 75553 658302 75573
rect 658302 75553 658305 75573
rect 658391 75553 658426 75573
rect 658426 75553 658447 75573
rect 658533 75553 658550 75573
rect 658550 75553 658589 75573
rect 658675 75553 658730 75573
rect 658730 75553 658731 75573
rect 658817 75553 658854 75573
rect 658854 75553 658873 75573
rect 658959 75553 658978 75573
rect 658978 75553 659015 75573
rect 659101 75553 659102 75573
rect 659102 75553 659157 75573
rect 659243 75553 659294 75573
rect 659294 75553 659299 75573
rect 659385 75553 659418 75573
rect 659418 75553 659441 75573
rect 659527 75553 659542 75573
rect 659542 75553 659583 75573
rect 659669 75553 659722 75573
rect 659722 75553 659725 75573
rect 657823 75449 657879 75467
rect 657965 75449 658021 75467
rect 658107 75449 658163 75467
rect 658249 75449 658305 75467
rect 658391 75449 658447 75467
rect 658533 75449 658589 75467
rect 658675 75449 658731 75467
rect 658817 75449 658873 75467
rect 658959 75449 659015 75467
rect 659101 75449 659157 75467
rect 659243 75449 659299 75467
rect 659385 75449 659441 75467
rect 659527 75449 659583 75467
rect 659669 75449 659725 75467
rect 657823 75411 657862 75449
rect 657862 75411 657879 75449
rect 657965 75411 657986 75449
rect 657986 75411 658021 75449
rect 658107 75411 658110 75449
rect 658110 75411 658163 75449
rect 658249 75411 658302 75449
rect 658302 75411 658305 75449
rect 658391 75411 658426 75449
rect 658426 75411 658447 75449
rect 658533 75411 658550 75449
rect 658550 75411 658589 75449
rect 658675 75411 658730 75449
rect 658730 75411 658731 75449
rect 658817 75411 658854 75449
rect 658854 75411 658873 75449
rect 658959 75411 658978 75449
rect 658978 75411 659015 75449
rect 659101 75411 659102 75449
rect 659102 75411 659157 75449
rect 659243 75411 659294 75449
rect 659294 75411 659299 75449
rect 659385 75411 659418 75449
rect 659418 75411 659441 75449
rect 659527 75411 659542 75449
rect 659542 75411 659583 75449
rect 659669 75411 659722 75449
rect 659722 75411 659725 75449
rect 657823 75269 657862 75325
rect 657862 75269 657879 75325
rect 657965 75269 657986 75325
rect 657986 75269 658021 75325
rect 658107 75269 658110 75325
rect 658110 75269 658163 75325
rect 658249 75269 658302 75325
rect 658302 75269 658305 75325
rect 658391 75269 658426 75325
rect 658426 75269 658447 75325
rect 658533 75269 658550 75325
rect 658550 75269 658589 75325
rect 658675 75269 658730 75325
rect 658730 75269 658731 75325
rect 658817 75269 658854 75325
rect 658854 75269 658873 75325
rect 658959 75269 658978 75325
rect 658978 75269 659015 75325
rect 659101 75269 659102 75325
rect 659102 75269 659157 75325
rect 659243 75269 659294 75325
rect 659294 75269 659299 75325
rect 659385 75269 659418 75325
rect 659418 75269 659441 75325
rect 659527 75269 659542 75325
rect 659542 75269 659583 75325
rect 659669 75269 659722 75325
rect 659722 75269 659725 75325
rect 657823 75145 657862 75183
rect 657862 75145 657879 75183
rect 657965 75145 657986 75183
rect 657986 75145 658021 75183
rect 658107 75145 658110 75183
rect 658110 75145 658163 75183
rect 658249 75145 658302 75183
rect 658302 75145 658305 75183
rect 658391 75145 658426 75183
rect 658426 75145 658447 75183
rect 658533 75145 658550 75183
rect 658550 75145 658589 75183
rect 658675 75145 658730 75183
rect 658730 75145 658731 75183
rect 658817 75145 658854 75183
rect 658854 75145 658873 75183
rect 658959 75145 658978 75183
rect 658978 75145 659015 75183
rect 659101 75145 659102 75183
rect 659102 75145 659157 75183
rect 659243 75145 659294 75183
rect 659294 75145 659299 75183
rect 659385 75145 659418 75183
rect 659418 75145 659441 75183
rect 659527 75145 659542 75183
rect 659542 75145 659583 75183
rect 659669 75145 659722 75183
rect 659722 75145 659725 75183
rect 657823 75127 657879 75145
rect 657965 75127 658021 75145
rect 658107 75127 658163 75145
rect 658249 75127 658305 75145
rect 658391 75127 658447 75145
rect 658533 75127 658589 75145
rect 658675 75127 658731 75145
rect 658817 75127 658873 75145
rect 658959 75127 659015 75145
rect 659101 75127 659157 75145
rect 659243 75127 659299 75145
rect 659385 75127 659441 75145
rect 659527 75127 659583 75145
rect 659669 75127 659725 75145
rect 657823 75021 657862 75041
rect 657862 75021 657879 75041
rect 657965 75021 657986 75041
rect 657986 75021 658021 75041
rect 658107 75021 658110 75041
rect 658110 75021 658163 75041
rect 658249 75021 658302 75041
rect 658302 75021 658305 75041
rect 658391 75021 658426 75041
rect 658426 75021 658447 75041
rect 658533 75021 658550 75041
rect 658550 75021 658589 75041
rect 658675 75021 658730 75041
rect 658730 75021 658731 75041
rect 658817 75021 658854 75041
rect 658854 75021 658873 75041
rect 658959 75021 658978 75041
rect 658978 75021 659015 75041
rect 659101 75021 659102 75041
rect 659102 75021 659157 75041
rect 659243 75021 659294 75041
rect 659294 75021 659299 75041
rect 659385 75021 659418 75041
rect 659418 75021 659441 75041
rect 659527 75021 659542 75041
rect 659542 75021 659583 75041
rect 659669 75021 659722 75041
rect 659722 75021 659725 75041
rect 657823 74985 657879 75021
rect 657965 74985 658021 75021
rect 658107 74985 658163 75021
rect 658249 74985 658305 75021
rect 658391 74985 658447 75021
rect 658533 74985 658589 75021
rect 658675 74985 658731 75021
rect 658817 74985 658873 75021
rect 658959 74985 659015 75021
rect 659101 74985 659157 75021
rect 659243 74985 659299 75021
rect 659385 74985 659441 75021
rect 659527 74985 659583 75021
rect 659669 74985 659725 75021
rect 657823 74897 657862 74899
rect 657862 74897 657879 74899
rect 657965 74897 657986 74899
rect 657986 74897 658021 74899
rect 658107 74897 658110 74899
rect 658110 74897 658163 74899
rect 658249 74897 658302 74899
rect 658302 74897 658305 74899
rect 658391 74897 658426 74899
rect 658426 74897 658447 74899
rect 658533 74897 658550 74899
rect 658550 74897 658589 74899
rect 658675 74897 658730 74899
rect 658730 74897 658731 74899
rect 658817 74897 658854 74899
rect 658854 74897 658873 74899
rect 658959 74897 658978 74899
rect 658978 74897 659015 74899
rect 659101 74897 659102 74899
rect 659102 74897 659157 74899
rect 659243 74897 659294 74899
rect 659294 74897 659299 74899
rect 659385 74897 659418 74899
rect 659418 74897 659441 74899
rect 659527 74897 659542 74899
rect 659542 74897 659583 74899
rect 659669 74897 659722 74899
rect 659722 74897 659725 74899
rect 657823 74843 657879 74897
rect 657965 74843 658021 74897
rect 658107 74843 658163 74897
rect 658249 74843 658305 74897
rect 658391 74843 658447 74897
rect 658533 74843 658589 74897
rect 658675 74843 658731 74897
rect 658817 74843 658873 74897
rect 658959 74843 659015 74897
rect 659101 74843 659157 74897
rect 659243 74843 659299 74897
rect 659385 74843 659441 74897
rect 659527 74843 659583 74897
rect 659669 74843 659725 74897
rect 657823 74705 657879 74757
rect 657965 74705 658021 74757
rect 658107 74705 658163 74757
rect 658249 74705 658305 74757
rect 658391 74705 658447 74757
rect 658533 74705 658589 74757
rect 658675 74705 658731 74757
rect 658817 74705 658873 74757
rect 658959 74705 659015 74757
rect 659101 74705 659157 74757
rect 659243 74705 659299 74757
rect 659385 74705 659441 74757
rect 659527 74705 659583 74757
rect 659669 74705 659725 74757
rect 657823 74701 657862 74705
rect 657862 74701 657879 74705
rect 657965 74701 657986 74705
rect 657986 74701 658021 74705
rect 658107 74701 658110 74705
rect 658110 74701 658163 74705
rect 658249 74701 658302 74705
rect 658302 74701 658305 74705
rect 658391 74701 658426 74705
rect 658426 74701 658447 74705
rect 658533 74701 658550 74705
rect 658550 74701 658589 74705
rect 658675 74701 658730 74705
rect 658730 74701 658731 74705
rect 658817 74701 658854 74705
rect 658854 74701 658873 74705
rect 658959 74701 658978 74705
rect 658978 74701 659015 74705
rect 659101 74701 659102 74705
rect 659102 74701 659157 74705
rect 659243 74701 659294 74705
rect 659294 74701 659299 74705
rect 659385 74701 659418 74705
rect 659418 74701 659441 74705
rect 659527 74701 659542 74705
rect 659542 74701 659583 74705
rect 659669 74701 659722 74705
rect 659722 74701 659725 74705
rect 657823 74581 657879 74615
rect 657965 74581 658021 74615
rect 658107 74581 658163 74615
rect 658249 74581 658305 74615
rect 658391 74581 658447 74615
rect 658533 74581 658589 74615
rect 658675 74581 658731 74615
rect 658817 74581 658873 74615
rect 658959 74581 659015 74615
rect 659101 74581 659157 74615
rect 659243 74581 659299 74615
rect 659385 74581 659441 74615
rect 659527 74581 659583 74615
rect 659669 74581 659725 74615
rect 657823 74559 657862 74581
rect 657862 74559 657879 74581
rect 657965 74559 657986 74581
rect 657986 74559 658021 74581
rect 658107 74559 658110 74581
rect 658110 74559 658163 74581
rect 658249 74559 658302 74581
rect 658302 74559 658305 74581
rect 658391 74559 658426 74581
rect 658426 74559 658447 74581
rect 658533 74559 658550 74581
rect 658550 74559 658589 74581
rect 658675 74559 658730 74581
rect 658730 74559 658731 74581
rect 658817 74559 658854 74581
rect 658854 74559 658873 74581
rect 658959 74559 658978 74581
rect 658978 74559 659015 74581
rect 659101 74559 659102 74581
rect 659102 74559 659157 74581
rect 659243 74559 659294 74581
rect 659294 74559 659299 74581
rect 659385 74559 659418 74581
rect 659418 74559 659441 74581
rect 659527 74559 659542 74581
rect 659542 74559 659583 74581
rect 659669 74559 659722 74581
rect 659722 74559 659725 74581
rect 660193 75979 660249 76035
rect 660335 75979 660391 76035
rect 660477 75979 660533 76035
rect 660619 75979 660675 76035
rect 660761 75979 660817 76035
rect 660903 75979 660959 76035
rect 661045 75979 661101 76035
rect 661187 75979 661243 76035
rect 661329 75979 661385 76035
rect 661471 75979 661527 76035
rect 661613 75979 661669 76035
rect 661755 75979 661811 76035
rect 661897 75979 661953 76035
rect 662039 75979 662095 76035
rect 660193 75889 660232 75893
rect 660232 75889 660249 75893
rect 660335 75889 660356 75893
rect 660356 75889 660391 75893
rect 660477 75889 660480 75893
rect 660480 75889 660533 75893
rect 660619 75889 660672 75893
rect 660672 75889 660675 75893
rect 660761 75889 660796 75893
rect 660796 75889 660817 75893
rect 660903 75889 660920 75893
rect 660920 75889 660959 75893
rect 661045 75889 661100 75893
rect 661100 75889 661101 75893
rect 661187 75889 661224 75893
rect 661224 75889 661243 75893
rect 661329 75889 661348 75893
rect 661348 75889 661385 75893
rect 661471 75889 661472 75893
rect 661472 75889 661527 75893
rect 661613 75889 661664 75893
rect 661664 75889 661669 75893
rect 661755 75889 661788 75893
rect 661788 75889 661811 75893
rect 661897 75889 661912 75893
rect 661912 75889 661953 75893
rect 662039 75889 662092 75893
rect 662092 75889 662095 75893
rect 660193 75837 660249 75889
rect 660335 75837 660391 75889
rect 660477 75837 660533 75889
rect 660619 75837 660675 75889
rect 660761 75837 660817 75889
rect 660903 75837 660959 75889
rect 661045 75837 661101 75889
rect 661187 75837 661243 75889
rect 661329 75837 661385 75889
rect 661471 75837 661527 75889
rect 661613 75837 661669 75889
rect 661755 75837 661811 75889
rect 661897 75837 661953 75889
rect 662039 75837 662095 75889
rect 660193 75697 660249 75751
rect 660335 75697 660391 75751
rect 660477 75697 660533 75751
rect 660619 75697 660675 75751
rect 660761 75697 660817 75751
rect 660903 75697 660959 75751
rect 661045 75697 661101 75751
rect 661187 75697 661243 75751
rect 661329 75697 661385 75751
rect 661471 75697 661527 75751
rect 661613 75697 661669 75751
rect 661755 75697 661811 75751
rect 661897 75697 661953 75751
rect 662039 75697 662095 75751
rect 660193 75695 660232 75697
rect 660232 75695 660249 75697
rect 660335 75695 660356 75697
rect 660356 75695 660391 75697
rect 660477 75695 660480 75697
rect 660480 75695 660533 75697
rect 660619 75695 660672 75697
rect 660672 75695 660675 75697
rect 660761 75695 660796 75697
rect 660796 75695 660817 75697
rect 660903 75695 660920 75697
rect 660920 75695 660959 75697
rect 661045 75695 661100 75697
rect 661100 75695 661101 75697
rect 661187 75695 661224 75697
rect 661224 75695 661243 75697
rect 661329 75695 661348 75697
rect 661348 75695 661385 75697
rect 661471 75695 661472 75697
rect 661472 75695 661527 75697
rect 661613 75695 661664 75697
rect 661664 75695 661669 75697
rect 661755 75695 661788 75697
rect 661788 75695 661811 75697
rect 661897 75695 661912 75697
rect 661912 75695 661953 75697
rect 662039 75695 662092 75697
rect 662092 75695 662095 75697
rect 660193 75573 660249 75609
rect 660335 75573 660391 75609
rect 660477 75573 660533 75609
rect 660619 75573 660675 75609
rect 660761 75573 660817 75609
rect 660903 75573 660959 75609
rect 661045 75573 661101 75609
rect 661187 75573 661243 75609
rect 661329 75573 661385 75609
rect 661471 75573 661527 75609
rect 661613 75573 661669 75609
rect 661755 75573 661811 75609
rect 661897 75573 661953 75609
rect 662039 75573 662095 75609
rect 660193 75553 660232 75573
rect 660232 75553 660249 75573
rect 660335 75553 660356 75573
rect 660356 75553 660391 75573
rect 660477 75553 660480 75573
rect 660480 75553 660533 75573
rect 660619 75553 660672 75573
rect 660672 75553 660675 75573
rect 660761 75553 660796 75573
rect 660796 75553 660817 75573
rect 660903 75553 660920 75573
rect 660920 75553 660959 75573
rect 661045 75553 661100 75573
rect 661100 75553 661101 75573
rect 661187 75553 661224 75573
rect 661224 75553 661243 75573
rect 661329 75553 661348 75573
rect 661348 75553 661385 75573
rect 661471 75553 661472 75573
rect 661472 75553 661527 75573
rect 661613 75553 661664 75573
rect 661664 75553 661669 75573
rect 661755 75553 661788 75573
rect 661788 75553 661811 75573
rect 661897 75553 661912 75573
rect 661912 75553 661953 75573
rect 662039 75553 662092 75573
rect 662092 75553 662095 75573
rect 660193 75449 660249 75467
rect 660335 75449 660391 75467
rect 660477 75449 660533 75467
rect 660619 75449 660675 75467
rect 660761 75449 660817 75467
rect 660903 75449 660959 75467
rect 661045 75449 661101 75467
rect 661187 75449 661243 75467
rect 661329 75449 661385 75467
rect 661471 75449 661527 75467
rect 661613 75449 661669 75467
rect 661755 75449 661811 75467
rect 661897 75449 661953 75467
rect 662039 75449 662095 75467
rect 660193 75411 660232 75449
rect 660232 75411 660249 75449
rect 660335 75411 660356 75449
rect 660356 75411 660391 75449
rect 660477 75411 660480 75449
rect 660480 75411 660533 75449
rect 660619 75411 660672 75449
rect 660672 75411 660675 75449
rect 660761 75411 660796 75449
rect 660796 75411 660817 75449
rect 660903 75411 660920 75449
rect 660920 75411 660959 75449
rect 661045 75411 661100 75449
rect 661100 75411 661101 75449
rect 661187 75411 661224 75449
rect 661224 75411 661243 75449
rect 661329 75411 661348 75449
rect 661348 75411 661385 75449
rect 661471 75411 661472 75449
rect 661472 75411 661527 75449
rect 661613 75411 661664 75449
rect 661664 75411 661669 75449
rect 661755 75411 661788 75449
rect 661788 75411 661811 75449
rect 661897 75411 661912 75449
rect 661912 75411 661953 75449
rect 662039 75411 662092 75449
rect 662092 75411 662095 75449
rect 660193 75269 660232 75325
rect 660232 75269 660249 75325
rect 660335 75269 660356 75325
rect 660356 75269 660391 75325
rect 660477 75269 660480 75325
rect 660480 75269 660533 75325
rect 660619 75269 660672 75325
rect 660672 75269 660675 75325
rect 660761 75269 660796 75325
rect 660796 75269 660817 75325
rect 660903 75269 660920 75325
rect 660920 75269 660959 75325
rect 661045 75269 661100 75325
rect 661100 75269 661101 75325
rect 661187 75269 661224 75325
rect 661224 75269 661243 75325
rect 661329 75269 661348 75325
rect 661348 75269 661385 75325
rect 661471 75269 661472 75325
rect 661472 75269 661527 75325
rect 661613 75269 661664 75325
rect 661664 75269 661669 75325
rect 661755 75269 661788 75325
rect 661788 75269 661811 75325
rect 661897 75269 661912 75325
rect 661912 75269 661953 75325
rect 662039 75269 662092 75325
rect 662092 75269 662095 75325
rect 660193 75145 660232 75183
rect 660232 75145 660249 75183
rect 660335 75145 660356 75183
rect 660356 75145 660391 75183
rect 660477 75145 660480 75183
rect 660480 75145 660533 75183
rect 660619 75145 660672 75183
rect 660672 75145 660675 75183
rect 660761 75145 660796 75183
rect 660796 75145 660817 75183
rect 660903 75145 660920 75183
rect 660920 75145 660959 75183
rect 661045 75145 661100 75183
rect 661100 75145 661101 75183
rect 661187 75145 661224 75183
rect 661224 75145 661243 75183
rect 661329 75145 661348 75183
rect 661348 75145 661385 75183
rect 661471 75145 661472 75183
rect 661472 75145 661527 75183
rect 661613 75145 661664 75183
rect 661664 75145 661669 75183
rect 661755 75145 661788 75183
rect 661788 75145 661811 75183
rect 661897 75145 661912 75183
rect 661912 75145 661953 75183
rect 662039 75145 662092 75183
rect 662092 75145 662095 75183
rect 660193 75127 660249 75145
rect 660335 75127 660391 75145
rect 660477 75127 660533 75145
rect 660619 75127 660675 75145
rect 660761 75127 660817 75145
rect 660903 75127 660959 75145
rect 661045 75127 661101 75145
rect 661187 75127 661243 75145
rect 661329 75127 661385 75145
rect 661471 75127 661527 75145
rect 661613 75127 661669 75145
rect 661755 75127 661811 75145
rect 661897 75127 661953 75145
rect 662039 75127 662095 75145
rect 660193 75021 660232 75041
rect 660232 75021 660249 75041
rect 660335 75021 660356 75041
rect 660356 75021 660391 75041
rect 660477 75021 660480 75041
rect 660480 75021 660533 75041
rect 660619 75021 660672 75041
rect 660672 75021 660675 75041
rect 660761 75021 660796 75041
rect 660796 75021 660817 75041
rect 660903 75021 660920 75041
rect 660920 75021 660959 75041
rect 661045 75021 661100 75041
rect 661100 75021 661101 75041
rect 661187 75021 661224 75041
rect 661224 75021 661243 75041
rect 661329 75021 661348 75041
rect 661348 75021 661385 75041
rect 661471 75021 661472 75041
rect 661472 75021 661527 75041
rect 661613 75021 661664 75041
rect 661664 75021 661669 75041
rect 661755 75021 661788 75041
rect 661788 75021 661811 75041
rect 661897 75021 661912 75041
rect 661912 75021 661953 75041
rect 662039 75021 662092 75041
rect 662092 75021 662095 75041
rect 660193 74985 660249 75021
rect 660335 74985 660391 75021
rect 660477 74985 660533 75021
rect 660619 74985 660675 75021
rect 660761 74985 660817 75021
rect 660903 74985 660959 75021
rect 661045 74985 661101 75021
rect 661187 74985 661243 75021
rect 661329 74985 661385 75021
rect 661471 74985 661527 75021
rect 661613 74985 661669 75021
rect 661755 74985 661811 75021
rect 661897 74985 661953 75021
rect 662039 74985 662095 75021
rect 660193 74897 660232 74899
rect 660232 74897 660249 74899
rect 660335 74897 660356 74899
rect 660356 74897 660391 74899
rect 660477 74897 660480 74899
rect 660480 74897 660533 74899
rect 660619 74897 660672 74899
rect 660672 74897 660675 74899
rect 660761 74897 660796 74899
rect 660796 74897 660817 74899
rect 660903 74897 660920 74899
rect 660920 74897 660959 74899
rect 661045 74897 661100 74899
rect 661100 74897 661101 74899
rect 661187 74897 661224 74899
rect 661224 74897 661243 74899
rect 661329 74897 661348 74899
rect 661348 74897 661385 74899
rect 661471 74897 661472 74899
rect 661472 74897 661527 74899
rect 661613 74897 661664 74899
rect 661664 74897 661669 74899
rect 661755 74897 661788 74899
rect 661788 74897 661811 74899
rect 661897 74897 661912 74899
rect 661912 74897 661953 74899
rect 662039 74897 662092 74899
rect 662092 74897 662095 74899
rect 660193 74843 660249 74897
rect 660335 74843 660391 74897
rect 660477 74843 660533 74897
rect 660619 74843 660675 74897
rect 660761 74843 660817 74897
rect 660903 74843 660959 74897
rect 661045 74843 661101 74897
rect 661187 74843 661243 74897
rect 661329 74843 661385 74897
rect 661471 74843 661527 74897
rect 661613 74843 661669 74897
rect 661755 74843 661811 74897
rect 661897 74843 661953 74897
rect 662039 74843 662095 74897
rect 660193 74705 660249 74757
rect 660335 74705 660391 74757
rect 660477 74705 660533 74757
rect 660619 74705 660675 74757
rect 660761 74705 660817 74757
rect 660903 74705 660959 74757
rect 661045 74705 661101 74757
rect 661187 74705 661243 74757
rect 661329 74705 661385 74757
rect 661471 74705 661527 74757
rect 661613 74705 661669 74757
rect 661755 74705 661811 74757
rect 661897 74705 661953 74757
rect 662039 74705 662095 74757
rect 660193 74701 660232 74705
rect 660232 74701 660249 74705
rect 660335 74701 660356 74705
rect 660356 74701 660391 74705
rect 660477 74701 660480 74705
rect 660480 74701 660533 74705
rect 660619 74701 660672 74705
rect 660672 74701 660675 74705
rect 660761 74701 660796 74705
rect 660796 74701 660817 74705
rect 660903 74701 660920 74705
rect 660920 74701 660959 74705
rect 661045 74701 661100 74705
rect 661100 74701 661101 74705
rect 661187 74701 661224 74705
rect 661224 74701 661243 74705
rect 661329 74701 661348 74705
rect 661348 74701 661385 74705
rect 661471 74701 661472 74705
rect 661472 74701 661527 74705
rect 661613 74701 661664 74705
rect 661664 74701 661669 74705
rect 661755 74701 661788 74705
rect 661788 74701 661811 74705
rect 661897 74701 661912 74705
rect 661912 74701 661953 74705
rect 662039 74701 662092 74705
rect 662092 74701 662095 74705
rect 660193 74581 660249 74615
rect 660335 74581 660391 74615
rect 660477 74581 660533 74615
rect 660619 74581 660675 74615
rect 660761 74581 660817 74615
rect 660903 74581 660959 74615
rect 661045 74581 661101 74615
rect 661187 74581 661243 74615
rect 661329 74581 661385 74615
rect 661471 74581 661527 74615
rect 661613 74581 661669 74615
rect 661755 74581 661811 74615
rect 661897 74581 661953 74615
rect 662039 74581 662095 74615
rect 660193 74559 660232 74581
rect 660232 74559 660249 74581
rect 660335 74559 660356 74581
rect 660356 74559 660391 74581
rect 660477 74559 660480 74581
rect 660480 74559 660533 74581
rect 660619 74559 660672 74581
rect 660672 74559 660675 74581
rect 660761 74559 660796 74581
rect 660796 74559 660817 74581
rect 660903 74559 660920 74581
rect 660920 74559 660959 74581
rect 661045 74559 661100 74581
rect 661100 74559 661101 74581
rect 661187 74559 661224 74581
rect 661224 74559 661243 74581
rect 661329 74559 661348 74581
rect 661348 74559 661385 74581
rect 661471 74559 661472 74581
rect 661472 74559 661527 74581
rect 661613 74559 661664 74581
rect 661664 74559 661669 74581
rect 661755 74559 661788 74581
rect 661788 74559 661811 74581
rect 661897 74559 661912 74581
rect 661912 74559 661953 74581
rect 662039 74559 662092 74581
rect 662092 74559 662095 74581
rect 662899 75979 662955 76035
rect 663041 75979 663097 76035
rect 663183 75979 663239 76035
rect 663325 75979 663381 76035
rect 663467 75979 663523 76035
rect 663609 75979 663665 76035
rect 663751 75979 663807 76035
rect 663893 75979 663949 76035
rect 664035 75979 664091 76035
rect 664177 75979 664233 76035
rect 664319 75979 664375 76035
rect 664461 75979 664517 76035
rect 664603 75979 664659 76035
rect 664745 75979 664801 76035
rect 662899 75889 662938 75893
rect 662938 75889 662955 75893
rect 663041 75889 663062 75893
rect 663062 75889 663097 75893
rect 663183 75889 663186 75893
rect 663186 75889 663239 75893
rect 663325 75889 663378 75893
rect 663378 75889 663381 75893
rect 663467 75889 663502 75893
rect 663502 75889 663523 75893
rect 663609 75889 663626 75893
rect 663626 75889 663665 75893
rect 663751 75889 663806 75893
rect 663806 75889 663807 75893
rect 663893 75889 663930 75893
rect 663930 75889 663949 75893
rect 664035 75889 664054 75893
rect 664054 75889 664091 75893
rect 664177 75889 664178 75893
rect 664178 75889 664233 75893
rect 664319 75889 664370 75893
rect 664370 75889 664375 75893
rect 664461 75889 664494 75893
rect 664494 75889 664517 75893
rect 664603 75889 664618 75893
rect 664618 75889 664659 75893
rect 664745 75889 664798 75893
rect 664798 75889 664801 75893
rect 662899 75837 662955 75889
rect 663041 75837 663097 75889
rect 663183 75837 663239 75889
rect 663325 75837 663381 75889
rect 663467 75837 663523 75889
rect 663609 75837 663665 75889
rect 663751 75837 663807 75889
rect 663893 75837 663949 75889
rect 664035 75837 664091 75889
rect 664177 75837 664233 75889
rect 664319 75837 664375 75889
rect 664461 75837 664517 75889
rect 664603 75837 664659 75889
rect 664745 75837 664801 75889
rect 662899 75697 662955 75751
rect 663041 75697 663097 75751
rect 663183 75697 663239 75751
rect 663325 75697 663381 75751
rect 663467 75697 663523 75751
rect 663609 75697 663665 75751
rect 663751 75697 663807 75751
rect 663893 75697 663949 75751
rect 664035 75697 664091 75751
rect 664177 75697 664233 75751
rect 664319 75697 664375 75751
rect 664461 75697 664517 75751
rect 664603 75697 664659 75751
rect 664745 75697 664801 75751
rect 662899 75695 662938 75697
rect 662938 75695 662955 75697
rect 663041 75695 663062 75697
rect 663062 75695 663097 75697
rect 663183 75695 663186 75697
rect 663186 75695 663239 75697
rect 663325 75695 663378 75697
rect 663378 75695 663381 75697
rect 663467 75695 663502 75697
rect 663502 75695 663523 75697
rect 663609 75695 663626 75697
rect 663626 75695 663665 75697
rect 663751 75695 663806 75697
rect 663806 75695 663807 75697
rect 663893 75695 663930 75697
rect 663930 75695 663949 75697
rect 664035 75695 664054 75697
rect 664054 75695 664091 75697
rect 664177 75695 664178 75697
rect 664178 75695 664233 75697
rect 664319 75695 664370 75697
rect 664370 75695 664375 75697
rect 664461 75695 664494 75697
rect 664494 75695 664517 75697
rect 664603 75695 664618 75697
rect 664618 75695 664659 75697
rect 664745 75695 664798 75697
rect 664798 75695 664801 75697
rect 662899 75573 662955 75609
rect 663041 75573 663097 75609
rect 663183 75573 663239 75609
rect 663325 75573 663381 75609
rect 663467 75573 663523 75609
rect 663609 75573 663665 75609
rect 663751 75573 663807 75609
rect 663893 75573 663949 75609
rect 664035 75573 664091 75609
rect 664177 75573 664233 75609
rect 664319 75573 664375 75609
rect 664461 75573 664517 75609
rect 664603 75573 664659 75609
rect 664745 75573 664801 75609
rect 662899 75553 662938 75573
rect 662938 75553 662955 75573
rect 663041 75553 663062 75573
rect 663062 75553 663097 75573
rect 663183 75553 663186 75573
rect 663186 75553 663239 75573
rect 663325 75553 663378 75573
rect 663378 75553 663381 75573
rect 663467 75553 663502 75573
rect 663502 75553 663523 75573
rect 663609 75553 663626 75573
rect 663626 75553 663665 75573
rect 663751 75553 663806 75573
rect 663806 75553 663807 75573
rect 663893 75553 663930 75573
rect 663930 75553 663949 75573
rect 664035 75553 664054 75573
rect 664054 75553 664091 75573
rect 664177 75553 664178 75573
rect 664178 75553 664233 75573
rect 664319 75553 664370 75573
rect 664370 75553 664375 75573
rect 664461 75553 664494 75573
rect 664494 75553 664517 75573
rect 664603 75553 664618 75573
rect 664618 75553 664659 75573
rect 664745 75553 664798 75573
rect 664798 75553 664801 75573
rect 662899 75449 662955 75467
rect 663041 75449 663097 75467
rect 663183 75449 663239 75467
rect 663325 75449 663381 75467
rect 663467 75449 663523 75467
rect 663609 75449 663665 75467
rect 663751 75449 663807 75467
rect 663893 75449 663949 75467
rect 664035 75449 664091 75467
rect 664177 75449 664233 75467
rect 664319 75449 664375 75467
rect 664461 75449 664517 75467
rect 664603 75449 664659 75467
rect 664745 75449 664801 75467
rect 662899 75411 662938 75449
rect 662938 75411 662955 75449
rect 663041 75411 663062 75449
rect 663062 75411 663097 75449
rect 663183 75411 663186 75449
rect 663186 75411 663239 75449
rect 663325 75411 663378 75449
rect 663378 75411 663381 75449
rect 663467 75411 663502 75449
rect 663502 75411 663523 75449
rect 663609 75411 663626 75449
rect 663626 75411 663665 75449
rect 663751 75411 663806 75449
rect 663806 75411 663807 75449
rect 663893 75411 663930 75449
rect 663930 75411 663949 75449
rect 664035 75411 664054 75449
rect 664054 75411 664091 75449
rect 664177 75411 664178 75449
rect 664178 75411 664233 75449
rect 664319 75411 664370 75449
rect 664370 75411 664375 75449
rect 664461 75411 664494 75449
rect 664494 75411 664517 75449
rect 664603 75411 664618 75449
rect 664618 75411 664659 75449
rect 664745 75411 664798 75449
rect 664798 75411 664801 75449
rect 662899 75269 662938 75325
rect 662938 75269 662955 75325
rect 663041 75269 663062 75325
rect 663062 75269 663097 75325
rect 663183 75269 663186 75325
rect 663186 75269 663239 75325
rect 663325 75269 663378 75325
rect 663378 75269 663381 75325
rect 663467 75269 663502 75325
rect 663502 75269 663523 75325
rect 663609 75269 663626 75325
rect 663626 75269 663665 75325
rect 663751 75269 663806 75325
rect 663806 75269 663807 75325
rect 663893 75269 663930 75325
rect 663930 75269 663949 75325
rect 664035 75269 664054 75325
rect 664054 75269 664091 75325
rect 664177 75269 664178 75325
rect 664178 75269 664233 75325
rect 664319 75269 664370 75325
rect 664370 75269 664375 75325
rect 664461 75269 664494 75325
rect 664494 75269 664517 75325
rect 664603 75269 664618 75325
rect 664618 75269 664659 75325
rect 664745 75269 664798 75325
rect 664798 75269 664801 75325
rect 662899 75145 662938 75183
rect 662938 75145 662955 75183
rect 663041 75145 663062 75183
rect 663062 75145 663097 75183
rect 663183 75145 663186 75183
rect 663186 75145 663239 75183
rect 663325 75145 663378 75183
rect 663378 75145 663381 75183
rect 663467 75145 663502 75183
rect 663502 75145 663523 75183
rect 663609 75145 663626 75183
rect 663626 75145 663665 75183
rect 663751 75145 663806 75183
rect 663806 75145 663807 75183
rect 663893 75145 663930 75183
rect 663930 75145 663949 75183
rect 664035 75145 664054 75183
rect 664054 75145 664091 75183
rect 664177 75145 664178 75183
rect 664178 75145 664233 75183
rect 664319 75145 664370 75183
rect 664370 75145 664375 75183
rect 664461 75145 664494 75183
rect 664494 75145 664517 75183
rect 664603 75145 664618 75183
rect 664618 75145 664659 75183
rect 664745 75145 664798 75183
rect 664798 75145 664801 75183
rect 662899 75127 662955 75145
rect 663041 75127 663097 75145
rect 663183 75127 663239 75145
rect 663325 75127 663381 75145
rect 663467 75127 663523 75145
rect 663609 75127 663665 75145
rect 663751 75127 663807 75145
rect 663893 75127 663949 75145
rect 664035 75127 664091 75145
rect 664177 75127 664233 75145
rect 664319 75127 664375 75145
rect 664461 75127 664517 75145
rect 664603 75127 664659 75145
rect 664745 75127 664801 75145
rect 662899 75021 662938 75041
rect 662938 75021 662955 75041
rect 663041 75021 663062 75041
rect 663062 75021 663097 75041
rect 663183 75021 663186 75041
rect 663186 75021 663239 75041
rect 663325 75021 663378 75041
rect 663378 75021 663381 75041
rect 663467 75021 663502 75041
rect 663502 75021 663523 75041
rect 663609 75021 663626 75041
rect 663626 75021 663665 75041
rect 663751 75021 663806 75041
rect 663806 75021 663807 75041
rect 663893 75021 663930 75041
rect 663930 75021 663949 75041
rect 664035 75021 664054 75041
rect 664054 75021 664091 75041
rect 664177 75021 664178 75041
rect 664178 75021 664233 75041
rect 664319 75021 664370 75041
rect 664370 75021 664375 75041
rect 664461 75021 664494 75041
rect 664494 75021 664517 75041
rect 664603 75021 664618 75041
rect 664618 75021 664659 75041
rect 664745 75021 664798 75041
rect 664798 75021 664801 75041
rect 662899 74985 662955 75021
rect 663041 74985 663097 75021
rect 663183 74985 663239 75021
rect 663325 74985 663381 75021
rect 663467 74985 663523 75021
rect 663609 74985 663665 75021
rect 663751 74985 663807 75021
rect 663893 74985 663949 75021
rect 664035 74985 664091 75021
rect 664177 74985 664233 75021
rect 664319 74985 664375 75021
rect 664461 74985 664517 75021
rect 664603 74985 664659 75021
rect 664745 74985 664801 75021
rect 662899 74897 662938 74899
rect 662938 74897 662955 74899
rect 663041 74897 663062 74899
rect 663062 74897 663097 74899
rect 663183 74897 663186 74899
rect 663186 74897 663239 74899
rect 663325 74897 663378 74899
rect 663378 74897 663381 74899
rect 663467 74897 663502 74899
rect 663502 74897 663523 74899
rect 663609 74897 663626 74899
rect 663626 74897 663665 74899
rect 663751 74897 663806 74899
rect 663806 74897 663807 74899
rect 663893 74897 663930 74899
rect 663930 74897 663949 74899
rect 664035 74897 664054 74899
rect 664054 74897 664091 74899
rect 664177 74897 664178 74899
rect 664178 74897 664233 74899
rect 664319 74897 664370 74899
rect 664370 74897 664375 74899
rect 664461 74897 664494 74899
rect 664494 74897 664517 74899
rect 664603 74897 664618 74899
rect 664618 74897 664659 74899
rect 664745 74897 664798 74899
rect 664798 74897 664801 74899
rect 662899 74843 662955 74897
rect 663041 74843 663097 74897
rect 663183 74843 663239 74897
rect 663325 74843 663381 74897
rect 663467 74843 663523 74897
rect 663609 74843 663665 74897
rect 663751 74843 663807 74897
rect 663893 74843 663949 74897
rect 664035 74843 664091 74897
rect 664177 74843 664233 74897
rect 664319 74843 664375 74897
rect 664461 74843 664517 74897
rect 664603 74843 664659 74897
rect 664745 74843 664801 74897
rect 662899 74705 662955 74757
rect 663041 74705 663097 74757
rect 663183 74705 663239 74757
rect 663325 74705 663381 74757
rect 663467 74705 663523 74757
rect 663609 74705 663665 74757
rect 663751 74705 663807 74757
rect 663893 74705 663949 74757
rect 664035 74705 664091 74757
rect 664177 74705 664233 74757
rect 664319 74705 664375 74757
rect 664461 74705 664517 74757
rect 664603 74705 664659 74757
rect 664745 74705 664801 74757
rect 662899 74701 662938 74705
rect 662938 74701 662955 74705
rect 663041 74701 663062 74705
rect 663062 74701 663097 74705
rect 663183 74701 663186 74705
rect 663186 74701 663239 74705
rect 663325 74701 663378 74705
rect 663378 74701 663381 74705
rect 663467 74701 663502 74705
rect 663502 74701 663523 74705
rect 663609 74701 663626 74705
rect 663626 74701 663665 74705
rect 663751 74701 663806 74705
rect 663806 74701 663807 74705
rect 663893 74701 663930 74705
rect 663930 74701 663949 74705
rect 664035 74701 664054 74705
rect 664054 74701 664091 74705
rect 664177 74701 664178 74705
rect 664178 74701 664233 74705
rect 664319 74701 664370 74705
rect 664370 74701 664375 74705
rect 664461 74701 664494 74705
rect 664494 74701 664517 74705
rect 664603 74701 664618 74705
rect 664618 74701 664659 74705
rect 664745 74701 664798 74705
rect 664798 74701 664801 74705
rect 662899 74581 662955 74615
rect 663041 74581 663097 74615
rect 663183 74581 663239 74615
rect 663325 74581 663381 74615
rect 663467 74581 663523 74615
rect 663609 74581 663665 74615
rect 663751 74581 663807 74615
rect 663893 74581 663949 74615
rect 664035 74581 664091 74615
rect 664177 74581 664233 74615
rect 664319 74581 664375 74615
rect 664461 74581 664517 74615
rect 664603 74581 664659 74615
rect 664745 74581 664801 74615
rect 662899 74559 662938 74581
rect 662938 74559 662955 74581
rect 663041 74559 663062 74581
rect 663062 74559 663097 74581
rect 663183 74559 663186 74581
rect 663186 74559 663239 74581
rect 663325 74559 663378 74581
rect 663378 74559 663381 74581
rect 663467 74559 663502 74581
rect 663502 74559 663523 74581
rect 663609 74559 663626 74581
rect 663626 74559 663665 74581
rect 663751 74559 663806 74581
rect 663806 74559 663807 74581
rect 663893 74559 663930 74581
rect 663930 74559 663949 74581
rect 664035 74559 664054 74581
rect 664054 74559 664091 74581
rect 664177 74559 664178 74581
rect 664178 74559 664233 74581
rect 664319 74559 664370 74581
rect 664370 74559 664375 74581
rect 664461 74559 664494 74581
rect 664494 74559 664517 74581
rect 664603 74559 664618 74581
rect 664618 74559 664659 74581
rect 664745 74559 664798 74581
rect 664798 74559 664801 74581
rect 665269 75979 665325 76035
rect 665411 75979 665467 76035
rect 665553 75979 665609 76035
rect 665695 75979 665751 76035
rect 665837 75979 665893 76035
rect 665979 75979 666035 76035
rect 666121 75979 666177 76035
rect 666263 75979 666319 76035
rect 666405 75979 666461 76035
rect 666547 75979 666603 76035
rect 666689 75979 666745 76035
rect 666831 75979 666887 76035
rect 666973 75979 667029 76035
rect 667115 75979 667171 76035
rect 665269 75889 665308 75893
rect 665308 75889 665325 75893
rect 665411 75889 665432 75893
rect 665432 75889 665467 75893
rect 665553 75889 665556 75893
rect 665556 75889 665609 75893
rect 665695 75889 665748 75893
rect 665748 75889 665751 75893
rect 665837 75889 665872 75893
rect 665872 75889 665893 75893
rect 665979 75889 665996 75893
rect 665996 75889 666035 75893
rect 666121 75889 666176 75893
rect 666176 75889 666177 75893
rect 666263 75889 666300 75893
rect 666300 75889 666319 75893
rect 666405 75889 666424 75893
rect 666424 75889 666461 75893
rect 666547 75889 666548 75893
rect 666548 75889 666603 75893
rect 666689 75889 666740 75893
rect 666740 75889 666745 75893
rect 666831 75889 666864 75893
rect 666864 75889 666887 75893
rect 666973 75889 666988 75893
rect 666988 75889 667029 75893
rect 667115 75889 667168 75893
rect 667168 75889 667171 75893
rect 665269 75837 665325 75889
rect 665411 75837 665467 75889
rect 665553 75837 665609 75889
rect 665695 75837 665751 75889
rect 665837 75837 665893 75889
rect 665979 75837 666035 75889
rect 666121 75837 666177 75889
rect 666263 75837 666319 75889
rect 666405 75837 666461 75889
rect 666547 75837 666603 75889
rect 666689 75837 666745 75889
rect 666831 75837 666887 75889
rect 666973 75837 667029 75889
rect 667115 75837 667171 75889
rect 665269 75697 665325 75751
rect 665411 75697 665467 75751
rect 665553 75697 665609 75751
rect 665695 75697 665751 75751
rect 665837 75697 665893 75751
rect 665979 75697 666035 75751
rect 666121 75697 666177 75751
rect 666263 75697 666319 75751
rect 666405 75697 666461 75751
rect 666547 75697 666603 75751
rect 666689 75697 666745 75751
rect 666831 75697 666887 75751
rect 666973 75697 667029 75751
rect 667115 75697 667171 75751
rect 665269 75695 665308 75697
rect 665308 75695 665325 75697
rect 665411 75695 665432 75697
rect 665432 75695 665467 75697
rect 665553 75695 665556 75697
rect 665556 75695 665609 75697
rect 665695 75695 665748 75697
rect 665748 75695 665751 75697
rect 665837 75695 665872 75697
rect 665872 75695 665893 75697
rect 665979 75695 665996 75697
rect 665996 75695 666035 75697
rect 666121 75695 666176 75697
rect 666176 75695 666177 75697
rect 666263 75695 666300 75697
rect 666300 75695 666319 75697
rect 666405 75695 666424 75697
rect 666424 75695 666461 75697
rect 666547 75695 666548 75697
rect 666548 75695 666603 75697
rect 666689 75695 666740 75697
rect 666740 75695 666745 75697
rect 666831 75695 666864 75697
rect 666864 75695 666887 75697
rect 666973 75695 666988 75697
rect 666988 75695 667029 75697
rect 667115 75695 667168 75697
rect 667168 75695 667171 75697
rect 665269 75573 665325 75609
rect 665411 75573 665467 75609
rect 665553 75573 665609 75609
rect 665695 75573 665751 75609
rect 665837 75573 665893 75609
rect 665979 75573 666035 75609
rect 666121 75573 666177 75609
rect 666263 75573 666319 75609
rect 666405 75573 666461 75609
rect 666547 75573 666603 75609
rect 666689 75573 666745 75609
rect 666831 75573 666887 75609
rect 666973 75573 667029 75609
rect 667115 75573 667171 75609
rect 665269 75553 665308 75573
rect 665308 75553 665325 75573
rect 665411 75553 665432 75573
rect 665432 75553 665467 75573
rect 665553 75553 665556 75573
rect 665556 75553 665609 75573
rect 665695 75553 665748 75573
rect 665748 75553 665751 75573
rect 665837 75553 665872 75573
rect 665872 75553 665893 75573
rect 665979 75553 665996 75573
rect 665996 75553 666035 75573
rect 666121 75553 666176 75573
rect 666176 75553 666177 75573
rect 666263 75553 666300 75573
rect 666300 75553 666319 75573
rect 666405 75553 666424 75573
rect 666424 75553 666461 75573
rect 666547 75553 666548 75573
rect 666548 75553 666603 75573
rect 666689 75553 666740 75573
rect 666740 75553 666745 75573
rect 666831 75553 666864 75573
rect 666864 75553 666887 75573
rect 666973 75553 666988 75573
rect 666988 75553 667029 75573
rect 667115 75553 667168 75573
rect 667168 75553 667171 75573
rect 665269 75449 665325 75467
rect 665411 75449 665467 75467
rect 665553 75449 665609 75467
rect 665695 75449 665751 75467
rect 665837 75449 665893 75467
rect 665979 75449 666035 75467
rect 666121 75449 666177 75467
rect 666263 75449 666319 75467
rect 666405 75449 666461 75467
rect 666547 75449 666603 75467
rect 666689 75449 666745 75467
rect 666831 75449 666887 75467
rect 666973 75449 667029 75467
rect 667115 75449 667171 75467
rect 665269 75411 665308 75449
rect 665308 75411 665325 75449
rect 665411 75411 665432 75449
rect 665432 75411 665467 75449
rect 665553 75411 665556 75449
rect 665556 75411 665609 75449
rect 665695 75411 665748 75449
rect 665748 75411 665751 75449
rect 665837 75411 665872 75449
rect 665872 75411 665893 75449
rect 665979 75411 665996 75449
rect 665996 75411 666035 75449
rect 666121 75411 666176 75449
rect 666176 75411 666177 75449
rect 666263 75411 666300 75449
rect 666300 75411 666319 75449
rect 666405 75411 666424 75449
rect 666424 75411 666461 75449
rect 666547 75411 666548 75449
rect 666548 75411 666603 75449
rect 666689 75411 666740 75449
rect 666740 75411 666745 75449
rect 666831 75411 666864 75449
rect 666864 75411 666887 75449
rect 666973 75411 666988 75449
rect 666988 75411 667029 75449
rect 667115 75411 667168 75449
rect 667168 75411 667171 75449
rect 665269 75269 665308 75325
rect 665308 75269 665325 75325
rect 665411 75269 665432 75325
rect 665432 75269 665467 75325
rect 665553 75269 665556 75325
rect 665556 75269 665609 75325
rect 665695 75269 665748 75325
rect 665748 75269 665751 75325
rect 665837 75269 665872 75325
rect 665872 75269 665893 75325
rect 665979 75269 665996 75325
rect 665996 75269 666035 75325
rect 666121 75269 666176 75325
rect 666176 75269 666177 75325
rect 666263 75269 666300 75325
rect 666300 75269 666319 75325
rect 666405 75269 666424 75325
rect 666424 75269 666461 75325
rect 666547 75269 666548 75325
rect 666548 75269 666603 75325
rect 666689 75269 666740 75325
rect 666740 75269 666745 75325
rect 666831 75269 666864 75325
rect 666864 75269 666887 75325
rect 666973 75269 666988 75325
rect 666988 75269 667029 75325
rect 667115 75269 667168 75325
rect 667168 75269 667171 75325
rect 665269 75145 665308 75183
rect 665308 75145 665325 75183
rect 665411 75145 665432 75183
rect 665432 75145 665467 75183
rect 665553 75145 665556 75183
rect 665556 75145 665609 75183
rect 665695 75145 665748 75183
rect 665748 75145 665751 75183
rect 665837 75145 665872 75183
rect 665872 75145 665893 75183
rect 665979 75145 665996 75183
rect 665996 75145 666035 75183
rect 666121 75145 666176 75183
rect 666176 75145 666177 75183
rect 666263 75145 666300 75183
rect 666300 75145 666319 75183
rect 666405 75145 666424 75183
rect 666424 75145 666461 75183
rect 666547 75145 666548 75183
rect 666548 75145 666603 75183
rect 666689 75145 666740 75183
rect 666740 75145 666745 75183
rect 666831 75145 666864 75183
rect 666864 75145 666887 75183
rect 666973 75145 666988 75183
rect 666988 75145 667029 75183
rect 667115 75145 667168 75183
rect 667168 75145 667171 75183
rect 665269 75127 665325 75145
rect 665411 75127 665467 75145
rect 665553 75127 665609 75145
rect 665695 75127 665751 75145
rect 665837 75127 665893 75145
rect 665979 75127 666035 75145
rect 666121 75127 666177 75145
rect 666263 75127 666319 75145
rect 666405 75127 666461 75145
rect 666547 75127 666603 75145
rect 666689 75127 666745 75145
rect 666831 75127 666887 75145
rect 666973 75127 667029 75145
rect 667115 75127 667171 75145
rect 665269 75021 665308 75041
rect 665308 75021 665325 75041
rect 665411 75021 665432 75041
rect 665432 75021 665467 75041
rect 665553 75021 665556 75041
rect 665556 75021 665609 75041
rect 665695 75021 665748 75041
rect 665748 75021 665751 75041
rect 665837 75021 665872 75041
rect 665872 75021 665893 75041
rect 665979 75021 665996 75041
rect 665996 75021 666035 75041
rect 666121 75021 666176 75041
rect 666176 75021 666177 75041
rect 666263 75021 666300 75041
rect 666300 75021 666319 75041
rect 666405 75021 666424 75041
rect 666424 75021 666461 75041
rect 666547 75021 666548 75041
rect 666548 75021 666603 75041
rect 666689 75021 666740 75041
rect 666740 75021 666745 75041
rect 666831 75021 666864 75041
rect 666864 75021 666887 75041
rect 666973 75021 666988 75041
rect 666988 75021 667029 75041
rect 667115 75021 667168 75041
rect 667168 75021 667171 75041
rect 665269 74985 665325 75021
rect 665411 74985 665467 75021
rect 665553 74985 665609 75021
rect 665695 74985 665751 75021
rect 665837 74985 665893 75021
rect 665979 74985 666035 75021
rect 666121 74985 666177 75021
rect 666263 74985 666319 75021
rect 666405 74985 666461 75021
rect 666547 74985 666603 75021
rect 666689 74985 666745 75021
rect 666831 74985 666887 75021
rect 666973 74985 667029 75021
rect 667115 74985 667171 75021
rect 665269 74897 665308 74899
rect 665308 74897 665325 74899
rect 665411 74897 665432 74899
rect 665432 74897 665467 74899
rect 665553 74897 665556 74899
rect 665556 74897 665609 74899
rect 665695 74897 665748 74899
rect 665748 74897 665751 74899
rect 665837 74897 665872 74899
rect 665872 74897 665893 74899
rect 665979 74897 665996 74899
rect 665996 74897 666035 74899
rect 666121 74897 666176 74899
rect 666176 74897 666177 74899
rect 666263 74897 666300 74899
rect 666300 74897 666319 74899
rect 666405 74897 666424 74899
rect 666424 74897 666461 74899
rect 666547 74897 666548 74899
rect 666548 74897 666603 74899
rect 666689 74897 666740 74899
rect 666740 74897 666745 74899
rect 666831 74897 666864 74899
rect 666864 74897 666887 74899
rect 666973 74897 666988 74899
rect 666988 74897 667029 74899
rect 667115 74897 667168 74899
rect 667168 74897 667171 74899
rect 665269 74843 665325 74897
rect 665411 74843 665467 74897
rect 665553 74843 665609 74897
rect 665695 74843 665751 74897
rect 665837 74843 665893 74897
rect 665979 74843 666035 74897
rect 666121 74843 666177 74897
rect 666263 74843 666319 74897
rect 666405 74843 666461 74897
rect 666547 74843 666603 74897
rect 666689 74843 666745 74897
rect 666831 74843 666887 74897
rect 666973 74843 667029 74897
rect 667115 74843 667171 74897
rect 665269 74705 665325 74757
rect 665411 74705 665467 74757
rect 665553 74705 665609 74757
rect 665695 74705 665751 74757
rect 665837 74705 665893 74757
rect 665979 74705 666035 74757
rect 666121 74705 666177 74757
rect 666263 74705 666319 74757
rect 666405 74705 666461 74757
rect 666547 74705 666603 74757
rect 666689 74705 666745 74757
rect 666831 74705 666887 74757
rect 666973 74705 667029 74757
rect 667115 74705 667171 74757
rect 665269 74701 665308 74705
rect 665308 74701 665325 74705
rect 665411 74701 665432 74705
rect 665432 74701 665467 74705
rect 665553 74701 665556 74705
rect 665556 74701 665609 74705
rect 665695 74701 665748 74705
rect 665748 74701 665751 74705
rect 665837 74701 665872 74705
rect 665872 74701 665893 74705
rect 665979 74701 665996 74705
rect 665996 74701 666035 74705
rect 666121 74701 666176 74705
rect 666176 74701 666177 74705
rect 666263 74701 666300 74705
rect 666300 74701 666319 74705
rect 666405 74701 666424 74705
rect 666424 74701 666461 74705
rect 666547 74701 666548 74705
rect 666548 74701 666603 74705
rect 666689 74701 666740 74705
rect 666740 74701 666745 74705
rect 666831 74701 666864 74705
rect 666864 74701 666887 74705
rect 666973 74701 666988 74705
rect 666988 74701 667029 74705
rect 667115 74701 667168 74705
rect 667168 74701 667171 74705
rect 665269 74581 665325 74615
rect 665411 74581 665467 74615
rect 665553 74581 665609 74615
rect 665695 74581 665751 74615
rect 665837 74581 665893 74615
rect 665979 74581 666035 74615
rect 666121 74581 666177 74615
rect 666263 74581 666319 74615
rect 666405 74581 666461 74615
rect 666547 74581 666603 74615
rect 666689 74581 666745 74615
rect 666831 74581 666887 74615
rect 666973 74581 667029 74615
rect 667115 74581 667171 74615
rect 665269 74559 665308 74581
rect 665308 74559 665325 74581
rect 665411 74559 665432 74581
rect 665432 74559 665467 74581
rect 665553 74559 665556 74581
rect 665556 74559 665609 74581
rect 665695 74559 665748 74581
rect 665748 74559 665751 74581
rect 665837 74559 665872 74581
rect 665872 74559 665893 74581
rect 665979 74559 665996 74581
rect 665996 74559 666035 74581
rect 666121 74559 666176 74581
rect 666176 74559 666177 74581
rect 666263 74559 666300 74581
rect 666300 74559 666319 74581
rect 666405 74559 666424 74581
rect 666424 74559 666461 74581
rect 666547 74559 666548 74581
rect 666548 74559 666603 74581
rect 666689 74559 666740 74581
rect 666740 74559 666745 74581
rect 666831 74559 666864 74581
rect 666864 74559 666887 74581
rect 666973 74559 666988 74581
rect 666988 74559 667029 74581
rect 667115 74559 667168 74581
rect 667168 74559 667171 74581
rect 667899 75979 667955 76035
rect 668041 75979 668097 76035
rect 668183 75979 668239 76035
rect 668325 75979 668381 76035
rect 668467 75979 668523 76035
rect 668609 75979 668665 76035
rect 668751 75979 668807 76035
rect 668893 75979 668949 76035
rect 669035 75979 669091 76035
rect 669177 75979 669233 76035
rect 669319 75979 669375 76035
rect 669461 75979 669517 76035
rect 669603 75979 669659 76035
rect 667899 75889 667938 75893
rect 667938 75889 667955 75893
rect 668041 75889 668062 75893
rect 668062 75889 668097 75893
rect 668183 75889 668186 75893
rect 668186 75889 668239 75893
rect 668325 75889 668378 75893
rect 668378 75889 668381 75893
rect 668467 75889 668502 75893
rect 668502 75889 668523 75893
rect 668609 75889 668626 75893
rect 668626 75889 668665 75893
rect 668751 75889 668806 75893
rect 668806 75889 668807 75893
rect 668893 75889 668930 75893
rect 668930 75889 668949 75893
rect 669035 75889 669054 75893
rect 669054 75889 669091 75893
rect 669177 75889 669178 75893
rect 669178 75889 669233 75893
rect 669319 75889 669370 75893
rect 669370 75889 669375 75893
rect 669461 75889 669494 75893
rect 669494 75889 669517 75893
rect 669603 75889 669618 75893
rect 669618 75889 669659 75893
rect 667899 75837 667955 75889
rect 668041 75837 668097 75889
rect 668183 75837 668239 75889
rect 668325 75837 668381 75889
rect 668467 75837 668523 75889
rect 668609 75837 668665 75889
rect 668751 75837 668807 75889
rect 668893 75837 668949 75889
rect 669035 75837 669091 75889
rect 669177 75837 669233 75889
rect 669319 75837 669375 75889
rect 669461 75837 669517 75889
rect 669603 75837 669659 75889
rect 667899 75697 667955 75751
rect 668041 75697 668097 75751
rect 668183 75697 668239 75751
rect 668325 75697 668381 75751
rect 668467 75697 668523 75751
rect 668609 75697 668665 75751
rect 668751 75697 668807 75751
rect 668893 75697 668949 75751
rect 669035 75697 669091 75751
rect 669177 75697 669233 75751
rect 669319 75697 669375 75751
rect 669461 75697 669517 75751
rect 669603 75697 669659 75751
rect 667899 75695 667938 75697
rect 667938 75695 667955 75697
rect 668041 75695 668062 75697
rect 668062 75695 668097 75697
rect 668183 75695 668186 75697
rect 668186 75695 668239 75697
rect 668325 75695 668378 75697
rect 668378 75695 668381 75697
rect 668467 75695 668502 75697
rect 668502 75695 668523 75697
rect 668609 75695 668626 75697
rect 668626 75695 668665 75697
rect 668751 75695 668806 75697
rect 668806 75695 668807 75697
rect 668893 75695 668930 75697
rect 668930 75695 668949 75697
rect 669035 75695 669054 75697
rect 669054 75695 669091 75697
rect 669177 75695 669178 75697
rect 669178 75695 669233 75697
rect 669319 75695 669370 75697
rect 669370 75695 669375 75697
rect 669461 75695 669494 75697
rect 669494 75695 669517 75697
rect 669603 75695 669618 75697
rect 669618 75695 669659 75697
rect 667899 75573 667955 75609
rect 668041 75573 668097 75609
rect 668183 75573 668239 75609
rect 668325 75573 668381 75609
rect 668467 75573 668523 75609
rect 668609 75573 668665 75609
rect 668751 75573 668807 75609
rect 668893 75573 668949 75609
rect 669035 75573 669091 75609
rect 669177 75573 669233 75609
rect 669319 75573 669375 75609
rect 669461 75573 669517 75609
rect 669603 75573 669659 75609
rect 667899 75553 667938 75573
rect 667938 75553 667955 75573
rect 668041 75553 668062 75573
rect 668062 75553 668097 75573
rect 668183 75553 668186 75573
rect 668186 75553 668239 75573
rect 668325 75553 668378 75573
rect 668378 75553 668381 75573
rect 668467 75553 668502 75573
rect 668502 75553 668523 75573
rect 668609 75553 668626 75573
rect 668626 75553 668665 75573
rect 668751 75553 668806 75573
rect 668806 75553 668807 75573
rect 668893 75553 668930 75573
rect 668930 75553 668949 75573
rect 669035 75553 669054 75573
rect 669054 75553 669091 75573
rect 669177 75553 669178 75573
rect 669178 75553 669233 75573
rect 669319 75553 669370 75573
rect 669370 75553 669375 75573
rect 669461 75553 669494 75573
rect 669494 75553 669517 75573
rect 669603 75553 669618 75573
rect 669618 75553 669659 75573
rect 667899 75449 667955 75467
rect 668041 75449 668097 75467
rect 668183 75449 668239 75467
rect 668325 75449 668381 75467
rect 668467 75449 668523 75467
rect 668609 75449 668665 75467
rect 668751 75449 668807 75467
rect 668893 75449 668949 75467
rect 669035 75449 669091 75467
rect 669177 75449 669233 75467
rect 669319 75449 669375 75467
rect 669461 75449 669517 75467
rect 669603 75449 669659 75467
rect 667899 75411 667938 75449
rect 667938 75411 667955 75449
rect 668041 75411 668062 75449
rect 668062 75411 668097 75449
rect 668183 75411 668186 75449
rect 668186 75411 668239 75449
rect 668325 75411 668378 75449
rect 668378 75411 668381 75449
rect 668467 75411 668502 75449
rect 668502 75411 668523 75449
rect 668609 75411 668626 75449
rect 668626 75411 668665 75449
rect 668751 75411 668806 75449
rect 668806 75411 668807 75449
rect 668893 75411 668930 75449
rect 668930 75411 668949 75449
rect 669035 75411 669054 75449
rect 669054 75411 669091 75449
rect 669177 75411 669178 75449
rect 669178 75411 669233 75449
rect 669319 75411 669370 75449
rect 669370 75411 669375 75449
rect 669461 75411 669494 75449
rect 669494 75411 669517 75449
rect 669603 75411 669618 75449
rect 669618 75411 669659 75449
rect 667899 75269 667938 75325
rect 667938 75269 667955 75325
rect 668041 75269 668062 75325
rect 668062 75269 668097 75325
rect 668183 75269 668186 75325
rect 668186 75269 668239 75325
rect 668325 75269 668378 75325
rect 668378 75269 668381 75325
rect 668467 75269 668502 75325
rect 668502 75269 668523 75325
rect 668609 75269 668626 75325
rect 668626 75269 668665 75325
rect 668751 75269 668806 75325
rect 668806 75269 668807 75325
rect 668893 75269 668930 75325
rect 668930 75269 668949 75325
rect 669035 75269 669054 75325
rect 669054 75269 669091 75325
rect 669177 75269 669178 75325
rect 669178 75269 669233 75325
rect 669319 75269 669370 75325
rect 669370 75269 669375 75325
rect 669461 75269 669494 75325
rect 669494 75269 669517 75325
rect 669603 75269 669618 75325
rect 669618 75269 669659 75325
rect 667899 75145 667938 75183
rect 667938 75145 667955 75183
rect 668041 75145 668062 75183
rect 668062 75145 668097 75183
rect 668183 75145 668186 75183
rect 668186 75145 668239 75183
rect 668325 75145 668378 75183
rect 668378 75145 668381 75183
rect 668467 75145 668502 75183
rect 668502 75145 668523 75183
rect 668609 75145 668626 75183
rect 668626 75145 668665 75183
rect 668751 75145 668806 75183
rect 668806 75145 668807 75183
rect 668893 75145 668930 75183
rect 668930 75145 668949 75183
rect 669035 75145 669054 75183
rect 669054 75145 669091 75183
rect 669177 75145 669178 75183
rect 669178 75145 669233 75183
rect 669319 75145 669370 75183
rect 669370 75145 669375 75183
rect 669461 75145 669494 75183
rect 669494 75145 669517 75183
rect 669603 75145 669618 75183
rect 669618 75145 669659 75183
rect 667899 75127 667955 75145
rect 668041 75127 668097 75145
rect 668183 75127 668239 75145
rect 668325 75127 668381 75145
rect 668467 75127 668523 75145
rect 668609 75127 668665 75145
rect 668751 75127 668807 75145
rect 668893 75127 668949 75145
rect 669035 75127 669091 75145
rect 669177 75127 669233 75145
rect 669319 75127 669375 75145
rect 669461 75127 669517 75145
rect 669603 75127 669659 75145
rect 667899 75021 667938 75041
rect 667938 75021 667955 75041
rect 668041 75021 668062 75041
rect 668062 75021 668097 75041
rect 668183 75021 668186 75041
rect 668186 75021 668239 75041
rect 668325 75021 668378 75041
rect 668378 75021 668381 75041
rect 668467 75021 668502 75041
rect 668502 75021 668523 75041
rect 668609 75021 668626 75041
rect 668626 75021 668665 75041
rect 668751 75021 668806 75041
rect 668806 75021 668807 75041
rect 668893 75021 668930 75041
rect 668930 75021 668949 75041
rect 669035 75021 669054 75041
rect 669054 75021 669091 75041
rect 669177 75021 669178 75041
rect 669178 75021 669233 75041
rect 669319 75021 669370 75041
rect 669370 75021 669375 75041
rect 669461 75021 669494 75041
rect 669494 75021 669517 75041
rect 669603 75021 669618 75041
rect 669618 75021 669659 75041
rect 667899 74985 667955 75021
rect 668041 74985 668097 75021
rect 668183 74985 668239 75021
rect 668325 74985 668381 75021
rect 668467 74985 668523 75021
rect 668609 74985 668665 75021
rect 668751 74985 668807 75021
rect 668893 74985 668949 75021
rect 669035 74985 669091 75021
rect 669177 74985 669233 75021
rect 669319 74985 669375 75021
rect 669461 74985 669517 75021
rect 669603 74985 669659 75021
rect 667899 74897 667938 74899
rect 667938 74897 667955 74899
rect 668041 74897 668062 74899
rect 668062 74897 668097 74899
rect 668183 74897 668186 74899
rect 668186 74897 668239 74899
rect 668325 74897 668378 74899
rect 668378 74897 668381 74899
rect 668467 74897 668502 74899
rect 668502 74897 668523 74899
rect 668609 74897 668626 74899
rect 668626 74897 668665 74899
rect 668751 74897 668806 74899
rect 668806 74897 668807 74899
rect 668893 74897 668930 74899
rect 668930 74897 668949 74899
rect 669035 74897 669054 74899
rect 669054 74897 669091 74899
rect 669177 74897 669178 74899
rect 669178 74897 669233 74899
rect 669319 74897 669370 74899
rect 669370 74897 669375 74899
rect 669461 74897 669494 74899
rect 669494 74897 669517 74899
rect 669603 74897 669618 74899
rect 669618 74897 669659 74899
rect 667899 74843 667955 74897
rect 668041 74843 668097 74897
rect 668183 74843 668239 74897
rect 668325 74843 668381 74897
rect 668467 74843 668523 74897
rect 668609 74843 668665 74897
rect 668751 74843 668807 74897
rect 668893 74843 668949 74897
rect 669035 74843 669091 74897
rect 669177 74843 669233 74897
rect 669319 74843 669375 74897
rect 669461 74843 669517 74897
rect 669603 74843 669659 74897
rect 667899 74705 667955 74757
rect 668041 74705 668097 74757
rect 668183 74705 668239 74757
rect 668325 74705 668381 74757
rect 668467 74705 668523 74757
rect 668609 74705 668665 74757
rect 668751 74705 668807 74757
rect 668893 74705 668949 74757
rect 669035 74705 669091 74757
rect 669177 74705 669233 74757
rect 669319 74705 669375 74757
rect 669461 74705 669517 74757
rect 669603 74705 669659 74757
rect 667899 74701 667938 74705
rect 667938 74701 667955 74705
rect 668041 74701 668062 74705
rect 668062 74701 668097 74705
rect 668183 74701 668186 74705
rect 668186 74701 668239 74705
rect 668325 74701 668378 74705
rect 668378 74701 668381 74705
rect 668467 74701 668502 74705
rect 668502 74701 668523 74705
rect 668609 74701 668626 74705
rect 668626 74701 668665 74705
rect 668751 74701 668806 74705
rect 668806 74701 668807 74705
rect 668893 74701 668930 74705
rect 668930 74701 668949 74705
rect 669035 74701 669054 74705
rect 669054 74701 669091 74705
rect 669177 74701 669178 74705
rect 669178 74701 669233 74705
rect 669319 74701 669370 74705
rect 669370 74701 669375 74705
rect 669461 74701 669494 74705
rect 669494 74701 669517 74705
rect 669603 74701 669618 74705
rect 669618 74701 669659 74705
rect 667899 74581 667955 74615
rect 668041 74581 668097 74615
rect 668183 74581 668239 74615
rect 668325 74581 668381 74615
rect 668467 74581 668523 74615
rect 668609 74581 668665 74615
rect 668751 74581 668807 74615
rect 668893 74581 668949 74615
rect 669035 74581 669091 74615
rect 669177 74581 669233 74615
rect 669319 74581 669375 74615
rect 669461 74581 669517 74615
rect 669603 74581 669659 74615
rect 667899 74559 667938 74581
rect 667938 74559 667955 74581
rect 668041 74559 668062 74581
rect 668062 74559 668097 74581
rect 668183 74559 668186 74581
rect 668186 74559 668239 74581
rect 668325 74559 668378 74581
rect 668378 74559 668381 74581
rect 668467 74559 668502 74581
rect 668502 74559 668523 74581
rect 668609 74559 668626 74581
rect 668626 74559 668665 74581
rect 668751 74559 668806 74581
rect 668806 74559 668807 74581
rect 668893 74559 668930 74581
rect 668930 74559 668949 74581
rect 669035 74559 669054 74581
rect 669054 74559 669091 74581
rect 669177 74559 669178 74581
rect 669178 74559 669233 74581
rect 669319 74559 669370 74581
rect 669370 74559 669375 74581
rect 669461 74559 669494 74581
rect 669494 74559 669517 74581
rect 669603 74559 669618 74581
rect 669618 74559 669659 74581
rect 105343 73979 105399 74035
rect 105485 73979 105541 74035
rect 105627 73979 105683 74035
rect 105769 73979 105825 74035
rect 105911 73979 105967 74035
rect 106053 73979 106109 74035
rect 106195 73979 106251 74035
rect 106337 73979 106393 74035
rect 106479 73979 106535 74035
rect 106621 73979 106677 74035
rect 106763 73979 106819 74035
rect 106905 73979 106961 74035
rect 107047 73979 107103 74035
rect 105343 73889 105382 73893
rect 105382 73889 105399 73893
rect 105485 73889 105506 73893
rect 105506 73889 105541 73893
rect 105627 73889 105630 73893
rect 105630 73889 105683 73893
rect 105769 73889 105822 73893
rect 105822 73889 105825 73893
rect 105911 73889 105946 73893
rect 105946 73889 105967 73893
rect 106053 73889 106070 73893
rect 106070 73889 106109 73893
rect 106195 73889 106250 73893
rect 106250 73889 106251 73893
rect 106337 73889 106374 73893
rect 106374 73889 106393 73893
rect 106479 73889 106498 73893
rect 106498 73889 106535 73893
rect 106621 73889 106622 73893
rect 106622 73889 106677 73893
rect 106763 73889 106814 73893
rect 106814 73889 106819 73893
rect 106905 73889 106938 73893
rect 106938 73889 106961 73893
rect 107047 73889 107062 73893
rect 107062 73889 107103 73893
rect 105343 73837 105399 73889
rect 105485 73837 105541 73889
rect 105627 73837 105683 73889
rect 105769 73837 105825 73889
rect 105911 73837 105967 73889
rect 106053 73837 106109 73889
rect 106195 73837 106251 73889
rect 106337 73837 106393 73889
rect 106479 73837 106535 73889
rect 106621 73837 106677 73889
rect 106763 73837 106819 73889
rect 106905 73837 106961 73889
rect 107047 73837 107103 73889
rect 105343 73697 105399 73751
rect 105485 73697 105541 73751
rect 105627 73697 105683 73751
rect 105769 73697 105825 73751
rect 105911 73697 105967 73751
rect 106053 73697 106109 73751
rect 106195 73697 106251 73751
rect 106337 73697 106393 73751
rect 106479 73697 106535 73751
rect 106621 73697 106677 73751
rect 106763 73697 106819 73751
rect 106905 73697 106961 73751
rect 107047 73697 107103 73751
rect 105343 73695 105382 73697
rect 105382 73695 105399 73697
rect 105485 73695 105506 73697
rect 105506 73695 105541 73697
rect 105627 73695 105630 73697
rect 105630 73695 105683 73697
rect 105769 73695 105822 73697
rect 105822 73695 105825 73697
rect 105911 73695 105946 73697
rect 105946 73695 105967 73697
rect 106053 73695 106070 73697
rect 106070 73695 106109 73697
rect 106195 73695 106250 73697
rect 106250 73695 106251 73697
rect 106337 73695 106374 73697
rect 106374 73695 106393 73697
rect 106479 73695 106498 73697
rect 106498 73695 106535 73697
rect 106621 73695 106622 73697
rect 106622 73695 106677 73697
rect 106763 73695 106814 73697
rect 106814 73695 106819 73697
rect 106905 73695 106938 73697
rect 106938 73695 106961 73697
rect 107047 73695 107062 73697
rect 107062 73695 107103 73697
rect 105343 73573 105399 73609
rect 105485 73573 105541 73609
rect 105627 73573 105683 73609
rect 105769 73573 105825 73609
rect 105911 73573 105967 73609
rect 106053 73573 106109 73609
rect 106195 73573 106251 73609
rect 106337 73573 106393 73609
rect 106479 73573 106535 73609
rect 106621 73573 106677 73609
rect 106763 73573 106819 73609
rect 106905 73573 106961 73609
rect 107047 73573 107103 73609
rect 105343 73553 105382 73573
rect 105382 73553 105399 73573
rect 105485 73553 105506 73573
rect 105506 73553 105541 73573
rect 105627 73553 105630 73573
rect 105630 73553 105683 73573
rect 105769 73553 105822 73573
rect 105822 73553 105825 73573
rect 105911 73553 105946 73573
rect 105946 73553 105967 73573
rect 106053 73553 106070 73573
rect 106070 73553 106109 73573
rect 106195 73553 106250 73573
rect 106250 73553 106251 73573
rect 106337 73553 106374 73573
rect 106374 73553 106393 73573
rect 106479 73553 106498 73573
rect 106498 73553 106535 73573
rect 106621 73553 106622 73573
rect 106622 73553 106677 73573
rect 106763 73553 106814 73573
rect 106814 73553 106819 73573
rect 106905 73553 106938 73573
rect 106938 73553 106961 73573
rect 107047 73553 107062 73573
rect 107062 73553 107103 73573
rect 105343 73449 105399 73467
rect 105485 73449 105541 73467
rect 105627 73449 105683 73467
rect 105769 73449 105825 73467
rect 105911 73449 105967 73467
rect 106053 73449 106109 73467
rect 106195 73449 106251 73467
rect 106337 73449 106393 73467
rect 106479 73449 106535 73467
rect 106621 73449 106677 73467
rect 106763 73449 106819 73467
rect 106905 73449 106961 73467
rect 107047 73449 107103 73467
rect 105343 73411 105382 73449
rect 105382 73411 105399 73449
rect 105485 73411 105506 73449
rect 105506 73411 105541 73449
rect 105627 73411 105630 73449
rect 105630 73411 105683 73449
rect 105769 73411 105822 73449
rect 105822 73411 105825 73449
rect 105911 73411 105946 73449
rect 105946 73411 105967 73449
rect 106053 73411 106070 73449
rect 106070 73411 106109 73449
rect 106195 73411 106250 73449
rect 106250 73411 106251 73449
rect 106337 73411 106374 73449
rect 106374 73411 106393 73449
rect 106479 73411 106498 73449
rect 106498 73411 106535 73449
rect 106621 73411 106622 73449
rect 106622 73411 106677 73449
rect 106763 73411 106814 73449
rect 106814 73411 106819 73449
rect 106905 73411 106938 73449
rect 106938 73411 106961 73449
rect 107047 73411 107062 73449
rect 107062 73411 107103 73449
rect 105343 73269 105382 73325
rect 105382 73269 105399 73325
rect 105485 73269 105506 73325
rect 105506 73269 105541 73325
rect 105627 73269 105630 73325
rect 105630 73269 105683 73325
rect 105769 73269 105822 73325
rect 105822 73269 105825 73325
rect 105911 73269 105946 73325
rect 105946 73269 105967 73325
rect 106053 73269 106070 73325
rect 106070 73269 106109 73325
rect 106195 73269 106250 73325
rect 106250 73269 106251 73325
rect 106337 73269 106374 73325
rect 106374 73269 106393 73325
rect 106479 73269 106498 73325
rect 106498 73269 106535 73325
rect 106621 73269 106622 73325
rect 106622 73269 106677 73325
rect 106763 73269 106814 73325
rect 106814 73269 106819 73325
rect 106905 73269 106938 73325
rect 106938 73269 106961 73325
rect 107047 73269 107062 73325
rect 107062 73269 107103 73325
rect 105343 73145 105382 73183
rect 105382 73145 105399 73183
rect 105485 73145 105506 73183
rect 105506 73145 105541 73183
rect 105627 73145 105630 73183
rect 105630 73145 105683 73183
rect 105769 73145 105822 73183
rect 105822 73145 105825 73183
rect 105911 73145 105946 73183
rect 105946 73145 105967 73183
rect 106053 73145 106070 73183
rect 106070 73145 106109 73183
rect 106195 73145 106250 73183
rect 106250 73145 106251 73183
rect 106337 73145 106374 73183
rect 106374 73145 106393 73183
rect 106479 73145 106498 73183
rect 106498 73145 106535 73183
rect 106621 73145 106622 73183
rect 106622 73145 106677 73183
rect 106763 73145 106814 73183
rect 106814 73145 106819 73183
rect 106905 73145 106938 73183
rect 106938 73145 106961 73183
rect 107047 73145 107062 73183
rect 107062 73145 107103 73183
rect 105343 73127 105399 73145
rect 105485 73127 105541 73145
rect 105627 73127 105683 73145
rect 105769 73127 105825 73145
rect 105911 73127 105967 73145
rect 106053 73127 106109 73145
rect 106195 73127 106251 73145
rect 106337 73127 106393 73145
rect 106479 73127 106535 73145
rect 106621 73127 106677 73145
rect 106763 73127 106819 73145
rect 106905 73127 106961 73145
rect 107047 73127 107103 73145
rect 105343 73021 105382 73041
rect 105382 73021 105399 73041
rect 105485 73021 105506 73041
rect 105506 73021 105541 73041
rect 105627 73021 105630 73041
rect 105630 73021 105683 73041
rect 105769 73021 105822 73041
rect 105822 73021 105825 73041
rect 105911 73021 105946 73041
rect 105946 73021 105967 73041
rect 106053 73021 106070 73041
rect 106070 73021 106109 73041
rect 106195 73021 106250 73041
rect 106250 73021 106251 73041
rect 106337 73021 106374 73041
rect 106374 73021 106393 73041
rect 106479 73021 106498 73041
rect 106498 73021 106535 73041
rect 106621 73021 106622 73041
rect 106622 73021 106677 73041
rect 106763 73021 106814 73041
rect 106814 73021 106819 73041
rect 106905 73021 106938 73041
rect 106938 73021 106961 73041
rect 107047 73021 107062 73041
rect 107062 73021 107103 73041
rect 105343 72985 105399 73021
rect 105485 72985 105541 73021
rect 105627 72985 105683 73021
rect 105769 72985 105825 73021
rect 105911 72985 105967 73021
rect 106053 72985 106109 73021
rect 106195 72985 106251 73021
rect 106337 72985 106393 73021
rect 106479 72985 106535 73021
rect 106621 72985 106677 73021
rect 106763 72985 106819 73021
rect 106905 72985 106961 73021
rect 107047 72985 107103 73021
rect 105343 72897 105382 72899
rect 105382 72897 105399 72899
rect 105485 72897 105506 72899
rect 105506 72897 105541 72899
rect 105627 72897 105630 72899
rect 105630 72897 105683 72899
rect 105769 72897 105822 72899
rect 105822 72897 105825 72899
rect 105911 72897 105946 72899
rect 105946 72897 105967 72899
rect 106053 72897 106070 72899
rect 106070 72897 106109 72899
rect 106195 72897 106250 72899
rect 106250 72897 106251 72899
rect 106337 72897 106374 72899
rect 106374 72897 106393 72899
rect 106479 72897 106498 72899
rect 106498 72897 106535 72899
rect 106621 72897 106622 72899
rect 106622 72897 106677 72899
rect 106763 72897 106814 72899
rect 106814 72897 106819 72899
rect 106905 72897 106938 72899
rect 106938 72897 106961 72899
rect 107047 72897 107062 72899
rect 107062 72897 107103 72899
rect 105343 72843 105399 72897
rect 105485 72843 105541 72897
rect 105627 72843 105683 72897
rect 105769 72843 105825 72897
rect 105911 72843 105967 72897
rect 106053 72843 106109 72897
rect 106195 72843 106251 72897
rect 106337 72843 106393 72897
rect 106479 72843 106535 72897
rect 106621 72843 106677 72897
rect 106763 72843 106819 72897
rect 106905 72843 106961 72897
rect 107047 72843 107103 72897
rect 105343 72705 105399 72757
rect 105485 72705 105541 72757
rect 105627 72705 105683 72757
rect 105769 72705 105825 72757
rect 105911 72705 105967 72757
rect 106053 72705 106109 72757
rect 106195 72705 106251 72757
rect 106337 72705 106393 72757
rect 106479 72705 106535 72757
rect 106621 72705 106677 72757
rect 106763 72705 106819 72757
rect 106905 72705 106961 72757
rect 107047 72705 107103 72757
rect 105343 72701 105382 72705
rect 105382 72701 105399 72705
rect 105485 72701 105506 72705
rect 105506 72701 105541 72705
rect 105627 72701 105630 72705
rect 105630 72701 105683 72705
rect 105769 72701 105822 72705
rect 105822 72701 105825 72705
rect 105911 72701 105946 72705
rect 105946 72701 105967 72705
rect 106053 72701 106070 72705
rect 106070 72701 106109 72705
rect 106195 72701 106250 72705
rect 106250 72701 106251 72705
rect 106337 72701 106374 72705
rect 106374 72701 106393 72705
rect 106479 72701 106498 72705
rect 106498 72701 106535 72705
rect 106621 72701 106622 72705
rect 106622 72701 106677 72705
rect 106763 72701 106814 72705
rect 106814 72701 106819 72705
rect 106905 72701 106938 72705
rect 106938 72701 106961 72705
rect 107047 72701 107062 72705
rect 107062 72701 107103 72705
rect 105343 72581 105399 72615
rect 105485 72581 105541 72615
rect 105627 72581 105683 72615
rect 105769 72581 105825 72615
rect 105911 72581 105967 72615
rect 106053 72581 106109 72615
rect 106195 72581 106251 72615
rect 106337 72581 106393 72615
rect 106479 72581 106535 72615
rect 106621 72581 106677 72615
rect 106763 72581 106819 72615
rect 106905 72581 106961 72615
rect 107047 72581 107103 72615
rect 105343 72559 105382 72581
rect 105382 72559 105399 72581
rect 105485 72559 105506 72581
rect 105506 72559 105541 72581
rect 105627 72559 105630 72581
rect 105630 72559 105683 72581
rect 105769 72559 105822 72581
rect 105822 72559 105825 72581
rect 105911 72559 105946 72581
rect 105946 72559 105967 72581
rect 106053 72559 106070 72581
rect 106070 72559 106109 72581
rect 106195 72559 106250 72581
rect 106250 72559 106251 72581
rect 106337 72559 106374 72581
rect 106374 72559 106393 72581
rect 106479 72559 106498 72581
rect 106498 72559 106535 72581
rect 106621 72559 106622 72581
rect 106622 72559 106677 72581
rect 106763 72559 106814 72581
rect 106814 72559 106819 72581
rect 106905 72559 106938 72581
rect 106938 72559 106961 72581
rect 107047 72559 107062 72581
rect 107062 72559 107103 72581
rect 105343 72457 105399 72473
rect 105485 72457 105541 72473
rect 105627 72457 105683 72473
rect 105769 72457 105825 72473
rect 105911 72457 105967 72473
rect 106053 72457 106109 72473
rect 106195 72457 106251 72473
rect 106337 72457 106393 72473
rect 106479 72457 106535 72473
rect 106621 72457 106677 72473
rect 106763 72457 106819 72473
rect 106905 72457 106961 72473
rect 107047 72457 107103 72473
rect 105343 72417 105382 72457
rect 105382 72417 105399 72457
rect 105485 72417 105506 72457
rect 105506 72417 105541 72457
rect 105627 72417 105630 72457
rect 105630 72417 105683 72457
rect 105769 72417 105822 72457
rect 105822 72417 105825 72457
rect 105911 72417 105946 72457
rect 105946 72417 105967 72457
rect 106053 72417 106070 72457
rect 106070 72417 106109 72457
rect 106195 72417 106250 72457
rect 106250 72417 106251 72457
rect 106337 72417 106374 72457
rect 106374 72417 106393 72457
rect 106479 72417 106498 72457
rect 106498 72417 106535 72457
rect 106621 72417 106622 72457
rect 106622 72417 106677 72457
rect 106763 72417 106814 72457
rect 106814 72417 106819 72457
rect 106905 72417 106938 72457
rect 106938 72417 106961 72457
rect 107047 72417 107062 72457
rect 107062 72417 107103 72457
rect 105343 72277 105382 72331
rect 105382 72277 105399 72331
rect 105485 72277 105506 72331
rect 105506 72277 105541 72331
rect 105627 72277 105630 72331
rect 105630 72277 105683 72331
rect 105769 72277 105822 72331
rect 105822 72277 105825 72331
rect 105911 72277 105946 72331
rect 105946 72277 105967 72331
rect 106053 72277 106070 72331
rect 106070 72277 106109 72331
rect 106195 72277 106250 72331
rect 106250 72277 106251 72331
rect 106337 72277 106374 72331
rect 106374 72277 106393 72331
rect 106479 72277 106498 72331
rect 106498 72277 106535 72331
rect 106621 72277 106622 72331
rect 106622 72277 106677 72331
rect 106763 72277 106814 72331
rect 106814 72277 106819 72331
rect 106905 72277 106938 72331
rect 106938 72277 106961 72331
rect 107047 72277 107062 72331
rect 107062 72277 107103 72331
rect 105343 72275 105399 72277
rect 105485 72275 105541 72277
rect 105627 72275 105683 72277
rect 105769 72275 105825 72277
rect 105911 72275 105967 72277
rect 106053 72275 106109 72277
rect 106195 72275 106251 72277
rect 106337 72275 106393 72277
rect 106479 72275 106535 72277
rect 106621 72275 106677 72277
rect 106763 72275 106819 72277
rect 106905 72275 106961 72277
rect 107047 72275 107103 72277
rect 105343 72153 105382 72189
rect 105382 72153 105399 72189
rect 105485 72153 105506 72189
rect 105506 72153 105541 72189
rect 105627 72153 105630 72189
rect 105630 72153 105683 72189
rect 105769 72153 105822 72189
rect 105822 72153 105825 72189
rect 105911 72153 105946 72189
rect 105946 72153 105967 72189
rect 106053 72153 106070 72189
rect 106070 72153 106109 72189
rect 106195 72153 106250 72189
rect 106250 72153 106251 72189
rect 106337 72153 106374 72189
rect 106374 72153 106393 72189
rect 106479 72153 106498 72189
rect 106498 72153 106535 72189
rect 106621 72153 106622 72189
rect 106622 72153 106677 72189
rect 106763 72153 106814 72189
rect 106814 72153 106819 72189
rect 106905 72153 106938 72189
rect 106938 72153 106961 72189
rect 107047 72153 107062 72189
rect 107062 72153 107103 72189
rect 105343 72133 105399 72153
rect 105485 72133 105541 72153
rect 105627 72133 105683 72153
rect 105769 72133 105825 72153
rect 105911 72133 105967 72153
rect 106053 72133 106109 72153
rect 106195 72133 106251 72153
rect 106337 72133 106393 72153
rect 106479 72133 106535 72153
rect 106621 72133 106677 72153
rect 106763 72133 106819 72153
rect 106905 72133 106961 72153
rect 107047 72133 107103 72153
rect 108995 73979 109051 74035
rect 109137 73979 109193 74035
rect 109279 73979 109335 74035
rect 109421 73979 109477 74035
rect 109563 73979 109619 74035
rect 109705 73979 109761 74035
rect 108995 73889 109046 73893
rect 109046 73889 109051 73893
rect 109137 73889 109170 73893
rect 109170 73889 109193 73893
rect 109279 73889 109294 73893
rect 109294 73889 109335 73893
rect 109421 73889 109474 73893
rect 109474 73889 109477 73893
rect 109563 73889 109598 73893
rect 109598 73889 109619 73893
rect 109705 73889 109722 73893
rect 109722 73889 109761 73893
rect 108995 73837 109051 73889
rect 109137 73837 109193 73889
rect 109279 73837 109335 73889
rect 109421 73837 109477 73889
rect 109563 73837 109619 73889
rect 109705 73837 109761 73889
rect 108995 73697 109051 73751
rect 109137 73697 109193 73751
rect 109279 73697 109335 73751
rect 109421 73697 109477 73751
rect 109563 73697 109619 73751
rect 109705 73697 109761 73751
rect 108995 73695 109046 73697
rect 109046 73695 109051 73697
rect 109137 73695 109170 73697
rect 109170 73695 109193 73697
rect 109279 73695 109294 73697
rect 109294 73695 109335 73697
rect 109421 73695 109474 73697
rect 109474 73695 109477 73697
rect 109563 73695 109598 73697
rect 109598 73695 109619 73697
rect 109705 73695 109722 73697
rect 109722 73695 109761 73697
rect 108995 73573 109051 73609
rect 109137 73573 109193 73609
rect 109279 73573 109335 73609
rect 109421 73573 109477 73609
rect 109563 73573 109619 73609
rect 109705 73573 109761 73609
rect 108995 73553 109046 73573
rect 109046 73553 109051 73573
rect 109137 73553 109170 73573
rect 109170 73553 109193 73573
rect 109279 73553 109294 73573
rect 109294 73553 109335 73573
rect 109421 73553 109474 73573
rect 109474 73553 109477 73573
rect 109563 73553 109598 73573
rect 109598 73553 109619 73573
rect 109705 73553 109722 73573
rect 109722 73553 109761 73573
rect 108995 73449 109051 73467
rect 109137 73449 109193 73467
rect 109279 73449 109335 73467
rect 109421 73449 109477 73467
rect 109563 73449 109619 73467
rect 109705 73449 109761 73467
rect 108995 73411 109046 73449
rect 109046 73411 109051 73449
rect 109137 73411 109170 73449
rect 109170 73411 109193 73449
rect 109279 73411 109294 73449
rect 109294 73411 109335 73449
rect 109421 73411 109474 73449
rect 109474 73411 109477 73449
rect 109563 73411 109598 73449
rect 109598 73411 109619 73449
rect 109705 73411 109722 73449
rect 109722 73411 109761 73449
rect 108995 73269 109046 73325
rect 109046 73269 109051 73325
rect 109137 73269 109170 73325
rect 109170 73269 109193 73325
rect 109279 73269 109294 73325
rect 109294 73269 109335 73325
rect 109421 73269 109474 73325
rect 109474 73269 109477 73325
rect 109563 73269 109598 73325
rect 109598 73269 109619 73325
rect 109705 73269 109722 73325
rect 109722 73269 109761 73325
rect 108995 73145 109046 73183
rect 109046 73145 109051 73183
rect 109137 73145 109170 73183
rect 109170 73145 109193 73183
rect 109279 73145 109294 73183
rect 109294 73145 109335 73183
rect 109421 73145 109474 73183
rect 109474 73145 109477 73183
rect 109563 73145 109598 73183
rect 109598 73145 109619 73183
rect 109705 73145 109722 73183
rect 109722 73145 109761 73183
rect 108995 73127 109051 73145
rect 109137 73127 109193 73145
rect 109279 73127 109335 73145
rect 109421 73127 109477 73145
rect 109563 73127 109619 73145
rect 109705 73127 109761 73145
rect 108995 73021 109046 73041
rect 109046 73021 109051 73041
rect 109137 73021 109170 73041
rect 109170 73021 109193 73041
rect 109279 73021 109294 73041
rect 109294 73021 109335 73041
rect 109421 73021 109474 73041
rect 109474 73021 109477 73041
rect 109563 73021 109598 73041
rect 109598 73021 109619 73041
rect 109705 73021 109722 73041
rect 109722 73021 109761 73041
rect 108995 72985 109051 73021
rect 109137 72985 109193 73021
rect 109279 72985 109335 73021
rect 109421 72985 109477 73021
rect 109563 72985 109619 73021
rect 109705 72985 109761 73021
rect 108995 72897 109046 72899
rect 109046 72897 109051 72899
rect 109137 72897 109170 72899
rect 109170 72897 109193 72899
rect 109279 72897 109294 72899
rect 109294 72897 109335 72899
rect 109421 72897 109474 72899
rect 109474 72897 109477 72899
rect 109563 72897 109598 72899
rect 109598 72897 109619 72899
rect 109705 72897 109722 72899
rect 109722 72897 109761 72899
rect 108995 72843 109051 72897
rect 109137 72843 109193 72897
rect 109279 72843 109335 72897
rect 109421 72843 109477 72897
rect 109563 72843 109619 72897
rect 109705 72843 109761 72897
rect 108995 72705 109051 72757
rect 109137 72705 109193 72757
rect 109279 72705 109335 72757
rect 109421 72705 109477 72757
rect 109563 72705 109619 72757
rect 109705 72705 109761 72757
rect 108995 72701 109046 72705
rect 109046 72701 109051 72705
rect 109137 72701 109170 72705
rect 109170 72701 109193 72705
rect 109279 72701 109294 72705
rect 109294 72701 109335 72705
rect 109421 72701 109474 72705
rect 109474 72701 109477 72705
rect 109563 72701 109598 72705
rect 109598 72701 109619 72705
rect 109705 72701 109722 72705
rect 109722 72701 109761 72705
rect 108995 72581 109051 72615
rect 109137 72581 109193 72615
rect 109279 72581 109335 72615
rect 109421 72581 109477 72615
rect 109563 72581 109619 72615
rect 109705 72581 109761 72615
rect 108995 72559 109046 72581
rect 109046 72559 109051 72581
rect 109137 72559 109170 72581
rect 109170 72559 109193 72581
rect 109279 72559 109294 72581
rect 109294 72559 109335 72581
rect 109421 72559 109474 72581
rect 109474 72559 109477 72581
rect 109563 72559 109598 72581
rect 109598 72559 109619 72581
rect 109705 72559 109722 72581
rect 109722 72559 109761 72581
rect 108995 72457 109051 72473
rect 109137 72457 109193 72473
rect 109279 72457 109335 72473
rect 109421 72457 109477 72473
rect 109563 72457 109619 72473
rect 109705 72457 109761 72473
rect 108995 72417 109046 72457
rect 109046 72417 109051 72457
rect 109137 72417 109170 72457
rect 109170 72417 109193 72457
rect 109279 72417 109294 72457
rect 109294 72417 109335 72457
rect 109421 72417 109474 72457
rect 109474 72417 109477 72457
rect 109563 72417 109598 72457
rect 109598 72417 109619 72457
rect 109705 72417 109722 72457
rect 109722 72417 109761 72457
rect 108995 72277 109046 72331
rect 109046 72277 109051 72331
rect 109137 72277 109170 72331
rect 109170 72277 109193 72331
rect 109279 72277 109294 72331
rect 109294 72277 109335 72331
rect 109421 72277 109474 72331
rect 109474 72277 109477 72331
rect 109563 72277 109598 72331
rect 109598 72277 109619 72331
rect 109705 72277 109722 72331
rect 109722 72277 109761 72331
rect 108995 72275 109051 72277
rect 109137 72275 109193 72277
rect 109279 72275 109335 72277
rect 109421 72275 109477 72277
rect 109563 72275 109619 72277
rect 109705 72275 109761 72277
rect 108995 72153 109046 72189
rect 109046 72153 109051 72189
rect 109137 72153 109170 72189
rect 109170 72153 109193 72189
rect 109279 72153 109294 72189
rect 109294 72153 109335 72189
rect 109421 72153 109474 72189
rect 109474 72153 109477 72189
rect 109563 72153 109598 72189
rect 109598 72153 109619 72189
rect 109705 72153 109722 72189
rect 109722 72153 109761 72189
rect 108995 72133 109051 72153
rect 109137 72133 109193 72153
rect 109279 72133 109335 72153
rect 109421 72133 109477 72153
rect 109563 72133 109619 72153
rect 109705 72133 109761 72153
rect 110193 73979 110249 74035
rect 110335 73979 110391 74035
rect 110477 73979 110533 74035
rect 110619 73979 110675 74035
rect 110761 73979 110817 74035
rect 110903 73979 110959 74035
rect 111045 73979 111101 74035
rect 111187 73979 111243 74035
rect 111329 73979 111385 74035
rect 111471 73979 111527 74035
rect 111613 73979 111669 74035
rect 111755 73979 111811 74035
rect 111897 73979 111953 74035
rect 112039 73979 112095 74035
rect 110193 73889 110232 73893
rect 110232 73889 110249 73893
rect 110335 73889 110356 73893
rect 110356 73889 110391 73893
rect 110477 73889 110480 73893
rect 110480 73889 110533 73893
rect 110619 73889 110672 73893
rect 110672 73889 110675 73893
rect 110761 73889 110796 73893
rect 110796 73889 110817 73893
rect 110903 73889 110920 73893
rect 110920 73889 110959 73893
rect 111045 73889 111100 73893
rect 111100 73889 111101 73893
rect 111187 73889 111224 73893
rect 111224 73889 111243 73893
rect 111329 73889 111348 73893
rect 111348 73889 111385 73893
rect 111471 73889 111472 73893
rect 111472 73889 111527 73893
rect 111613 73889 111664 73893
rect 111664 73889 111669 73893
rect 111755 73889 111788 73893
rect 111788 73889 111811 73893
rect 111897 73889 111912 73893
rect 111912 73889 111953 73893
rect 112039 73889 112092 73893
rect 112092 73889 112095 73893
rect 110193 73837 110249 73889
rect 110335 73837 110391 73889
rect 110477 73837 110533 73889
rect 110619 73837 110675 73889
rect 110761 73837 110817 73889
rect 110903 73837 110959 73889
rect 111045 73837 111101 73889
rect 111187 73837 111243 73889
rect 111329 73837 111385 73889
rect 111471 73837 111527 73889
rect 111613 73837 111669 73889
rect 111755 73837 111811 73889
rect 111897 73837 111953 73889
rect 112039 73837 112095 73889
rect 110193 73697 110249 73751
rect 110335 73697 110391 73751
rect 110477 73697 110533 73751
rect 110619 73697 110675 73751
rect 110761 73697 110817 73751
rect 110903 73697 110959 73751
rect 111045 73697 111101 73751
rect 111187 73697 111243 73751
rect 111329 73697 111385 73751
rect 111471 73697 111527 73751
rect 111613 73697 111669 73751
rect 111755 73697 111811 73751
rect 111897 73697 111953 73751
rect 112039 73697 112095 73751
rect 110193 73695 110232 73697
rect 110232 73695 110249 73697
rect 110335 73695 110356 73697
rect 110356 73695 110391 73697
rect 110477 73695 110480 73697
rect 110480 73695 110533 73697
rect 110619 73695 110672 73697
rect 110672 73695 110675 73697
rect 110761 73695 110796 73697
rect 110796 73695 110817 73697
rect 110903 73695 110920 73697
rect 110920 73695 110959 73697
rect 111045 73695 111100 73697
rect 111100 73695 111101 73697
rect 111187 73695 111224 73697
rect 111224 73695 111243 73697
rect 111329 73695 111348 73697
rect 111348 73695 111385 73697
rect 111471 73695 111472 73697
rect 111472 73695 111527 73697
rect 111613 73695 111664 73697
rect 111664 73695 111669 73697
rect 111755 73695 111788 73697
rect 111788 73695 111811 73697
rect 111897 73695 111912 73697
rect 111912 73695 111953 73697
rect 112039 73695 112092 73697
rect 112092 73695 112095 73697
rect 110193 73573 110249 73609
rect 110335 73573 110391 73609
rect 110477 73573 110533 73609
rect 110619 73573 110675 73609
rect 110761 73573 110817 73609
rect 110903 73573 110959 73609
rect 111045 73573 111101 73609
rect 111187 73573 111243 73609
rect 111329 73573 111385 73609
rect 111471 73573 111527 73609
rect 111613 73573 111669 73609
rect 111755 73573 111811 73609
rect 111897 73573 111953 73609
rect 112039 73573 112095 73609
rect 110193 73553 110232 73573
rect 110232 73553 110249 73573
rect 110335 73553 110356 73573
rect 110356 73553 110391 73573
rect 110477 73553 110480 73573
rect 110480 73553 110533 73573
rect 110619 73553 110672 73573
rect 110672 73553 110675 73573
rect 110761 73553 110796 73573
rect 110796 73553 110817 73573
rect 110903 73553 110920 73573
rect 110920 73553 110959 73573
rect 111045 73553 111100 73573
rect 111100 73553 111101 73573
rect 111187 73553 111224 73573
rect 111224 73553 111243 73573
rect 111329 73553 111348 73573
rect 111348 73553 111385 73573
rect 111471 73553 111472 73573
rect 111472 73553 111527 73573
rect 111613 73553 111664 73573
rect 111664 73553 111669 73573
rect 111755 73553 111788 73573
rect 111788 73553 111811 73573
rect 111897 73553 111912 73573
rect 111912 73553 111953 73573
rect 112039 73553 112092 73573
rect 112092 73553 112095 73573
rect 110193 73449 110249 73467
rect 110335 73449 110391 73467
rect 110477 73449 110533 73467
rect 110619 73449 110675 73467
rect 110761 73449 110817 73467
rect 110903 73449 110959 73467
rect 111045 73449 111101 73467
rect 111187 73449 111243 73467
rect 111329 73449 111385 73467
rect 111471 73449 111527 73467
rect 111613 73449 111669 73467
rect 111755 73449 111811 73467
rect 111897 73449 111953 73467
rect 112039 73449 112095 73467
rect 110193 73411 110232 73449
rect 110232 73411 110249 73449
rect 110335 73411 110356 73449
rect 110356 73411 110391 73449
rect 110477 73411 110480 73449
rect 110480 73411 110533 73449
rect 110619 73411 110672 73449
rect 110672 73411 110675 73449
rect 110761 73411 110796 73449
rect 110796 73411 110817 73449
rect 110903 73411 110920 73449
rect 110920 73411 110959 73449
rect 111045 73411 111100 73449
rect 111100 73411 111101 73449
rect 111187 73411 111224 73449
rect 111224 73411 111243 73449
rect 111329 73411 111348 73449
rect 111348 73411 111385 73449
rect 111471 73411 111472 73449
rect 111472 73411 111527 73449
rect 111613 73411 111664 73449
rect 111664 73411 111669 73449
rect 111755 73411 111788 73449
rect 111788 73411 111811 73449
rect 111897 73411 111912 73449
rect 111912 73411 111953 73449
rect 112039 73411 112092 73449
rect 112092 73411 112095 73449
rect 110193 73269 110232 73325
rect 110232 73269 110249 73325
rect 110335 73269 110356 73325
rect 110356 73269 110391 73325
rect 110477 73269 110480 73325
rect 110480 73269 110533 73325
rect 110619 73269 110672 73325
rect 110672 73269 110675 73325
rect 110761 73269 110796 73325
rect 110796 73269 110817 73325
rect 110903 73269 110920 73325
rect 110920 73269 110959 73325
rect 111045 73269 111100 73325
rect 111100 73269 111101 73325
rect 111187 73269 111224 73325
rect 111224 73269 111243 73325
rect 111329 73269 111348 73325
rect 111348 73269 111385 73325
rect 111471 73269 111472 73325
rect 111472 73269 111527 73325
rect 111613 73269 111664 73325
rect 111664 73269 111669 73325
rect 111755 73269 111788 73325
rect 111788 73269 111811 73325
rect 111897 73269 111912 73325
rect 111912 73269 111953 73325
rect 112039 73269 112092 73325
rect 112092 73269 112095 73325
rect 110193 73145 110232 73183
rect 110232 73145 110249 73183
rect 110335 73145 110356 73183
rect 110356 73145 110391 73183
rect 110477 73145 110480 73183
rect 110480 73145 110533 73183
rect 110619 73145 110672 73183
rect 110672 73145 110675 73183
rect 110761 73145 110796 73183
rect 110796 73145 110817 73183
rect 110903 73145 110920 73183
rect 110920 73145 110959 73183
rect 111045 73145 111100 73183
rect 111100 73145 111101 73183
rect 111187 73145 111224 73183
rect 111224 73145 111243 73183
rect 111329 73145 111348 73183
rect 111348 73145 111385 73183
rect 111471 73145 111472 73183
rect 111472 73145 111527 73183
rect 111613 73145 111664 73183
rect 111664 73145 111669 73183
rect 111755 73145 111788 73183
rect 111788 73145 111811 73183
rect 111897 73145 111912 73183
rect 111912 73145 111953 73183
rect 112039 73145 112092 73183
rect 112092 73145 112095 73183
rect 110193 73127 110249 73145
rect 110335 73127 110391 73145
rect 110477 73127 110533 73145
rect 110619 73127 110675 73145
rect 110761 73127 110817 73145
rect 110903 73127 110959 73145
rect 111045 73127 111101 73145
rect 111187 73127 111243 73145
rect 111329 73127 111385 73145
rect 111471 73127 111527 73145
rect 111613 73127 111669 73145
rect 111755 73127 111811 73145
rect 111897 73127 111953 73145
rect 112039 73127 112095 73145
rect 110193 73021 110232 73041
rect 110232 73021 110249 73041
rect 110335 73021 110356 73041
rect 110356 73021 110391 73041
rect 110477 73021 110480 73041
rect 110480 73021 110533 73041
rect 110619 73021 110672 73041
rect 110672 73021 110675 73041
rect 110761 73021 110796 73041
rect 110796 73021 110817 73041
rect 110903 73021 110920 73041
rect 110920 73021 110959 73041
rect 111045 73021 111100 73041
rect 111100 73021 111101 73041
rect 111187 73021 111224 73041
rect 111224 73021 111243 73041
rect 111329 73021 111348 73041
rect 111348 73021 111385 73041
rect 111471 73021 111472 73041
rect 111472 73021 111527 73041
rect 111613 73021 111664 73041
rect 111664 73021 111669 73041
rect 111755 73021 111788 73041
rect 111788 73021 111811 73041
rect 111897 73021 111912 73041
rect 111912 73021 111953 73041
rect 112039 73021 112092 73041
rect 112092 73021 112095 73041
rect 110193 72985 110249 73021
rect 110335 72985 110391 73021
rect 110477 72985 110533 73021
rect 110619 72985 110675 73021
rect 110761 72985 110817 73021
rect 110903 72985 110959 73021
rect 111045 72985 111101 73021
rect 111187 72985 111243 73021
rect 111329 72985 111385 73021
rect 111471 72985 111527 73021
rect 111613 72985 111669 73021
rect 111755 72985 111811 73021
rect 111897 72985 111953 73021
rect 112039 72985 112095 73021
rect 110193 72897 110232 72899
rect 110232 72897 110249 72899
rect 110335 72897 110356 72899
rect 110356 72897 110391 72899
rect 110477 72897 110480 72899
rect 110480 72897 110533 72899
rect 110619 72897 110672 72899
rect 110672 72897 110675 72899
rect 110761 72897 110796 72899
rect 110796 72897 110817 72899
rect 110903 72897 110920 72899
rect 110920 72897 110959 72899
rect 111045 72897 111100 72899
rect 111100 72897 111101 72899
rect 111187 72897 111224 72899
rect 111224 72897 111243 72899
rect 111329 72897 111348 72899
rect 111348 72897 111385 72899
rect 111471 72897 111472 72899
rect 111472 72897 111527 72899
rect 111613 72897 111664 72899
rect 111664 72897 111669 72899
rect 111755 72897 111788 72899
rect 111788 72897 111811 72899
rect 111897 72897 111912 72899
rect 111912 72897 111953 72899
rect 112039 72897 112092 72899
rect 112092 72897 112095 72899
rect 110193 72843 110249 72897
rect 110335 72843 110391 72897
rect 110477 72843 110533 72897
rect 110619 72843 110675 72897
rect 110761 72843 110817 72897
rect 110903 72843 110959 72897
rect 111045 72843 111101 72897
rect 111187 72843 111243 72897
rect 111329 72843 111385 72897
rect 111471 72843 111527 72897
rect 111613 72843 111669 72897
rect 111755 72843 111811 72897
rect 111897 72843 111953 72897
rect 112039 72843 112095 72897
rect 110193 72705 110249 72757
rect 110335 72705 110391 72757
rect 110477 72705 110533 72757
rect 110619 72705 110675 72757
rect 110761 72705 110817 72757
rect 110903 72705 110959 72757
rect 111045 72705 111101 72757
rect 111187 72705 111243 72757
rect 111329 72705 111385 72757
rect 111471 72705 111527 72757
rect 111613 72705 111669 72757
rect 111755 72705 111811 72757
rect 111897 72705 111953 72757
rect 112039 72705 112095 72757
rect 110193 72701 110232 72705
rect 110232 72701 110249 72705
rect 110335 72701 110356 72705
rect 110356 72701 110391 72705
rect 110477 72701 110480 72705
rect 110480 72701 110533 72705
rect 110619 72701 110672 72705
rect 110672 72701 110675 72705
rect 110761 72701 110796 72705
rect 110796 72701 110817 72705
rect 110903 72701 110920 72705
rect 110920 72701 110959 72705
rect 111045 72701 111100 72705
rect 111100 72701 111101 72705
rect 111187 72701 111224 72705
rect 111224 72701 111243 72705
rect 111329 72701 111348 72705
rect 111348 72701 111385 72705
rect 111471 72701 111472 72705
rect 111472 72701 111527 72705
rect 111613 72701 111664 72705
rect 111664 72701 111669 72705
rect 111755 72701 111788 72705
rect 111788 72701 111811 72705
rect 111897 72701 111912 72705
rect 111912 72701 111953 72705
rect 112039 72701 112092 72705
rect 112092 72701 112095 72705
rect 110193 72581 110249 72615
rect 110335 72581 110391 72615
rect 110477 72581 110533 72615
rect 110619 72581 110675 72615
rect 110761 72581 110817 72615
rect 110903 72581 110959 72615
rect 111045 72581 111101 72615
rect 111187 72581 111243 72615
rect 111329 72581 111385 72615
rect 111471 72581 111527 72615
rect 111613 72581 111669 72615
rect 111755 72581 111811 72615
rect 111897 72581 111953 72615
rect 112039 72581 112095 72615
rect 110193 72559 110232 72581
rect 110232 72559 110249 72581
rect 110335 72559 110356 72581
rect 110356 72559 110391 72581
rect 110477 72559 110480 72581
rect 110480 72559 110533 72581
rect 110619 72559 110672 72581
rect 110672 72559 110675 72581
rect 110761 72559 110796 72581
rect 110796 72559 110817 72581
rect 110903 72559 110920 72581
rect 110920 72559 110959 72581
rect 111045 72559 111100 72581
rect 111100 72559 111101 72581
rect 111187 72559 111224 72581
rect 111224 72559 111243 72581
rect 111329 72559 111348 72581
rect 111348 72559 111385 72581
rect 111471 72559 111472 72581
rect 111472 72559 111527 72581
rect 111613 72559 111664 72581
rect 111664 72559 111669 72581
rect 111755 72559 111788 72581
rect 111788 72559 111811 72581
rect 111897 72559 111912 72581
rect 111912 72559 111953 72581
rect 112039 72559 112092 72581
rect 112092 72559 112095 72581
rect 110193 72457 110249 72473
rect 110335 72457 110391 72473
rect 110477 72457 110533 72473
rect 110619 72457 110675 72473
rect 110761 72457 110817 72473
rect 110903 72457 110959 72473
rect 111045 72457 111101 72473
rect 111187 72457 111243 72473
rect 111329 72457 111385 72473
rect 111471 72457 111527 72473
rect 111613 72457 111669 72473
rect 111755 72457 111811 72473
rect 111897 72457 111953 72473
rect 112039 72457 112095 72473
rect 110193 72417 110232 72457
rect 110232 72417 110249 72457
rect 110335 72417 110356 72457
rect 110356 72417 110391 72457
rect 110477 72417 110480 72457
rect 110480 72417 110533 72457
rect 110619 72417 110672 72457
rect 110672 72417 110675 72457
rect 110761 72417 110796 72457
rect 110796 72417 110817 72457
rect 110903 72417 110920 72457
rect 110920 72417 110959 72457
rect 111045 72417 111100 72457
rect 111100 72417 111101 72457
rect 111187 72417 111224 72457
rect 111224 72417 111243 72457
rect 111329 72417 111348 72457
rect 111348 72417 111385 72457
rect 111471 72417 111472 72457
rect 111472 72417 111527 72457
rect 111613 72417 111664 72457
rect 111664 72417 111669 72457
rect 111755 72417 111788 72457
rect 111788 72417 111811 72457
rect 111897 72417 111912 72457
rect 111912 72417 111953 72457
rect 112039 72417 112092 72457
rect 112092 72417 112095 72457
rect 110193 72277 110232 72331
rect 110232 72277 110249 72331
rect 110335 72277 110356 72331
rect 110356 72277 110391 72331
rect 110477 72277 110480 72331
rect 110480 72277 110533 72331
rect 110619 72277 110672 72331
rect 110672 72277 110675 72331
rect 110761 72277 110796 72331
rect 110796 72277 110817 72331
rect 110903 72277 110920 72331
rect 110920 72277 110959 72331
rect 111045 72277 111100 72331
rect 111100 72277 111101 72331
rect 111187 72277 111224 72331
rect 111224 72277 111243 72331
rect 111329 72277 111348 72331
rect 111348 72277 111385 72331
rect 111471 72277 111472 72331
rect 111472 72277 111527 72331
rect 111613 72277 111664 72331
rect 111664 72277 111669 72331
rect 111755 72277 111788 72331
rect 111788 72277 111811 72331
rect 111897 72277 111912 72331
rect 111912 72277 111953 72331
rect 112039 72277 112092 72331
rect 112092 72277 112095 72331
rect 110193 72275 110249 72277
rect 110335 72275 110391 72277
rect 110477 72275 110533 72277
rect 110619 72275 110675 72277
rect 110761 72275 110817 72277
rect 110903 72275 110959 72277
rect 111045 72275 111101 72277
rect 111187 72275 111243 72277
rect 111329 72275 111385 72277
rect 111471 72275 111527 72277
rect 111613 72275 111669 72277
rect 111755 72275 111811 72277
rect 111897 72275 111953 72277
rect 112039 72275 112095 72277
rect 110193 72153 110232 72189
rect 110232 72153 110249 72189
rect 110335 72153 110356 72189
rect 110356 72153 110391 72189
rect 110477 72153 110480 72189
rect 110480 72153 110533 72189
rect 110619 72153 110672 72189
rect 110672 72153 110675 72189
rect 110761 72153 110796 72189
rect 110796 72153 110817 72189
rect 110903 72153 110920 72189
rect 110920 72153 110959 72189
rect 111045 72153 111100 72189
rect 111100 72153 111101 72189
rect 111187 72153 111224 72189
rect 111224 72153 111243 72189
rect 111329 72153 111348 72189
rect 111348 72153 111385 72189
rect 111471 72153 111472 72189
rect 111472 72153 111527 72189
rect 111613 72153 111664 72189
rect 111664 72153 111669 72189
rect 111755 72153 111788 72189
rect 111788 72153 111811 72189
rect 111897 72153 111912 72189
rect 111912 72153 111953 72189
rect 112039 72153 112092 72189
rect 112092 72153 112095 72189
rect 110193 72133 110249 72153
rect 110335 72133 110391 72153
rect 110477 72133 110533 72153
rect 110619 72133 110675 72153
rect 110761 72133 110817 72153
rect 110903 72133 110959 72153
rect 111045 72133 111101 72153
rect 111187 72133 111243 72153
rect 111329 72133 111385 72153
rect 111471 72133 111527 72153
rect 111613 72133 111669 72153
rect 111755 72133 111811 72153
rect 111897 72133 111953 72153
rect 112039 72133 112095 72153
rect 113325 73979 113381 74035
rect 113467 73979 113523 74035
rect 113609 73979 113665 74035
rect 113751 73979 113807 74035
rect 113893 73979 113949 74035
rect 114035 73979 114091 74035
rect 114177 73979 114233 74035
rect 114319 73979 114375 74035
rect 114461 73979 114517 74035
rect 114603 73979 114659 74035
rect 114745 73979 114801 74035
rect 113325 73889 113378 73893
rect 113378 73889 113381 73893
rect 113467 73889 113502 73893
rect 113502 73889 113523 73893
rect 113609 73889 113626 73893
rect 113626 73889 113665 73893
rect 113751 73889 113806 73893
rect 113806 73889 113807 73893
rect 113893 73889 113930 73893
rect 113930 73889 113949 73893
rect 114035 73889 114054 73893
rect 114054 73889 114091 73893
rect 114177 73889 114178 73893
rect 114178 73889 114233 73893
rect 114319 73889 114370 73893
rect 114370 73889 114375 73893
rect 114461 73889 114494 73893
rect 114494 73889 114517 73893
rect 114603 73889 114618 73893
rect 114618 73889 114659 73893
rect 114745 73889 114798 73893
rect 114798 73889 114801 73893
rect 113325 73837 113381 73889
rect 113467 73837 113523 73889
rect 113609 73837 113665 73889
rect 113751 73837 113807 73889
rect 113893 73837 113949 73889
rect 114035 73837 114091 73889
rect 114177 73837 114233 73889
rect 114319 73837 114375 73889
rect 114461 73837 114517 73889
rect 114603 73837 114659 73889
rect 114745 73837 114801 73889
rect 113325 73697 113381 73751
rect 113467 73697 113523 73751
rect 113609 73697 113665 73751
rect 113751 73697 113807 73751
rect 113893 73697 113949 73751
rect 114035 73697 114091 73751
rect 114177 73697 114233 73751
rect 114319 73697 114375 73751
rect 114461 73697 114517 73751
rect 114603 73697 114659 73751
rect 114745 73697 114801 73751
rect 113325 73695 113378 73697
rect 113378 73695 113381 73697
rect 113467 73695 113502 73697
rect 113502 73695 113523 73697
rect 113609 73695 113626 73697
rect 113626 73695 113665 73697
rect 113751 73695 113806 73697
rect 113806 73695 113807 73697
rect 113893 73695 113930 73697
rect 113930 73695 113949 73697
rect 114035 73695 114054 73697
rect 114054 73695 114091 73697
rect 114177 73695 114178 73697
rect 114178 73695 114233 73697
rect 114319 73695 114370 73697
rect 114370 73695 114375 73697
rect 114461 73695 114494 73697
rect 114494 73695 114517 73697
rect 114603 73695 114618 73697
rect 114618 73695 114659 73697
rect 114745 73695 114798 73697
rect 114798 73695 114801 73697
rect 113325 73573 113381 73609
rect 113467 73573 113523 73609
rect 113609 73573 113665 73609
rect 113751 73573 113807 73609
rect 113893 73573 113949 73609
rect 114035 73573 114091 73609
rect 114177 73573 114233 73609
rect 114319 73573 114375 73609
rect 114461 73573 114517 73609
rect 114603 73573 114659 73609
rect 114745 73573 114801 73609
rect 113325 73553 113378 73573
rect 113378 73553 113381 73573
rect 113467 73553 113502 73573
rect 113502 73553 113523 73573
rect 113609 73553 113626 73573
rect 113626 73553 113665 73573
rect 113751 73553 113806 73573
rect 113806 73553 113807 73573
rect 113893 73553 113930 73573
rect 113930 73553 113949 73573
rect 114035 73553 114054 73573
rect 114054 73553 114091 73573
rect 114177 73553 114178 73573
rect 114178 73553 114233 73573
rect 114319 73553 114370 73573
rect 114370 73553 114375 73573
rect 114461 73553 114494 73573
rect 114494 73553 114517 73573
rect 114603 73553 114618 73573
rect 114618 73553 114659 73573
rect 114745 73553 114798 73573
rect 114798 73553 114801 73573
rect 113325 73449 113381 73467
rect 113467 73449 113523 73467
rect 113609 73449 113665 73467
rect 113751 73449 113807 73467
rect 113893 73449 113949 73467
rect 114035 73449 114091 73467
rect 114177 73449 114233 73467
rect 114319 73449 114375 73467
rect 114461 73449 114517 73467
rect 114603 73449 114659 73467
rect 114745 73449 114801 73467
rect 113325 73411 113378 73449
rect 113378 73411 113381 73449
rect 113467 73411 113502 73449
rect 113502 73411 113523 73449
rect 113609 73411 113626 73449
rect 113626 73411 113665 73449
rect 113751 73411 113806 73449
rect 113806 73411 113807 73449
rect 113893 73411 113930 73449
rect 113930 73411 113949 73449
rect 114035 73411 114054 73449
rect 114054 73411 114091 73449
rect 114177 73411 114178 73449
rect 114178 73411 114233 73449
rect 114319 73411 114370 73449
rect 114370 73411 114375 73449
rect 114461 73411 114494 73449
rect 114494 73411 114517 73449
rect 114603 73411 114618 73449
rect 114618 73411 114659 73449
rect 114745 73411 114798 73449
rect 114798 73411 114801 73449
rect 113325 73269 113378 73325
rect 113378 73269 113381 73325
rect 113467 73269 113502 73325
rect 113502 73269 113523 73325
rect 113609 73269 113626 73325
rect 113626 73269 113665 73325
rect 113751 73269 113806 73325
rect 113806 73269 113807 73325
rect 113893 73269 113930 73325
rect 113930 73269 113949 73325
rect 114035 73269 114054 73325
rect 114054 73269 114091 73325
rect 114177 73269 114178 73325
rect 114178 73269 114233 73325
rect 114319 73269 114370 73325
rect 114370 73269 114375 73325
rect 114461 73269 114494 73325
rect 114494 73269 114517 73325
rect 114603 73269 114618 73325
rect 114618 73269 114659 73325
rect 114745 73269 114798 73325
rect 114798 73269 114801 73325
rect 113325 73145 113378 73183
rect 113378 73145 113381 73183
rect 113467 73145 113502 73183
rect 113502 73145 113523 73183
rect 113609 73145 113626 73183
rect 113626 73145 113665 73183
rect 113751 73145 113806 73183
rect 113806 73145 113807 73183
rect 113893 73145 113930 73183
rect 113930 73145 113949 73183
rect 114035 73145 114054 73183
rect 114054 73145 114091 73183
rect 114177 73145 114178 73183
rect 114178 73145 114233 73183
rect 114319 73145 114370 73183
rect 114370 73145 114375 73183
rect 114461 73145 114494 73183
rect 114494 73145 114517 73183
rect 114603 73145 114618 73183
rect 114618 73145 114659 73183
rect 114745 73145 114798 73183
rect 114798 73145 114801 73183
rect 113325 73127 113381 73145
rect 113467 73127 113523 73145
rect 113609 73127 113665 73145
rect 113751 73127 113807 73145
rect 113893 73127 113949 73145
rect 114035 73127 114091 73145
rect 114177 73127 114233 73145
rect 114319 73127 114375 73145
rect 114461 73127 114517 73145
rect 114603 73127 114659 73145
rect 114745 73127 114801 73145
rect 113325 73021 113378 73041
rect 113378 73021 113381 73041
rect 113467 73021 113502 73041
rect 113502 73021 113523 73041
rect 113609 73021 113626 73041
rect 113626 73021 113665 73041
rect 113751 73021 113806 73041
rect 113806 73021 113807 73041
rect 113893 73021 113930 73041
rect 113930 73021 113949 73041
rect 114035 73021 114054 73041
rect 114054 73021 114091 73041
rect 114177 73021 114178 73041
rect 114178 73021 114233 73041
rect 114319 73021 114370 73041
rect 114370 73021 114375 73041
rect 114461 73021 114494 73041
rect 114494 73021 114517 73041
rect 114603 73021 114618 73041
rect 114618 73021 114659 73041
rect 114745 73021 114798 73041
rect 114798 73021 114801 73041
rect 113325 72985 113381 73021
rect 113467 72985 113523 73021
rect 113609 72985 113665 73021
rect 113751 72985 113807 73021
rect 113893 72985 113949 73021
rect 114035 72985 114091 73021
rect 114177 72985 114233 73021
rect 114319 72985 114375 73021
rect 114461 72985 114517 73021
rect 114603 72985 114659 73021
rect 114745 72985 114801 73021
rect 113325 72897 113378 72899
rect 113378 72897 113381 72899
rect 113467 72897 113502 72899
rect 113502 72897 113523 72899
rect 113609 72897 113626 72899
rect 113626 72897 113665 72899
rect 113751 72897 113806 72899
rect 113806 72897 113807 72899
rect 113893 72897 113930 72899
rect 113930 72897 113949 72899
rect 114035 72897 114054 72899
rect 114054 72897 114091 72899
rect 114177 72897 114178 72899
rect 114178 72897 114233 72899
rect 114319 72897 114370 72899
rect 114370 72897 114375 72899
rect 114461 72897 114494 72899
rect 114494 72897 114517 72899
rect 114603 72897 114618 72899
rect 114618 72897 114659 72899
rect 114745 72897 114798 72899
rect 114798 72897 114801 72899
rect 113325 72843 113381 72897
rect 113467 72843 113523 72897
rect 113609 72843 113665 72897
rect 113751 72843 113807 72897
rect 113893 72843 113949 72897
rect 114035 72843 114091 72897
rect 114177 72843 114233 72897
rect 114319 72843 114375 72897
rect 114461 72843 114517 72897
rect 114603 72843 114659 72897
rect 114745 72843 114801 72897
rect 113325 72705 113381 72757
rect 113467 72705 113523 72757
rect 113609 72705 113665 72757
rect 113751 72705 113807 72757
rect 113893 72705 113949 72757
rect 114035 72705 114091 72757
rect 114177 72705 114233 72757
rect 114319 72705 114375 72757
rect 114461 72705 114517 72757
rect 114603 72705 114659 72757
rect 114745 72705 114801 72757
rect 113325 72701 113378 72705
rect 113378 72701 113381 72705
rect 113467 72701 113502 72705
rect 113502 72701 113523 72705
rect 113609 72701 113626 72705
rect 113626 72701 113665 72705
rect 113751 72701 113806 72705
rect 113806 72701 113807 72705
rect 113893 72701 113930 72705
rect 113930 72701 113949 72705
rect 114035 72701 114054 72705
rect 114054 72701 114091 72705
rect 114177 72701 114178 72705
rect 114178 72701 114233 72705
rect 114319 72701 114370 72705
rect 114370 72701 114375 72705
rect 114461 72701 114494 72705
rect 114494 72701 114517 72705
rect 114603 72701 114618 72705
rect 114618 72701 114659 72705
rect 114745 72701 114798 72705
rect 114798 72701 114801 72705
rect 113325 72581 113381 72615
rect 113467 72581 113523 72615
rect 113609 72581 113665 72615
rect 113751 72581 113807 72615
rect 113893 72581 113949 72615
rect 114035 72581 114091 72615
rect 114177 72581 114233 72615
rect 114319 72581 114375 72615
rect 114461 72581 114517 72615
rect 114603 72581 114659 72615
rect 114745 72581 114801 72615
rect 113325 72559 113378 72581
rect 113378 72559 113381 72581
rect 113467 72559 113502 72581
rect 113502 72559 113523 72581
rect 113609 72559 113626 72581
rect 113626 72559 113665 72581
rect 113751 72559 113806 72581
rect 113806 72559 113807 72581
rect 113893 72559 113930 72581
rect 113930 72559 113949 72581
rect 114035 72559 114054 72581
rect 114054 72559 114091 72581
rect 114177 72559 114178 72581
rect 114178 72559 114233 72581
rect 114319 72559 114370 72581
rect 114370 72559 114375 72581
rect 114461 72559 114494 72581
rect 114494 72559 114517 72581
rect 114603 72559 114618 72581
rect 114618 72559 114659 72581
rect 114745 72559 114798 72581
rect 114798 72559 114801 72581
rect 113325 72457 113381 72473
rect 113467 72457 113523 72473
rect 113609 72457 113665 72473
rect 113751 72457 113807 72473
rect 113893 72457 113949 72473
rect 114035 72457 114091 72473
rect 114177 72457 114233 72473
rect 114319 72457 114375 72473
rect 114461 72457 114517 72473
rect 114603 72457 114659 72473
rect 114745 72457 114801 72473
rect 113325 72417 113378 72457
rect 113378 72417 113381 72457
rect 113467 72417 113502 72457
rect 113502 72417 113523 72457
rect 113609 72417 113626 72457
rect 113626 72417 113665 72457
rect 113751 72417 113806 72457
rect 113806 72417 113807 72457
rect 113893 72417 113930 72457
rect 113930 72417 113949 72457
rect 114035 72417 114054 72457
rect 114054 72417 114091 72457
rect 114177 72417 114178 72457
rect 114178 72417 114233 72457
rect 114319 72417 114370 72457
rect 114370 72417 114375 72457
rect 114461 72417 114494 72457
rect 114494 72417 114517 72457
rect 114603 72417 114618 72457
rect 114618 72417 114659 72457
rect 114745 72417 114798 72457
rect 114798 72417 114801 72457
rect 113325 72277 113378 72331
rect 113378 72277 113381 72331
rect 113467 72277 113502 72331
rect 113502 72277 113523 72331
rect 113609 72277 113626 72331
rect 113626 72277 113665 72331
rect 113751 72277 113806 72331
rect 113806 72277 113807 72331
rect 113893 72277 113930 72331
rect 113930 72277 113949 72331
rect 114035 72277 114054 72331
rect 114054 72277 114091 72331
rect 114177 72277 114178 72331
rect 114178 72277 114233 72331
rect 114319 72277 114370 72331
rect 114370 72277 114375 72331
rect 114461 72277 114494 72331
rect 114494 72277 114517 72331
rect 114603 72277 114618 72331
rect 114618 72277 114659 72331
rect 114745 72277 114798 72331
rect 114798 72277 114801 72331
rect 113325 72275 113381 72277
rect 113467 72275 113523 72277
rect 113609 72275 113665 72277
rect 113751 72275 113807 72277
rect 113893 72275 113949 72277
rect 114035 72275 114091 72277
rect 114177 72275 114233 72277
rect 114319 72275 114375 72277
rect 114461 72275 114517 72277
rect 114603 72275 114659 72277
rect 114745 72275 114801 72277
rect 113325 72153 113378 72189
rect 113378 72153 113381 72189
rect 113467 72153 113502 72189
rect 113502 72153 113523 72189
rect 113609 72153 113626 72189
rect 113626 72153 113665 72189
rect 113751 72153 113806 72189
rect 113806 72153 113807 72189
rect 113893 72153 113930 72189
rect 113930 72153 113949 72189
rect 114035 72153 114054 72189
rect 114054 72153 114091 72189
rect 114177 72153 114178 72189
rect 114178 72153 114233 72189
rect 114319 72153 114370 72189
rect 114370 72153 114375 72189
rect 114461 72153 114494 72189
rect 114494 72153 114517 72189
rect 114603 72153 114618 72189
rect 114618 72153 114659 72189
rect 114745 72153 114798 72189
rect 114798 72153 114801 72189
rect 113325 72133 113381 72153
rect 113467 72133 113523 72153
rect 113609 72133 113665 72153
rect 113751 72133 113807 72153
rect 113893 72133 113949 72153
rect 114035 72133 114091 72153
rect 114177 72133 114233 72153
rect 114319 72133 114375 72153
rect 114461 72133 114517 72153
rect 114603 72133 114659 72153
rect 114745 72133 114801 72153
rect 115269 73979 115325 74035
rect 115411 73979 115467 74035
rect 115553 73979 115609 74035
rect 115695 73979 115751 74035
rect 115837 73979 115893 74035
rect 115979 73979 116035 74035
rect 116121 73979 116177 74035
rect 116263 73979 116319 74035
rect 116405 73979 116461 74035
rect 116547 73979 116603 74035
rect 116689 73979 116745 74035
rect 116831 73979 116887 74035
rect 116973 73979 117029 74035
rect 117115 73979 117171 74035
rect 115269 73889 115308 73893
rect 115308 73889 115325 73893
rect 115411 73889 115432 73893
rect 115432 73889 115467 73893
rect 115553 73889 115556 73893
rect 115556 73889 115609 73893
rect 115695 73889 115748 73893
rect 115748 73889 115751 73893
rect 115837 73889 115872 73893
rect 115872 73889 115893 73893
rect 115979 73889 115996 73893
rect 115996 73889 116035 73893
rect 116121 73889 116176 73893
rect 116176 73889 116177 73893
rect 116263 73889 116300 73893
rect 116300 73889 116319 73893
rect 116405 73889 116424 73893
rect 116424 73889 116461 73893
rect 116547 73889 116548 73893
rect 116548 73889 116603 73893
rect 116689 73889 116740 73893
rect 116740 73889 116745 73893
rect 116831 73889 116864 73893
rect 116864 73889 116887 73893
rect 116973 73889 116988 73893
rect 116988 73889 117029 73893
rect 117115 73889 117168 73893
rect 117168 73889 117171 73893
rect 115269 73837 115325 73889
rect 115411 73837 115467 73889
rect 115553 73837 115609 73889
rect 115695 73837 115751 73889
rect 115837 73837 115893 73889
rect 115979 73837 116035 73889
rect 116121 73837 116177 73889
rect 116263 73837 116319 73889
rect 116405 73837 116461 73889
rect 116547 73837 116603 73889
rect 116689 73837 116745 73889
rect 116831 73837 116887 73889
rect 116973 73837 117029 73889
rect 117115 73837 117171 73889
rect 115269 73697 115325 73751
rect 115411 73697 115467 73751
rect 115553 73697 115609 73751
rect 115695 73697 115751 73751
rect 115837 73697 115893 73751
rect 115979 73697 116035 73751
rect 116121 73697 116177 73751
rect 116263 73697 116319 73751
rect 116405 73697 116461 73751
rect 116547 73697 116603 73751
rect 116689 73697 116745 73751
rect 116831 73697 116887 73751
rect 116973 73697 117029 73751
rect 117115 73697 117171 73751
rect 115269 73695 115308 73697
rect 115308 73695 115325 73697
rect 115411 73695 115432 73697
rect 115432 73695 115467 73697
rect 115553 73695 115556 73697
rect 115556 73695 115609 73697
rect 115695 73695 115748 73697
rect 115748 73695 115751 73697
rect 115837 73695 115872 73697
rect 115872 73695 115893 73697
rect 115979 73695 115996 73697
rect 115996 73695 116035 73697
rect 116121 73695 116176 73697
rect 116176 73695 116177 73697
rect 116263 73695 116300 73697
rect 116300 73695 116319 73697
rect 116405 73695 116424 73697
rect 116424 73695 116461 73697
rect 116547 73695 116548 73697
rect 116548 73695 116603 73697
rect 116689 73695 116740 73697
rect 116740 73695 116745 73697
rect 116831 73695 116864 73697
rect 116864 73695 116887 73697
rect 116973 73695 116988 73697
rect 116988 73695 117029 73697
rect 117115 73695 117168 73697
rect 117168 73695 117171 73697
rect 115269 73573 115325 73609
rect 115411 73573 115467 73609
rect 115553 73573 115609 73609
rect 115695 73573 115751 73609
rect 115837 73573 115893 73609
rect 115979 73573 116035 73609
rect 116121 73573 116177 73609
rect 116263 73573 116319 73609
rect 116405 73573 116461 73609
rect 116547 73573 116603 73609
rect 116689 73573 116745 73609
rect 116831 73573 116887 73609
rect 116973 73573 117029 73609
rect 117115 73573 117171 73609
rect 115269 73553 115308 73573
rect 115308 73553 115325 73573
rect 115411 73553 115432 73573
rect 115432 73553 115467 73573
rect 115553 73553 115556 73573
rect 115556 73553 115609 73573
rect 115695 73553 115748 73573
rect 115748 73553 115751 73573
rect 115837 73553 115872 73573
rect 115872 73553 115893 73573
rect 115979 73553 115996 73573
rect 115996 73553 116035 73573
rect 116121 73553 116176 73573
rect 116176 73553 116177 73573
rect 116263 73553 116300 73573
rect 116300 73553 116319 73573
rect 116405 73553 116424 73573
rect 116424 73553 116461 73573
rect 116547 73553 116548 73573
rect 116548 73553 116603 73573
rect 116689 73553 116740 73573
rect 116740 73553 116745 73573
rect 116831 73553 116864 73573
rect 116864 73553 116887 73573
rect 116973 73553 116988 73573
rect 116988 73553 117029 73573
rect 117115 73553 117168 73573
rect 117168 73553 117171 73573
rect 115269 73449 115325 73467
rect 115411 73449 115467 73467
rect 115553 73449 115609 73467
rect 115695 73449 115751 73467
rect 115837 73449 115893 73467
rect 115979 73449 116035 73467
rect 116121 73449 116177 73467
rect 116263 73449 116319 73467
rect 116405 73449 116461 73467
rect 116547 73449 116603 73467
rect 116689 73449 116745 73467
rect 116831 73449 116887 73467
rect 116973 73449 117029 73467
rect 117115 73449 117171 73467
rect 115269 73411 115308 73449
rect 115308 73411 115325 73449
rect 115411 73411 115432 73449
rect 115432 73411 115467 73449
rect 115553 73411 115556 73449
rect 115556 73411 115609 73449
rect 115695 73411 115748 73449
rect 115748 73411 115751 73449
rect 115837 73411 115872 73449
rect 115872 73411 115893 73449
rect 115979 73411 115996 73449
rect 115996 73411 116035 73449
rect 116121 73411 116176 73449
rect 116176 73411 116177 73449
rect 116263 73411 116300 73449
rect 116300 73411 116319 73449
rect 116405 73411 116424 73449
rect 116424 73411 116461 73449
rect 116547 73411 116548 73449
rect 116548 73411 116603 73449
rect 116689 73411 116740 73449
rect 116740 73411 116745 73449
rect 116831 73411 116864 73449
rect 116864 73411 116887 73449
rect 116973 73411 116988 73449
rect 116988 73411 117029 73449
rect 117115 73411 117168 73449
rect 117168 73411 117171 73449
rect 115269 73269 115308 73325
rect 115308 73269 115325 73325
rect 115411 73269 115432 73325
rect 115432 73269 115467 73325
rect 115553 73269 115556 73325
rect 115556 73269 115609 73325
rect 115695 73269 115748 73325
rect 115748 73269 115751 73325
rect 115837 73269 115872 73325
rect 115872 73269 115893 73325
rect 115979 73269 115996 73325
rect 115996 73269 116035 73325
rect 116121 73269 116176 73325
rect 116176 73269 116177 73325
rect 116263 73269 116300 73325
rect 116300 73269 116319 73325
rect 116405 73269 116424 73325
rect 116424 73269 116461 73325
rect 116547 73269 116548 73325
rect 116548 73269 116603 73325
rect 116689 73269 116740 73325
rect 116740 73269 116745 73325
rect 116831 73269 116864 73325
rect 116864 73269 116887 73325
rect 116973 73269 116988 73325
rect 116988 73269 117029 73325
rect 117115 73269 117168 73325
rect 117168 73269 117171 73325
rect 115269 73145 115308 73183
rect 115308 73145 115325 73183
rect 115411 73145 115432 73183
rect 115432 73145 115467 73183
rect 115553 73145 115556 73183
rect 115556 73145 115609 73183
rect 115695 73145 115748 73183
rect 115748 73145 115751 73183
rect 115837 73145 115872 73183
rect 115872 73145 115893 73183
rect 115979 73145 115996 73183
rect 115996 73145 116035 73183
rect 116121 73145 116176 73183
rect 116176 73145 116177 73183
rect 116263 73145 116300 73183
rect 116300 73145 116319 73183
rect 116405 73145 116424 73183
rect 116424 73145 116461 73183
rect 116547 73145 116548 73183
rect 116548 73145 116603 73183
rect 116689 73145 116740 73183
rect 116740 73145 116745 73183
rect 116831 73145 116864 73183
rect 116864 73145 116887 73183
rect 116973 73145 116988 73183
rect 116988 73145 117029 73183
rect 117115 73145 117168 73183
rect 117168 73145 117171 73183
rect 115269 73127 115325 73145
rect 115411 73127 115467 73145
rect 115553 73127 115609 73145
rect 115695 73127 115751 73145
rect 115837 73127 115893 73145
rect 115979 73127 116035 73145
rect 116121 73127 116177 73145
rect 116263 73127 116319 73145
rect 116405 73127 116461 73145
rect 116547 73127 116603 73145
rect 116689 73127 116745 73145
rect 116831 73127 116887 73145
rect 116973 73127 117029 73145
rect 117115 73127 117171 73145
rect 115269 73021 115308 73041
rect 115308 73021 115325 73041
rect 115411 73021 115432 73041
rect 115432 73021 115467 73041
rect 115553 73021 115556 73041
rect 115556 73021 115609 73041
rect 115695 73021 115748 73041
rect 115748 73021 115751 73041
rect 115837 73021 115872 73041
rect 115872 73021 115893 73041
rect 115979 73021 115996 73041
rect 115996 73021 116035 73041
rect 116121 73021 116176 73041
rect 116176 73021 116177 73041
rect 116263 73021 116300 73041
rect 116300 73021 116319 73041
rect 116405 73021 116424 73041
rect 116424 73021 116461 73041
rect 116547 73021 116548 73041
rect 116548 73021 116603 73041
rect 116689 73021 116740 73041
rect 116740 73021 116745 73041
rect 116831 73021 116864 73041
rect 116864 73021 116887 73041
rect 116973 73021 116988 73041
rect 116988 73021 117029 73041
rect 117115 73021 117168 73041
rect 117168 73021 117171 73041
rect 115269 72985 115325 73021
rect 115411 72985 115467 73021
rect 115553 72985 115609 73021
rect 115695 72985 115751 73021
rect 115837 72985 115893 73021
rect 115979 72985 116035 73021
rect 116121 72985 116177 73021
rect 116263 72985 116319 73021
rect 116405 72985 116461 73021
rect 116547 72985 116603 73021
rect 116689 72985 116745 73021
rect 116831 72985 116887 73021
rect 116973 72985 117029 73021
rect 117115 72985 117171 73021
rect 115269 72897 115308 72899
rect 115308 72897 115325 72899
rect 115411 72897 115432 72899
rect 115432 72897 115467 72899
rect 115553 72897 115556 72899
rect 115556 72897 115609 72899
rect 115695 72897 115748 72899
rect 115748 72897 115751 72899
rect 115837 72897 115872 72899
rect 115872 72897 115893 72899
rect 115979 72897 115996 72899
rect 115996 72897 116035 72899
rect 116121 72897 116176 72899
rect 116176 72897 116177 72899
rect 116263 72897 116300 72899
rect 116300 72897 116319 72899
rect 116405 72897 116424 72899
rect 116424 72897 116461 72899
rect 116547 72897 116548 72899
rect 116548 72897 116603 72899
rect 116689 72897 116740 72899
rect 116740 72897 116745 72899
rect 116831 72897 116864 72899
rect 116864 72897 116887 72899
rect 116973 72897 116988 72899
rect 116988 72897 117029 72899
rect 117115 72897 117168 72899
rect 117168 72897 117171 72899
rect 115269 72843 115325 72897
rect 115411 72843 115467 72897
rect 115553 72843 115609 72897
rect 115695 72843 115751 72897
rect 115837 72843 115893 72897
rect 115979 72843 116035 72897
rect 116121 72843 116177 72897
rect 116263 72843 116319 72897
rect 116405 72843 116461 72897
rect 116547 72843 116603 72897
rect 116689 72843 116745 72897
rect 116831 72843 116887 72897
rect 116973 72843 117029 72897
rect 117115 72843 117171 72897
rect 115269 72705 115325 72757
rect 115411 72705 115467 72757
rect 115553 72705 115609 72757
rect 115695 72705 115751 72757
rect 115837 72705 115893 72757
rect 115979 72705 116035 72757
rect 116121 72705 116177 72757
rect 116263 72705 116319 72757
rect 116405 72705 116461 72757
rect 116547 72705 116603 72757
rect 116689 72705 116745 72757
rect 116831 72705 116887 72757
rect 116973 72705 117029 72757
rect 117115 72705 117171 72757
rect 115269 72701 115308 72705
rect 115308 72701 115325 72705
rect 115411 72701 115432 72705
rect 115432 72701 115467 72705
rect 115553 72701 115556 72705
rect 115556 72701 115609 72705
rect 115695 72701 115748 72705
rect 115748 72701 115751 72705
rect 115837 72701 115872 72705
rect 115872 72701 115893 72705
rect 115979 72701 115996 72705
rect 115996 72701 116035 72705
rect 116121 72701 116176 72705
rect 116176 72701 116177 72705
rect 116263 72701 116300 72705
rect 116300 72701 116319 72705
rect 116405 72701 116424 72705
rect 116424 72701 116461 72705
rect 116547 72701 116548 72705
rect 116548 72701 116603 72705
rect 116689 72701 116740 72705
rect 116740 72701 116745 72705
rect 116831 72701 116864 72705
rect 116864 72701 116887 72705
rect 116973 72701 116988 72705
rect 116988 72701 117029 72705
rect 117115 72701 117168 72705
rect 117168 72701 117171 72705
rect 115269 72581 115325 72615
rect 115411 72581 115467 72615
rect 115553 72581 115609 72615
rect 115695 72581 115751 72615
rect 115837 72581 115893 72615
rect 115979 72581 116035 72615
rect 116121 72581 116177 72615
rect 116263 72581 116319 72615
rect 116405 72581 116461 72615
rect 116547 72581 116603 72615
rect 116689 72581 116745 72615
rect 116831 72581 116887 72615
rect 116973 72581 117029 72615
rect 117115 72581 117171 72615
rect 115269 72559 115308 72581
rect 115308 72559 115325 72581
rect 115411 72559 115432 72581
rect 115432 72559 115467 72581
rect 115553 72559 115556 72581
rect 115556 72559 115609 72581
rect 115695 72559 115748 72581
rect 115748 72559 115751 72581
rect 115837 72559 115872 72581
rect 115872 72559 115893 72581
rect 115979 72559 115996 72581
rect 115996 72559 116035 72581
rect 116121 72559 116176 72581
rect 116176 72559 116177 72581
rect 116263 72559 116300 72581
rect 116300 72559 116319 72581
rect 116405 72559 116424 72581
rect 116424 72559 116461 72581
rect 116547 72559 116548 72581
rect 116548 72559 116603 72581
rect 116689 72559 116740 72581
rect 116740 72559 116745 72581
rect 116831 72559 116864 72581
rect 116864 72559 116887 72581
rect 116973 72559 116988 72581
rect 116988 72559 117029 72581
rect 117115 72559 117168 72581
rect 117168 72559 117171 72581
rect 115269 72457 115325 72473
rect 115411 72457 115467 72473
rect 115553 72457 115609 72473
rect 115695 72457 115751 72473
rect 115837 72457 115893 72473
rect 115979 72457 116035 72473
rect 116121 72457 116177 72473
rect 116263 72457 116319 72473
rect 116405 72457 116461 72473
rect 116547 72457 116603 72473
rect 116689 72457 116745 72473
rect 116831 72457 116887 72473
rect 116973 72457 117029 72473
rect 117115 72457 117171 72473
rect 115269 72417 115308 72457
rect 115308 72417 115325 72457
rect 115411 72417 115432 72457
rect 115432 72417 115467 72457
rect 115553 72417 115556 72457
rect 115556 72417 115609 72457
rect 115695 72417 115748 72457
rect 115748 72417 115751 72457
rect 115837 72417 115872 72457
rect 115872 72417 115893 72457
rect 115979 72417 115996 72457
rect 115996 72417 116035 72457
rect 116121 72417 116176 72457
rect 116176 72417 116177 72457
rect 116263 72417 116300 72457
rect 116300 72417 116319 72457
rect 116405 72417 116424 72457
rect 116424 72417 116461 72457
rect 116547 72417 116548 72457
rect 116548 72417 116603 72457
rect 116689 72417 116740 72457
rect 116740 72417 116745 72457
rect 116831 72417 116864 72457
rect 116864 72417 116887 72457
rect 116973 72417 116988 72457
rect 116988 72417 117029 72457
rect 117115 72417 117168 72457
rect 117168 72417 117171 72457
rect 115269 72277 115308 72331
rect 115308 72277 115325 72331
rect 115411 72277 115432 72331
rect 115432 72277 115467 72331
rect 115553 72277 115556 72331
rect 115556 72277 115609 72331
rect 115695 72277 115748 72331
rect 115748 72277 115751 72331
rect 115837 72277 115872 72331
rect 115872 72277 115893 72331
rect 115979 72277 115996 72331
rect 115996 72277 116035 72331
rect 116121 72277 116176 72331
rect 116176 72277 116177 72331
rect 116263 72277 116300 72331
rect 116300 72277 116319 72331
rect 116405 72277 116424 72331
rect 116424 72277 116461 72331
rect 116547 72277 116548 72331
rect 116548 72277 116603 72331
rect 116689 72277 116740 72331
rect 116740 72277 116745 72331
rect 116831 72277 116864 72331
rect 116864 72277 116887 72331
rect 116973 72277 116988 72331
rect 116988 72277 117029 72331
rect 117115 72277 117168 72331
rect 117168 72277 117171 72331
rect 115269 72275 115325 72277
rect 115411 72275 115467 72277
rect 115553 72275 115609 72277
rect 115695 72275 115751 72277
rect 115837 72275 115893 72277
rect 115979 72275 116035 72277
rect 116121 72275 116177 72277
rect 116263 72275 116319 72277
rect 116405 72275 116461 72277
rect 116547 72275 116603 72277
rect 116689 72275 116745 72277
rect 116831 72275 116887 72277
rect 116973 72275 117029 72277
rect 117115 72275 117171 72277
rect 115269 72153 115308 72189
rect 115308 72153 115325 72189
rect 115411 72153 115432 72189
rect 115432 72153 115467 72189
rect 115553 72153 115556 72189
rect 115556 72153 115609 72189
rect 115695 72153 115748 72189
rect 115748 72153 115751 72189
rect 115837 72153 115872 72189
rect 115872 72153 115893 72189
rect 115979 72153 115996 72189
rect 115996 72153 116035 72189
rect 116121 72153 116176 72189
rect 116176 72153 116177 72189
rect 116263 72153 116300 72189
rect 116300 72153 116319 72189
rect 116405 72153 116424 72189
rect 116424 72153 116461 72189
rect 116547 72153 116548 72189
rect 116548 72153 116603 72189
rect 116689 72153 116740 72189
rect 116740 72153 116745 72189
rect 116831 72153 116864 72189
rect 116864 72153 116887 72189
rect 116973 72153 116988 72189
rect 116988 72153 117029 72189
rect 117115 72153 117168 72189
rect 117168 72153 117171 72189
rect 115269 72133 115325 72153
rect 115411 72133 115467 72153
rect 115553 72133 115609 72153
rect 115695 72133 115751 72153
rect 115837 72133 115893 72153
rect 115979 72133 116035 72153
rect 116121 72133 116177 72153
rect 116263 72133 116319 72153
rect 116405 72133 116461 72153
rect 116547 72133 116603 72153
rect 116689 72133 116745 72153
rect 116831 72133 116887 72153
rect 116973 72133 117029 72153
rect 117115 72133 117171 72153
rect 117899 73979 117955 74035
rect 118041 73979 118097 74035
rect 118183 73979 118239 74035
rect 118325 73979 118381 74035
rect 118467 73979 118523 74035
rect 118609 73979 118665 74035
rect 118751 73979 118807 74035
rect 118893 73979 118949 74035
rect 119035 73979 119091 74035
rect 119177 73979 119233 74035
rect 119319 73979 119375 74035
rect 119461 73979 119517 74035
rect 119603 73979 119659 74035
rect 117899 73889 117938 73893
rect 117938 73889 117955 73893
rect 118041 73889 118062 73893
rect 118062 73889 118097 73893
rect 118183 73889 118186 73893
rect 118186 73889 118239 73893
rect 118325 73889 118378 73893
rect 118378 73889 118381 73893
rect 118467 73889 118502 73893
rect 118502 73889 118523 73893
rect 118609 73889 118626 73893
rect 118626 73889 118665 73893
rect 118751 73889 118806 73893
rect 118806 73889 118807 73893
rect 118893 73889 118930 73893
rect 118930 73889 118949 73893
rect 119035 73889 119054 73893
rect 119054 73889 119091 73893
rect 119177 73889 119178 73893
rect 119178 73889 119233 73893
rect 119319 73889 119370 73893
rect 119370 73889 119375 73893
rect 119461 73889 119494 73893
rect 119494 73889 119517 73893
rect 119603 73889 119618 73893
rect 119618 73889 119659 73893
rect 117899 73837 117955 73889
rect 118041 73837 118097 73889
rect 118183 73837 118239 73889
rect 118325 73837 118381 73889
rect 118467 73837 118523 73889
rect 118609 73837 118665 73889
rect 118751 73837 118807 73889
rect 118893 73837 118949 73889
rect 119035 73837 119091 73889
rect 119177 73837 119233 73889
rect 119319 73837 119375 73889
rect 119461 73837 119517 73889
rect 119603 73837 119659 73889
rect 117899 73697 117955 73751
rect 118041 73697 118097 73751
rect 118183 73697 118239 73751
rect 118325 73697 118381 73751
rect 118467 73697 118523 73751
rect 118609 73697 118665 73751
rect 118751 73697 118807 73751
rect 118893 73697 118949 73751
rect 119035 73697 119091 73751
rect 119177 73697 119233 73751
rect 119319 73697 119375 73751
rect 119461 73697 119517 73751
rect 119603 73697 119659 73751
rect 117899 73695 117938 73697
rect 117938 73695 117955 73697
rect 118041 73695 118062 73697
rect 118062 73695 118097 73697
rect 118183 73695 118186 73697
rect 118186 73695 118239 73697
rect 118325 73695 118378 73697
rect 118378 73695 118381 73697
rect 118467 73695 118502 73697
rect 118502 73695 118523 73697
rect 118609 73695 118626 73697
rect 118626 73695 118665 73697
rect 118751 73695 118806 73697
rect 118806 73695 118807 73697
rect 118893 73695 118930 73697
rect 118930 73695 118949 73697
rect 119035 73695 119054 73697
rect 119054 73695 119091 73697
rect 119177 73695 119178 73697
rect 119178 73695 119233 73697
rect 119319 73695 119370 73697
rect 119370 73695 119375 73697
rect 119461 73695 119494 73697
rect 119494 73695 119517 73697
rect 119603 73695 119618 73697
rect 119618 73695 119659 73697
rect 117899 73573 117955 73609
rect 118041 73573 118097 73609
rect 118183 73573 118239 73609
rect 118325 73573 118381 73609
rect 118467 73573 118523 73609
rect 118609 73573 118665 73609
rect 118751 73573 118807 73609
rect 118893 73573 118949 73609
rect 119035 73573 119091 73609
rect 119177 73573 119233 73609
rect 119319 73573 119375 73609
rect 119461 73573 119517 73609
rect 119603 73573 119659 73609
rect 117899 73553 117938 73573
rect 117938 73553 117955 73573
rect 118041 73553 118062 73573
rect 118062 73553 118097 73573
rect 118183 73553 118186 73573
rect 118186 73553 118239 73573
rect 118325 73553 118378 73573
rect 118378 73553 118381 73573
rect 118467 73553 118502 73573
rect 118502 73553 118523 73573
rect 118609 73553 118626 73573
rect 118626 73553 118665 73573
rect 118751 73553 118806 73573
rect 118806 73553 118807 73573
rect 118893 73553 118930 73573
rect 118930 73553 118949 73573
rect 119035 73553 119054 73573
rect 119054 73553 119091 73573
rect 119177 73553 119178 73573
rect 119178 73553 119233 73573
rect 119319 73553 119370 73573
rect 119370 73553 119375 73573
rect 119461 73553 119494 73573
rect 119494 73553 119517 73573
rect 119603 73553 119618 73573
rect 119618 73553 119659 73573
rect 117899 73449 117955 73467
rect 118041 73449 118097 73467
rect 118183 73449 118239 73467
rect 118325 73449 118381 73467
rect 118467 73449 118523 73467
rect 118609 73449 118665 73467
rect 118751 73449 118807 73467
rect 118893 73449 118949 73467
rect 119035 73449 119091 73467
rect 119177 73449 119233 73467
rect 119319 73449 119375 73467
rect 119461 73449 119517 73467
rect 119603 73449 119659 73467
rect 117899 73411 117938 73449
rect 117938 73411 117955 73449
rect 118041 73411 118062 73449
rect 118062 73411 118097 73449
rect 118183 73411 118186 73449
rect 118186 73411 118239 73449
rect 118325 73411 118378 73449
rect 118378 73411 118381 73449
rect 118467 73411 118502 73449
rect 118502 73411 118523 73449
rect 118609 73411 118626 73449
rect 118626 73411 118665 73449
rect 118751 73411 118806 73449
rect 118806 73411 118807 73449
rect 118893 73411 118930 73449
rect 118930 73411 118949 73449
rect 119035 73411 119054 73449
rect 119054 73411 119091 73449
rect 119177 73411 119178 73449
rect 119178 73411 119233 73449
rect 119319 73411 119370 73449
rect 119370 73411 119375 73449
rect 119461 73411 119494 73449
rect 119494 73411 119517 73449
rect 119603 73411 119618 73449
rect 119618 73411 119659 73449
rect 117899 73269 117938 73325
rect 117938 73269 117955 73325
rect 118041 73269 118062 73325
rect 118062 73269 118097 73325
rect 118183 73269 118186 73325
rect 118186 73269 118239 73325
rect 118325 73269 118378 73325
rect 118378 73269 118381 73325
rect 118467 73269 118502 73325
rect 118502 73269 118523 73325
rect 118609 73269 118626 73325
rect 118626 73269 118665 73325
rect 118751 73269 118806 73325
rect 118806 73269 118807 73325
rect 118893 73269 118930 73325
rect 118930 73269 118949 73325
rect 119035 73269 119054 73325
rect 119054 73269 119091 73325
rect 119177 73269 119178 73325
rect 119178 73269 119233 73325
rect 119319 73269 119370 73325
rect 119370 73269 119375 73325
rect 119461 73269 119494 73325
rect 119494 73269 119517 73325
rect 119603 73269 119618 73325
rect 119618 73269 119659 73325
rect 117899 73145 117938 73183
rect 117938 73145 117955 73183
rect 118041 73145 118062 73183
rect 118062 73145 118097 73183
rect 118183 73145 118186 73183
rect 118186 73145 118239 73183
rect 118325 73145 118378 73183
rect 118378 73145 118381 73183
rect 118467 73145 118502 73183
rect 118502 73145 118523 73183
rect 118609 73145 118626 73183
rect 118626 73145 118665 73183
rect 118751 73145 118806 73183
rect 118806 73145 118807 73183
rect 118893 73145 118930 73183
rect 118930 73145 118949 73183
rect 119035 73145 119054 73183
rect 119054 73145 119091 73183
rect 119177 73145 119178 73183
rect 119178 73145 119233 73183
rect 119319 73145 119370 73183
rect 119370 73145 119375 73183
rect 119461 73145 119494 73183
rect 119494 73145 119517 73183
rect 119603 73145 119618 73183
rect 119618 73145 119659 73183
rect 117899 73127 117955 73145
rect 118041 73127 118097 73145
rect 118183 73127 118239 73145
rect 118325 73127 118381 73145
rect 118467 73127 118523 73145
rect 118609 73127 118665 73145
rect 118751 73127 118807 73145
rect 118893 73127 118949 73145
rect 119035 73127 119091 73145
rect 119177 73127 119233 73145
rect 119319 73127 119375 73145
rect 119461 73127 119517 73145
rect 119603 73127 119659 73145
rect 117899 73021 117938 73041
rect 117938 73021 117955 73041
rect 118041 73021 118062 73041
rect 118062 73021 118097 73041
rect 118183 73021 118186 73041
rect 118186 73021 118239 73041
rect 118325 73021 118378 73041
rect 118378 73021 118381 73041
rect 118467 73021 118502 73041
rect 118502 73021 118523 73041
rect 118609 73021 118626 73041
rect 118626 73021 118665 73041
rect 118751 73021 118806 73041
rect 118806 73021 118807 73041
rect 118893 73021 118930 73041
rect 118930 73021 118949 73041
rect 119035 73021 119054 73041
rect 119054 73021 119091 73041
rect 119177 73021 119178 73041
rect 119178 73021 119233 73041
rect 119319 73021 119370 73041
rect 119370 73021 119375 73041
rect 119461 73021 119494 73041
rect 119494 73021 119517 73041
rect 119603 73021 119618 73041
rect 119618 73021 119659 73041
rect 117899 72985 117955 73021
rect 118041 72985 118097 73021
rect 118183 72985 118239 73021
rect 118325 72985 118381 73021
rect 118467 72985 118523 73021
rect 118609 72985 118665 73021
rect 118751 72985 118807 73021
rect 118893 72985 118949 73021
rect 119035 72985 119091 73021
rect 119177 72985 119233 73021
rect 119319 72985 119375 73021
rect 119461 72985 119517 73021
rect 119603 72985 119659 73021
rect 117899 72897 117938 72899
rect 117938 72897 117955 72899
rect 118041 72897 118062 72899
rect 118062 72897 118097 72899
rect 118183 72897 118186 72899
rect 118186 72897 118239 72899
rect 118325 72897 118378 72899
rect 118378 72897 118381 72899
rect 118467 72897 118502 72899
rect 118502 72897 118523 72899
rect 118609 72897 118626 72899
rect 118626 72897 118665 72899
rect 118751 72897 118806 72899
rect 118806 72897 118807 72899
rect 118893 72897 118930 72899
rect 118930 72897 118949 72899
rect 119035 72897 119054 72899
rect 119054 72897 119091 72899
rect 119177 72897 119178 72899
rect 119178 72897 119233 72899
rect 119319 72897 119370 72899
rect 119370 72897 119375 72899
rect 119461 72897 119494 72899
rect 119494 72897 119517 72899
rect 119603 72897 119618 72899
rect 119618 72897 119659 72899
rect 117899 72843 117955 72897
rect 118041 72843 118097 72897
rect 118183 72843 118239 72897
rect 118325 72843 118381 72897
rect 118467 72843 118523 72897
rect 118609 72843 118665 72897
rect 118751 72843 118807 72897
rect 118893 72843 118949 72897
rect 119035 72843 119091 72897
rect 119177 72843 119233 72897
rect 119319 72843 119375 72897
rect 119461 72843 119517 72897
rect 119603 72843 119659 72897
rect 117899 72705 117955 72757
rect 118041 72705 118097 72757
rect 118183 72705 118239 72757
rect 118325 72705 118381 72757
rect 118467 72705 118523 72757
rect 118609 72705 118665 72757
rect 118751 72705 118807 72757
rect 118893 72705 118949 72757
rect 119035 72705 119091 72757
rect 119177 72705 119233 72757
rect 119319 72705 119375 72757
rect 119461 72705 119517 72757
rect 119603 72705 119659 72757
rect 117899 72701 117938 72705
rect 117938 72701 117955 72705
rect 118041 72701 118062 72705
rect 118062 72701 118097 72705
rect 118183 72701 118186 72705
rect 118186 72701 118239 72705
rect 118325 72701 118378 72705
rect 118378 72701 118381 72705
rect 118467 72701 118502 72705
rect 118502 72701 118523 72705
rect 118609 72701 118626 72705
rect 118626 72701 118665 72705
rect 118751 72701 118806 72705
rect 118806 72701 118807 72705
rect 118893 72701 118930 72705
rect 118930 72701 118949 72705
rect 119035 72701 119054 72705
rect 119054 72701 119091 72705
rect 119177 72701 119178 72705
rect 119178 72701 119233 72705
rect 119319 72701 119370 72705
rect 119370 72701 119375 72705
rect 119461 72701 119494 72705
rect 119494 72701 119517 72705
rect 119603 72701 119618 72705
rect 119618 72701 119659 72705
rect 117899 72581 117955 72615
rect 118041 72581 118097 72615
rect 118183 72581 118239 72615
rect 118325 72581 118381 72615
rect 118467 72581 118523 72615
rect 118609 72581 118665 72615
rect 118751 72581 118807 72615
rect 118893 72581 118949 72615
rect 119035 72581 119091 72615
rect 119177 72581 119233 72615
rect 119319 72581 119375 72615
rect 119461 72581 119517 72615
rect 119603 72581 119659 72615
rect 117899 72559 117938 72581
rect 117938 72559 117955 72581
rect 118041 72559 118062 72581
rect 118062 72559 118097 72581
rect 118183 72559 118186 72581
rect 118186 72559 118239 72581
rect 118325 72559 118378 72581
rect 118378 72559 118381 72581
rect 118467 72559 118502 72581
rect 118502 72559 118523 72581
rect 118609 72559 118626 72581
rect 118626 72559 118665 72581
rect 118751 72559 118806 72581
rect 118806 72559 118807 72581
rect 118893 72559 118930 72581
rect 118930 72559 118949 72581
rect 119035 72559 119054 72581
rect 119054 72559 119091 72581
rect 119177 72559 119178 72581
rect 119178 72559 119233 72581
rect 119319 72559 119370 72581
rect 119370 72559 119375 72581
rect 119461 72559 119494 72581
rect 119494 72559 119517 72581
rect 119603 72559 119618 72581
rect 119618 72559 119659 72581
rect 117899 72457 117955 72473
rect 118041 72457 118097 72473
rect 118183 72457 118239 72473
rect 118325 72457 118381 72473
rect 118467 72457 118523 72473
rect 118609 72457 118665 72473
rect 118751 72457 118807 72473
rect 118893 72457 118949 72473
rect 119035 72457 119091 72473
rect 119177 72457 119233 72473
rect 119319 72457 119375 72473
rect 119461 72457 119517 72473
rect 119603 72457 119659 72473
rect 117899 72417 117938 72457
rect 117938 72417 117955 72457
rect 118041 72417 118062 72457
rect 118062 72417 118097 72457
rect 118183 72417 118186 72457
rect 118186 72417 118239 72457
rect 118325 72417 118378 72457
rect 118378 72417 118381 72457
rect 118467 72417 118502 72457
rect 118502 72417 118523 72457
rect 118609 72417 118626 72457
rect 118626 72417 118665 72457
rect 118751 72417 118806 72457
rect 118806 72417 118807 72457
rect 118893 72417 118930 72457
rect 118930 72417 118949 72457
rect 119035 72417 119054 72457
rect 119054 72417 119091 72457
rect 119177 72417 119178 72457
rect 119178 72417 119233 72457
rect 119319 72417 119370 72457
rect 119370 72417 119375 72457
rect 119461 72417 119494 72457
rect 119494 72417 119517 72457
rect 119603 72417 119618 72457
rect 119618 72417 119659 72457
rect 117899 72277 117938 72331
rect 117938 72277 117955 72331
rect 118041 72277 118062 72331
rect 118062 72277 118097 72331
rect 118183 72277 118186 72331
rect 118186 72277 118239 72331
rect 118325 72277 118378 72331
rect 118378 72277 118381 72331
rect 118467 72277 118502 72331
rect 118502 72277 118523 72331
rect 118609 72277 118626 72331
rect 118626 72277 118665 72331
rect 118751 72277 118806 72331
rect 118806 72277 118807 72331
rect 118893 72277 118930 72331
rect 118930 72277 118949 72331
rect 119035 72277 119054 72331
rect 119054 72277 119091 72331
rect 119177 72277 119178 72331
rect 119178 72277 119233 72331
rect 119319 72277 119370 72331
rect 119370 72277 119375 72331
rect 119461 72277 119494 72331
rect 119494 72277 119517 72331
rect 119603 72277 119618 72331
rect 119618 72277 119659 72331
rect 117899 72275 117955 72277
rect 118041 72275 118097 72277
rect 118183 72275 118239 72277
rect 118325 72275 118381 72277
rect 118467 72275 118523 72277
rect 118609 72275 118665 72277
rect 118751 72275 118807 72277
rect 118893 72275 118949 72277
rect 119035 72275 119091 72277
rect 119177 72275 119233 72277
rect 119319 72275 119375 72277
rect 119461 72275 119517 72277
rect 119603 72275 119659 72277
rect 117899 72153 117938 72189
rect 117938 72153 117955 72189
rect 118041 72153 118062 72189
rect 118062 72153 118097 72189
rect 118183 72153 118186 72189
rect 118186 72153 118239 72189
rect 118325 72153 118378 72189
rect 118378 72153 118381 72189
rect 118467 72153 118502 72189
rect 118502 72153 118523 72189
rect 118609 72153 118626 72189
rect 118626 72153 118665 72189
rect 118751 72153 118806 72189
rect 118806 72153 118807 72189
rect 118893 72153 118930 72189
rect 118930 72153 118949 72189
rect 119035 72153 119054 72189
rect 119054 72153 119091 72189
rect 119177 72153 119178 72189
rect 119178 72153 119233 72189
rect 119319 72153 119370 72189
rect 119370 72153 119375 72189
rect 119461 72153 119494 72189
rect 119494 72153 119517 72189
rect 119603 72153 119618 72189
rect 119618 72153 119659 72189
rect 117899 72133 117955 72153
rect 118041 72133 118097 72153
rect 118183 72133 118239 72153
rect 118325 72133 118381 72153
rect 118467 72133 118523 72153
rect 118609 72133 118665 72153
rect 118751 72133 118807 72153
rect 118893 72133 118949 72153
rect 119035 72133 119091 72153
rect 119177 72133 119233 72153
rect 119319 72133 119375 72153
rect 119461 72133 119517 72153
rect 119603 72133 119659 72153
rect 270343 73979 270399 74035
rect 270485 73979 270541 74035
rect 270627 73979 270683 74035
rect 270769 73979 270825 74035
rect 270911 73979 270967 74035
rect 271053 73979 271109 74035
rect 271195 73979 271251 74035
rect 271337 73979 271393 74035
rect 271479 73979 271535 74035
rect 271621 73979 271677 74035
rect 271763 73979 271819 74035
rect 271905 73979 271961 74035
rect 272047 73979 272103 74035
rect 270343 73889 270382 73893
rect 270382 73889 270399 73893
rect 270485 73889 270506 73893
rect 270506 73889 270541 73893
rect 270627 73889 270630 73893
rect 270630 73889 270683 73893
rect 270769 73889 270822 73893
rect 270822 73889 270825 73893
rect 270911 73889 270946 73893
rect 270946 73889 270967 73893
rect 271053 73889 271070 73893
rect 271070 73889 271109 73893
rect 271195 73889 271250 73893
rect 271250 73889 271251 73893
rect 271337 73889 271374 73893
rect 271374 73889 271393 73893
rect 271479 73889 271498 73893
rect 271498 73889 271535 73893
rect 271621 73889 271622 73893
rect 271622 73889 271677 73893
rect 271763 73889 271814 73893
rect 271814 73889 271819 73893
rect 271905 73889 271938 73893
rect 271938 73889 271961 73893
rect 272047 73889 272062 73893
rect 272062 73889 272103 73893
rect 270343 73837 270399 73889
rect 270485 73837 270541 73889
rect 270627 73837 270683 73889
rect 270769 73837 270825 73889
rect 270911 73837 270967 73889
rect 271053 73837 271109 73889
rect 271195 73837 271251 73889
rect 271337 73837 271393 73889
rect 271479 73837 271535 73889
rect 271621 73837 271677 73889
rect 271763 73837 271819 73889
rect 271905 73837 271961 73889
rect 272047 73837 272103 73889
rect 270343 73697 270399 73751
rect 270485 73697 270541 73751
rect 270627 73697 270683 73751
rect 270769 73697 270825 73751
rect 270911 73697 270967 73751
rect 271053 73697 271109 73751
rect 271195 73697 271251 73751
rect 271337 73697 271393 73751
rect 271479 73697 271535 73751
rect 271621 73697 271677 73751
rect 271763 73697 271819 73751
rect 271905 73697 271961 73751
rect 272047 73697 272103 73751
rect 270343 73695 270382 73697
rect 270382 73695 270399 73697
rect 270485 73695 270506 73697
rect 270506 73695 270541 73697
rect 270627 73695 270630 73697
rect 270630 73695 270683 73697
rect 270769 73695 270822 73697
rect 270822 73695 270825 73697
rect 270911 73695 270946 73697
rect 270946 73695 270967 73697
rect 271053 73695 271070 73697
rect 271070 73695 271109 73697
rect 271195 73695 271250 73697
rect 271250 73695 271251 73697
rect 271337 73695 271374 73697
rect 271374 73695 271393 73697
rect 271479 73695 271498 73697
rect 271498 73695 271535 73697
rect 271621 73695 271622 73697
rect 271622 73695 271677 73697
rect 271763 73695 271814 73697
rect 271814 73695 271819 73697
rect 271905 73695 271938 73697
rect 271938 73695 271961 73697
rect 272047 73695 272062 73697
rect 272062 73695 272103 73697
rect 270343 73573 270399 73609
rect 270485 73573 270541 73609
rect 270627 73573 270683 73609
rect 270769 73573 270825 73609
rect 270911 73573 270967 73609
rect 271053 73573 271109 73609
rect 271195 73573 271251 73609
rect 271337 73573 271393 73609
rect 271479 73573 271535 73609
rect 271621 73573 271677 73609
rect 271763 73573 271819 73609
rect 271905 73573 271961 73609
rect 272047 73573 272103 73609
rect 270343 73553 270382 73573
rect 270382 73553 270399 73573
rect 270485 73553 270506 73573
rect 270506 73553 270541 73573
rect 270627 73553 270630 73573
rect 270630 73553 270683 73573
rect 270769 73553 270822 73573
rect 270822 73553 270825 73573
rect 270911 73553 270946 73573
rect 270946 73553 270967 73573
rect 271053 73553 271070 73573
rect 271070 73553 271109 73573
rect 271195 73553 271250 73573
rect 271250 73553 271251 73573
rect 271337 73553 271374 73573
rect 271374 73553 271393 73573
rect 271479 73553 271498 73573
rect 271498 73553 271535 73573
rect 271621 73553 271622 73573
rect 271622 73553 271677 73573
rect 271763 73553 271814 73573
rect 271814 73553 271819 73573
rect 271905 73553 271938 73573
rect 271938 73553 271961 73573
rect 272047 73553 272062 73573
rect 272062 73553 272103 73573
rect 270343 73449 270399 73467
rect 270485 73449 270541 73467
rect 270627 73449 270683 73467
rect 270769 73449 270825 73467
rect 270911 73449 270967 73467
rect 271053 73449 271109 73467
rect 271195 73449 271251 73467
rect 271337 73449 271393 73467
rect 271479 73449 271535 73467
rect 271621 73449 271677 73467
rect 271763 73449 271819 73467
rect 271905 73449 271961 73467
rect 272047 73449 272103 73467
rect 270343 73411 270382 73449
rect 270382 73411 270399 73449
rect 270485 73411 270506 73449
rect 270506 73411 270541 73449
rect 270627 73411 270630 73449
rect 270630 73411 270683 73449
rect 270769 73411 270822 73449
rect 270822 73411 270825 73449
rect 270911 73411 270946 73449
rect 270946 73411 270967 73449
rect 271053 73411 271070 73449
rect 271070 73411 271109 73449
rect 271195 73411 271250 73449
rect 271250 73411 271251 73449
rect 271337 73411 271374 73449
rect 271374 73411 271393 73449
rect 271479 73411 271498 73449
rect 271498 73411 271535 73449
rect 271621 73411 271622 73449
rect 271622 73411 271677 73449
rect 271763 73411 271814 73449
rect 271814 73411 271819 73449
rect 271905 73411 271938 73449
rect 271938 73411 271961 73449
rect 272047 73411 272062 73449
rect 272062 73411 272103 73449
rect 270343 73269 270382 73325
rect 270382 73269 270399 73325
rect 270485 73269 270506 73325
rect 270506 73269 270541 73325
rect 270627 73269 270630 73325
rect 270630 73269 270683 73325
rect 270769 73269 270822 73325
rect 270822 73269 270825 73325
rect 270911 73269 270946 73325
rect 270946 73269 270967 73325
rect 271053 73269 271070 73325
rect 271070 73269 271109 73325
rect 271195 73269 271250 73325
rect 271250 73269 271251 73325
rect 271337 73269 271374 73325
rect 271374 73269 271393 73325
rect 271479 73269 271498 73325
rect 271498 73269 271535 73325
rect 271621 73269 271622 73325
rect 271622 73269 271677 73325
rect 271763 73269 271814 73325
rect 271814 73269 271819 73325
rect 271905 73269 271938 73325
rect 271938 73269 271961 73325
rect 272047 73269 272062 73325
rect 272062 73269 272103 73325
rect 270343 73145 270382 73183
rect 270382 73145 270399 73183
rect 270485 73145 270506 73183
rect 270506 73145 270541 73183
rect 270627 73145 270630 73183
rect 270630 73145 270683 73183
rect 270769 73145 270822 73183
rect 270822 73145 270825 73183
rect 270911 73145 270946 73183
rect 270946 73145 270967 73183
rect 271053 73145 271070 73183
rect 271070 73145 271109 73183
rect 271195 73145 271250 73183
rect 271250 73145 271251 73183
rect 271337 73145 271374 73183
rect 271374 73145 271393 73183
rect 271479 73145 271498 73183
rect 271498 73145 271535 73183
rect 271621 73145 271622 73183
rect 271622 73145 271677 73183
rect 271763 73145 271814 73183
rect 271814 73145 271819 73183
rect 271905 73145 271938 73183
rect 271938 73145 271961 73183
rect 272047 73145 272062 73183
rect 272062 73145 272103 73183
rect 270343 73127 270399 73145
rect 270485 73127 270541 73145
rect 270627 73127 270683 73145
rect 270769 73127 270825 73145
rect 270911 73127 270967 73145
rect 271053 73127 271109 73145
rect 271195 73127 271251 73145
rect 271337 73127 271393 73145
rect 271479 73127 271535 73145
rect 271621 73127 271677 73145
rect 271763 73127 271819 73145
rect 271905 73127 271961 73145
rect 272047 73127 272103 73145
rect 270343 73021 270382 73041
rect 270382 73021 270399 73041
rect 270485 73021 270506 73041
rect 270506 73021 270541 73041
rect 270627 73021 270630 73041
rect 270630 73021 270683 73041
rect 270769 73021 270822 73041
rect 270822 73021 270825 73041
rect 270911 73021 270946 73041
rect 270946 73021 270967 73041
rect 271053 73021 271070 73041
rect 271070 73021 271109 73041
rect 271195 73021 271250 73041
rect 271250 73021 271251 73041
rect 271337 73021 271374 73041
rect 271374 73021 271393 73041
rect 271479 73021 271498 73041
rect 271498 73021 271535 73041
rect 271621 73021 271622 73041
rect 271622 73021 271677 73041
rect 271763 73021 271814 73041
rect 271814 73021 271819 73041
rect 271905 73021 271938 73041
rect 271938 73021 271961 73041
rect 272047 73021 272062 73041
rect 272062 73021 272103 73041
rect 270343 72985 270399 73021
rect 270485 72985 270541 73021
rect 270627 72985 270683 73021
rect 270769 72985 270825 73021
rect 270911 72985 270967 73021
rect 271053 72985 271109 73021
rect 271195 72985 271251 73021
rect 271337 72985 271393 73021
rect 271479 72985 271535 73021
rect 271621 72985 271677 73021
rect 271763 72985 271819 73021
rect 271905 72985 271961 73021
rect 272047 72985 272103 73021
rect 270343 72897 270382 72899
rect 270382 72897 270399 72899
rect 270485 72897 270506 72899
rect 270506 72897 270541 72899
rect 270627 72897 270630 72899
rect 270630 72897 270683 72899
rect 270769 72897 270822 72899
rect 270822 72897 270825 72899
rect 270911 72897 270946 72899
rect 270946 72897 270967 72899
rect 271053 72897 271070 72899
rect 271070 72897 271109 72899
rect 271195 72897 271250 72899
rect 271250 72897 271251 72899
rect 271337 72897 271374 72899
rect 271374 72897 271393 72899
rect 271479 72897 271498 72899
rect 271498 72897 271535 72899
rect 271621 72897 271622 72899
rect 271622 72897 271677 72899
rect 271763 72897 271814 72899
rect 271814 72897 271819 72899
rect 271905 72897 271938 72899
rect 271938 72897 271961 72899
rect 272047 72897 272062 72899
rect 272062 72897 272103 72899
rect 270343 72843 270399 72897
rect 270485 72843 270541 72897
rect 270627 72843 270683 72897
rect 270769 72843 270825 72897
rect 270911 72843 270967 72897
rect 271053 72843 271109 72897
rect 271195 72843 271251 72897
rect 271337 72843 271393 72897
rect 271479 72843 271535 72897
rect 271621 72843 271677 72897
rect 271763 72843 271819 72897
rect 271905 72843 271961 72897
rect 272047 72843 272103 72897
rect 270343 72705 270399 72757
rect 270485 72705 270541 72757
rect 270627 72705 270683 72757
rect 270769 72705 270825 72757
rect 270911 72705 270967 72757
rect 271053 72705 271109 72757
rect 271195 72705 271251 72757
rect 271337 72705 271393 72757
rect 271479 72705 271535 72757
rect 271621 72705 271677 72757
rect 271763 72705 271819 72757
rect 271905 72705 271961 72757
rect 272047 72705 272103 72757
rect 270343 72701 270382 72705
rect 270382 72701 270399 72705
rect 270485 72701 270506 72705
rect 270506 72701 270541 72705
rect 270627 72701 270630 72705
rect 270630 72701 270683 72705
rect 270769 72701 270822 72705
rect 270822 72701 270825 72705
rect 270911 72701 270946 72705
rect 270946 72701 270967 72705
rect 271053 72701 271070 72705
rect 271070 72701 271109 72705
rect 271195 72701 271250 72705
rect 271250 72701 271251 72705
rect 271337 72701 271374 72705
rect 271374 72701 271393 72705
rect 271479 72701 271498 72705
rect 271498 72701 271535 72705
rect 271621 72701 271622 72705
rect 271622 72701 271677 72705
rect 271763 72701 271814 72705
rect 271814 72701 271819 72705
rect 271905 72701 271938 72705
rect 271938 72701 271961 72705
rect 272047 72701 272062 72705
rect 272062 72701 272103 72705
rect 270343 72581 270399 72615
rect 270485 72581 270541 72615
rect 270627 72581 270683 72615
rect 270769 72581 270825 72615
rect 270911 72581 270967 72615
rect 271053 72581 271109 72615
rect 271195 72581 271251 72615
rect 271337 72581 271393 72615
rect 271479 72581 271535 72615
rect 271621 72581 271677 72615
rect 271763 72581 271819 72615
rect 271905 72581 271961 72615
rect 272047 72581 272103 72615
rect 270343 72559 270382 72581
rect 270382 72559 270399 72581
rect 270485 72559 270506 72581
rect 270506 72559 270541 72581
rect 270627 72559 270630 72581
rect 270630 72559 270683 72581
rect 270769 72559 270822 72581
rect 270822 72559 270825 72581
rect 270911 72559 270946 72581
rect 270946 72559 270967 72581
rect 271053 72559 271070 72581
rect 271070 72559 271109 72581
rect 271195 72559 271250 72581
rect 271250 72559 271251 72581
rect 271337 72559 271374 72581
rect 271374 72559 271393 72581
rect 271479 72559 271498 72581
rect 271498 72559 271535 72581
rect 271621 72559 271622 72581
rect 271622 72559 271677 72581
rect 271763 72559 271814 72581
rect 271814 72559 271819 72581
rect 271905 72559 271938 72581
rect 271938 72559 271961 72581
rect 272047 72559 272062 72581
rect 272062 72559 272103 72581
rect 270343 72457 270399 72473
rect 270485 72457 270541 72473
rect 270627 72457 270683 72473
rect 270769 72457 270825 72473
rect 270911 72457 270967 72473
rect 271053 72457 271109 72473
rect 271195 72457 271251 72473
rect 271337 72457 271393 72473
rect 271479 72457 271535 72473
rect 271621 72457 271677 72473
rect 271763 72457 271819 72473
rect 271905 72457 271961 72473
rect 272047 72457 272103 72473
rect 270343 72417 270382 72457
rect 270382 72417 270399 72457
rect 270485 72417 270506 72457
rect 270506 72417 270541 72457
rect 270627 72417 270630 72457
rect 270630 72417 270683 72457
rect 270769 72417 270822 72457
rect 270822 72417 270825 72457
rect 270911 72417 270946 72457
rect 270946 72417 270967 72457
rect 271053 72417 271070 72457
rect 271070 72417 271109 72457
rect 271195 72417 271250 72457
rect 271250 72417 271251 72457
rect 271337 72417 271374 72457
rect 271374 72417 271393 72457
rect 271479 72417 271498 72457
rect 271498 72417 271535 72457
rect 271621 72417 271622 72457
rect 271622 72417 271677 72457
rect 271763 72417 271814 72457
rect 271814 72417 271819 72457
rect 271905 72417 271938 72457
rect 271938 72417 271961 72457
rect 272047 72417 272062 72457
rect 272062 72417 272103 72457
rect 270343 72277 270382 72331
rect 270382 72277 270399 72331
rect 270485 72277 270506 72331
rect 270506 72277 270541 72331
rect 270627 72277 270630 72331
rect 270630 72277 270683 72331
rect 270769 72277 270822 72331
rect 270822 72277 270825 72331
rect 270911 72277 270946 72331
rect 270946 72277 270967 72331
rect 271053 72277 271070 72331
rect 271070 72277 271109 72331
rect 271195 72277 271250 72331
rect 271250 72277 271251 72331
rect 271337 72277 271374 72331
rect 271374 72277 271393 72331
rect 271479 72277 271498 72331
rect 271498 72277 271535 72331
rect 271621 72277 271622 72331
rect 271622 72277 271677 72331
rect 271763 72277 271814 72331
rect 271814 72277 271819 72331
rect 271905 72277 271938 72331
rect 271938 72277 271961 72331
rect 272047 72277 272062 72331
rect 272062 72277 272103 72331
rect 270343 72275 270399 72277
rect 270485 72275 270541 72277
rect 270627 72275 270683 72277
rect 270769 72275 270825 72277
rect 270911 72275 270967 72277
rect 271053 72275 271109 72277
rect 271195 72275 271251 72277
rect 271337 72275 271393 72277
rect 271479 72275 271535 72277
rect 271621 72275 271677 72277
rect 271763 72275 271819 72277
rect 271905 72275 271961 72277
rect 272047 72275 272103 72277
rect 270343 72153 270382 72189
rect 270382 72153 270399 72189
rect 270485 72153 270506 72189
rect 270506 72153 270541 72189
rect 270627 72153 270630 72189
rect 270630 72153 270683 72189
rect 270769 72153 270822 72189
rect 270822 72153 270825 72189
rect 270911 72153 270946 72189
rect 270946 72153 270967 72189
rect 271053 72153 271070 72189
rect 271070 72153 271109 72189
rect 271195 72153 271250 72189
rect 271250 72153 271251 72189
rect 271337 72153 271374 72189
rect 271374 72153 271393 72189
rect 271479 72153 271498 72189
rect 271498 72153 271535 72189
rect 271621 72153 271622 72189
rect 271622 72153 271677 72189
rect 271763 72153 271814 72189
rect 271814 72153 271819 72189
rect 271905 72153 271938 72189
rect 271938 72153 271961 72189
rect 272047 72153 272062 72189
rect 272062 72153 272103 72189
rect 270343 72133 270399 72153
rect 270485 72133 270541 72153
rect 270627 72133 270683 72153
rect 270769 72133 270825 72153
rect 270911 72133 270967 72153
rect 271053 72133 271109 72153
rect 271195 72133 271251 72153
rect 271337 72133 271393 72153
rect 271479 72133 271535 72153
rect 271621 72133 271677 72153
rect 271763 72133 271819 72153
rect 271905 72133 271961 72153
rect 272047 72133 272103 72153
rect 272823 73979 272879 74035
rect 272965 73979 273021 74035
rect 273107 73979 273163 74035
rect 273249 73979 273305 74035
rect 273391 73979 273447 74035
rect 273533 73979 273589 74035
rect 273675 73979 273731 74035
rect 273817 73979 273873 74035
rect 273959 73979 274015 74035
rect 274101 73979 274157 74035
rect 274243 73979 274299 74035
rect 274385 73979 274441 74035
rect 274527 73979 274583 74035
rect 274669 73979 274725 74035
rect 272823 73889 272862 73893
rect 272862 73889 272879 73893
rect 272965 73889 272986 73893
rect 272986 73889 273021 73893
rect 273107 73889 273110 73893
rect 273110 73889 273163 73893
rect 273249 73889 273302 73893
rect 273302 73889 273305 73893
rect 273391 73889 273426 73893
rect 273426 73889 273447 73893
rect 273533 73889 273550 73893
rect 273550 73889 273589 73893
rect 273675 73889 273730 73893
rect 273730 73889 273731 73893
rect 273817 73889 273854 73893
rect 273854 73889 273873 73893
rect 273959 73889 273978 73893
rect 273978 73889 274015 73893
rect 274101 73889 274102 73893
rect 274102 73889 274157 73893
rect 274243 73889 274294 73893
rect 274294 73889 274299 73893
rect 274385 73889 274418 73893
rect 274418 73889 274441 73893
rect 274527 73889 274542 73893
rect 274542 73889 274583 73893
rect 274669 73889 274722 73893
rect 274722 73889 274725 73893
rect 272823 73837 272879 73889
rect 272965 73837 273021 73889
rect 273107 73837 273163 73889
rect 273249 73837 273305 73889
rect 273391 73837 273447 73889
rect 273533 73837 273589 73889
rect 273675 73837 273731 73889
rect 273817 73837 273873 73889
rect 273959 73837 274015 73889
rect 274101 73837 274157 73889
rect 274243 73837 274299 73889
rect 274385 73837 274441 73889
rect 274527 73837 274583 73889
rect 274669 73837 274725 73889
rect 272823 73697 272879 73751
rect 272965 73697 273021 73751
rect 273107 73697 273163 73751
rect 273249 73697 273305 73751
rect 273391 73697 273447 73751
rect 273533 73697 273589 73751
rect 273675 73697 273731 73751
rect 273817 73697 273873 73751
rect 273959 73697 274015 73751
rect 274101 73697 274157 73751
rect 274243 73697 274299 73751
rect 274385 73697 274441 73751
rect 274527 73697 274583 73751
rect 274669 73697 274725 73751
rect 272823 73695 272862 73697
rect 272862 73695 272879 73697
rect 272965 73695 272986 73697
rect 272986 73695 273021 73697
rect 273107 73695 273110 73697
rect 273110 73695 273163 73697
rect 273249 73695 273302 73697
rect 273302 73695 273305 73697
rect 273391 73695 273426 73697
rect 273426 73695 273447 73697
rect 273533 73695 273550 73697
rect 273550 73695 273589 73697
rect 273675 73695 273730 73697
rect 273730 73695 273731 73697
rect 273817 73695 273854 73697
rect 273854 73695 273873 73697
rect 273959 73695 273978 73697
rect 273978 73695 274015 73697
rect 274101 73695 274102 73697
rect 274102 73695 274157 73697
rect 274243 73695 274294 73697
rect 274294 73695 274299 73697
rect 274385 73695 274418 73697
rect 274418 73695 274441 73697
rect 274527 73695 274542 73697
rect 274542 73695 274583 73697
rect 274669 73695 274722 73697
rect 274722 73695 274725 73697
rect 272823 73573 272879 73609
rect 272965 73573 273021 73609
rect 273107 73573 273163 73609
rect 273249 73573 273305 73609
rect 273391 73573 273447 73609
rect 273533 73573 273589 73609
rect 273675 73573 273731 73609
rect 273817 73573 273873 73609
rect 273959 73573 274015 73609
rect 274101 73573 274157 73609
rect 274243 73573 274299 73609
rect 274385 73573 274441 73609
rect 274527 73573 274583 73609
rect 274669 73573 274725 73609
rect 272823 73553 272862 73573
rect 272862 73553 272879 73573
rect 272965 73553 272986 73573
rect 272986 73553 273021 73573
rect 273107 73553 273110 73573
rect 273110 73553 273163 73573
rect 273249 73553 273302 73573
rect 273302 73553 273305 73573
rect 273391 73553 273426 73573
rect 273426 73553 273447 73573
rect 273533 73553 273550 73573
rect 273550 73553 273589 73573
rect 273675 73553 273730 73573
rect 273730 73553 273731 73573
rect 273817 73553 273854 73573
rect 273854 73553 273873 73573
rect 273959 73553 273978 73573
rect 273978 73553 274015 73573
rect 274101 73553 274102 73573
rect 274102 73553 274157 73573
rect 274243 73553 274294 73573
rect 274294 73553 274299 73573
rect 274385 73553 274418 73573
rect 274418 73553 274441 73573
rect 274527 73553 274542 73573
rect 274542 73553 274583 73573
rect 274669 73553 274722 73573
rect 274722 73553 274725 73573
rect 272823 73449 272879 73467
rect 272965 73449 273021 73467
rect 273107 73449 273163 73467
rect 273249 73449 273305 73467
rect 273391 73449 273447 73467
rect 273533 73449 273589 73467
rect 273675 73449 273731 73467
rect 273817 73449 273873 73467
rect 273959 73449 274015 73467
rect 274101 73449 274157 73467
rect 274243 73449 274299 73467
rect 274385 73449 274441 73467
rect 274527 73449 274583 73467
rect 274669 73449 274725 73467
rect 272823 73411 272862 73449
rect 272862 73411 272879 73449
rect 272965 73411 272986 73449
rect 272986 73411 273021 73449
rect 273107 73411 273110 73449
rect 273110 73411 273163 73449
rect 273249 73411 273302 73449
rect 273302 73411 273305 73449
rect 273391 73411 273426 73449
rect 273426 73411 273447 73449
rect 273533 73411 273550 73449
rect 273550 73411 273589 73449
rect 273675 73411 273730 73449
rect 273730 73411 273731 73449
rect 273817 73411 273854 73449
rect 273854 73411 273873 73449
rect 273959 73411 273978 73449
rect 273978 73411 274015 73449
rect 274101 73411 274102 73449
rect 274102 73411 274157 73449
rect 274243 73411 274294 73449
rect 274294 73411 274299 73449
rect 274385 73411 274418 73449
rect 274418 73411 274441 73449
rect 274527 73411 274542 73449
rect 274542 73411 274583 73449
rect 274669 73411 274722 73449
rect 274722 73411 274725 73449
rect 272823 73269 272862 73325
rect 272862 73269 272879 73325
rect 272965 73269 272986 73325
rect 272986 73269 273021 73325
rect 273107 73269 273110 73325
rect 273110 73269 273163 73325
rect 273249 73269 273302 73325
rect 273302 73269 273305 73325
rect 273391 73269 273426 73325
rect 273426 73269 273447 73325
rect 273533 73269 273550 73325
rect 273550 73269 273589 73325
rect 273675 73269 273730 73325
rect 273730 73269 273731 73325
rect 273817 73269 273854 73325
rect 273854 73269 273873 73325
rect 273959 73269 273978 73325
rect 273978 73269 274015 73325
rect 274101 73269 274102 73325
rect 274102 73269 274157 73325
rect 274243 73269 274294 73325
rect 274294 73269 274299 73325
rect 274385 73269 274418 73325
rect 274418 73269 274441 73325
rect 274527 73269 274542 73325
rect 274542 73269 274583 73325
rect 274669 73269 274722 73325
rect 274722 73269 274725 73325
rect 272823 73145 272862 73183
rect 272862 73145 272879 73183
rect 272965 73145 272986 73183
rect 272986 73145 273021 73183
rect 273107 73145 273110 73183
rect 273110 73145 273163 73183
rect 273249 73145 273302 73183
rect 273302 73145 273305 73183
rect 273391 73145 273426 73183
rect 273426 73145 273447 73183
rect 273533 73145 273550 73183
rect 273550 73145 273589 73183
rect 273675 73145 273730 73183
rect 273730 73145 273731 73183
rect 273817 73145 273854 73183
rect 273854 73145 273873 73183
rect 273959 73145 273978 73183
rect 273978 73145 274015 73183
rect 274101 73145 274102 73183
rect 274102 73145 274157 73183
rect 274243 73145 274294 73183
rect 274294 73145 274299 73183
rect 274385 73145 274418 73183
rect 274418 73145 274441 73183
rect 274527 73145 274542 73183
rect 274542 73145 274583 73183
rect 274669 73145 274722 73183
rect 274722 73145 274725 73183
rect 272823 73127 272879 73145
rect 272965 73127 273021 73145
rect 273107 73127 273163 73145
rect 273249 73127 273305 73145
rect 273391 73127 273447 73145
rect 273533 73127 273589 73145
rect 273675 73127 273731 73145
rect 273817 73127 273873 73145
rect 273959 73127 274015 73145
rect 274101 73127 274157 73145
rect 274243 73127 274299 73145
rect 274385 73127 274441 73145
rect 274527 73127 274583 73145
rect 274669 73127 274725 73145
rect 272823 73021 272862 73041
rect 272862 73021 272879 73041
rect 272965 73021 272986 73041
rect 272986 73021 273021 73041
rect 273107 73021 273110 73041
rect 273110 73021 273163 73041
rect 273249 73021 273302 73041
rect 273302 73021 273305 73041
rect 273391 73021 273426 73041
rect 273426 73021 273447 73041
rect 273533 73021 273550 73041
rect 273550 73021 273589 73041
rect 273675 73021 273730 73041
rect 273730 73021 273731 73041
rect 273817 73021 273854 73041
rect 273854 73021 273873 73041
rect 273959 73021 273978 73041
rect 273978 73021 274015 73041
rect 274101 73021 274102 73041
rect 274102 73021 274157 73041
rect 274243 73021 274294 73041
rect 274294 73021 274299 73041
rect 274385 73021 274418 73041
rect 274418 73021 274441 73041
rect 274527 73021 274542 73041
rect 274542 73021 274583 73041
rect 274669 73021 274722 73041
rect 274722 73021 274725 73041
rect 272823 72985 272879 73021
rect 272965 72985 273021 73021
rect 273107 72985 273163 73021
rect 273249 72985 273305 73021
rect 273391 72985 273447 73021
rect 273533 72985 273589 73021
rect 273675 72985 273731 73021
rect 273817 72985 273873 73021
rect 273959 72985 274015 73021
rect 274101 72985 274157 73021
rect 274243 72985 274299 73021
rect 274385 72985 274441 73021
rect 274527 72985 274583 73021
rect 274669 72985 274725 73021
rect 272823 72897 272862 72899
rect 272862 72897 272879 72899
rect 272965 72897 272986 72899
rect 272986 72897 273021 72899
rect 273107 72897 273110 72899
rect 273110 72897 273163 72899
rect 273249 72897 273302 72899
rect 273302 72897 273305 72899
rect 273391 72897 273426 72899
rect 273426 72897 273447 72899
rect 273533 72897 273550 72899
rect 273550 72897 273589 72899
rect 273675 72897 273730 72899
rect 273730 72897 273731 72899
rect 273817 72897 273854 72899
rect 273854 72897 273873 72899
rect 273959 72897 273978 72899
rect 273978 72897 274015 72899
rect 274101 72897 274102 72899
rect 274102 72897 274157 72899
rect 274243 72897 274294 72899
rect 274294 72897 274299 72899
rect 274385 72897 274418 72899
rect 274418 72897 274441 72899
rect 274527 72897 274542 72899
rect 274542 72897 274583 72899
rect 274669 72897 274722 72899
rect 274722 72897 274725 72899
rect 272823 72843 272879 72897
rect 272965 72843 273021 72897
rect 273107 72843 273163 72897
rect 273249 72843 273305 72897
rect 273391 72843 273447 72897
rect 273533 72843 273589 72897
rect 273675 72843 273731 72897
rect 273817 72843 273873 72897
rect 273959 72843 274015 72897
rect 274101 72843 274157 72897
rect 274243 72843 274299 72897
rect 274385 72843 274441 72897
rect 274527 72843 274583 72897
rect 274669 72843 274725 72897
rect 272823 72705 272879 72757
rect 272965 72705 273021 72757
rect 273107 72705 273163 72757
rect 273249 72705 273305 72757
rect 273391 72705 273447 72757
rect 273533 72705 273589 72757
rect 273675 72705 273731 72757
rect 273817 72705 273873 72757
rect 273959 72705 274015 72757
rect 274101 72705 274157 72757
rect 274243 72705 274299 72757
rect 274385 72705 274441 72757
rect 274527 72705 274583 72757
rect 274669 72705 274725 72757
rect 272823 72701 272862 72705
rect 272862 72701 272879 72705
rect 272965 72701 272986 72705
rect 272986 72701 273021 72705
rect 273107 72701 273110 72705
rect 273110 72701 273163 72705
rect 273249 72701 273302 72705
rect 273302 72701 273305 72705
rect 273391 72701 273426 72705
rect 273426 72701 273447 72705
rect 273533 72701 273550 72705
rect 273550 72701 273589 72705
rect 273675 72701 273730 72705
rect 273730 72701 273731 72705
rect 273817 72701 273854 72705
rect 273854 72701 273873 72705
rect 273959 72701 273978 72705
rect 273978 72701 274015 72705
rect 274101 72701 274102 72705
rect 274102 72701 274157 72705
rect 274243 72701 274294 72705
rect 274294 72701 274299 72705
rect 274385 72701 274418 72705
rect 274418 72701 274441 72705
rect 274527 72701 274542 72705
rect 274542 72701 274583 72705
rect 274669 72701 274722 72705
rect 274722 72701 274725 72705
rect 272823 72581 272879 72615
rect 272965 72581 273021 72615
rect 273107 72581 273163 72615
rect 273249 72581 273305 72615
rect 273391 72581 273447 72615
rect 273533 72581 273589 72615
rect 273675 72581 273731 72615
rect 273817 72581 273873 72615
rect 273959 72581 274015 72615
rect 274101 72581 274157 72615
rect 274243 72581 274299 72615
rect 274385 72581 274441 72615
rect 274527 72581 274583 72615
rect 274669 72581 274725 72615
rect 272823 72559 272862 72581
rect 272862 72559 272879 72581
rect 272965 72559 272986 72581
rect 272986 72559 273021 72581
rect 273107 72559 273110 72581
rect 273110 72559 273163 72581
rect 273249 72559 273302 72581
rect 273302 72559 273305 72581
rect 273391 72559 273426 72581
rect 273426 72559 273447 72581
rect 273533 72559 273550 72581
rect 273550 72559 273589 72581
rect 273675 72559 273730 72581
rect 273730 72559 273731 72581
rect 273817 72559 273854 72581
rect 273854 72559 273873 72581
rect 273959 72559 273978 72581
rect 273978 72559 274015 72581
rect 274101 72559 274102 72581
rect 274102 72559 274157 72581
rect 274243 72559 274294 72581
rect 274294 72559 274299 72581
rect 274385 72559 274418 72581
rect 274418 72559 274441 72581
rect 274527 72559 274542 72581
rect 274542 72559 274583 72581
rect 274669 72559 274722 72581
rect 274722 72559 274725 72581
rect 272823 72457 272879 72473
rect 272965 72457 273021 72473
rect 273107 72457 273163 72473
rect 273249 72457 273305 72473
rect 273391 72457 273447 72473
rect 273533 72457 273589 72473
rect 273675 72457 273731 72473
rect 273817 72457 273873 72473
rect 273959 72457 274015 72473
rect 274101 72457 274157 72473
rect 274243 72457 274299 72473
rect 274385 72457 274441 72473
rect 274527 72457 274583 72473
rect 274669 72457 274725 72473
rect 272823 72417 272862 72457
rect 272862 72417 272879 72457
rect 272965 72417 272986 72457
rect 272986 72417 273021 72457
rect 273107 72417 273110 72457
rect 273110 72417 273163 72457
rect 273249 72417 273302 72457
rect 273302 72417 273305 72457
rect 273391 72417 273426 72457
rect 273426 72417 273447 72457
rect 273533 72417 273550 72457
rect 273550 72417 273589 72457
rect 273675 72417 273730 72457
rect 273730 72417 273731 72457
rect 273817 72417 273854 72457
rect 273854 72417 273873 72457
rect 273959 72417 273978 72457
rect 273978 72417 274015 72457
rect 274101 72417 274102 72457
rect 274102 72417 274157 72457
rect 274243 72417 274294 72457
rect 274294 72417 274299 72457
rect 274385 72417 274418 72457
rect 274418 72417 274441 72457
rect 274527 72417 274542 72457
rect 274542 72417 274583 72457
rect 274669 72417 274722 72457
rect 274722 72417 274725 72457
rect 272823 72277 272862 72331
rect 272862 72277 272879 72331
rect 272965 72277 272986 72331
rect 272986 72277 273021 72331
rect 273107 72277 273110 72331
rect 273110 72277 273163 72331
rect 273249 72277 273302 72331
rect 273302 72277 273305 72331
rect 273391 72277 273426 72331
rect 273426 72277 273447 72331
rect 273533 72277 273550 72331
rect 273550 72277 273589 72331
rect 273675 72277 273730 72331
rect 273730 72277 273731 72331
rect 273817 72277 273854 72331
rect 273854 72277 273873 72331
rect 273959 72277 273978 72331
rect 273978 72277 274015 72331
rect 274101 72277 274102 72331
rect 274102 72277 274157 72331
rect 274243 72277 274294 72331
rect 274294 72277 274299 72331
rect 274385 72277 274418 72331
rect 274418 72277 274441 72331
rect 274527 72277 274542 72331
rect 274542 72277 274583 72331
rect 274669 72277 274722 72331
rect 274722 72277 274725 72331
rect 272823 72275 272879 72277
rect 272965 72275 273021 72277
rect 273107 72275 273163 72277
rect 273249 72275 273305 72277
rect 273391 72275 273447 72277
rect 273533 72275 273589 72277
rect 273675 72275 273731 72277
rect 273817 72275 273873 72277
rect 273959 72275 274015 72277
rect 274101 72275 274157 72277
rect 274243 72275 274299 72277
rect 274385 72275 274441 72277
rect 274527 72275 274583 72277
rect 274669 72275 274725 72277
rect 272823 72153 272862 72189
rect 272862 72153 272879 72189
rect 272965 72153 272986 72189
rect 272986 72153 273021 72189
rect 273107 72153 273110 72189
rect 273110 72153 273163 72189
rect 273249 72153 273302 72189
rect 273302 72153 273305 72189
rect 273391 72153 273426 72189
rect 273426 72153 273447 72189
rect 273533 72153 273550 72189
rect 273550 72153 273589 72189
rect 273675 72153 273730 72189
rect 273730 72153 273731 72189
rect 273817 72153 273854 72189
rect 273854 72153 273873 72189
rect 273959 72153 273978 72189
rect 273978 72153 274015 72189
rect 274101 72153 274102 72189
rect 274102 72153 274157 72189
rect 274243 72153 274294 72189
rect 274294 72153 274299 72189
rect 274385 72153 274418 72189
rect 274418 72153 274441 72189
rect 274527 72153 274542 72189
rect 274542 72153 274583 72189
rect 274669 72153 274722 72189
rect 274722 72153 274725 72189
rect 272823 72133 272879 72153
rect 272965 72133 273021 72153
rect 273107 72133 273163 72153
rect 273249 72133 273305 72153
rect 273391 72133 273447 72153
rect 273533 72133 273589 72153
rect 273675 72133 273731 72153
rect 273817 72133 273873 72153
rect 273959 72133 274015 72153
rect 274101 72133 274157 72153
rect 274243 72133 274299 72153
rect 274385 72133 274441 72153
rect 274527 72133 274583 72153
rect 274669 72133 274725 72153
rect 275193 73979 275249 74035
rect 275335 73979 275391 74035
rect 275477 73979 275533 74035
rect 275619 73979 275675 74035
rect 275761 73979 275817 74035
rect 275903 73979 275959 74035
rect 276045 73979 276101 74035
rect 276187 73979 276243 74035
rect 276329 73979 276385 74035
rect 276471 73979 276527 74035
rect 276613 73979 276669 74035
rect 276755 73979 276811 74035
rect 276897 73979 276953 74035
rect 277039 73979 277095 74035
rect 275193 73889 275232 73893
rect 275232 73889 275249 73893
rect 275335 73889 275356 73893
rect 275356 73889 275391 73893
rect 275477 73889 275480 73893
rect 275480 73889 275533 73893
rect 275619 73889 275672 73893
rect 275672 73889 275675 73893
rect 275761 73889 275796 73893
rect 275796 73889 275817 73893
rect 275903 73889 275920 73893
rect 275920 73889 275959 73893
rect 276045 73889 276100 73893
rect 276100 73889 276101 73893
rect 276187 73889 276224 73893
rect 276224 73889 276243 73893
rect 276329 73889 276348 73893
rect 276348 73889 276385 73893
rect 276471 73889 276472 73893
rect 276472 73889 276527 73893
rect 276613 73889 276664 73893
rect 276664 73889 276669 73893
rect 276755 73889 276788 73893
rect 276788 73889 276811 73893
rect 276897 73889 276912 73893
rect 276912 73889 276953 73893
rect 277039 73889 277092 73893
rect 277092 73889 277095 73893
rect 275193 73837 275249 73889
rect 275335 73837 275391 73889
rect 275477 73837 275533 73889
rect 275619 73837 275675 73889
rect 275761 73837 275817 73889
rect 275903 73837 275959 73889
rect 276045 73837 276101 73889
rect 276187 73837 276243 73889
rect 276329 73837 276385 73889
rect 276471 73837 276527 73889
rect 276613 73837 276669 73889
rect 276755 73837 276811 73889
rect 276897 73837 276953 73889
rect 277039 73837 277095 73889
rect 275193 73697 275249 73751
rect 275335 73697 275391 73751
rect 275477 73697 275533 73751
rect 275619 73697 275675 73751
rect 275761 73697 275817 73751
rect 275903 73697 275959 73751
rect 276045 73697 276101 73751
rect 276187 73697 276243 73751
rect 276329 73697 276385 73751
rect 276471 73697 276527 73751
rect 276613 73697 276669 73751
rect 276755 73697 276811 73751
rect 276897 73697 276953 73751
rect 277039 73697 277095 73751
rect 275193 73695 275232 73697
rect 275232 73695 275249 73697
rect 275335 73695 275356 73697
rect 275356 73695 275391 73697
rect 275477 73695 275480 73697
rect 275480 73695 275533 73697
rect 275619 73695 275672 73697
rect 275672 73695 275675 73697
rect 275761 73695 275796 73697
rect 275796 73695 275817 73697
rect 275903 73695 275920 73697
rect 275920 73695 275959 73697
rect 276045 73695 276100 73697
rect 276100 73695 276101 73697
rect 276187 73695 276224 73697
rect 276224 73695 276243 73697
rect 276329 73695 276348 73697
rect 276348 73695 276385 73697
rect 276471 73695 276472 73697
rect 276472 73695 276527 73697
rect 276613 73695 276664 73697
rect 276664 73695 276669 73697
rect 276755 73695 276788 73697
rect 276788 73695 276811 73697
rect 276897 73695 276912 73697
rect 276912 73695 276953 73697
rect 277039 73695 277092 73697
rect 277092 73695 277095 73697
rect 275193 73573 275249 73609
rect 275335 73573 275391 73609
rect 275477 73573 275533 73609
rect 275619 73573 275675 73609
rect 275761 73573 275817 73609
rect 275903 73573 275959 73609
rect 276045 73573 276101 73609
rect 276187 73573 276243 73609
rect 276329 73573 276385 73609
rect 276471 73573 276527 73609
rect 276613 73573 276669 73609
rect 276755 73573 276811 73609
rect 276897 73573 276953 73609
rect 277039 73573 277095 73609
rect 275193 73553 275232 73573
rect 275232 73553 275249 73573
rect 275335 73553 275356 73573
rect 275356 73553 275391 73573
rect 275477 73553 275480 73573
rect 275480 73553 275533 73573
rect 275619 73553 275672 73573
rect 275672 73553 275675 73573
rect 275761 73553 275796 73573
rect 275796 73553 275817 73573
rect 275903 73553 275920 73573
rect 275920 73553 275959 73573
rect 276045 73553 276100 73573
rect 276100 73553 276101 73573
rect 276187 73553 276224 73573
rect 276224 73553 276243 73573
rect 276329 73553 276348 73573
rect 276348 73553 276385 73573
rect 276471 73553 276472 73573
rect 276472 73553 276527 73573
rect 276613 73553 276664 73573
rect 276664 73553 276669 73573
rect 276755 73553 276788 73573
rect 276788 73553 276811 73573
rect 276897 73553 276912 73573
rect 276912 73553 276953 73573
rect 277039 73553 277092 73573
rect 277092 73553 277095 73573
rect 275193 73449 275249 73467
rect 275335 73449 275391 73467
rect 275477 73449 275533 73467
rect 275619 73449 275675 73467
rect 275761 73449 275817 73467
rect 275903 73449 275959 73467
rect 276045 73449 276101 73467
rect 276187 73449 276243 73467
rect 276329 73449 276385 73467
rect 276471 73449 276527 73467
rect 276613 73449 276669 73467
rect 276755 73449 276811 73467
rect 276897 73449 276953 73467
rect 277039 73449 277095 73467
rect 275193 73411 275232 73449
rect 275232 73411 275249 73449
rect 275335 73411 275356 73449
rect 275356 73411 275391 73449
rect 275477 73411 275480 73449
rect 275480 73411 275533 73449
rect 275619 73411 275672 73449
rect 275672 73411 275675 73449
rect 275761 73411 275796 73449
rect 275796 73411 275817 73449
rect 275903 73411 275920 73449
rect 275920 73411 275959 73449
rect 276045 73411 276100 73449
rect 276100 73411 276101 73449
rect 276187 73411 276224 73449
rect 276224 73411 276243 73449
rect 276329 73411 276348 73449
rect 276348 73411 276385 73449
rect 276471 73411 276472 73449
rect 276472 73411 276527 73449
rect 276613 73411 276664 73449
rect 276664 73411 276669 73449
rect 276755 73411 276788 73449
rect 276788 73411 276811 73449
rect 276897 73411 276912 73449
rect 276912 73411 276953 73449
rect 277039 73411 277092 73449
rect 277092 73411 277095 73449
rect 275193 73269 275232 73325
rect 275232 73269 275249 73325
rect 275335 73269 275356 73325
rect 275356 73269 275391 73325
rect 275477 73269 275480 73325
rect 275480 73269 275533 73325
rect 275619 73269 275672 73325
rect 275672 73269 275675 73325
rect 275761 73269 275796 73325
rect 275796 73269 275817 73325
rect 275903 73269 275920 73325
rect 275920 73269 275959 73325
rect 276045 73269 276100 73325
rect 276100 73269 276101 73325
rect 276187 73269 276224 73325
rect 276224 73269 276243 73325
rect 276329 73269 276348 73325
rect 276348 73269 276385 73325
rect 276471 73269 276472 73325
rect 276472 73269 276527 73325
rect 276613 73269 276664 73325
rect 276664 73269 276669 73325
rect 276755 73269 276788 73325
rect 276788 73269 276811 73325
rect 276897 73269 276912 73325
rect 276912 73269 276953 73325
rect 277039 73269 277092 73325
rect 277092 73269 277095 73325
rect 275193 73145 275232 73183
rect 275232 73145 275249 73183
rect 275335 73145 275356 73183
rect 275356 73145 275391 73183
rect 275477 73145 275480 73183
rect 275480 73145 275533 73183
rect 275619 73145 275672 73183
rect 275672 73145 275675 73183
rect 275761 73145 275796 73183
rect 275796 73145 275817 73183
rect 275903 73145 275920 73183
rect 275920 73145 275959 73183
rect 276045 73145 276100 73183
rect 276100 73145 276101 73183
rect 276187 73145 276224 73183
rect 276224 73145 276243 73183
rect 276329 73145 276348 73183
rect 276348 73145 276385 73183
rect 276471 73145 276472 73183
rect 276472 73145 276527 73183
rect 276613 73145 276664 73183
rect 276664 73145 276669 73183
rect 276755 73145 276788 73183
rect 276788 73145 276811 73183
rect 276897 73145 276912 73183
rect 276912 73145 276953 73183
rect 277039 73145 277092 73183
rect 277092 73145 277095 73183
rect 275193 73127 275249 73145
rect 275335 73127 275391 73145
rect 275477 73127 275533 73145
rect 275619 73127 275675 73145
rect 275761 73127 275817 73145
rect 275903 73127 275959 73145
rect 276045 73127 276101 73145
rect 276187 73127 276243 73145
rect 276329 73127 276385 73145
rect 276471 73127 276527 73145
rect 276613 73127 276669 73145
rect 276755 73127 276811 73145
rect 276897 73127 276953 73145
rect 277039 73127 277095 73145
rect 275193 73021 275232 73041
rect 275232 73021 275249 73041
rect 275335 73021 275356 73041
rect 275356 73021 275391 73041
rect 275477 73021 275480 73041
rect 275480 73021 275533 73041
rect 275619 73021 275672 73041
rect 275672 73021 275675 73041
rect 275761 73021 275796 73041
rect 275796 73021 275817 73041
rect 275903 73021 275920 73041
rect 275920 73021 275959 73041
rect 276045 73021 276100 73041
rect 276100 73021 276101 73041
rect 276187 73021 276224 73041
rect 276224 73021 276243 73041
rect 276329 73021 276348 73041
rect 276348 73021 276385 73041
rect 276471 73021 276472 73041
rect 276472 73021 276527 73041
rect 276613 73021 276664 73041
rect 276664 73021 276669 73041
rect 276755 73021 276788 73041
rect 276788 73021 276811 73041
rect 276897 73021 276912 73041
rect 276912 73021 276953 73041
rect 277039 73021 277092 73041
rect 277092 73021 277095 73041
rect 275193 72985 275249 73021
rect 275335 72985 275391 73021
rect 275477 72985 275533 73021
rect 275619 72985 275675 73021
rect 275761 72985 275817 73021
rect 275903 72985 275959 73021
rect 276045 72985 276101 73021
rect 276187 72985 276243 73021
rect 276329 72985 276385 73021
rect 276471 72985 276527 73021
rect 276613 72985 276669 73021
rect 276755 72985 276811 73021
rect 276897 72985 276953 73021
rect 277039 72985 277095 73021
rect 275193 72897 275232 72899
rect 275232 72897 275249 72899
rect 275335 72897 275356 72899
rect 275356 72897 275391 72899
rect 275477 72897 275480 72899
rect 275480 72897 275533 72899
rect 275619 72897 275672 72899
rect 275672 72897 275675 72899
rect 275761 72897 275796 72899
rect 275796 72897 275817 72899
rect 275903 72897 275920 72899
rect 275920 72897 275959 72899
rect 276045 72897 276100 72899
rect 276100 72897 276101 72899
rect 276187 72897 276224 72899
rect 276224 72897 276243 72899
rect 276329 72897 276348 72899
rect 276348 72897 276385 72899
rect 276471 72897 276472 72899
rect 276472 72897 276527 72899
rect 276613 72897 276664 72899
rect 276664 72897 276669 72899
rect 276755 72897 276788 72899
rect 276788 72897 276811 72899
rect 276897 72897 276912 72899
rect 276912 72897 276953 72899
rect 277039 72897 277092 72899
rect 277092 72897 277095 72899
rect 275193 72843 275249 72897
rect 275335 72843 275391 72897
rect 275477 72843 275533 72897
rect 275619 72843 275675 72897
rect 275761 72843 275817 72897
rect 275903 72843 275959 72897
rect 276045 72843 276101 72897
rect 276187 72843 276243 72897
rect 276329 72843 276385 72897
rect 276471 72843 276527 72897
rect 276613 72843 276669 72897
rect 276755 72843 276811 72897
rect 276897 72843 276953 72897
rect 277039 72843 277095 72897
rect 275193 72705 275249 72757
rect 275335 72705 275391 72757
rect 275477 72705 275533 72757
rect 275619 72705 275675 72757
rect 275761 72705 275817 72757
rect 275903 72705 275959 72757
rect 276045 72705 276101 72757
rect 276187 72705 276243 72757
rect 276329 72705 276385 72757
rect 276471 72705 276527 72757
rect 276613 72705 276669 72757
rect 276755 72705 276811 72757
rect 276897 72705 276953 72757
rect 277039 72705 277095 72757
rect 275193 72701 275232 72705
rect 275232 72701 275249 72705
rect 275335 72701 275356 72705
rect 275356 72701 275391 72705
rect 275477 72701 275480 72705
rect 275480 72701 275533 72705
rect 275619 72701 275672 72705
rect 275672 72701 275675 72705
rect 275761 72701 275796 72705
rect 275796 72701 275817 72705
rect 275903 72701 275920 72705
rect 275920 72701 275959 72705
rect 276045 72701 276100 72705
rect 276100 72701 276101 72705
rect 276187 72701 276224 72705
rect 276224 72701 276243 72705
rect 276329 72701 276348 72705
rect 276348 72701 276385 72705
rect 276471 72701 276472 72705
rect 276472 72701 276527 72705
rect 276613 72701 276664 72705
rect 276664 72701 276669 72705
rect 276755 72701 276788 72705
rect 276788 72701 276811 72705
rect 276897 72701 276912 72705
rect 276912 72701 276953 72705
rect 277039 72701 277092 72705
rect 277092 72701 277095 72705
rect 275193 72581 275249 72615
rect 275335 72581 275391 72615
rect 275477 72581 275533 72615
rect 275619 72581 275675 72615
rect 275761 72581 275817 72615
rect 275903 72581 275959 72615
rect 276045 72581 276101 72615
rect 276187 72581 276243 72615
rect 276329 72581 276385 72615
rect 276471 72581 276527 72615
rect 276613 72581 276669 72615
rect 276755 72581 276811 72615
rect 276897 72581 276953 72615
rect 277039 72581 277095 72615
rect 275193 72559 275232 72581
rect 275232 72559 275249 72581
rect 275335 72559 275356 72581
rect 275356 72559 275391 72581
rect 275477 72559 275480 72581
rect 275480 72559 275533 72581
rect 275619 72559 275672 72581
rect 275672 72559 275675 72581
rect 275761 72559 275796 72581
rect 275796 72559 275817 72581
rect 275903 72559 275920 72581
rect 275920 72559 275959 72581
rect 276045 72559 276100 72581
rect 276100 72559 276101 72581
rect 276187 72559 276224 72581
rect 276224 72559 276243 72581
rect 276329 72559 276348 72581
rect 276348 72559 276385 72581
rect 276471 72559 276472 72581
rect 276472 72559 276527 72581
rect 276613 72559 276664 72581
rect 276664 72559 276669 72581
rect 276755 72559 276788 72581
rect 276788 72559 276811 72581
rect 276897 72559 276912 72581
rect 276912 72559 276953 72581
rect 277039 72559 277092 72581
rect 277092 72559 277095 72581
rect 275193 72457 275249 72473
rect 275335 72457 275391 72473
rect 275477 72457 275533 72473
rect 275619 72457 275675 72473
rect 275761 72457 275817 72473
rect 275903 72457 275959 72473
rect 276045 72457 276101 72473
rect 276187 72457 276243 72473
rect 276329 72457 276385 72473
rect 276471 72457 276527 72473
rect 276613 72457 276669 72473
rect 276755 72457 276811 72473
rect 276897 72457 276953 72473
rect 277039 72457 277095 72473
rect 275193 72417 275232 72457
rect 275232 72417 275249 72457
rect 275335 72417 275356 72457
rect 275356 72417 275391 72457
rect 275477 72417 275480 72457
rect 275480 72417 275533 72457
rect 275619 72417 275672 72457
rect 275672 72417 275675 72457
rect 275761 72417 275796 72457
rect 275796 72417 275817 72457
rect 275903 72417 275920 72457
rect 275920 72417 275959 72457
rect 276045 72417 276100 72457
rect 276100 72417 276101 72457
rect 276187 72417 276224 72457
rect 276224 72417 276243 72457
rect 276329 72417 276348 72457
rect 276348 72417 276385 72457
rect 276471 72417 276472 72457
rect 276472 72417 276527 72457
rect 276613 72417 276664 72457
rect 276664 72417 276669 72457
rect 276755 72417 276788 72457
rect 276788 72417 276811 72457
rect 276897 72417 276912 72457
rect 276912 72417 276953 72457
rect 277039 72417 277092 72457
rect 277092 72417 277095 72457
rect 275193 72277 275232 72331
rect 275232 72277 275249 72331
rect 275335 72277 275356 72331
rect 275356 72277 275391 72331
rect 275477 72277 275480 72331
rect 275480 72277 275533 72331
rect 275619 72277 275672 72331
rect 275672 72277 275675 72331
rect 275761 72277 275796 72331
rect 275796 72277 275817 72331
rect 275903 72277 275920 72331
rect 275920 72277 275959 72331
rect 276045 72277 276100 72331
rect 276100 72277 276101 72331
rect 276187 72277 276224 72331
rect 276224 72277 276243 72331
rect 276329 72277 276348 72331
rect 276348 72277 276385 72331
rect 276471 72277 276472 72331
rect 276472 72277 276527 72331
rect 276613 72277 276664 72331
rect 276664 72277 276669 72331
rect 276755 72277 276788 72331
rect 276788 72277 276811 72331
rect 276897 72277 276912 72331
rect 276912 72277 276953 72331
rect 277039 72277 277092 72331
rect 277092 72277 277095 72331
rect 275193 72275 275249 72277
rect 275335 72275 275391 72277
rect 275477 72275 275533 72277
rect 275619 72275 275675 72277
rect 275761 72275 275817 72277
rect 275903 72275 275959 72277
rect 276045 72275 276101 72277
rect 276187 72275 276243 72277
rect 276329 72275 276385 72277
rect 276471 72275 276527 72277
rect 276613 72275 276669 72277
rect 276755 72275 276811 72277
rect 276897 72275 276953 72277
rect 277039 72275 277095 72277
rect 275193 72153 275232 72189
rect 275232 72153 275249 72189
rect 275335 72153 275356 72189
rect 275356 72153 275391 72189
rect 275477 72153 275480 72189
rect 275480 72153 275533 72189
rect 275619 72153 275672 72189
rect 275672 72153 275675 72189
rect 275761 72153 275796 72189
rect 275796 72153 275817 72189
rect 275903 72153 275920 72189
rect 275920 72153 275959 72189
rect 276045 72153 276100 72189
rect 276100 72153 276101 72189
rect 276187 72153 276224 72189
rect 276224 72153 276243 72189
rect 276329 72153 276348 72189
rect 276348 72153 276385 72189
rect 276471 72153 276472 72189
rect 276472 72153 276527 72189
rect 276613 72153 276664 72189
rect 276664 72153 276669 72189
rect 276755 72153 276788 72189
rect 276788 72153 276811 72189
rect 276897 72153 276912 72189
rect 276912 72153 276953 72189
rect 277039 72153 277092 72189
rect 277092 72153 277095 72189
rect 275193 72133 275249 72153
rect 275335 72133 275391 72153
rect 275477 72133 275533 72153
rect 275619 72133 275675 72153
rect 275761 72133 275817 72153
rect 275903 72133 275959 72153
rect 276045 72133 276101 72153
rect 276187 72133 276243 72153
rect 276329 72133 276385 72153
rect 276471 72133 276527 72153
rect 276613 72133 276669 72153
rect 276755 72133 276811 72153
rect 276897 72133 276953 72153
rect 277039 72133 277095 72153
rect 277899 73979 277955 74035
rect 278041 73979 278097 74035
rect 278183 73979 278239 74035
rect 278325 73979 278381 74035
rect 278467 73979 278523 74035
rect 278609 73979 278665 74035
rect 278751 73979 278807 74035
rect 278893 73979 278949 74035
rect 279035 73979 279091 74035
rect 279177 73979 279233 74035
rect 279319 73979 279375 74035
rect 279461 73979 279517 74035
rect 279603 73979 279659 74035
rect 279745 73979 279801 74035
rect 277899 73889 277938 73893
rect 277938 73889 277955 73893
rect 278041 73889 278062 73893
rect 278062 73889 278097 73893
rect 278183 73889 278186 73893
rect 278186 73889 278239 73893
rect 278325 73889 278378 73893
rect 278378 73889 278381 73893
rect 278467 73889 278502 73893
rect 278502 73889 278523 73893
rect 278609 73889 278626 73893
rect 278626 73889 278665 73893
rect 278751 73889 278806 73893
rect 278806 73889 278807 73893
rect 278893 73889 278930 73893
rect 278930 73889 278949 73893
rect 279035 73889 279054 73893
rect 279054 73889 279091 73893
rect 279177 73889 279178 73893
rect 279178 73889 279233 73893
rect 279319 73889 279370 73893
rect 279370 73889 279375 73893
rect 279461 73889 279494 73893
rect 279494 73889 279517 73893
rect 279603 73889 279618 73893
rect 279618 73889 279659 73893
rect 279745 73889 279798 73893
rect 279798 73889 279801 73893
rect 277899 73837 277955 73889
rect 278041 73837 278097 73889
rect 278183 73837 278239 73889
rect 278325 73837 278381 73889
rect 278467 73837 278523 73889
rect 278609 73837 278665 73889
rect 278751 73837 278807 73889
rect 278893 73837 278949 73889
rect 279035 73837 279091 73889
rect 279177 73837 279233 73889
rect 279319 73837 279375 73889
rect 279461 73837 279517 73889
rect 279603 73837 279659 73889
rect 279745 73837 279801 73889
rect 277899 73697 277955 73751
rect 278041 73697 278097 73751
rect 278183 73697 278239 73751
rect 278325 73697 278381 73751
rect 278467 73697 278523 73751
rect 278609 73697 278665 73751
rect 278751 73697 278807 73751
rect 278893 73697 278949 73751
rect 279035 73697 279091 73751
rect 279177 73697 279233 73751
rect 279319 73697 279375 73751
rect 279461 73697 279517 73751
rect 279603 73697 279659 73751
rect 279745 73697 279801 73751
rect 277899 73695 277938 73697
rect 277938 73695 277955 73697
rect 278041 73695 278062 73697
rect 278062 73695 278097 73697
rect 278183 73695 278186 73697
rect 278186 73695 278239 73697
rect 278325 73695 278378 73697
rect 278378 73695 278381 73697
rect 278467 73695 278502 73697
rect 278502 73695 278523 73697
rect 278609 73695 278626 73697
rect 278626 73695 278665 73697
rect 278751 73695 278806 73697
rect 278806 73695 278807 73697
rect 278893 73695 278930 73697
rect 278930 73695 278949 73697
rect 279035 73695 279054 73697
rect 279054 73695 279091 73697
rect 279177 73695 279178 73697
rect 279178 73695 279233 73697
rect 279319 73695 279370 73697
rect 279370 73695 279375 73697
rect 279461 73695 279494 73697
rect 279494 73695 279517 73697
rect 279603 73695 279618 73697
rect 279618 73695 279659 73697
rect 279745 73695 279798 73697
rect 279798 73695 279801 73697
rect 277899 73573 277955 73609
rect 278041 73573 278097 73609
rect 278183 73573 278239 73609
rect 278325 73573 278381 73609
rect 278467 73573 278523 73609
rect 278609 73573 278665 73609
rect 278751 73573 278807 73609
rect 278893 73573 278949 73609
rect 279035 73573 279091 73609
rect 279177 73573 279233 73609
rect 279319 73573 279375 73609
rect 279461 73573 279517 73609
rect 279603 73573 279659 73609
rect 279745 73573 279801 73609
rect 277899 73553 277938 73573
rect 277938 73553 277955 73573
rect 278041 73553 278062 73573
rect 278062 73553 278097 73573
rect 278183 73553 278186 73573
rect 278186 73553 278239 73573
rect 278325 73553 278378 73573
rect 278378 73553 278381 73573
rect 278467 73553 278502 73573
rect 278502 73553 278523 73573
rect 278609 73553 278626 73573
rect 278626 73553 278665 73573
rect 278751 73553 278806 73573
rect 278806 73553 278807 73573
rect 278893 73553 278930 73573
rect 278930 73553 278949 73573
rect 279035 73553 279054 73573
rect 279054 73553 279091 73573
rect 279177 73553 279178 73573
rect 279178 73553 279233 73573
rect 279319 73553 279370 73573
rect 279370 73553 279375 73573
rect 279461 73553 279494 73573
rect 279494 73553 279517 73573
rect 279603 73553 279618 73573
rect 279618 73553 279659 73573
rect 279745 73553 279798 73573
rect 279798 73553 279801 73573
rect 277899 73449 277955 73467
rect 278041 73449 278097 73467
rect 278183 73449 278239 73467
rect 278325 73449 278381 73467
rect 278467 73449 278523 73467
rect 278609 73449 278665 73467
rect 278751 73449 278807 73467
rect 278893 73449 278949 73467
rect 279035 73449 279091 73467
rect 279177 73449 279233 73467
rect 279319 73449 279375 73467
rect 279461 73449 279517 73467
rect 279603 73449 279659 73467
rect 279745 73449 279801 73467
rect 277899 73411 277938 73449
rect 277938 73411 277955 73449
rect 278041 73411 278062 73449
rect 278062 73411 278097 73449
rect 278183 73411 278186 73449
rect 278186 73411 278239 73449
rect 278325 73411 278378 73449
rect 278378 73411 278381 73449
rect 278467 73411 278502 73449
rect 278502 73411 278523 73449
rect 278609 73411 278626 73449
rect 278626 73411 278665 73449
rect 278751 73411 278806 73449
rect 278806 73411 278807 73449
rect 278893 73411 278930 73449
rect 278930 73411 278949 73449
rect 279035 73411 279054 73449
rect 279054 73411 279091 73449
rect 279177 73411 279178 73449
rect 279178 73411 279233 73449
rect 279319 73411 279370 73449
rect 279370 73411 279375 73449
rect 279461 73411 279494 73449
rect 279494 73411 279517 73449
rect 279603 73411 279618 73449
rect 279618 73411 279659 73449
rect 279745 73411 279798 73449
rect 279798 73411 279801 73449
rect 277899 73269 277938 73325
rect 277938 73269 277955 73325
rect 278041 73269 278062 73325
rect 278062 73269 278097 73325
rect 278183 73269 278186 73325
rect 278186 73269 278239 73325
rect 278325 73269 278378 73325
rect 278378 73269 278381 73325
rect 278467 73269 278502 73325
rect 278502 73269 278523 73325
rect 278609 73269 278626 73325
rect 278626 73269 278665 73325
rect 278751 73269 278806 73325
rect 278806 73269 278807 73325
rect 278893 73269 278930 73325
rect 278930 73269 278949 73325
rect 279035 73269 279054 73325
rect 279054 73269 279091 73325
rect 279177 73269 279178 73325
rect 279178 73269 279233 73325
rect 279319 73269 279370 73325
rect 279370 73269 279375 73325
rect 279461 73269 279494 73325
rect 279494 73269 279517 73325
rect 279603 73269 279618 73325
rect 279618 73269 279659 73325
rect 279745 73269 279798 73325
rect 279798 73269 279801 73325
rect 277899 73145 277938 73183
rect 277938 73145 277955 73183
rect 278041 73145 278062 73183
rect 278062 73145 278097 73183
rect 278183 73145 278186 73183
rect 278186 73145 278239 73183
rect 278325 73145 278378 73183
rect 278378 73145 278381 73183
rect 278467 73145 278502 73183
rect 278502 73145 278523 73183
rect 278609 73145 278626 73183
rect 278626 73145 278665 73183
rect 278751 73145 278806 73183
rect 278806 73145 278807 73183
rect 278893 73145 278930 73183
rect 278930 73145 278949 73183
rect 279035 73145 279054 73183
rect 279054 73145 279091 73183
rect 279177 73145 279178 73183
rect 279178 73145 279233 73183
rect 279319 73145 279370 73183
rect 279370 73145 279375 73183
rect 279461 73145 279494 73183
rect 279494 73145 279517 73183
rect 279603 73145 279618 73183
rect 279618 73145 279659 73183
rect 279745 73145 279798 73183
rect 279798 73145 279801 73183
rect 277899 73127 277955 73145
rect 278041 73127 278097 73145
rect 278183 73127 278239 73145
rect 278325 73127 278381 73145
rect 278467 73127 278523 73145
rect 278609 73127 278665 73145
rect 278751 73127 278807 73145
rect 278893 73127 278949 73145
rect 279035 73127 279091 73145
rect 279177 73127 279233 73145
rect 279319 73127 279375 73145
rect 279461 73127 279517 73145
rect 279603 73127 279659 73145
rect 279745 73127 279801 73145
rect 277899 73021 277938 73041
rect 277938 73021 277955 73041
rect 278041 73021 278062 73041
rect 278062 73021 278097 73041
rect 278183 73021 278186 73041
rect 278186 73021 278239 73041
rect 278325 73021 278378 73041
rect 278378 73021 278381 73041
rect 278467 73021 278502 73041
rect 278502 73021 278523 73041
rect 278609 73021 278626 73041
rect 278626 73021 278665 73041
rect 278751 73021 278806 73041
rect 278806 73021 278807 73041
rect 278893 73021 278930 73041
rect 278930 73021 278949 73041
rect 279035 73021 279054 73041
rect 279054 73021 279091 73041
rect 279177 73021 279178 73041
rect 279178 73021 279233 73041
rect 279319 73021 279370 73041
rect 279370 73021 279375 73041
rect 279461 73021 279494 73041
rect 279494 73021 279517 73041
rect 279603 73021 279618 73041
rect 279618 73021 279659 73041
rect 279745 73021 279798 73041
rect 279798 73021 279801 73041
rect 277899 72985 277955 73021
rect 278041 72985 278097 73021
rect 278183 72985 278239 73021
rect 278325 72985 278381 73021
rect 278467 72985 278523 73021
rect 278609 72985 278665 73021
rect 278751 72985 278807 73021
rect 278893 72985 278949 73021
rect 279035 72985 279091 73021
rect 279177 72985 279233 73021
rect 279319 72985 279375 73021
rect 279461 72985 279517 73021
rect 279603 72985 279659 73021
rect 279745 72985 279801 73021
rect 277899 72897 277938 72899
rect 277938 72897 277955 72899
rect 278041 72897 278062 72899
rect 278062 72897 278097 72899
rect 278183 72897 278186 72899
rect 278186 72897 278239 72899
rect 278325 72897 278378 72899
rect 278378 72897 278381 72899
rect 278467 72897 278502 72899
rect 278502 72897 278523 72899
rect 278609 72897 278626 72899
rect 278626 72897 278665 72899
rect 278751 72897 278806 72899
rect 278806 72897 278807 72899
rect 278893 72897 278930 72899
rect 278930 72897 278949 72899
rect 279035 72897 279054 72899
rect 279054 72897 279091 72899
rect 279177 72897 279178 72899
rect 279178 72897 279233 72899
rect 279319 72897 279370 72899
rect 279370 72897 279375 72899
rect 279461 72897 279494 72899
rect 279494 72897 279517 72899
rect 279603 72897 279618 72899
rect 279618 72897 279659 72899
rect 279745 72897 279798 72899
rect 279798 72897 279801 72899
rect 277899 72843 277955 72897
rect 278041 72843 278097 72897
rect 278183 72843 278239 72897
rect 278325 72843 278381 72897
rect 278467 72843 278523 72897
rect 278609 72843 278665 72897
rect 278751 72843 278807 72897
rect 278893 72843 278949 72897
rect 279035 72843 279091 72897
rect 279177 72843 279233 72897
rect 279319 72843 279375 72897
rect 279461 72843 279517 72897
rect 279603 72843 279659 72897
rect 279745 72843 279801 72897
rect 277899 72705 277955 72757
rect 278041 72705 278097 72757
rect 278183 72705 278239 72757
rect 278325 72705 278381 72757
rect 278467 72705 278523 72757
rect 278609 72705 278665 72757
rect 278751 72705 278807 72757
rect 278893 72705 278949 72757
rect 279035 72705 279091 72757
rect 279177 72705 279233 72757
rect 279319 72705 279375 72757
rect 279461 72705 279517 72757
rect 279603 72705 279659 72757
rect 279745 72705 279801 72757
rect 277899 72701 277938 72705
rect 277938 72701 277955 72705
rect 278041 72701 278062 72705
rect 278062 72701 278097 72705
rect 278183 72701 278186 72705
rect 278186 72701 278239 72705
rect 278325 72701 278378 72705
rect 278378 72701 278381 72705
rect 278467 72701 278502 72705
rect 278502 72701 278523 72705
rect 278609 72701 278626 72705
rect 278626 72701 278665 72705
rect 278751 72701 278806 72705
rect 278806 72701 278807 72705
rect 278893 72701 278930 72705
rect 278930 72701 278949 72705
rect 279035 72701 279054 72705
rect 279054 72701 279091 72705
rect 279177 72701 279178 72705
rect 279178 72701 279233 72705
rect 279319 72701 279370 72705
rect 279370 72701 279375 72705
rect 279461 72701 279494 72705
rect 279494 72701 279517 72705
rect 279603 72701 279618 72705
rect 279618 72701 279659 72705
rect 279745 72701 279798 72705
rect 279798 72701 279801 72705
rect 277899 72581 277955 72615
rect 278041 72581 278097 72615
rect 278183 72581 278239 72615
rect 278325 72581 278381 72615
rect 278467 72581 278523 72615
rect 278609 72581 278665 72615
rect 278751 72581 278807 72615
rect 278893 72581 278949 72615
rect 279035 72581 279091 72615
rect 279177 72581 279233 72615
rect 279319 72581 279375 72615
rect 279461 72581 279517 72615
rect 279603 72581 279659 72615
rect 279745 72581 279801 72615
rect 277899 72559 277938 72581
rect 277938 72559 277955 72581
rect 278041 72559 278062 72581
rect 278062 72559 278097 72581
rect 278183 72559 278186 72581
rect 278186 72559 278239 72581
rect 278325 72559 278378 72581
rect 278378 72559 278381 72581
rect 278467 72559 278502 72581
rect 278502 72559 278523 72581
rect 278609 72559 278626 72581
rect 278626 72559 278665 72581
rect 278751 72559 278806 72581
rect 278806 72559 278807 72581
rect 278893 72559 278930 72581
rect 278930 72559 278949 72581
rect 279035 72559 279054 72581
rect 279054 72559 279091 72581
rect 279177 72559 279178 72581
rect 279178 72559 279233 72581
rect 279319 72559 279370 72581
rect 279370 72559 279375 72581
rect 279461 72559 279494 72581
rect 279494 72559 279517 72581
rect 279603 72559 279618 72581
rect 279618 72559 279659 72581
rect 279745 72559 279798 72581
rect 279798 72559 279801 72581
rect 277899 72457 277955 72473
rect 278041 72457 278097 72473
rect 278183 72457 278239 72473
rect 278325 72457 278381 72473
rect 278467 72457 278523 72473
rect 278609 72457 278665 72473
rect 278751 72457 278807 72473
rect 278893 72457 278949 72473
rect 279035 72457 279091 72473
rect 279177 72457 279233 72473
rect 279319 72457 279375 72473
rect 279461 72457 279517 72473
rect 279603 72457 279659 72473
rect 279745 72457 279801 72473
rect 277899 72417 277938 72457
rect 277938 72417 277955 72457
rect 278041 72417 278062 72457
rect 278062 72417 278097 72457
rect 278183 72417 278186 72457
rect 278186 72417 278239 72457
rect 278325 72417 278378 72457
rect 278378 72417 278381 72457
rect 278467 72417 278502 72457
rect 278502 72417 278523 72457
rect 278609 72417 278626 72457
rect 278626 72417 278665 72457
rect 278751 72417 278806 72457
rect 278806 72417 278807 72457
rect 278893 72417 278930 72457
rect 278930 72417 278949 72457
rect 279035 72417 279054 72457
rect 279054 72417 279091 72457
rect 279177 72417 279178 72457
rect 279178 72417 279233 72457
rect 279319 72417 279370 72457
rect 279370 72417 279375 72457
rect 279461 72417 279494 72457
rect 279494 72417 279517 72457
rect 279603 72417 279618 72457
rect 279618 72417 279659 72457
rect 279745 72417 279798 72457
rect 279798 72417 279801 72457
rect 277899 72277 277938 72331
rect 277938 72277 277955 72331
rect 278041 72277 278062 72331
rect 278062 72277 278097 72331
rect 278183 72277 278186 72331
rect 278186 72277 278239 72331
rect 278325 72277 278378 72331
rect 278378 72277 278381 72331
rect 278467 72277 278502 72331
rect 278502 72277 278523 72331
rect 278609 72277 278626 72331
rect 278626 72277 278665 72331
rect 278751 72277 278806 72331
rect 278806 72277 278807 72331
rect 278893 72277 278930 72331
rect 278930 72277 278949 72331
rect 279035 72277 279054 72331
rect 279054 72277 279091 72331
rect 279177 72277 279178 72331
rect 279178 72277 279233 72331
rect 279319 72277 279370 72331
rect 279370 72277 279375 72331
rect 279461 72277 279494 72331
rect 279494 72277 279517 72331
rect 279603 72277 279618 72331
rect 279618 72277 279659 72331
rect 279745 72277 279798 72331
rect 279798 72277 279801 72331
rect 277899 72275 277955 72277
rect 278041 72275 278097 72277
rect 278183 72275 278239 72277
rect 278325 72275 278381 72277
rect 278467 72275 278523 72277
rect 278609 72275 278665 72277
rect 278751 72275 278807 72277
rect 278893 72275 278949 72277
rect 279035 72275 279091 72277
rect 279177 72275 279233 72277
rect 279319 72275 279375 72277
rect 279461 72275 279517 72277
rect 279603 72275 279659 72277
rect 279745 72275 279801 72277
rect 277899 72153 277938 72189
rect 277938 72153 277955 72189
rect 278041 72153 278062 72189
rect 278062 72153 278097 72189
rect 278183 72153 278186 72189
rect 278186 72153 278239 72189
rect 278325 72153 278378 72189
rect 278378 72153 278381 72189
rect 278467 72153 278502 72189
rect 278502 72153 278523 72189
rect 278609 72153 278626 72189
rect 278626 72153 278665 72189
rect 278751 72153 278806 72189
rect 278806 72153 278807 72189
rect 278893 72153 278930 72189
rect 278930 72153 278949 72189
rect 279035 72153 279054 72189
rect 279054 72153 279091 72189
rect 279177 72153 279178 72189
rect 279178 72153 279233 72189
rect 279319 72153 279370 72189
rect 279370 72153 279375 72189
rect 279461 72153 279494 72189
rect 279494 72153 279517 72189
rect 279603 72153 279618 72189
rect 279618 72153 279659 72189
rect 279745 72153 279798 72189
rect 279798 72153 279801 72189
rect 277899 72133 277955 72153
rect 278041 72133 278097 72153
rect 278183 72133 278239 72153
rect 278325 72133 278381 72153
rect 278467 72133 278523 72153
rect 278609 72133 278665 72153
rect 278751 72133 278807 72153
rect 278893 72133 278949 72153
rect 279035 72133 279091 72153
rect 279177 72133 279233 72153
rect 279319 72133 279375 72153
rect 279461 72133 279517 72153
rect 279603 72133 279659 72153
rect 279745 72133 279801 72153
rect 280269 73979 280325 74035
rect 280411 73979 280467 74035
rect 280553 73979 280609 74035
rect 280695 73979 280751 74035
rect 280837 73979 280893 74035
rect 280979 73979 281035 74035
rect 281121 73979 281177 74035
rect 281263 73979 281319 74035
rect 281405 73979 281461 74035
rect 281547 73979 281603 74035
rect 281689 73979 281745 74035
rect 281831 73979 281887 74035
rect 281973 73979 282029 74035
rect 282115 73979 282171 74035
rect 280269 73889 280308 73893
rect 280308 73889 280325 73893
rect 280411 73889 280432 73893
rect 280432 73889 280467 73893
rect 280553 73889 280556 73893
rect 280556 73889 280609 73893
rect 280695 73889 280748 73893
rect 280748 73889 280751 73893
rect 280837 73889 280872 73893
rect 280872 73889 280893 73893
rect 280979 73889 280996 73893
rect 280996 73889 281035 73893
rect 281121 73889 281176 73893
rect 281176 73889 281177 73893
rect 281263 73889 281300 73893
rect 281300 73889 281319 73893
rect 281405 73889 281424 73893
rect 281424 73889 281461 73893
rect 281547 73889 281548 73893
rect 281548 73889 281603 73893
rect 281689 73889 281740 73893
rect 281740 73889 281745 73893
rect 281831 73889 281864 73893
rect 281864 73889 281887 73893
rect 281973 73889 281988 73893
rect 281988 73889 282029 73893
rect 282115 73889 282168 73893
rect 282168 73889 282171 73893
rect 280269 73837 280325 73889
rect 280411 73837 280467 73889
rect 280553 73837 280609 73889
rect 280695 73837 280751 73889
rect 280837 73837 280893 73889
rect 280979 73837 281035 73889
rect 281121 73837 281177 73889
rect 281263 73837 281319 73889
rect 281405 73837 281461 73889
rect 281547 73837 281603 73889
rect 281689 73837 281745 73889
rect 281831 73837 281887 73889
rect 281973 73837 282029 73889
rect 282115 73837 282171 73889
rect 280269 73697 280325 73751
rect 280411 73697 280467 73751
rect 280553 73697 280609 73751
rect 280695 73697 280751 73751
rect 280837 73697 280893 73751
rect 280979 73697 281035 73751
rect 281121 73697 281177 73751
rect 281263 73697 281319 73751
rect 281405 73697 281461 73751
rect 281547 73697 281603 73751
rect 281689 73697 281745 73751
rect 281831 73697 281887 73751
rect 281973 73697 282029 73751
rect 282115 73697 282171 73751
rect 280269 73695 280308 73697
rect 280308 73695 280325 73697
rect 280411 73695 280432 73697
rect 280432 73695 280467 73697
rect 280553 73695 280556 73697
rect 280556 73695 280609 73697
rect 280695 73695 280748 73697
rect 280748 73695 280751 73697
rect 280837 73695 280872 73697
rect 280872 73695 280893 73697
rect 280979 73695 280996 73697
rect 280996 73695 281035 73697
rect 281121 73695 281176 73697
rect 281176 73695 281177 73697
rect 281263 73695 281300 73697
rect 281300 73695 281319 73697
rect 281405 73695 281424 73697
rect 281424 73695 281461 73697
rect 281547 73695 281548 73697
rect 281548 73695 281603 73697
rect 281689 73695 281740 73697
rect 281740 73695 281745 73697
rect 281831 73695 281864 73697
rect 281864 73695 281887 73697
rect 281973 73695 281988 73697
rect 281988 73695 282029 73697
rect 282115 73695 282168 73697
rect 282168 73695 282171 73697
rect 280269 73573 280325 73609
rect 280411 73573 280467 73609
rect 280553 73573 280609 73609
rect 280695 73573 280751 73609
rect 280837 73573 280893 73609
rect 280979 73573 281035 73609
rect 281121 73573 281177 73609
rect 281263 73573 281319 73609
rect 281405 73573 281461 73609
rect 281547 73573 281603 73609
rect 281689 73573 281745 73609
rect 281831 73573 281887 73609
rect 281973 73573 282029 73609
rect 282115 73573 282171 73609
rect 280269 73553 280308 73573
rect 280308 73553 280325 73573
rect 280411 73553 280432 73573
rect 280432 73553 280467 73573
rect 280553 73553 280556 73573
rect 280556 73553 280609 73573
rect 280695 73553 280748 73573
rect 280748 73553 280751 73573
rect 280837 73553 280872 73573
rect 280872 73553 280893 73573
rect 280979 73553 280996 73573
rect 280996 73553 281035 73573
rect 281121 73553 281176 73573
rect 281176 73553 281177 73573
rect 281263 73553 281300 73573
rect 281300 73553 281319 73573
rect 281405 73553 281424 73573
rect 281424 73553 281461 73573
rect 281547 73553 281548 73573
rect 281548 73553 281603 73573
rect 281689 73553 281740 73573
rect 281740 73553 281745 73573
rect 281831 73553 281864 73573
rect 281864 73553 281887 73573
rect 281973 73553 281988 73573
rect 281988 73553 282029 73573
rect 282115 73553 282168 73573
rect 282168 73553 282171 73573
rect 280269 73449 280325 73467
rect 280411 73449 280467 73467
rect 280553 73449 280609 73467
rect 280695 73449 280751 73467
rect 280837 73449 280893 73467
rect 280979 73449 281035 73467
rect 281121 73449 281177 73467
rect 281263 73449 281319 73467
rect 281405 73449 281461 73467
rect 281547 73449 281603 73467
rect 281689 73449 281745 73467
rect 281831 73449 281887 73467
rect 281973 73449 282029 73467
rect 282115 73449 282171 73467
rect 280269 73411 280308 73449
rect 280308 73411 280325 73449
rect 280411 73411 280432 73449
rect 280432 73411 280467 73449
rect 280553 73411 280556 73449
rect 280556 73411 280609 73449
rect 280695 73411 280748 73449
rect 280748 73411 280751 73449
rect 280837 73411 280872 73449
rect 280872 73411 280893 73449
rect 280979 73411 280996 73449
rect 280996 73411 281035 73449
rect 281121 73411 281176 73449
rect 281176 73411 281177 73449
rect 281263 73411 281300 73449
rect 281300 73411 281319 73449
rect 281405 73411 281424 73449
rect 281424 73411 281461 73449
rect 281547 73411 281548 73449
rect 281548 73411 281603 73449
rect 281689 73411 281740 73449
rect 281740 73411 281745 73449
rect 281831 73411 281864 73449
rect 281864 73411 281887 73449
rect 281973 73411 281988 73449
rect 281988 73411 282029 73449
rect 282115 73411 282168 73449
rect 282168 73411 282171 73449
rect 280269 73269 280308 73325
rect 280308 73269 280325 73325
rect 280411 73269 280432 73325
rect 280432 73269 280467 73325
rect 280553 73269 280556 73325
rect 280556 73269 280609 73325
rect 280695 73269 280748 73325
rect 280748 73269 280751 73325
rect 280837 73269 280872 73325
rect 280872 73269 280893 73325
rect 280979 73269 280996 73325
rect 280996 73269 281035 73325
rect 281121 73269 281176 73325
rect 281176 73269 281177 73325
rect 281263 73269 281300 73325
rect 281300 73269 281319 73325
rect 281405 73269 281424 73325
rect 281424 73269 281461 73325
rect 281547 73269 281548 73325
rect 281548 73269 281603 73325
rect 281689 73269 281740 73325
rect 281740 73269 281745 73325
rect 281831 73269 281864 73325
rect 281864 73269 281887 73325
rect 281973 73269 281988 73325
rect 281988 73269 282029 73325
rect 282115 73269 282168 73325
rect 282168 73269 282171 73325
rect 280269 73145 280308 73183
rect 280308 73145 280325 73183
rect 280411 73145 280432 73183
rect 280432 73145 280467 73183
rect 280553 73145 280556 73183
rect 280556 73145 280609 73183
rect 280695 73145 280748 73183
rect 280748 73145 280751 73183
rect 280837 73145 280872 73183
rect 280872 73145 280893 73183
rect 280979 73145 280996 73183
rect 280996 73145 281035 73183
rect 281121 73145 281176 73183
rect 281176 73145 281177 73183
rect 281263 73145 281300 73183
rect 281300 73145 281319 73183
rect 281405 73145 281424 73183
rect 281424 73145 281461 73183
rect 281547 73145 281548 73183
rect 281548 73145 281603 73183
rect 281689 73145 281740 73183
rect 281740 73145 281745 73183
rect 281831 73145 281864 73183
rect 281864 73145 281887 73183
rect 281973 73145 281988 73183
rect 281988 73145 282029 73183
rect 282115 73145 282168 73183
rect 282168 73145 282171 73183
rect 280269 73127 280325 73145
rect 280411 73127 280467 73145
rect 280553 73127 280609 73145
rect 280695 73127 280751 73145
rect 280837 73127 280893 73145
rect 280979 73127 281035 73145
rect 281121 73127 281177 73145
rect 281263 73127 281319 73145
rect 281405 73127 281461 73145
rect 281547 73127 281603 73145
rect 281689 73127 281745 73145
rect 281831 73127 281887 73145
rect 281973 73127 282029 73145
rect 282115 73127 282171 73145
rect 280269 73021 280308 73041
rect 280308 73021 280325 73041
rect 280411 73021 280432 73041
rect 280432 73021 280467 73041
rect 280553 73021 280556 73041
rect 280556 73021 280609 73041
rect 280695 73021 280748 73041
rect 280748 73021 280751 73041
rect 280837 73021 280872 73041
rect 280872 73021 280893 73041
rect 280979 73021 280996 73041
rect 280996 73021 281035 73041
rect 281121 73021 281176 73041
rect 281176 73021 281177 73041
rect 281263 73021 281300 73041
rect 281300 73021 281319 73041
rect 281405 73021 281424 73041
rect 281424 73021 281461 73041
rect 281547 73021 281548 73041
rect 281548 73021 281603 73041
rect 281689 73021 281740 73041
rect 281740 73021 281745 73041
rect 281831 73021 281864 73041
rect 281864 73021 281887 73041
rect 281973 73021 281988 73041
rect 281988 73021 282029 73041
rect 282115 73021 282168 73041
rect 282168 73021 282171 73041
rect 280269 72985 280325 73021
rect 280411 72985 280467 73021
rect 280553 72985 280609 73021
rect 280695 72985 280751 73021
rect 280837 72985 280893 73021
rect 280979 72985 281035 73021
rect 281121 72985 281177 73021
rect 281263 72985 281319 73021
rect 281405 72985 281461 73021
rect 281547 72985 281603 73021
rect 281689 72985 281745 73021
rect 281831 72985 281887 73021
rect 281973 72985 282029 73021
rect 282115 72985 282171 73021
rect 280269 72897 280308 72899
rect 280308 72897 280325 72899
rect 280411 72897 280432 72899
rect 280432 72897 280467 72899
rect 280553 72897 280556 72899
rect 280556 72897 280609 72899
rect 280695 72897 280748 72899
rect 280748 72897 280751 72899
rect 280837 72897 280872 72899
rect 280872 72897 280893 72899
rect 280979 72897 280996 72899
rect 280996 72897 281035 72899
rect 281121 72897 281176 72899
rect 281176 72897 281177 72899
rect 281263 72897 281300 72899
rect 281300 72897 281319 72899
rect 281405 72897 281424 72899
rect 281424 72897 281461 72899
rect 281547 72897 281548 72899
rect 281548 72897 281603 72899
rect 281689 72897 281740 72899
rect 281740 72897 281745 72899
rect 281831 72897 281864 72899
rect 281864 72897 281887 72899
rect 281973 72897 281988 72899
rect 281988 72897 282029 72899
rect 282115 72897 282168 72899
rect 282168 72897 282171 72899
rect 280269 72843 280325 72897
rect 280411 72843 280467 72897
rect 280553 72843 280609 72897
rect 280695 72843 280751 72897
rect 280837 72843 280893 72897
rect 280979 72843 281035 72897
rect 281121 72843 281177 72897
rect 281263 72843 281319 72897
rect 281405 72843 281461 72897
rect 281547 72843 281603 72897
rect 281689 72843 281745 72897
rect 281831 72843 281887 72897
rect 281973 72843 282029 72897
rect 282115 72843 282171 72897
rect 280269 72705 280325 72757
rect 280411 72705 280467 72757
rect 280553 72705 280609 72757
rect 280695 72705 280751 72757
rect 280837 72705 280893 72757
rect 280979 72705 281035 72757
rect 281121 72705 281177 72757
rect 281263 72705 281319 72757
rect 281405 72705 281461 72757
rect 281547 72705 281603 72757
rect 281689 72705 281745 72757
rect 281831 72705 281887 72757
rect 281973 72705 282029 72757
rect 282115 72705 282171 72757
rect 280269 72701 280308 72705
rect 280308 72701 280325 72705
rect 280411 72701 280432 72705
rect 280432 72701 280467 72705
rect 280553 72701 280556 72705
rect 280556 72701 280609 72705
rect 280695 72701 280748 72705
rect 280748 72701 280751 72705
rect 280837 72701 280872 72705
rect 280872 72701 280893 72705
rect 280979 72701 280996 72705
rect 280996 72701 281035 72705
rect 281121 72701 281176 72705
rect 281176 72701 281177 72705
rect 281263 72701 281300 72705
rect 281300 72701 281319 72705
rect 281405 72701 281424 72705
rect 281424 72701 281461 72705
rect 281547 72701 281548 72705
rect 281548 72701 281603 72705
rect 281689 72701 281740 72705
rect 281740 72701 281745 72705
rect 281831 72701 281864 72705
rect 281864 72701 281887 72705
rect 281973 72701 281988 72705
rect 281988 72701 282029 72705
rect 282115 72701 282168 72705
rect 282168 72701 282171 72705
rect 280269 72581 280325 72615
rect 280411 72581 280467 72615
rect 280553 72581 280609 72615
rect 280695 72581 280751 72615
rect 280837 72581 280893 72615
rect 280979 72581 281035 72615
rect 281121 72581 281177 72615
rect 281263 72581 281319 72615
rect 281405 72581 281461 72615
rect 281547 72581 281603 72615
rect 281689 72581 281745 72615
rect 281831 72581 281887 72615
rect 281973 72581 282029 72615
rect 282115 72581 282171 72615
rect 280269 72559 280308 72581
rect 280308 72559 280325 72581
rect 280411 72559 280432 72581
rect 280432 72559 280467 72581
rect 280553 72559 280556 72581
rect 280556 72559 280609 72581
rect 280695 72559 280748 72581
rect 280748 72559 280751 72581
rect 280837 72559 280872 72581
rect 280872 72559 280893 72581
rect 280979 72559 280996 72581
rect 280996 72559 281035 72581
rect 281121 72559 281176 72581
rect 281176 72559 281177 72581
rect 281263 72559 281300 72581
rect 281300 72559 281319 72581
rect 281405 72559 281424 72581
rect 281424 72559 281461 72581
rect 281547 72559 281548 72581
rect 281548 72559 281603 72581
rect 281689 72559 281740 72581
rect 281740 72559 281745 72581
rect 281831 72559 281864 72581
rect 281864 72559 281887 72581
rect 281973 72559 281988 72581
rect 281988 72559 282029 72581
rect 282115 72559 282168 72581
rect 282168 72559 282171 72581
rect 280269 72457 280325 72473
rect 280411 72457 280467 72473
rect 280553 72457 280609 72473
rect 280695 72457 280751 72473
rect 280837 72457 280893 72473
rect 280979 72457 281035 72473
rect 281121 72457 281177 72473
rect 281263 72457 281319 72473
rect 281405 72457 281461 72473
rect 281547 72457 281603 72473
rect 281689 72457 281745 72473
rect 281831 72457 281887 72473
rect 281973 72457 282029 72473
rect 282115 72457 282171 72473
rect 280269 72417 280308 72457
rect 280308 72417 280325 72457
rect 280411 72417 280432 72457
rect 280432 72417 280467 72457
rect 280553 72417 280556 72457
rect 280556 72417 280609 72457
rect 280695 72417 280748 72457
rect 280748 72417 280751 72457
rect 280837 72417 280872 72457
rect 280872 72417 280893 72457
rect 280979 72417 280996 72457
rect 280996 72417 281035 72457
rect 281121 72417 281176 72457
rect 281176 72417 281177 72457
rect 281263 72417 281300 72457
rect 281300 72417 281319 72457
rect 281405 72417 281424 72457
rect 281424 72417 281461 72457
rect 281547 72417 281548 72457
rect 281548 72417 281603 72457
rect 281689 72417 281740 72457
rect 281740 72417 281745 72457
rect 281831 72417 281864 72457
rect 281864 72417 281887 72457
rect 281973 72417 281988 72457
rect 281988 72417 282029 72457
rect 282115 72417 282168 72457
rect 282168 72417 282171 72457
rect 280269 72277 280308 72331
rect 280308 72277 280325 72331
rect 280411 72277 280432 72331
rect 280432 72277 280467 72331
rect 280553 72277 280556 72331
rect 280556 72277 280609 72331
rect 280695 72277 280748 72331
rect 280748 72277 280751 72331
rect 280837 72277 280872 72331
rect 280872 72277 280893 72331
rect 280979 72277 280996 72331
rect 280996 72277 281035 72331
rect 281121 72277 281176 72331
rect 281176 72277 281177 72331
rect 281263 72277 281300 72331
rect 281300 72277 281319 72331
rect 281405 72277 281424 72331
rect 281424 72277 281461 72331
rect 281547 72277 281548 72331
rect 281548 72277 281603 72331
rect 281689 72277 281740 72331
rect 281740 72277 281745 72331
rect 281831 72277 281864 72331
rect 281864 72277 281887 72331
rect 281973 72277 281988 72331
rect 281988 72277 282029 72331
rect 282115 72277 282168 72331
rect 282168 72277 282171 72331
rect 280269 72275 280325 72277
rect 280411 72275 280467 72277
rect 280553 72275 280609 72277
rect 280695 72275 280751 72277
rect 280837 72275 280893 72277
rect 280979 72275 281035 72277
rect 281121 72275 281177 72277
rect 281263 72275 281319 72277
rect 281405 72275 281461 72277
rect 281547 72275 281603 72277
rect 281689 72275 281745 72277
rect 281831 72275 281887 72277
rect 281973 72275 282029 72277
rect 282115 72275 282171 72277
rect 280269 72153 280308 72189
rect 280308 72153 280325 72189
rect 280411 72153 280432 72189
rect 280432 72153 280467 72189
rect 280553 72153 280556 72189
rect 280556 72153 280609 72189
rect 280695 72153 280748 72189
rect 280748 72153 280751 72189
rect 280837 72153 280872 72189
rect 280872 72153 280893 72189
rect 280979 72153 280996 72189
rect 280996 72153 281035 72189
rect 281121 72153 281176 72189
rect 281176 72153 281177 72189
rect 281263 72153 281300 72189
rect 281300 72153 281319 72189
rect 281405 72153 281424 72189
rect 281424 72153 281461 72189
rect 281547 72153 281548 72189
rect 281548 72153 281603 72189
rect 281689 72153 281740 72189
rect 281740 72153 281745 72189
rect 281831 72153 281864 72189
rect 281864 72153 281887 72189
rect 281973 72153 281988 72189
rect 281988 72153 282029 72189
rect 282115 72153 282168 72189
rect 282168 72153 282171 72189
rect 280269 72133 280325 72153
rect 280411 72133 280467 72153
rect 280553 72133 280609 72153
rect 280695 72133 280751 72153
rect 280837 72133 280893 72153
rect 280979 72133 281035 72153
rect 281121 72133 281177 72153
rect 281263 72133 281319 72153
rect 281405 72133 281461 72153
rect 281547 72133 281603 72153
rect 281689 72133 281745 72153
rect 281831 72133 281887 72153
rect 281973 72133 282029 72153
rect 282115 72133 282171 72153
rect 282899 73979 282955 74035
rect 283041 73979 283097 74035
rect 283183 73979 283239 74035
rect 283325 73979 283381 74035
rect 283467 73979 283523 74035
rect 283609 73979 283665 74035
rect 283751 73979 283807 74035
rect 283893 73979 283949 74035
rect 282899 73889 282938 73893
rect 282938 73889 282955 73893
rect 283041 73889 283062 73893
rect 283062 73889 283097 73893
rect 283183 73889 283186 73893
rect 283186 73889 283239 73893
rect 283325 73889 283378 73893
rect 283378 73889 283381 73893
rect 283467 73889 283502 73893
rect 283502 73889 283523 73893
rect 283609 73889 283626 73893
rect 283626 73889 283665 73893
rect 283751 73889 283806 73893
rect 283806 73889 283807 73893
rect 283893 73889 283930 73893
rect 283930 73889 283949 73893
rect 282899 73837 282955 73889
rect 283041 73837 283097 73889
rect 283183 73837 283239 73889
rect 283325 73837 283381 73889
rect 283467 73837 283523 73889
rect 283609 73837 283665 73889
rect 283751 73837 283807 73889
rect 283893 73837 283949 73889
rect 282899 73697 282955 73751
rect 283041 73697 283097 73751
rect 283183 73697 283239 73751
rect 283325 73697 283381 73751
rect 283467 73697 283523 73751
rect 283609 73697 283665 73751
rect 283751 73697 283807 73751
rect 283893 73697 283949 73751
rect 282899 73695 282938 73697
rect 282938 73695 282955 73697
rect 283041 73695 283062 73697
rect 283062 73695 283097 73697
rect 283183 73695 283186 73697
rect 283186 73695 283239 73697
rect 283325 73695 283378 73697
rect 283378 73695 283381 73697
rect 283467 73695 283502 73697
rect 283502 73695 283523 73697
rect 283609 73695 283626 73697
rect 283626 73695 283665 73697
rect 283751 73695 283806 73697
rect 283806 73695 283807 73697
rect 283893 73695 283930 73697
rect 283930 73695 283949 73697
rect 282899 73573 282955 73609
rect 283041 73573 283097 73609
rect 283183 73573 283239 73609
rect 283325 73573 283381 73609
rect 283467 73573 283523 73609
rect 283609 73573 283665 73609
rect 283751 73573 283807 73609
rect 283893 73573 283949 73609
rect 282899 73553 282938 73573
rect 282938 73553 282955 73573
rect 283041 73553 283062 73573
rect 283062 73553 283097 73573
rect 283183 73553 283186 73573
rect 283186 73553 283239 73573
rect 283325 73553 283378 73573
rect 283378 73553 283381 73573
rect 283467 73553 283502 73573
rect 283502 73553 283523 73573
rect 283609 73553 283626 73573
rect 283626 73553 283665 73573
rect 283751 73553 283806 73573
rect 283806 73553 283807 73573
rect 283893 73553 283930 73573
rect 283930 73553 283949 73573
rect 282899 73449 282955 73467
rect 283041 73449 283097 73467
rect 283183 73449 283239 73467
rect 283325 73449 283381 73467
rect 283467 73449 283523 73467
rect 283609 73449 283665 73467
rect 283751 73449 283807 73467
rect 283893 73449 283949 73467
rect 282899 73411 282938 73449
rect 282938 73411 282955 73449
rect 283041 73411 283062 73449
rect 283062 73411 283097 73449
rect 283183 73411 283186 73449
rect 283186 73411 283239 73449
rect 283325 73411 283378 73449
rect 283378 73411 283381 73449
rect 283467 73411 283502 73449
rect 283502 73411 283523 73449
rect 283609 73411 283626 73449
rect 283626 73411 283665 73449
rect 283751 73411 283806 73449
rect 283806 73411 283807 73449
rect 283893 73411 283930 73449
rect 283930 73411 283949 73449
rect 282899 73269 282938 73325
rect 282938 73269 282955 73325
rect 283041 73269 283062 73325
rect 283062 73269 283097 73325
rect 283183 73269 283186 73325
rect 283186 73269 283239 73325
rect 283325 73269 283378 73325
rect 283378 73269 283381 73325
rect 283467 73269 283502 73325
rect 283502 73269 283523 73325
rect 283609 73269 283626 73325
rect 283626 73269 283665 73325
rect 283751 73269 283806 73325
rect 283806 73269 283807 73325
rect 283893 73269 283930 73325
rect 283930 73269 283949 73325
rect 282899 73145 282938 73183
rect 282938 73145 282955 73183
rect 283041 73145 283062 73183
rect 283062 73145 283097 73183
rect 283183 73145 283186 73183
rect 283186 73145 283239 73183
rect 283325 73145 283378 73183
rect 283378 73145 283381 73183
rect 283467 73145 283502 73183
rect 283502 73145 283523 73183
rect 283609 73145 283626 73183
rect 283626 73145 283665 73183
rect 283751 73145 283806 73183
rect 283806 73145 283807 73183
rect 283893 73145 283930 73183
rect 283930 73145 283949 73183
rect 282899 73127 282955 73145
rect 283041 73127 283097 73145
rect 283183 73127 283239 73145
rect 283325 73127 283381 73145
rect 283467 73127 283523 73145
rect 283609 73127 283665 73145
rect 283751 73127 283807 73145
rect 283893 73127 283949 73145
rect 282899 73021 282938 73041
rect 282938 73021 282955 73041
rect 283041 73021 283062 73041
rect 283062 73021 283097 73041
rect 283183 73021 283186 73041
rect 283186 73021 283239 73041
rect 283325 73021 283378 73041
rect 283378 73021 283381 73041
rect 283467 73021 283502 73041
rect 283502 73021 283523 73041
rect 283609 73021 283626 73041
rect 283626 73021 283665 73041
rect 283751 73021 283806 73041
rect 283806 73021 283807 73041
rect 283893 73021 283930 73041
rect 283930 73021 283949 73041
rect 282899 72985 282955 73021
rect 283041 72985 283097 73021
rect 283183 72985 283239 73021
rect 283325 72985 283381 73021
rect 283467 72985 283523 73021
rect 283609 72985 283665 73021
rect 283751 72985 283807 73021
rect 283893 72985 283949 73021
rect 282899 72897 282938 72899
rect 282938 72897 282955 72899
rect 283041 72897 283062 72899
rect 283062 72897 283097 72899
rect 283183 72897 283186 72899
rect 283186 72897 283239 72899
rect 283325 72897 283378 72899
rect 283378 72897 283381 72899
rect 283467 72897 283502 72899
rect 283502 72897 283523 72899
rect 283609 72897 283626 72899
rect 283626 72897 283665 72899
rect 283751 72897 283806 72899
rect 283806 72897 283807 72899
rect 283893 72897 283930 72899
rect 283930 72897 283949 72899
rect 282899 72843 282955 72897
rect 283041 72843 283097 72897
rect 283183 72843 283239 72897
rect 283325 72843 283381 72897
rect 283467 72843 283523 72897
rect 283609 72843 283665 72897
rect 283751 72843 283807 72897
rect 283893 72843 283949 72897
rect 282899 72705 282955 72757
rect 283041 72705 283097 72757
rect 283183 72705 283239 72757
rect 283325 72705 283381 72757
rect 283467 72705 283523 72757
rect 283609 72705 283665 72757
rect 283751 72705 283807 72757
rect 283893 72705 283949 72757
rect 282899 72701 282938 72705
rect 282938 72701 282955 72705
rect 283041 72701 283062 72705
rect 283062 72701 283097 72705
rect 283183 72701 283186 72705
rect 283186 72701 283239 72705
rect 283325 72701 283378 72705
rect 283378 72701 283381 72705
rect 283467 72701 283502 72705
rect 283502 72701 283523 72705
rect 283609 72701 283626 72705
rect 283626 72701 283665 72705
rect 283751 72701 283806 72705
rect 283806 72701 283807 72705
rect 283893 72701 283930 72705
rect 283930 72701 283949 72705
rect 282899 72581 282955 72615
rect 283041 72581 283097 72615
rect 283183 72581 283239 72615
rect 283325 72581 283381 72615
rect 283467 72581 283523 72615
rect 283609 72581 283665 72615
rect 283751 72581 283807 72615
rect 283893 72581 283949 72615
rect 282899 72559 282938 72581
rect 282938 72559 282955 72581
rect 283041 72559 283062 72581
rect 283062 72559 283097 72581
rect 283183 72559 283186 72581
rect 283186 72559 283239 72581
rect 283325 72559 283378 72581
rect 283378 72559 283381 72581
rect 283467 72559 283502 72581
rect 283502 72559 283523 72581
rect 283609 72559 283626 72581
rect 283626 72559 283665 72581
rect 283751 72559 283806 72581
rect 283806 72559 283807 72581
rect 283893 72559 283930 72581
rect 283930 72559 283949 72581
rect 282899 72457 282955 72473
rect 283041 72457 283097 72473
rect 283183 72457 283239 72473
rect 283325 72457 283381 72473
rect 283467 72457 283523 72473
rect 283609 72457 283665 72473
rect 283751 72457 283807 72473
rect 283893 72457 283949 72473
rect 282899 72417 282938 72457
rect 282938 72417 282955 72457
rect 283041 72417 283062 72457
rect 283062 72417 283097 72457
rect 283183 72417 283186 72457
rect 283186 72417 283239 72457
rect 283325 72417 283378 72457
rect 283378 72417 283381 72457
rect 283467 72417 283502 72457
rect 283502 72417 283523 72457
rect 283609 72417 283626 72457
rect 283626 72417 283665 72457
rect 283751 72417 283806 72457
rect 283806 72417 283807 72457
rect 283893 72417 283930 72457
rect 283930 72417 283949 72457
rect 282899 72277 282938 72331
rect 282938 72277 282955 72331
rect 283041 72277 283062 72331
rect 283062 72277 283097 72331
rect 283183 72277 283186 72331
rect 283186 72277 283239 72331
rect 283325 72277 283378 72331
rect 283378 72277 283381 72331
rect 283467 72277 283502 72331
rect 283502 72277 283523 72331
rect 283609 72277 283626 72331
rect 283626 72277 283665 72331
rect 283751 72277 283806 72331
rect 283806 72277 283807 72331
rect 283893 72277 283930 72331
rect 283930 72277 283949 72331
rect 282899 72275 282955 72277
rect 283041 72275 283097 72277
rect 283183 72275 283239 72277
rect 283325 72275 283381 72277
rect 283467 72275 283523 72277
rect 283609 72275 283665 72277
rect 283751 72275 283807 72277
rect 283893 72275 283949 72277
rect 282899 72153 282938 72189
rect 282938 72153 282955 72189
rect 283041 72153 283062 72189
rect 283062 72153 283097 72189
rect 283183 72153 283186 72189
rect 283186 72153 283239 72189
rect 283325 72153 283378 72189
rect 283378 72153 283381 72189
rect 283467 72153 283502 72189
rect 283502 72153 283523 72189
rect 283609 72153 283626 72189
rect 283626 72153 283665 72189
rect 283751 72153 283806 72189
rect 283806 72153 283807 72189
rect 283893 72153 283930 72189
rect 283930 72153 283949 72189
rect 282899 72133 282955 72153
rect 283041 72133 283097 72153
rect 283183 72133 283239 72153
rect 283325 72133 283381 72153
rect 283467 72133 283523 72153
rect 283609 72133 283665 72153
rect 283751 72133 283807 72153
rect 283893 72133 283949 72153
rect 600343 73979 600399 74035
rect 600485 73979 600541 74035
rect 600627 73979 600683 74035
rect 600769 73979 600825 74035
rect 600911 73979 600967 74035
rect 601053 73979 601109 74035
rect 601195 73979 601251 74035
rect 601337 73979 601393 74035
rect 601479 73979 601535 74035
rect 601621 73979 601677 74035
rect 601763 73979 601819 74035
rect 601905 73979 601961 74035
rect 602047 73979 602103 74035
rect 600343 73889 600382 73893
rect 600382 73889 600399 73893
rect 600485 73889 600506 73893
rect 600506 73889 600541 73893
rect 600627 73889 600630 73893
rect 600630 73889 600683 73893
rect 600769 73889 600822 73893
rect 600822 73889 600825 73893
rect 600911 73889 600946 73893
rect 600946 73889 600967 73893
rect 601053 73889 601070 73893
rect 601070 73889 601109 73893
rect 601195 73889 601250 73893
rect 601250 73889 601251 73893
rect 601337 73889 601374 73893
rect 601374 73889 601393 73893
rect 601479 73889 601498 73893
rect 601498 73889 601535 73893
rect 601621 73889 601622 73893
rect 601622 73889 601677 73893
rect 601763 73889 601814 73893
rect 601814 73889 601819 73893
rect 601905 73889 601938 73893
rect 601938 73889 601961 73893
rect 602047 73889 602062 73893
rect 602062 73889 602103 73893
rect 600343 73837 600399 73889
rect 600485 73837 600541 73889
rect 600627 73837 600683 73889
rect 600769 73837 600825 73889
rect 600911 73837 600967 73889
rect 601053 73837 601109 73889
rect 601195 73837 601251 73889
rect 601337 73837 601393 73889
rect 601479 73837 601535 73889
rect 601621 73837 601677 73889
rect 601763 73837 601819 73889
rect 601905 73837 601961 73889
rect 602047 73837 602103 73889
rect 600343 73697 600399 73751
rect 600485 73697 600541 73751
rect 600627 73697 600683 73751
rect 600769 73697 600825 73751
rect 600911 73697 600967 73751
rect 601053 73697 601109 73751
rect 601195 73697 601251 73751
rect 601337 73697 601393 73751
rect 601479 73697 601535 73751
rect 601621 73697 601677 73751
rect 601763 73697 601819 73751
rect 601905 73697 601961 73751
rect 602047 73697 602103 73751
rect 600343 73695 600382 73697
rect 600382 73695 600399 73697
rect 600485 73695 600506 73697
rect 600506 73695 600541 73697
rect 600627 73695 600630 73697
rect 600630 73695 600683 73697
rect 600769 73695 600822 73697
rect 600822 73695 600825 73697
rect 600911 73695 600946 73697
rect 600946 73695 600967 73697
rect 601053 73695 601070 73697
rect 601070 73695 601109 73697
rect 601195 73695 601250 73697
rect 601250 73695 601251 73697
rect 601337 73695 601374 73697
rect 601374 73695 601393 73697
rect 601479 73695 601498 73697
rect 601498 73695 601535 73697
rect 601621 73695 601622 73697
rect 601622 73695 601677 73697
rect 601763 73695 601814 73697
rect 601814 73695 601819 73697
rect 601905 73695 601938 73697
rect 601938 73695 601961 73697
rect 602047 73695 602062 73697
rect 602062 73695 602103 73697
rect 600343 73573 600399 73609
rect 600485 73573 600541 73609
rect 600627 73573 600683 73609
rect 600769 73573 600825 73609
rect 600911 73573 600967 73609
rect 601053 73573 601109 73609
rect 601195 73573 601251 73609
rect 601337 73573 601393 73609
rect 601479 73573 601535 73609
rect 601621 73573 601677 73609
rect 601763 73573 601819 73609
rect 601905 73573 601961 73609
rect 602047 73573 602103 73609
rect 600343 73553 600382 73573
rect 600382 73553 600399 73573
rect 600485 73553 600506 73573
rect 600506 73553 600541 73573
rect 600627 73553 600630 73573
rect 600630 73553 600683 73573
rect 600769 73553 600822 73573
rect 600822 73553 600825 73573
rect 600911 73553 600946 73573
rect 600946 73553 600967 73573
rect 601053 73553 601070 73573
rect 601070 73553 601109 73573
rect 601195 73553 601250 73573
rect 601250 73553 601251 73573
rect 601337 73553 601374 73573
rect 601374 73553 601393 73573
rect 601479 73553 601498 73573
rect 601498 73553 601535 73573
rect 601621 73553 601622 73573
rect 601622 73553 601677 73573
rect 601763 73553 601814 73573
rect 601814 73553 601819 73573
rect 601905 73553 601938 73573
rect 601938 73553 601961 73573
rect 602047 73553 602062 73573
rect 602062 73553 602103 73573
rect 600343 73449 600399 73467
rect 600485 73449 600541 73467
rect 600627 73449 600683 73467
rect 600769 73449 600825 73467
rect 600911 73449 600967 73467
rect 601053 73449 601109 73467
rect 601195 73449 601251 73467
rect 601337 73449 601393 73467
rect 601479 73449 601535 73467
rect 601621 73449 601677 73467
rect 601763 73449 601819 73467
rect 601905 73449 601961 73467
rect 602047 73449 602103 73467
rect 600343 73411 600382 73449
rect 600382 73411 600399 73449
rect 600485 73411 600506 73449
rect 600506 73411 600541 73449
rect 600627 73411 600630 73449
rect 600630 73411 600683 73449
rect 600769 73411 600822 73449
rect 600822 73411 600825 73449
rect 600911 73411 600946 73449
rect 600946 73411 600967 73449
rect 601053 73411 601070 73449
rect 601070 73411 601109 73449
rect 601195 73411 601250 73449
rect 601250 73411 601251 73449
rect 601337 73411 601374 73449
rect 601374 73411 601393 73449
rect 601479 73411 601498 73449
rect 601498 73411 601535 73449
rect 601621 73411 601622 73449
rect 601622 73411 601677 73449
rect 601763 73411 601814 73449
rect 601814 73411 601819 73449
rect 601905 73411 601938 73449
rect 601938 73411 601961 73449
rect 602047 73411 602062 73449
rect 602062 73411 602103 73449
rect 600343 73269 600382 73325
rect 600382 73269 600399 73325
rect 600485 73269 600506 73325
rect 600506 73269 600541 73325
rect 600627 73269 600630 73325
rect 600630 73269 600683 73325
rect 600769 73269 600822 73325
rect 600822 73269 600825 73325
rect 600911 73269 600946 73325
rect 600946 73269 600967 73325
rect 601053 73269 601070 73325
rect 601070 73269 601109 73325
rect 601195 73269 601250 73325
rect 601250 73269 601251 73325
rect 601337 73269 601374 73325
rect 601374 73269 601393 73325
rect 601479 73269 601498 73325
rect 601498 73269 601535 73325
rect 601621 73269 601622 73325
rect 601622 73269 601677 73325
rect 601763 73269 601814 73325
rect 601814 73269 601819 73325
rect 601905 73269 601938 73325
rect 601938 73269 601961 73325
rect 602047 73269 602062 73325
rect 602062 73269 602103 73325
rect 600343 73145 600382 73183
rect 600382 73145 600399 73183
rect 600485 73145 600506 73183
rect 600506 73145 600541 73183
rect 600627 73145 600630 73183
rect 600630 73145 600683 73183
rect 600769 73145 600822 73183
rect 600822 73145 600825 73183
rect 600911 73145 600946 73183
rect 600946 73145 600967 73183
rect 601053 73145 601070 73183
rect 601070 73145 601109 73183
rect 601195 73145 601250 73183
rect 601250 73145 601251 73183
rect 601337 73145 601374 73183
rect 601374 73145 601393 73183
rect 601479 73145 601498 73183
rect 601498 73145 601535 73183
rect 601621 73145 601622 73183
rect 601622 73145 601677 73183
rect 601763 73145 601814 73183
rect 601814 73145 601819 73183
rect 601905 73145 601938 73183
rect 601938 73145 601961 73183
rect 602047 73145 602062 73183
rect 602062 73145 602103 73183
rect 600343 73127 600399 73145
rect 600485 73127 600541 73145
rect 600627 73127 600683 73145
rect 600769 73127 600825 73145
rect 600911 73127 600967 73145
rect 601053 73127 601109 73145
rect 601195 73127 601251 73145
rect 601337 73127 601393 73145
rect 601479 73127 601535 73145
rect 601621 73127 601677 73145
rect 601763 73127 601819 73145
rect 601905 73127 601961 73145
rect 602047 73127 602103 73145
rect 600343 73021 600382 73041
rect 600382 73021 600399 73041
rect 600485 73021 600506 73041
rect 600506 73021 600541 73041
rect 600627 73021 600630 73041
rect 600630 73021 600683 73041
rect 600769 73021 600822 73041
rect 600822 73021 600825 73041
rect 600911 73021 600946 73041
rect 600946 73021 600967 73041
rect 601053 73021 601070 73041
rect 601070 73021 601109 73041
rect 601195 73021 601250 73041
rect 601250 73021 601251 73041
rect 601337 73021 601374 73041
rect 601374 73021 601393 73041
rect 601479 73021 601498 73041
rect 601498 73021 601535 73041
rect 601621 73021 601622 73041
rect 601622 73021 601677 73041
rect 601763 73021 601814 73041
rect 601814 73021 601819 73041
rect 601905 73021 601938 73041
rect 601938 73021 601961 73041
rect 602047 73021 602062 73041
rect 602062 73021 602103 73041
rect 600343 72985 600399 73021
rect 600485 72985 600541 73021
rect 600627 72985 600683 73021
rect 600769 72985 600825 73021
rect 600911 72985 600967 73021
rect 601053 72985 601109 73021
rect 601195 72985 601251 73021
rect 601337 72985 601393 73021
rect 601479 72985 601535 73021
rect 601621 72985 601677 73021
rect 601763 72985 601819 73021
rect 601905 72985 601961 73021
rect 602047 72985 602103 73021
rect 600343 72897 600382 72899
rect 600382 72897 600399 72899
rect 600485 72897 600506 72899
rect 600506 72897 600541 72899
rect 600627 72897 600630 72899
rect 600630 72897 600683 72899
rect 600769 72897 600822 72899
rect 600822 72897 600825 72899
rect 600911 72897 600946 72899
rect 600946 72897 600967 72899
rect 601053 72897 601070 72899
rect 601070 72897 601109 72899
rect 601195 72897 601250 72899
rect 601250 72897 601251 72899
rect 601337 72897 601374 72899
rect 601374 72897 601393 72899
rect 601479 72897 601498 72899
rect 601498 72897 601535 72899
rect 601621 72897 601622 72899
rect 601622 72897 601677 72899
rect 601763 72897 601814 72899
rect 601814 72897 601819 72899
rect 601905 72897 601938 72899
rect 601938 72897 601961 72899
rect 602047 72897 602062 72899
rect 602062 72897 602103 72899
rect 600343 72843 600399 72897
rect 600485 72843 600541 72897
rect 600627 72843 600683 72897
rect 600769 72843 600825 72897
rect 600911 72843 600967 72897
rect 601053 72843 601109 72897
rect 601195 72843 601251 72897
rect 601337 72843 601393 72897
rect 601479 72843 601535 72897
rect 601621 72843 601677 72897
rect 601763 72843 601819 72897
rect 601905 72843 601961 72897
rect 602047 72843 602103 72897
rect 600343 72705 600399 72757
rect 600485 72705 600541 72757
rect 600627 72705 600683 72757
rect 600769 72705 600825 72757
rect 600911 72705 600967 72757
rect 601053 72705 601109 72757
rect 601195 72705 601251 72757
rect 601337 72705 601393 72757
rect 601479 72705 601535 72757
rect 601621 72705 601677 72757
rect 601763 72705 601819 72757
rect 601905 72705 601961 72757
rect 602047 72705 602103 72757
rect 600343 72701 600382 72705
rect 600382 72701 600399 72705
rect 600485 72701 600506 72705
rect 600506 72701 600541 72705
rect 600627 72701 600630 72705
rect 600630 72701 600683 72705
rect 600769 72701 600822 72705
rect 600822 72701 600825 72705
rect 600911 72701 600946 72705
rect 600946 72701 600967 72705
rect 601053 72701 601070 72705
rect 601070 72701 601109 72705
rect 601195 72701 601250 72705
rect 601250 72701 601251 72705
rect 601337 72701 601374 72705
rect 601374 72701 601393 72705
rect 601479 72701 601498 72705
rect 601498 72701 601535 72705
rect 601621 72701 601622 72705
rect 601622 72701 601677 72705
rect 601763 72701 601814 72705
rect 601814 72701 601819 72705
rect 601905 72701 601938 72705
rect 601938 72701 601961 72705
rect 602047 72701 602062 72705
rect 602062 72701 602103 72705
rect 600343 72581 600399 72615
rect 600485 72581 600541 72615
rect 600627 72581 600683 72615
rect 600769 72581 600825 72615
rect 600911 72581 600967 72615
rect 601053 72581 601109 72615
rect 601195 72581 601251 72615
rect 601337 72581 601393 72615
rect 601479 72581 601535 72615
rect 601621 72581 601677 72615
rect 601763 72581 601819 72615
rect 601905 72581 601961 72615
rect 602047 72581 602103 72615
rect 600343 72559 600382 72581
rect 600382 72559 600399 72581
rect 600485 72559 600506 72581
rect 600506 72559 600541 72581
rect 600627 72559 600630 72581
rect 600630 72559 600683 72581
rect 600769 72559 600822 72581
rect 600822 72559 600825 72581
rect 600911 72559 600946 72581
rect 600946 72559 600967 72581
rect 601053 72559 601070 72581
rect 601070 72559 601109 72581
rect 601195 72559 601250 72581
rect 601250 72559 601251 72581
rect 601337 72559 601374 72581
rect 601374 72559 601393 72581
rect 601479 72559 601498 72581
rect 601498 72559 601535 72581
rect 601621 72559 601622 72581
rect 601622 72559 601677 72581
rect 601763 72559 601814 72581
rect 601814 72559 601819 72581
rect 601905 72559 601938 72581
rect 601938 72559 601961 72581
rect 602047 72559 602062 72581
rect 602062 72559 602103 72581
rect 600343 72457 600399 72473
rect 600485 72457 600541 72473
rect 600627 72457 600683 72473
rect 600769 72457 600825 72473
rect 600911 72457 600967 72473
rect 601053 72457 601109 72473
rect 601195 72457 601251 72473
rect 601337 72457 601393 72473
rect 601479 72457 601535 72473
rect 601621 72457 601677 72473
rect 601763 72457 601819 72473
rect 601905 72457 601961 72473
rect 602047 72457 602103 72473
rect 600343 72417 600382 72457
rect 600382 72417 600399 72457
rect 600485 72417 600506 72457
rect 600506 72417 600541 72457
rect 600627 72417 600630 72457
rect 600630 72417 600683 72457
rect 600769 72417 600822 72457
rect 600822 72417 600825 72457
rect 600911 72417 600946 72457
rect 600946 72417 600967 72457
rect 601053 72417 601070 72457
rect 601070 72417 601109 72457
rect 601195 72417 601250 72457
rect 601250 72417 601251 72457
rect 601337 72417 601374 72457
rect 601374 72417 601393 72457
rect 601479 72417 601498 72457
rect 601498 72417 601535 72457
rect 601621 72417 601622 72457
rect 601622 72417 601677 72457
rect 601763 72417 601814 72457
rect 601814 72417 601819 72457
rect 601905 72417 601938 72457
rect 601938 72417 601961 72457
rect 602047 72417 602062 72457
rect 602062 72417 602103 72457
rect 600343 72277 600382 72331
rect 600382 72277 600399 72331
rect 600485 72277 600506 72331
rect 600506 72277 600541 72331
rect 600627 72277 600630 72331
rect 600630 72277 600683 72331
rect 600769 72277 600822 72331
rect 600822 72277 600825 72331
rect 600911 72277 600946 72331
rect 600946 72277 600967 72331
rect 601053 72277 601070 72331
rect 601070 72277 601109 72331
rect 601195 72277 601250 72331
rect 601250 72277 601251 72331
rect 601337 72277 601374 72331
rect 601374 72277 601393 72331
rect 601479 72277 601498 72331
rect 601498 72277 601535 72331
rect 601621 72277 601622 72331
rect 601622 72277 601677 72331
rect 601763 72277 601814 72331
rect 601814 72277 601819 72331
rect 601905 72277 601938 72331
rect 601938 72277 601961 72331
rect 602047 72277 602062 72331
rect 602062 72277 602103 72331
rect 600343 72275 600399 72277
rect 600485 72275 600541 72277
rect 600627 72275 600683 72277
rect 600769 72275 600825 72277
rect 600911 72275 600967 72277
rect 601053 72275 601109 72277
rect 601195 72275 601251 72277
rect 601337 72275 601393 72277
rect 601479 72275 601535 72277
rect 601621 72275 601677 72277
rect 601763 72275 601819 72277
rect 601905 72275 601961 72277
rect 602047 72275 602103 72277
rect 600343 72153 600382 72189
rect 600382 72153 600399 72189
rect 600485 72153 600506 72189
rect 600506 72153 600541 72189
rect 600627 72153 600630 72189
rect 600630 72153 600683 72189
rect 600769 72153 600822 72189
rect 600822 72153 600825 72189
rect 600911 72153 600946 72189
rect 600946 72153 600967 72189
rect 601053 72153 601070 72189
rect 601070 72153 601109 72189
rect 601195 72153 601250 72189
rect 601250 72153 601251 72189
rect 601337 72153 601374 72189
rect 601374 72153 601393 72189
rect 601479 72153 601498 72189
rect 601498 72153 601535 72189
rect 601621 72153 601622 72189
rect 601622 72153 601677 72189
rect 601763 72153 601814 72189
rect 601814 72153 601819 72189
rect 601905 72153 601938 72189
rect 601938 72153 601961 72189
rect 602047 72153 602062 72189
rect 602062 72153 602103 72189
rect 600343 72133 600399 72153
rect 600485 72133 600541 72153
rect 600627 72133 600683 72153
rect 600769 72133 600825 72153
rect 600911 72133 600967 72153
rect 601053 72133 601109 72153
rect 601195 72133 601251 72153
rect 601337 72133 601393 72153
rect 601479 72133 601535 72153
rect 601621 72133 601677 72153
rect 601763 72133 601819 72153
rect 601905 72133 601961 72153
rect 602047 72133 602103 72153
rect 602823 73979 602879 74035
rect 602965 73979 603021 74035
rect 603107 73979 603163 74035
rect 603249 73979 603305 74035
rect 603391 73979 603447 74035
rect 603533 73979 603589 74035
rect 603675 73979 603731 74035
rect 603817 73979 603873 74035
rect 603959 73979 604015 74035
rect 602823 73889 602862 73893
rect 602862 73889 602879 73893
rect 602965 73889 602986 73893
rect 602986 73889 603021 73893
rect 603107 73889 603110 73893
rect 603110 73889 603163 73893
rect 603249 73889 603302 73893
rect 603302 73889 603305 73893
rect 603391 73889 603426 73893
rect 603426 73889 603447 73893
rect 603533 73889 603550 73893
rect 603550 73889 603589 73893
rect 603675 73889 603730 73893
rect 603730 73889 603731 73893
rect 603817 73889 603854 73893
rect 603854 73889 603873 73893
rect 603959 73889 603978 73893
rect 603978 73889 604015 73893
rect 602823 73837 602879 73889
rect 602965 73837 603021 73889
rect 603107 73837 603163 73889
rect 603249 73837 603305 73889
rect 603391 73837 603447 73889
rect 603533 73837 603589 73889
rect 603675 73837 603731 73889
rect 603817 73837 603873 73889
rect 603959 73837 604015 73889
rect 602823 73697 602879 73751
rect 602965 73697 603021 73751
rect 603107 73697 603163 73751
rect 603249 73697 603305 73751
rect 603391 73697 603447 73751
rect 603533 73697 603589 73751
rect 603675 73697 603731 73751
rect 603817 73697 603873 73751
rect 603959 73697 604015 73751
rect 602823 73695 602862 73697
rect 602862 73695 602879 73697
rect 602965 73695 602986 73697
rect 602986 73695 603021 73697
rect 603107 73695 603110 73697
rect 603110 73695 603163 73697
rect 603249 73695 603302 73697
rect 603302 73695 603305 73697
rect 603391 73695 603426 73697
rect 603426 73695 603447 73697
rect 603533 73695 603550 73697
rect 603550 73695 603589 73697
rect 603675 73695 603730 73697
rect 603730 73695 603731 73697
rect 603817 73695 603854 73697
rect 603854 73695 603873 73697
rect 603959 73695 603978 73697
rect 603978 73695 604015 73697
rect 602823 73573 602879 73609
rect 602965 73573 603021 73609
rect 603107 73573 603163 73609
rect 603249 73573 603305 73609
rect 603391 73573 603447 73609
rect 603533 73573 603589 73609
rect 603675 73573 603731 73609
rect 603817 73573 603873 73609
rect 603959 73573 604015 73609
rect 602823 73553 602862 73573
rect 602862 73553 602879 73573
rect 602965 73553 602986 73573
rect 602986 73553 603021 73573
rect 603107 73553 603110 73573
rect 603110 73553 603163 73573
rect 603249 73553 603302 73573
rect 603302 73553 603305 73573
rect 603391 73553 603426 73573
rect 603426 73553 603447 73573
rect 603533 73553 603550 73573
rect 603550 73553 603589 73573
rect 603675 73553 603730 73573
rect 603730 73553 603731 73573
rect 603817 73553 603854 73573
rect 603854 73553 603873 73573
rect 603959 73553 603978 73573
rect 603978 73553 604015 73573
rect 602823 73449 602879 73467
rect 602965 73449 603021 73467
rect 603107 73449 603163 73467
rect 603249 73449 603305 73467
rect 603391 73449 603447 73467
rect 603533 73449 603589 73467
rect 603675 73449 603731 73467
rect 603817 73449 603873 73467
rect 603959 73449 604015 73467
rect 602823 73411 602862 73449
rect 602862 73411 602879 73449
rect 602965 73411 602986 73449
rect 602986 73411 603021 73449
rect 603107 73411 603110 73449
rect 603110 73411 603163 73449
rect 603249 73411 603302 73449
rect 603302 73411 603305 73449
rect 603391 73411 603426 73449
rect 603426 73411 603447 73449
rect 603533 73411 603550 73449
rect 603550 73411 603589 73449
rect 603675 73411 603730 73449
rect 603730 73411 603731 73449
rect 603817 73411 603854 73449
rect 603854 73411 603873 73449
rect 603959 73411 603978 73449
rect 603978 73411 604015 73449
rect 602823 73269 602862 73325
rect 602862 73269 602879 73325
rect 602965 73269 602986 73325
rect 602986 73269 603021 73325
rect 603107 73269 603110 73325
rect 603110 73269 603163 73325
rect 603249 73269 603302 73325
rect 603302 73269 603305 73325
rect 603391 73269 603426 73325
rect 603426 73269 603447 73325
rect 603533 73269 603550 73325
rect 603550 73269 603589 73325
rect 603675 73269 603730 73325
rect 603730 73269 603731 73325
rect 603817 73269 603854 73325
rect 603854 73269 603873 73325
rect 603959 73269 603978 73325
rect 603978 73269 604015 73325
rect 602823 73145 602862 73183
rect 602862 73145 602879 73183
rect 602965 73145 602986 73183
rect 602986 73145 603021 73183
rect 603107 73145 603110 73183
rect 603110 73145 603163 73183
rect 603249 73145 603302 73183
rect 603302 73145 603305 73183
rect 603391 73145 603426 73183
rect 603426 73145 603447 73183
rect 603533 73145 603550 73183
rect 603550 73145 603589 73183
rect 603675 73145 603730 73183
rect 603730 73145 603731 73183
rect 603817 73145 603854 73183
rect 603854 73145 603873 73183
rect 603959 73145 603978 73183
rect 603978 73145 604015 73183
rect 602823 73127 602879 73145
rect 602965 73127 603021 73145
rect 603107 73127 603163 73145
rect 603249 73127 603305 73145
rect 603391 73127 603447 73145
rect 603533 73127 603589 73145
rect 603675 73127 603731 73145
rect 603817 73127 603873 73145
rect 603959 73127 604015 73145
rect 602823 73021 602862 73041
rect 602862 73021 602879 73041
rect 602965 73021 602986 73041
rect 602986 73021 603021 73041
rect 603107 73021 603110 73041
rect 603110 73021 603163 73041
rect 603249 73021 603302 73041
rect 603302 73021 603305 73041
rect 603391 73021 603426 73041
rect 603426 73021 603447 73041
rect 603533 73021 603550 73041
rect 603550 73021 603589 73041
rect 603675 73021 603730 73041
rect 603730 73021 603731 73041
rect 603817 73021 603854 73041
rect 603854 73021 603873 73041
rect 603959 73021 603978 73041
rect 603978 73021 604015 73041
rect 602823 72985 602879 73021
rect 602965 72985 603021 73021
rect 603107 72985 603163 73021
rect 603249 72985 603305 73021
rect 603391 72985 603447 73021
rect 603533 72985 603589 73021
rect 603675 72985 603731 73021
rect 603817 72985 603873 73021
rect 603959 72985 604015 73021
rect 602823 72897 602862 72899
rect 602862 72897 602879 72899
rect 602965 72897 602986 72899
rect 602986 72897 603021 72899
rect 603107 72897 603110 72899
rect 603110 72897 603163 72899
rect 603249 72897 603302 72899
rect 603302 72897 603305 72899
rect 603391 72897 603426 72899
rect 603426 72897 603447 72899
rect 603533 72897 603550 72899
rect 603550 72897 603589 72899
rect 603675 72897 603730 72899
rect 603730 72897 603731 72899
rect 603817 72897 603854 72899
rect 603854 72897 603873 72899
rect 603959 72897 603978 72899
rect 603978 72897 604015 72899
rect 602823 72843 602879 72897
rect 602965 72843 603021 72897
rect 603107 72843 603163 72897
rect 603249 72843 603305 72897
rect 603391 72843 603447 72897
rect 603533 72843 603589 72897
rect 603675 72843 603731 72897
rect 603817 72843 603873 72897
rect 603959 72843 604015 72897
rect 602823 72705 602879 72757
rect 602965 72705 603021 72757
rect 603107 72705 603163 72757
rect 603249 72705 603305 72757
rect 603391 72705 603447 72757
rect 603533 72705 603589 72757
rect 603675 72705 603731 72757
rect 603817 72705 603873 72757
rect 603959 72705 604015 72757
rect 602823 72701 602862 72705
rect 602862 72701 602879 72705
rect 602965 72701 602986 72705
rect 602986 72701 603021 72705
rect 603107 72701 603110 72705
rect 603110 72701 603163 72705
rect 603249 72701 603302 72705
rect 603302 72701 603305 72705
rect 603391 72701 603426 72705
rect 603426 72701 603447 72705
rect 603533 72701 603550 72705
rect 603550 72701 603589 72705
rect 603675 72701 603730 72705
rect 603730 72701 603731 72705
rect 603817 72701 603854 72705
rect 603854 72701 603873 72705
rect 603959 72701 603978 72705
rect 603978 72701 604015 72705
rect 602823 72581 602879 72615
rect 602965 72581 603021 72615
rect 603107 72581 603163 72615
rect 603249 72581 603305 72615
rect 603391 72581 603447 72615
rect 603533 72581 603589 72615
rect 603675 72581 603731 72615
rect 603817 72581 603873 72615
rect 603959 72581 604015 72615
rect 602823 72559 602862 72581
rect 602862 72559 602879 72581
rect 602965 72559 602986 72581
rect 602986 72559 603021 72581
rect 603107 72559 603110 72581
rect 603110 72559 603163 72581
rect 603249 72559 603302 72581
rect 603302 72559 603305 72581
rect 603391 72559 603426 72581
rect 603426 72559 603447 72581
rect 603533 72559 603550 72581
rect 603550 72559 603589 72581
rect 603675 72559 603730 72581
rect 603730 72559 603731 72581
rect 603817 72559 603854 72581
rect 603854 72559 603873 72581
rect 603959 72559 603978 72581
rect 603978 72559 604015 72581
rect 602823 72457 602879 72473
rect 602965 72457 603021 72473
rect 603107 72457 603163 72473
rect 603249 72457 603305 72473
rect 603391 72457 603447 72473
rect 603533 72457 603589 72473
rect 603675 72457 603731 72473
rect 603817 72457 603873 72473
rect 603959 72457 604015 72473
rect 602823 72417 602862 72457
rect 602862 72417 602879 72457
rect 602965 72417 602986 72457
rect 602986 72417 603021 72457
rect 603107 72417 603110 72457
rect 603110 72417 603163 72457
rect 603249 72417 603302 72457
rect 603302 72417 603305 72457
rect 603391 72417 603426 72457
rect 603426 72417 603447 72457
rect 603533 72417 603550 72457
rect 603550 72417 603589 72457
rect 603675 72417 603730 72457
rect 603730 72417 603731 72457
rect 603817 72417 603854 72457
rect 603854 72417 603873 72457
rect 603959 72417 603978 72457
rect 603978 72417 604015 72457
rect 602823 72277 602862 72331
rect 602862 72277 602879 72331
rect 602965 72277 602986 72331
rect 602986 72277 603021 72331
rect 603107 72277 603110 72331
rect 603110 72277 603163 72331
rect 603249 72277 603302 72331
rect 603302 72277 603305 72331
rect 603391 72277 603426 72331
rect 603426 72277 603447 72331
rect 603533 72277 603550 72331
rect 603550 72277 603589 72331
rect 603675 72277 603730 72331
rect 603730 72277 603731 72331
rect 603817 72277 603854 72331
rect 603854 72277 603873 72331
rect 603959 72277 603978 72331
rect 603978 72277 604015 72331
rect 602823 72275 602879 72277
rect 602965 72275 603021 72277
rect 603107 72275 603163 72277
rect 603249 72275 603305 72277
rect 603391 72275 603447 72277
rect 603533 72275 603589 72277
rect 603675 72275 603731 72277
rect 603817 72275 603873 72277
rect 603959 72275 604015 72277
rect 602823 72153 602862 72189
rect 602862 72153 602879 72189
rect 602965 72153 602986 72189
rect 602986 72153 603021 72189
rect 603107 72153 603110 72189
rect 603110 72153 603163 72189
rect 603249 72153 603302 72189
rect 603302 72153 603305 72189
rect 603391 72153 603426 72189
rect 603426 72153 603447 72189
rect 603533 72153 603550 72189
rect 603550 72153 603589 72189
rect 603675 72153 603730 72189
rect 603730 72153 603731 72189
rect 603817 72153 603854 72189
rect 603854 72153 603873 72189
rect 603959 72153 603978 72189
rect 603978 72153 604015 72189
rect 602823 72133 602879 72153
rect 602965 72133 603021 72153
rect 603107 72133 603163 72153
rect 603249 72133 603305 72153
rect 603391 72133 603447 72153
rect 603533 72133 603589 72153
rect 603675 72133 603731 72153
rect 603817 72133 603873 72153
rect 603959 72133 604015 72153
rect 605193 73979 605249 74035
rect 605335 73979 605391 74035
rect 605477 73979 605533 74035
rect 605619 73979 605675 74035
rect 605761 73979 605817 74035
rect 605903 73979 605959 74035
rect 606045 73979 606101 74035
rect 606187 73979 606243 74035
rect 606329 73979 606385 74035
rect 606471 73979 606527 74035
rect 606613 73979 606669 74035
rect 606755 73979 606811 74035
rect 606897 73979 606953 74035
rect 607039 73979 607095 74035
rect 605193 73889 605232 73893
rect 605232 73889 605249 73893
rect 605335 73889 605356 73893
rect 605356 73889 605391 73893
rect 605477 73889 605480 73893
rect 605480 73889 605533 73893
rect 605619 73889 605672 73893
rect 605672 73889 605675 73893
rect 605761 73889 605796 73893
rect 605796 73889 605817 73893
rect 605903 73889 605920 73893
rect 605920 73889 605959 73893
rect 606045 73889 606100 73893
rect 606100 73889 606101 73893
rect 606187 73889 606224 73893
rect 606224 73889 606243 73893
rect 606329 73889 606348 73893
rect 606348 73889 606385 73893
rect 606471 73889 606472 73893
rect 606472 73889 606527 73893
rect 606613 73889 606664 73893
rect 606664 73889 606669 73893
rect 606755 73889 606788 73893
rect 606788 73889 606811 73893
rect 606897 73889 606912 73893
rect 606912 73889 606953 73893
rect 607039 73889 607092 73893
rect 607092 73889 607095 73893
rect 605193 73837 605249 73889
rect 605335 73837 605391 73889
rect 605477 73837 605533 73889
rect 605619 73837 605675 73889
rect 605761 73837 605817 73889
rect 605903 73837 605959 73889
rect 606045 73837 606101 73889
rect 606187 73837 606243 73889
rect 606329 73837 606385 73889
rect 606471 73837 606527 73889
rect 606613 73837 606669 73889
rect 606755 73837 606811 73889
rect 606897 73837 606953 73889
rect 607039 73837 607095 73889
rect 605193 73697 605249 73751
rect 605335 73697 605391 73751
rect 605477 73697 605533 73751
rect 605619 73697 605675 73751
rect 605761 73697 605817 73751
rect 605903 73697 605959 73751
rect 606045 73697 606101 73751
rect 606187 73697 606243 73751
rect 606329 73697 606385 73751
rect 606471 73697 606527 73751
rect 606613 73697 606669 73751
rect 606755 73697 606811 73751
rect 606897 73697 606953 73751
rect 607039 73697 607095 73751
rect 605193 73695 605232 73697
rect 605232 73695 605249 73697
rect 605335 73695 605356 73697
rect 605356 73695 605391 73697
rect 605477 73695 605480 73697
rect 605480 73695 605533 73697
rect 605619 73695 605672 73697
rect 605672 73695 605675 73697
rect 605761 73695 605796 73697
rect 605796 73695 605817 73697
rect 605903 73695 605920 73697
rect 605920 73695 605959 73697
rect 606045 73695 606100 73697
rect 606100 73695 606101 73697
rect 606187 73695 606224 73697
rect 606224 73695 606243 73697
rect 606329 73695 606348 73697
rect 606348 73695 606385 73697
rect 606471 73695 606472 73697
rect 606472 73695 606527 73697
rect 606613 73695 606664 73697
rect 606664 73695 606669 73697
rect 606755 73695 606788 73697
rect 606788 73695 606811 73697
rect 606897 73695 606912 73697
rect 606912 73695 606953 73697
rect 607039 73695 607092 73697
rect 607092 73695 607095 73697
rect 605193 73573 605249 73609
rect 605335 73573 605391 73609
rect 605477 73573 605533 73609
rect 605619 73573 605675 73609
rect 605761 73573 605817 73609
rect 605903 73573 605959 73609
rect 606045 73573 606101 73609
rect 606187 73573 606243 73609
rect 606329 73573 606385 73609
rect 606471 73573 606527 73609
rect 606613 73573 606669 73609
rect 606755 73573 606811 73609
rect 606897 73573 606953 73609
rect 607039 73573 607095 73609
rect 605193 73553 605232 73573
rect 605232 73553 605249 73573
rect 605335 73553 605356 73573
rect 605356 73553 605391 73573
rect 605477 73553 605480 73573
rect 605480 73553 605533 73573
rect 605619 73553 605672 73573
rect 605672 73553 605675 73573
rect 605761 73553 605796 73573
rect 605796 73553 605817 73573
rect 605903 73553 605920 73573
rect 605920 73553 605959 73573
rect 606045 73553 606100 73573
rect 606100 73553 606101 73573
rect 606187 73553 606224 73573
rect 606224 73553 606243 73573
rect 606329 73553 606348 73573
rect 606348 73553 606385 73573
rect 606471 73553 606472 73573
rect 606472 73553 606527 73573
rect 606613 73553 606664 73573
rect 606664 73553 606669 73573
rect 606755 73553 606788 73573
rect 606788 73553 606811 73573
rect 606897 73553 606912 73573
rect 606912 73553 606953 73573
rect 607039 73553 607092 73573
rect 607092 73553 607095 73573
rect 605193 73449 605249 73467
rect 605335 73449 605391 73467
rect 605477 73449 605533 73467
rect 605619 73449 605675 73467
rect 605761 73449 605817 73467
rect 605903 73449 605959 73467
rect 606045 73449 606101 73467
rect 606187 73449 606243 73467
rect 606329 73449 606385 73467
rect 606471 73449 606527 73467
rect 606613 73449 606669 73467
rect 606755 73449 606811 73467
rect 606897 73449 606953 73467
rect 607039 73449 607095 73467
rect 605193 73411 605232 73449
rect 605232 73411 605249 73449
rect 605335 73411 605356 73449
rect 605356 73411 605391 73449
rect 605477 73411 605480 73449
rect 605480 73411 605533 73449
rect 605619 73411 605672 73449
rect 605672 73411 605675 73449
rect 605761 73411 605796 73449
rect 605796 73411 605817 73449
rect 605903 73411 605920 73449
rect 605920 73411 605959 73449
rect 606045 73411 606100 73449
rect 606100 73411 606101 73449
rect 606187 73411 606224 73449
rect 606224 73411 606243 73449
rect 606329 73411 606348 73449
rect 606348 73411 606385 73449
rect 606471 73411 606472 73449
rect 606472 73411 606527 73449
rect 606613 73411 606664 73449
rect 606664 73411 606669 73449
rect 606755 73411 606788 73449
rect 606788 73411 606811 73449
rect 606897 73411 606912 73449
rect 606912 73411 606953 73449
rect 607039 73411 607092 73449
rect 607092 73411 607095 73449
rect 605193 73269 605232 73325
rect 605232 73269 605249 73325
rect 605335 73269 605356 73325
rect 605356 73269 605391 73325
rect 605477 73269 605480 73325
rect 605480 73269 605533 73325
rect 605619 73269 605672 73325
rect 605672 73269 605675 73325
rect 605761 73269 605796 73325
rect 605796 73269 605817 73325
rect 605903 73269 605920 73325
rect 605920 73269 605959 73325
rect 606045 73269 606100 73325
rect 606100 73269 606101 73325
rect 606187 73269 606224 73325
rect 606224 73269 606243 73325
rect 606329 73269 606348 73325
rect 606348 73269 606385 73325
rect 606471 73269 606472 73325
rect 606472 73269 606527 73325
rect 606613 73269 606664 73325
rect 606664 73269 606669 73325
rect 606755 73269 606788 73325
rect 606788 73269 606811 73325
rect 606897 73269 606912 73325
rect 606912 73269 606953 73325
rect 607039 73269 607092 73325
rect 607092 73269 607095 73325
rect 605193 73145 605232 73183
rect 605232 73145 605249 73183
rect 605335 73145 605356 73183
rect 605356 73145 605391 73183
rect 605477 73145 605480 73183
rect 605480 73145 605533 73183
rect 605619 73145 605672 73183
rect 605672 73145 605675 73183
rect 605761 73145 605796 73183
rect 605796 73145 605817 73183
rect 605903 73145 605920 73183
rect 605920 73145 605959 73183
rect 606045 73145 606100 73183
rect 606100 73145 606101 73183
rect 606187 73145 606224 73183
rect 606224 73145 606243 73183
rect 606329 73145 606348 73183
rect 606348 73145 606385 73183
rect 606471 73145 606472 73183
rect 606472 73145 606527 73183
rect 606613 73145 606664 73183
rect 606664 73145 606669 73183
rect 606755 73145 606788 73183
rect 606788 73145 606811 73183
rect 606897 73145 606912 73183
rect 606912 73145 606953 73183
rect 607039 73145 607092 73183
rect 607092 73145 607095 73183
rect 605193 73127 605249 73145
rect 605335 73127 605391 73145
rect 605477 73127 605533 73145
rect 605619 73127 605675 73145
rect 605761 73127 605817 73145
rect 605903 73127 605959 73145
rect 606045 73127 606101 73145
rect 606187 73127 606243 73145
rect 606329 73127 606385 73145
rect 606471 73127 606527 73145
rect 606613 73127 606669 73145
rect 606755 73127 606811 73145
rect 606897 73127 606953 73145
rect 607039 73127 607095 73145
rect 605193 73021 605232 73041
rect 605232 73021 605249 73041
rect 605335 73021 605356 73041
rect 605356 73021 605391 73041
rect 605477 73021 605480 73041
rect 605480 73021 605533 73041
rect 605619 73021 605672 73041
rect 605672 73021 605675 73041
rect 605761 73021 605796 73041
rect 605796 73021 605817 73041
rect 605903 73021 605920 73041
rect 605920 73021 605959 73041
rect 606045 73021 606100 73041
rect 606100 73021 606101 73041
rect 606187 73021 606224 73041
rect 606224 73021 606243 73041
rect 606329 73021 606348 73041
rect 606348 73021 606385 73041
rect 606471 73021 606472 73041
rect 606472 73021 606527 73041
rect 606613 73021 606664 73041
rect 606664 73021 606669 73041
rect 606755 73021 606788 73041
rect 606788 73021 606811 73041
rect 606897 73021 606912 73041
rect 606912 73021 606953 73041
rect 607039 73021 607092 73041
rect 607092 73021 607095 73041
rect 605193 72985 605249 73021
rect 605335 72985 605391 73021
rect 605477 72985 605533 73021
rect 605619 72985 605675 73021
rect 605761 72985 605817 73021
rect 605903 72985 605959 73021
rect 606045 72985 606101 73021
rect 606187 72985 606243 73021
rect 606329 72985 606385 73021
rect 606471 72985 606527 73021
rect 606613 72985 606669 73021
rect 606755 72985 606811 73021
rect 606897 72985 606953 73021
rect 607039 72985 607095 73021
rect 605193 72897 605232 72899
rect 605232 72897 605249 72899
rect 605335 72897 605356 72899
rect 605356 72897 605391 72899
rect 605477 72897 605480 72899
rect 605480 72897 605533 72899
rect 605619 72897 605672 72899
rect 605672 72897 605675 72899
rect 605761 72897 605796 72899
rect 605796 72897 605817 72899
rect 605903 72897 605920 72899
rect 605920 72897 605959 72899
rect 606045 72897 606100 72899
rect 606100 72897 606101 72899
rect 606187 72897 606224 72899
rect 606224 72897 606243 72899
rect 606329 72897 606348 72899
rect 606348 72897 606385 72899
rect 606471 72897 606472 72899
rect 606472 72897 606527 72899
rect 606613 72897 606664 72899
rect 606664 72897 606669 72899
rect 606755 72897 606788 72899
rect 606788 72897 606811 72899
rect 606897 72897 606912 72899
rect 606912 72897 606953 72899
rect 607039 72897 607092 72899
rect 607092 72897 607095 72899
rect 605193 72843 605249 72897
rect 605335 72843 605391 72897
rect 605477 72843 605533 72897
rect 605619 72843 605675 72897
rect 605761 72843 605817 72897
rect 605903 72843 605959 72897
rect 606045 72843 606101 72897
rect 606187 72843 606243 72897
rect 606329 72843 606385 72897
rect 606471 72843 606527 72897
rect 606613 72843 606669 72897
rect 606755 72843 606811 72897
rect 606897 72843 606953 72897
rect 607039 72843 607095 72897
rect 605193 72705 605249 72757
rect 605335 72705 605391 72757
rect 605477 72705 605533 72757
rect 605619 72705 605675 72757
rect 605761 72705 605817 72757
rect 605903 72705 605959 72757
rect 606045 72705 606101 72757
rect 606187 72705 606243 72757
rect 606329 72705 606385 72757
rect 606471 72705 606527 72757
rect 606613 72705 606669 72757
rect 606755 72705 606811 72757
rect 606897 72705 606953 72757
rect 607039 72705 607095 72757
rect 605193 72701 605232 72705
rect 605232 72701 605249 72705
rect 605335 72701 605356 72705
rect 605356 72701 605391 72705
rect 605477 72701 605480 72705
rect 605480 72701 605533 72705
rect 605619 72701 605672 72705
rect 605672 72701 605675 72705
rect 605761 72701 605796 72705
rect 605796 72701 605817 72705
rect 605903 72701 605920 72705
rect 605920 72701 605959 72705
rect 606045 72701 606100 72705
rect 606100 72701 606101 72705
rect 606187 72701 606224 72705
rect 606224 72701 606243 72705
rect 606329 72701 606348 72705
rect 606348 72701 606385 72705
rect 606471 72701 606472 72705
rect 606472 72701 606527 72705
rect 606613 72701 606664 72705
rect 606664 72701 606669 72705
rect 606755 72701 606788 72705
rect 606788 72701 606811 72705
rect 606897 72701 606912 72705
rect 606912 72701 606953 72705
rect 607039 72701 607092 72705
rect 607092 72701 607095 72705
rect 605193 72581 605249 72615
rect 605335 72581 605391 72615
rect 605477 72581 605533 72615
rect 605619 72581 605675 72615
rect 605761 72581 605817 72615
rect 605903 72581 605959 72615
rect 606045 72581 606101 72615
rect 606187 72581 606243 72615
rect 606329 72581 606385 72615
rect 606471 72581 606527 72615
rect 606613 72581 606669 72615
rect 606755 72581 606811 72615
rect 606897 72581 606953 72615
rect 607039 72581 607095 72615
rect 605193 72559 605232 72581
rect 605232 72559 605249 72581
rect 605335 72559 605356 72581
rect 605356 72559 605391 72581
rect 605477 72559 605480 72581
rect 605480 72559 605533 72581
rect 605619 72559 605672 72581
rect 605672 72559 605675 72581
rect 605761 72559 605796 72581
rect 605796 72559 605817 72581
rect 605903 72559 605920 72581
rect 605920 72559 605959 72581
rect 606045 72559 606100 72581
rect 606100 72559 606101 72581
rect 606187 72559 606224 72581
rect 606224 72559 606243 72581
rect 606329 72559 606348 72581
rect 606348 72559 606385 72581
rect 606471 72559 606472 72581
rect 606472 72559 606527 72581
rect 606613 72559 606664 72581
rect 606664 72559 606669 72581
rect 606755 72559 606788 72581
rect 606788 72559 606811 72581
rect 606897 72559 606912 72581
rect 606912 72559 606953 72581
rect 607039 72559 607092 72581
rect 607092 72559 607095 72581
rect 605193 72457 605249 72473
rect 605335 72457 605391 72473
rect 605477 72457 605533 72473
rect 605619 72457 605675 72473
rect 605761 72457 605817 72473
rect 605903 72457 605959 72473
rect 606045 72457 606101 72473
rect 606187 72457 606243 72473
rect 606329 72457 606385 72473
rect 606471 72457 606527 72473
rect 606613 72457 606669 72473
rect 606755 72457 606811 72473
rect 606897 72457 606953 72473
rect 607039 72457 607095 72473
rect 605193 72417 605232 72457
rect 605232 72417 605249 72457
rect 605335 72417 605356 72457
rect 605356 72417 605391 72457
rect 605477 72417 605480 72457
rect 605480 72417 605533 72457
rect 605619 72417 605672 72457
rect 605672 72417 605675 72457
rect 605761 72417 605796 72457
rect 605796 72417 605817 72457
rect 605903 72417 605920 72457
rect 605920 72417 605959 72457
rect 606045 72417 606100 72457
rect 606100 72417 606101 72457
rect 606187 72417 606224 72457
rect 606224 72417 606243 72457
rect 606329 72417 606348 72457
rect 606348 72417 606385 72457
rect 606471 72417 606472 72457
rect 606472 72417 606527 72457
rect 606613 72417 606664 72457
rect 606664 72417 606669 72457
rect 606755 72417 606788 72457
rect 606788 72417 606811 72457
rect 606897 72417 606912 72457
rect 606912 72417 606953 72457
rect 607039 72417 607092 72457
rect 607092 72417 607095 72457
rect 605193 72277 605232 72331
rect 605232 72277 605249 72331
rect 605335 72277 605356 72331
rect 605356 72277 605391 72331
rect 605477 72277 605480 72331
rect 605480 72277 605533 72331
rect 605619 72277 605672 72331
rect 605672 72277 605675 72331
rect 605761 72277 605796 72331
rect 605796 72277 605817 72331
rect 605903 72277 605920 72331
rect 605920 72277 605959 72331
rect 606045 72277 606100 72331
rect 606100 72277 606101 72331
rect 606187 72277 606224 72331
rect 606224 72277 606243 72331
rect 606329 72277 606348 72331
rect 606348 72277 606385 72331
rect 606471 72277 606472 72331
rect 606472 72277 606527 72331
rect 606613 72277 606664 72331
rect 606664 72277 606669 72331
rect 606755 72277 606788 72331
rect 606788 72277 606811 72331
rect 606897 72277 606912 72331
rect 606912 72277 606953 72331
rect 607039 72277 607092 72331
rect 607092 72277 607095 72331
rect 605193 72275 605249 72277
rect 605335 72275 605391 72277
rect 605477 72275 605533 72277
rect 605619 72275 605675 72277
rect 605761 72275 605817 72277
rect 605903 72275 605959 72277
rect 606045 72275 606101 72277
rect 606187 72275 606243 72277
rect 606329 72275 606385 72277
rect 606471 72275 606527 72277
rect 606613 72275 606669 72277
rect 606755 72275 606811 72277
rect 606897 72275 606953 72277
rect 607039 72275 607095 72277
rect 605193 72153 605232 72189
rect 605232 72153 605249 72189
rect 605335 72153 605356 72189
rect 605356 72153 605391 72189
rect 605477 72153 605480 72189
rect 605480 72153 605533 72189
rect 605619 72153 605672 72189
rect 605672 72153 605675 72189
rect 605761 72153 605796 72189
rect 605796 72153 605817 72189
rect 605903 72153 605920 72189
rect 605920 72153 605959 72189
rect 606045 72153 606100 72189
rect 606100 72153 606101 72189
rect 606187 72153 606224 72189
rect 606224 72153 606243 72189
rect 606329 72153 606348 72189
rect 606348 72153 606385 72189
rect 606471 72153 606472 72189
rect 606472 72153 606527 72189
rect 606613 72153 606664 72189
rect 606664 72153 606669 72189
rect 606755 72153 606788 72189
rect 606788 72153 606811 72189
rect 606897 72153 606912 72189
rect 606912 72153 606953 72189
rect 607039 72153 607092 72189
rect 607092 72153 607095 72189
rect 605193 72133 605249 72153
rect 605335 72133 605391 72153
rect 605477 72133 605533 72153
rect 605619 72133 605675 72153
rect 605761 72133 605817 72153
rect 605903 72133 605959 72153
rect 606045 72133 606101 72153
rect 606187 72133 606243 72153
rect 606329 72133 606385 72153
rect 606471 72133 606527 72153
rect 606613 72133 606669 72153
rect 606755 72133 606811 72153
rect 606897 72133 606953 72153
rect 607039 72133 607095 72153
rect 607899 73979 607955 74035
rect 608041 73979 608097 74035
rect 608183 73979 608239 74035
rect 608325 73979 608381 74035
rect 608467 73979 608523 74035
rect 608609 73979 608665 74035
rect 608751 73979 608807 74035
rect 608893 73979 608949 74035
rect 609035 73979 609091 74035
rect 609177 73979 609233 74035
rect 609319 73979 609375 74035
rect 609461 73979 609517 74035
rect 609603 73979 609659 74035
rect 609745 73979 609801 74035
rect 607899 73889 607938 73893
rect 607938 73889 607955 73893
rect 608041 73889 608062 73893
rect 608062 73889 608097 73893
rect 608183 73889 608186 73893
rect 608186 73889 608239 73893
rect 608325 73889 608378 73893
rect 608378 73889 608381 73893
rect 608467 73889 608502 73893
rect 608502 73889 608523 73893
rect 608609 73889 608626 73893
rect 608626 73889 608665 73893
rect 608751 73889 608806 73893
rect 608806 73889 608807 73893
rect 608893 73889 608930 73893
rect 608930 73889 608949 73893
rect 609035 73889 609054 73893
rect 609054 73889 609091 73893
rect 609177 73889 609178 73893
rect 609178 73889 609233 73893
rect 609319 73889 609370 73893
rect 609370 73889 609375 73893
rect 609461 73889 609494 73893
rect 609494 73889 609517 73893
rect 609603 73889 609618 73893
rect 609618 73889 609659 73893
rect 609745 73889 609798 73893
rect 609798 73889 609801 73893
rect 607899 73837 607955 73889
rect 608041 73837 608097 73889
rect 608183 73837 608239 73889
rect 608325 73837 608381 73889
rect 608467 73837 608523 73889
rect 608609 73837 608665 73889
rect 608751 73837 608807 73889
rect 608893 73837 608949 73889
rect 609035 73837 609091 73889
rect 609177 73837 609233 73889
rect 609319 73837 609375 73889
rect 609461 73837 609517 73889
rect 609603 73837 609659 73889
rect 609745 73837 609801 73889
rect 607899 73697 607955 73751
rect 608041 73697 608097 73751
rect 608183 73697 608239 73751
rect 608325 73697 608381 73751
rect 608467 73697 608523 73751
rect 608609 73697 608665 73751
rect 608751 73697 608807 73751
rect 608893 73697 608949 73751
rect 609035 73697 609091 73751
rect 609177 73697 609233 73751
rect 609319 73697 609375 73751
rect 609461 73697 609517 73751
rect 609603 73697 609659 73751
rect 609745 73697 609801 73751
rect 607899 73695 607938 73697
rect 607938 73695 607955 73697
rect 608041 73695 608062 73697
rect 608062 73695 608097 73697
rect 608183 73695 608186 73697
rect 608186 73695 608239 73697
rect 608325 73695 608378 73697
rect 608378 73695 608381 73697
rect 608467 73695 608502 73697
rect 608502 73695 608523 73697
rect 608609 73695 608626 73697
rect 608626 73695 608665 73697
rect 608751 73695 608806 73697
rect 608806 73695 608807 73697
rect 608893 73695 608930 73697
rect 608930 73695 608949 73697
rect 609035 73695 609054 73697
rect 609054 73695 609091 73697
rect 609177 73695 609178 73697
rect 609178 73695 609233 73697
rect 609319 73695 609370 73697
rect 609370 73695 609375 73697
rect 609461 73695 609494 73697
rect 609494 73695 609517 73697
rect 609603 73695 609618 73697
rect 609618 73695 609659 73697
rect 609745 73695 609798 73697
rect 609798 73695 609801 73697
rect 607899 73573 607955 73609
rect 608041 73573 608097 73609
rect 608183 73573 608239 73609
rect 608325 73573 608381 73609
rect 608467 73573 608523 73609
rect 608609 73573 608665 73609
rect 608751 73573 608807 73609
rect 608893 73573 608949 73609
rect 609035 73573 609091 73609
rect 609177 73573 609233 73609
rect 609319 73573 609375 73609
rect 609461 73573 609517 73609
rect 609603 73573 609659 73609
rect 609745 73573 609801 73609
rect 607899 73553 607938 73573
rect 607938 73553 607955 73573
rect 608041 73553 608062 73573
rect 608062 73553 608097 73573
rect 608183 73553 608186 73573
rect 608186 73553 608239 73573
rect 608325 73553 608378 73573
rect 608378 73553 608381 73573
rect 608467 73553 608502 73573
rect 608502 73553 608523 73573
rect 608609 73553 608626 73573
rect 608626 73553 608665 73573
rect 608751 73553 608806 73573
rect 608806 73553 608807 73573
rect 608893 73553 608930 73573
rect 608930 73553 608949 73573
rect 609035 73553 609054 73573
rect 609054 73553 609091 73573
rect 609177 73553 609178 73573
rect 609178 73553 609233 73573
rect 609319 73553 609370 73573
rect 609370 73553 609375 73573
rect 609461 73553 609494 73573
rect 609494 73553 609517 73573
rect 609603 73553 609618 73573
rect 609618 73553 609659 73573
rect 609745 73553 609798 73573
rect 609798 73553 609801 73573
rect 607899 73449 607955 73467
rect 608041 73449 608097 73467
rect 608183 73449 608239 73467
rect 608325 73449 608381 73467
rect 608467 73449 608523 73467
rect 608609 73449 608665 73467
rect 608751 73449 608807 73467
rect 608893 73449 608949 73467
rect 609035 73449 609091 73467
rect 609177 73449 609233 73467
rect 609319 73449 609375 73467
rect 609461 73449 609517 73467
rect 609603 73449 609659 73467
rect 609745 73449 609801 73467
rect 607899 73411 607938 73449
rect 607938 73411 607955 73449
rect 608041 73411 608062 73449
rect 608062 73411 608097 73449
rect 608183 73411 608186 73449
rect 608186 73411 608239 73449
rect 608325 73411 608378 73449
rect 608378 73411 608381 73449
rect 608467 73411 608502 73449
rect 608502 73411 608523 73449
rect 608609 73411 608626 73449
rect 608626 73411 608665 73449
rect 608751 73411 608806 73449
rect 608806 73411 608807 73449
rect 608893 73411 608930 73449
rect 608930 73411 608949 73449
rect 609035 73411 609054 73449
rect 609054 73411 609091 73449
rect 609177 73411 609178 73449
rect 609178 73411 609233 73449
rect 609319 73411 609370 73449
rect 609370 73411 609375 73449
rect 609461 73411 609494 73449
rect 609494 73411 609517 73449
rect 609603 73411 609618 73449
rect 609618 73411 609659 73449
rect 609745 73411 609798 73449
rect 609798 73411 609801 73449
rect 607899 73269 607938 73325
rect 607938 73269 607955 73325
rect 608041 73269 608062 73325
rect 608062 73269 608097 73325
rect 608183 73269 608186 73325
rect 608186 73269 608239 73325
rect 608325 73269 608378 73325
rect 608378 73269 608381 73325
rect 608467 73269 608502 73325
rect 608502 73269 608523 73325
rect 608609 73269 608626 73325
rect 608626 73269 608665 73325
rect 608751 73269 608806 73325
rect 608806 73269 608807 73325
rect 608893 73269 608930 73325
rect 608930 73269 608949 73325
rect 609035 73269 609054 73325
rect 609054 73269 609091 73325
rect 609177 73269 609178 73325
rect 609178 73269 609233 73325
rect 609319 73269 609370 73325
rect 609370 73269 609375 73325
rect 609461 73269 609494 73325
rect 609494 73269 609517 73325
rect 609603 73269 609618 73325
rect 609618 73269 609659 73325
rect 609745 73269 609798 73325
rect 609798 73269 609801 73325
rect 607899 73145 607938 73183
rect 607938 73145 607955 73183
rect 608041 73145 608062 73183
rect 608062 73145 608097 73183
rect 608183 73145 608186 73183
rect 608186 73145 608239 73183
rect 608325 73145 608378 73183
rect 608378 73145 608381 73183
rect 608467 73145 608502 73183
rect 608502 73145 608523 73183
rect 608609 73145 608626 73183
rect 608626 73145 608665 73183
rect 608751 73145 608806 73183
rect 608806 73145 608807 73183
rect 608893 73145 608930 73183
rect 608930 73145 608949 73183
rect 609035 73145 609054 73183
rect 609054 73145 609091 73183
rect 609177 73145 609178 73183
rect 609178 73145 609233 73183
rect 609319 73145 609370 73183
rect 609370 73145 609375 73183
rect 609461 73145 609494 73183
rect 609494 73145 609517 73183
rect 609603 73145 609618 73183
rect 609618 73145 609659 73183
rect 609745 73145 609798 73183
rect 609798 73145 609801 73183
rect 607899 73127 607955 73145
rect 608041 73127 608097 73145
rect 608183 73127 608239 73145
rect 608325 73127 608381 73145
rect 608467 73127 608523 73145
rect 608609 73127 608665 73145
rect 608751 73127 608807 73145
rect 608893 73127 608949 73145
rect 609035 73127 609091 73145
rect 609177 73127 609233 73145
rect 609319 73127 609375 73145
rect 609461 73127 609517 73145
rect 609603 73127 609659 73145
rect 609745 73127 609801 73145
rect 607899 73021 607938 73041
rect 607938 73021 607955 73041
rect 608041 73021 608062 73041
rect 608062 73021 608097 73041
rect 608183 73021 608186 73041
rect 608186 73021 608239 73041
rect 608325 73021 608378 73041
rect 608378 73021 608381 73041
rect 608467 73021 608502 73041
rect 608502 73021 608523 73041
rect 608609 73021 608626 73041
rect 608626 73021 608665 73041
rect 608751 73021 608806 73041
rect 608806 73021 608807 73041
rect 608893 73021 608930 73041
rect 608930 73021 608949 73041
rect 609035 73021 609054 73041
rect 609054 73021 609091 73041
rect 609177 73021 609178 73041
rect 609178 73021 609233 73041
rect 609319 73021 609370 73041
rect 609370 73021 609375 73041
rect 609461 73021 609494 73041
rect 609494 73021 609517 73041
rect 609603 73021 609618 73041
rect 609618 73021 609659 73041
rect 609745 73021 609798 73041
rect 609798 73021 609801 73041
rect 607899 72985 607955 73021
rect 608041 72985 608097 73021
rect 608183 72985 608239 73021
rect 608325 72985 608381 73021
rect 608467 72985 608523 73021
rect 608609 72985 608665 73021
rect 608751 72985 608807 73021
rect 608893 72985 608949 73021
rect 609035 72985 609091 73021
rect 609177 72985 609233 73021
rect 609319 72985 609375 73021
rect 609461 72985 609517 73021
rect 609603 72985 609659 73021
rect 609745 72985 609801 73021
rect 607899 72897 607938 72899
rect 607938 72897 607955 72899
rect 608041 72897 608062 72899
rect 608062 72897 608097 72899
rect 608183 72897 608186 72899
rect 608186 72897 608239 72899
rect 608325 72897 608378 72899
rect 608378 72897 608381 72899
rect 608467 72897 608502 72899
rect 608502 72897 608523 72899
rect 608609 72897 608626 72899
rect 608626 72897 608665 72899
rect 608751 72897 608806 72899
rect 608806 72897 608807 72899
rect 608893 72897 608930 72899
rect 608930 72897 608949 72899
rect 609035 72897 609054 72899
rect 609054 72897 609091 72899
rect 609177 72897 609178 72899
rect 609178 72897 609233 72899
rect 609319 72897 609370 72899
rect 609370 72897 609375 72899
rect 609461 72897 609494 72899
rect 609494 72897 609517 72899
rect 609603 72897 609618 72899
rect 609618 72897 609659 72899
rect 609745 72897 609798 72899
rect 609798 72897 609801 72899
rect 607899 72843 607955 72897
rect 608041 72843 608097 72897
rect 608183 72843 608239 72897
rect 608325 72843 608381 72897
rect 608467 72843 608523 72897
rect 608609 72843 608665 72897
rect 608751 72843 608807 72897
rect 608893 72843 608949 72897
rect 609035 72843 609091 72897
rect 609177 72843 609233 72897
rect 609319 72843 609375 72897
rect 609461 72843 609517 72897
rect 609603 72843 609659 72897
rect 609745 72843 609801 72897
rect 607899 72705 607955 72757
rect 608041 72705 608097 72757
rect 608183 72705 608239 72757
rect 608325 72705 608381 72757
rect 608467 72705 608523 72757
rect 608609 72705 608665 72757
rect 608751 72705 608807 72757
rect 608893 72705 608949 72757
rect 609035 72705 609091 72757
rect 609177 72705 609233 72757
rect 609319 72705 609375 72757
rect 609461 72705 609517 72757
rect 609603 72705 609659 72757
rect 609745 72705 609801 72757
rect 607899 72701 607938 72705
rect 607938 72701 607955 72705
rect 608041 72701 608062 72705
rect 608062 72701 608097 72705
rect 608183 72701 608186 72705
rect 608186 72701 608239 72705
rect 608325 72701 608378 72705
rect 608378 72701 608381 72705
rect 608467 72701 608502 72705
rect 608502 72701 608523 72705
rect 608609 72701 608626 72705
rect 608626 72701 608665 72705
rect 608751 72701 608806 72705
rect 608806 72701 608807 72705
rect 608893 72701 608930 72705
rect 608930 72701 608949 72705
rect 609035 72701 609054 72705
rect 609054 72701 609091 72705
rect 609177 72701 609178 72705
rect 609178 72701 609233 72705
rect 609319 72701 609370 72705
rect 609370 72701 609375 72705
rect 609461 72701 609494 72705
rect 609494 72701 609517 72705
rect 609603 72701 609618 72705
rect 609618 72701 609659 72705
rect 609745 72701 609798 72705
rect 609798 72701 609801 72705
rect 607899 72581 607955 72615
rect 608041 72581 608097 72615
rect 608183 72581 608239 72615
rect 608325 72581 608381 72615
rect 608467 72581 608523 72615
rect 608609 72581 608665 72615
rect 608751 72581 608807 72615
rect 608893 72581 608949 72615
rect 609035 72581 609091 72615
rect 609177 72581 609233 72615
rect 609319 72581 609375 72615
rect 609461 72581 609517 72615
rect 609603 72581 609659 72615
rect 609745 72581 609801 72615
rect 607899 72559 607938 72581
rect 607938 72559 607955 72581
rect 608041 72559 608062 72581
rect 608062 72559 608097 72581
rect 608183 72559 608186 72581
rect 608186 72559 608239 72581
rect 608325 72559 608378 72581
rect 608378 72559 608381 72581
rect 608467 72559 608502 72581
rect 608502 72559 608523 72581
rect 608609 72559 608626 72581
rect 608626 72559 608665 72581
rect 608751 72559 608806 72581
rect 608806 72559 608807 72581
rect 608893 72559 608930 72581
rect 608930 72559 608949 72581
rect 609035 72559 609054 72581
rect 609054 72559 609091 72581
rect 609177 72559 609178 72581
rect 609178 72559 609233 72581
rect 609319 72559 609370 72581
rect 609370 72559 609375 72581
rect 609461 72559 609494 72581
rect 609494 72559 609517 72581
rect 609603 72559 609618 72581
rect 609618 72559 609659 72581
rect 609745 72559 609798 72581
rect 609798 72559 609801 72581
rect 607899 72457 607955 72473
rect 608041 72457 608097 72473
rect 608183 72457 608239 72473
rect 608325 72457 608381 72473
rect 608467 72457 608523 72473
rect 608609 72457 608665 72473
rect 608751 72457 608807 72473
rect 608893 72457 608949 72473
rect 609035 72457 609091 72473
rect 609177 72457 609233 72473
rect 609319 72457 609375 72473
rect 609461 72457 609517 72473
rect 609603 72457 609659 72473
rect 609745 72457 609801 72473
rect 607899 72417 607938 72457
rect 607938 72417 607955 72457
rect 608041 72417 608062 72457
rect 608062 72417 608097 72457
rect 608183 72417 608186 72457
rect 608186 72417 608239 72457
rect 608325 72417 608378 72457
rect 608378 72417 608381 72457
rect 608467 72417 608502 72457
rect 608502 72417 608523 72457
rect 608609 72417 608626 72457
rect 608626 72417 608665 72457
rect 608751 72417 608806 72457
rect 608806 72417 608807 72457
rect 608893 72417 608930 72457
rect 608930 72417 608949 72457
rect 609035 72417 609054 72457
rect 609054 72417 609091 72457
rect 609177 72417 609178 72457
rect 609178 72417 609233 72457
rect 609319 72417 609370 72457
rect 609370 72417 609375 72457
rect 609461 72417 609494 72457
rect 609494 72417 609517 72457
rect 609603 72417 609618 72457
rect 609618 72417 609659 72457
rect 609745 72417 609798 72457
rect 609798 72417 609801 72457
rect 607899 72277 607938 72331
rect 607938 72277 607955 72331
rect 608041 72277 608062 72331
rect 608062 72277 608097 72331
rect 608183 72277 608186 72331
rect 608186 72277 608239 72331
rect 608325 72277 608378 72331
rect 608378 72277 608381 72331
rect 608467 72277 608502 72331
rect 608502 72277 608523 72331
rect 608609 72277 608626 72331
rect 608626 72277 608665 72331
rect 608751 72277 608806 72331
rect 608806 72277 608807 72331
rect 608893 72277 608930 72331
rect 608930 72277 608949 72331
rect 609035 72277 609054 72331
rect 609054 72277 609091 72331
rect 609177 72277 609178 72331
rect 609178 72277 609233 72331
rect 609319 72277 609370 72331
rect 609370 72277 609375 72331
rect 609461 72277 609494 72331
rect 609494 72277 609517 72331
rect 609603 72277 609618 72331
rect 609618 72277 609659 72331
rect 609745 72277 609798 72331
rect 609798 72277 609801 72331
rect 607899 72275 607955 72277
rect 608041 72275 608097 72277
rect 608183 72275 608239 72277
rect 608325 72275 608381 72277
rect 608467 72275 608523 72277
rect 608609 72275 608665 72277
rect 608751 72275 608807 72277
rect 608893 72275 608949 72277
rect 609035 72275 609091 72277
rect 609177 72275 609233 72277
rect 609319 72275 609375 72277
rect 609461 72275 609517 72277
rect 609603 72275 609659 72277
rect 609745 72275 609801 72277
rect 607899 72153 607938 72189
rect 607938 72153 607955 72189
rect 608041 72153 608062 72189
rect 608062 72153 608097 72189
rect 608183 72153 608186 72189
rect 608186 72153 608239 72189
rect 608325 72153 608378 72189
rect 608378 72153 608381 72189
rect 608467 72153 608502 72189
rect 608502 72153 608523 72189
rect 608609 72153 608626 72189
rect 608626 72153 608665 72189
rect 608751 72153 608806 72189
rect 608806 72153 608807 72189
rect 608893 72153 608930 72189
rect 608930 72153 608949 72189
rect 609035 72153 609054 72189
rect 609054 72153 609091 72189
rect 609177 72153 609178 72189
rect 609178 72153 609233 72189
rect 609319 72153 609370 72189
rect 609370 72153 609375 72189
rect 609461 72153 609494 72189
rect 609494 72153 609517 72189
rect 609603 72153 609618 72189
rect 609618 72153 609659 72189
rect 609745 72153 609798 72189
rect 609798 72153 609801 72189
rect 607899 72133 607955 72153
rect 608041 72133 608097 72153
rect 608183 72133 608239 72153
rect 608325 72133 608381 72153
rect 608467 72133 608523 72153
rect 608609 72133 608665 72153
rect 608751 72133 608807 72153
rect 608893 72133 608949 72153
rect 609035 72133 609091 72153
rect 609177 72133 609233 72153
rect 609319 72133 609375 72153
rect 609461 72133 609517 72153
rect 609603 72133 609659 72153
rect 609745 72133 609801 72153
rect 610269 73979 610325 74035
rect 610411 73979 610467 74035
rect 610553 73979 610609 74035
rect 610695 73979 610751 74035
rect 610837 73979 610893 74035
rect 610979 73979 611035 74035
rect 611121 73979 611177 74035
rect 611263 73979 611319 74035
rect 611405 73979 611461 74035
rect 611547 73979 611603 74035
rect 611689 73979 611745 74035
rect 611831 73979 611887 74035
rect 611973 73979 612029 74035
rect 612115 73979 612171 74035
rect 610269 73889 610308 73893
rect 610308 73889 610325 73893
rect 610411 73889 610432 73893
rect 610432 73889 610467 73893
rect 610553 73889 610556 73893
rect 610556 73889 610609 73893
rect 610695 73889 610748 73893
rect 610748 73889 610751 73893
rect 610837 73889 610872 73893
rect 610872 73889 610893 73893
rect 610979 73889 610996 73893
rect 610996 73889 611035 73893
rect 611121 73889 611176 73893
rect 611176 73889 611177 73893
rect 611263 73889 611300 73893
rect 611300 73889 611319 73893
rect 611405 73889 611424 73893
rect 611424 73889 611461 73893
rect 611547 73889 611548 73893
rect 611548 73889 611603 73893
rect 611689 73889 611740 73893
rect 611740 73889 611745 73893
rect 611831 73889 611864 73893
rect 611864 73889 611887 73893
rect 611973 73889 611988 73893
rect 611988 73889 612029 73893
rect 612115 73889 612168 73893
rect 612168 73889 612171 73893
rect 610269 73837 610325 73889
rect 610411 73837 610467 73889
rect 610553 73837 610609 73889
rect 610695 73837 610751 73889
rect 610837 73837 610893 73889
rect 610979 73837 611035 73889
rect 611121 73837 611177 73889
rect 611263 73837 611319 73889
rect 611405 73837 611461 73889
rect 611547 73837 611603 73889
rect 611689 73837 611745 73889
rect 611831 73837 611887 73889
rect 611973 73837 612029 73889
rect 612115 73837 612171 73889
rect 610269 73697 610325 73751
rect 610411 73697 610467 73751
rect 610553 73697 610609 73751
rect 610695 73697 610751 73751
rect 610837 73697 610893 73751
rect 610979 73697 611035 73751
rect 611121 73697 611177 73751
rect 611263 73697 611319 73751
rect 611405 73697 611461 73751
rect 611547 73697 611603 73751
rect 611689 73697 611745 73751
rect 611831 73697 611887 73751
rect 611973 73697 612029 73751
rect 612115 73697 612171 73751
rect 610269 73695 610308 73697
rect 610308 73695 610325 73697
rect 610411 73695 610432 73697
rect 610432 73695 610467 73697
rect 610553 73695 610556 73697
rect 610556 73695 610609 73697
rect 610695 73695 610748 73697
rect 610748 73695 610751 73697
rect 610837 73695 610872 73697
rect 610872 73695 610893 73697
rect 610979 73695 610996 73697
rect 610996 73695 611035 73697
rect 611121 73695 611176 73697
rect 611176 73695 611177 73697
rect 611263 73695 611300 73697
rect 611300 73695 611319 73697
rect 611405 73695 611424 73697
rect 611424 73695 611461 73697
rect 611547 73695 611548 73697
rect 611548 73695 611603 73697
rect 611689 73695 611740 73697
rect 611740 73695 611745 73697
rect 611831 73695 611864 73697
rect 611864 73695 611887 73697
rect 611973 73695 611988 73697
rect 611988 73695 612029 73697
rect 612115 73695 612168 73697
rect 612168 73695 612171 73697
rect 610269 73573 610325 73609
rect 610411 73573 610467 73609
rect 610553 73573 610609 73609
rect 610695 73573 610751 73609
rect 610837 73573 610893 73609
rect 610979 73573 611035 73609
rect 611121 73573 611177 73609
rect 611263 73573 611319 73609
rect 611405 73573 611461 73609
rect 611547 73573 611603 73609
rect 611689 73573 611745 73609
rect 611831 73573 611887 73609
rect 611973 73573 612029 73609
rect 612115 73573 612171 73609
rect 610269 73553 610308 73573
rect 610308 73553 610325 73573
rect 610411 73553 610432 73573
rect 610432 73553 610467 73573
rect 610553 73553 610556 73573
rect 610556 73553 610609 73573
rect 610695 73553 610748 73573
rect 610748 73553 610751 73573
rect 610837 73553 610872 73573
rect 610872 73553 610893 73573
rect 610979 73553 610996 73573
rect 610996 73553 611035 73573
rect 611121 73553 611176 73573
rect 611176 73553 611177 73573
rect 611263 73553 611300 73573
rect 611300 73553 611319 73573
rect 611405 73553 611424 73573
rect 611424 73553 611461 73573
rect 611547 73553 611548 73573
rect 611548 73553 611603 73573
rect 611689 73553 611740 73573
rect 611740 73553 611745 73573
rect 611831 73553 611864 73573
rect 611864 73553 611887 73573
rect 611973 73553 611988 73573
rect 611988 73553 612029 73573
rect 612115 73553 612168 73573
rect 612168 73553 612171 73573
rect 610269 73449 610325 73467
rect 610411 73449 610467 73467
rect 610553 73449 610609 73467
rect 610695 73449 610751 73467
rect 610837 73449 610893 73467
rect 610979 73449 611035 73467
rect 611121 73449 611177 73467
rect 611263 73449 611319 73467
rect 611405 73449 611461 73467
rect 611547 73449 611603 73467
rect 611689 73449 611745 73467
rect 611831 73449 611887 73467
rect 611973 73449 612029 73467
rect 612115 73449 612171 73467
rect 610269 73411 610308 73449
rect 610308 73411 610325 73449
rect 610411 73411 610432 73449
rect 610432 73411 610467 73449
rect 610553 73411 610556 73449
rect 610556 73411 610609 73449
rect 610695 73411 610748 73449
rect 610748 73411 610751 73449
rect 610837 73411 610872 73449
rect 610872 73411 610893 73449
rect 610979 73411 610996 73449
rect 610996 73411 611035 73449
rect 611121 73411 611176 73449
rect 611176 73411 611177 73449
rect 611263 73411 611300 73449
rect 611300 73411 611319 73449
rect 611405 73411 611424 73449
rect 611424 73411 611461 73449
rect 611547 73411 611548 73449
rect 611548 73411 611603 73449
rect 611689 73411 611740 73449
rect 611740 73411 611745 73449
rect 611831 73411 611864 73449
rect 611864 73411 611887 73449
rect 611973 73411 611988 73449
rect 611988 73411 612029 73449
rect 612115 73411 612168 73449
rect 612168 73411 612171 73449
rect 610269 73269 610308 73325
rect 610308 73269 610325 73325
rect 610411 73269 610432 73325
rect 610432 73269 610467 73325
rect 610553 73269 610556 73325
rect 610556 73269 610609 73325
rect 610695 73269 610748 73325
rect 610748 73269 610751 73325
rect 610837 73269 610872 73325
rect 610872 73269 610893 73325
rect 610979 73269 610996 73325
rect 610996 73269 611035 73325
rect 611121 73269 611176 73325
rect 611176 73269 611177 73325
rect 611263 73269 611300 73325
rect 611300 73269 611319 73325
rect 611405 73269 611424 73325
rect 611424 73269 611461 73325
rect 611547 73269 611548 73325
rect 611548 73269 611603 73325
rect 611689 73269 611740 73325
rect 611740 73269 611745 73325
rect 611831 73269 611864 73325
rect 611864 73269 611887 73325
rect 611973 73269 611988 73325
rect 611988 73269 612029 73325
rect 612115 73269 612168 73325
rect 612168 73269 612171 73325
rect 610269 73145 610308 73183
rect 610308 73145 610325 73183
rect 610411 73145 610432 73183
rect 610432 73145 610467 73183
rect 610553 73145 610556 73183
rect 610556 73145 610609 73183
rect 610695 73145 610748 73183
rect 610748 73145 610751 73183
rect 610837 73145 610872 73183
rect 610872 73145 610893 73183
rect 610979 73145 610996 73183
rect 610996 73145 611035 73183
rect 611121 73145 611176 73183
rect 611176 73145 611177 73183
rect 611263 73145 611300 73183
rect 611300 73145 611319 73183
rect 611405 73145 611424 73183
rect 611424 73145 611461 73183
rect 611547 73145 611548 73183
rect 611548 73145 611603 73183
rect 611689 73145 611740 73183
rect 611740 73145 611745 73183
rect 611831 73145 611864 73183
rect 611864 73145 611887 73183
rect 611973 73145 611988 73183
rect 611988 73145 612029 73183
rect 612115 73145 612168 73183
rect 612168 73145 612171 73183
rect 610269 73127 610325 73145
rect 610411 73127 610467 73145
rect 610553 73127 610609 73145
rect 610695 73127 610751 73145
rect 610837 73127 610893 73145
rect 610979 73127 611035 73145
rect 611121 73127 611177 73145
rect 611263 73127 611319 73145
rect 611405 73127 611461 73145
rect 611547 73127 611603 73145
rect 611689 73127 611745 73145
rect 611831 73127 611887 73145
rect 611973 73127 612029 73145
rect 612115 73127 612171 73145
rect 610269 73021 610308 73041
rect 610308 73021 610325 73041
rect 610411 73021 610432 73041
rect 610432 73021 610467 73041
rect 610553 73021 610556 73041
rect 610556 73021 610609 73041
rect 610695 73021 610748 73041
rect 610748 73021 610751 73041
rect 610837 73021 610872 73041
rect 610872 73021 610893 73041
rect 610979 73021 610996 73041
rect 610996 73021 611035 73041
rect 611121 73021 611176 73041
rect 611176 73021 611177 73041
rect 611263 73021 611300 73041
rect 611300 73021 611319 73041
rect 611405 73021 611424 73041
rect 611424 73021 611461 73041
rect 611547 73021 611548 73041
rect 611548 73021 611603 73041
rect 611689 73021 611740 73041
rect 611740 73021 611745 73041
rect 611831 73021 611864 73041
rect 611864 73021 611887 73041
rect 611973 73021 611988 73041
rect 611988 73021 612029 73041
rect 612115 73021 612168 73041
rect 612168 73021 612171 73041
rect 610269 72985 610325 73021
rect 610411 72985 610467 73021
rect 610553 72985 610609 73021
rect 610695 72985 610751 73021
rect 610837 72985 610893 73021
rect 610979 72985 611035 73021
rect 611121 72985 611177 73021
rect 611263 72985 611319 73021
rect 611405 72985 611461 73021
rect 611547 72985 611603 73021
rect 611689 72985 611745 73021
rect 611831 72985 611887 73021
rect 611973 72985 612029 73021
rect 612115 72985 612171 73021
rect 610269 72897 610308 72899
rect 610308 72897 610325 72899
rect 610411 72897 610432 72899
rect 610432 72897 610467 72899
rect 610553 72897 610556 72899
rect 610556 72897 610609 72899
rect 610695 72897 610748 72899
rect 610748 72897 610751 72899
rect 610837 72897 610872 72899
rect 610872 72897 610893 72899
rect 610979 72897 610996 72899
rect 610996 72897 611035 72899
rect 611121 72897 611176 72899
rect 611176 72897 611177 72899
rect 611263 72897 611300 72899
rect 611300 72897 611319 72899
rect 611405 72897 611424 72899
rect 611424 72897 611461 72899
rect 611547 72897 611548 72899
rect 611548 72897 611603 72899
rect 611689 72897 611740 72899
rect 611740 72897 611745 72899
rect 611831 72897 611864 72899
rect 611864 72897 611887 72899
rect 611973 72897 611988 72899
rect 611988 72897 612029 72899
rect 612115 72897 612168 72899
rect 612168 72897 612171 72899
rect 610269 72843 610325 72897
rect 610411 72843 610467 72897
rect 610553 72843 610609 72897
rect 610695 72843 610751 72897
rect 610837 72843 610893 72897
rect 610979 72843 611035 72897
rect 611121 72843 611177 72897
rect 611263 72843 611319 72897
rect 611405 72843 611461 72897
rect 611547 72843 611603 72897
rect 611689 72843 611745 72897
rect 611831 72843 611887 72897
rect 611973 72843 612029 72897
rect 612115 72843 612171 72897
rect 610269 72705 610325 72757
rect 610411 72705 610467 72757
rect 610553 72705 610609 72757
rect 610695 72705 610751 72757
rect 610837 72705 610893 72757
rect 610979 72705 611035 72757
rect 611121 72705 611177 72757
rect 611263 72705 611319 72757
rect 611405 72705 611461 72757
rect 611547 72705 611603 72757
rect 611689 72705 611745 72757
rect 611831 72705 611887 72757
rect 611973 72705 612029 72757
rect 612115 72705 612171 72757
rect 610269 72701 610308 72705
rect 610308 72701 610325 72705
rect 610411 72701 610432 72705
rect 610432 72701 610467 72705
rect 610553 72701 610556 72705
rect 610556 72701 610609 72705
rect 610695 72701 610748 72705
rect 610748 72701 610751 72705
rect 610837 72701 610872 72705
rect 610872 72701 610893 72705
rect 610979 72701 610996 72705
rect 610996 72701 611035 72705
rect 611121 72701 611176 72705
rect 611176 72701 611177 72705
rect 611263 72701 611300 72705
rect 611300 72701 611319 72705
rect 611405 72701 611424 72705
rect 611424 72701 611461 72705
rect 611547 72701 611548 72705
rect 611548 72701 611603 72705
rect 611689 72701 611740 72705
rect 611740 72701 611745 72705
rect 611831 72701 611864 72705
rect 611864 72701 611887 72705
rect 611973 72701 611988 72705
rect 611988 72701 612029 72705
rect 612115 72701 612168 72705
rect 612168 72701 612171 72705
rect 610269 72581 610325 72615
rect 610411 72581 610467 72615
rect 610553 72581 610609 72615
rect 610695 72581 610751 72615
rect 610837 72581 610893 72615
rect 610979 72581 611035 72615
rect 611121 72581 611177 72615
rect 611263 72581 611319 72615
rect 611405 72581 611461 72615
rect 611547 72581 611603 72615
rect 611689 72581 611745 72615
rect 611831 72581 611887 72615
rect 611973 72581 612029 72615
rect 612115 72581 612171 72615
rect 610269 72559 610308 72581
rect 610308 72559 610325 72581
rect 610411 72559 610432 72581
rect 610432 72559 610467 72581
rect 610553 72559 610556 72581
rect 610556 72559 610609 72581
rect 610695 72559 610748 72581
rect 610748 72559 610751 72581
rect 610837 72559 610872 72581
rect 610872 72559 610893 72581
rect 610979 72559 610996 72581
rect 610996 72559 611035 72581
rect 611121 72559 611176 72581
rect 611176 72559 611177 72581
rect 611263 72559 611300 72581
rect 611300 72559 611319 72581
rect 611405 72559 611424 72581
rect 611424 72559 611461 72581
rect 611547 72559 611548 72581
rect 611548 72559 611603 72581
rect 611689 72559 611740 72581
rect 611740 72559 611745 72581
rect 611831 72559 611864 72581
rect 611864 72559 611887 72581
rect 611973 72559 611988 72581
rect 611988 72559 612029 72581
rect 612115 72559 612168 72581
rect 612168 72559 612171 72581
rect 610269 72457 610325 72473
rect 610411 72457 610467 72473
rect 610553 72457 610609 72473
rect 610695 72457 610751 72473
rect 610837 72457 610893 72473
rect 610979 72457 611035 72473
rect 611121 72457 611177 72473
rect 611263 72457 611319 72473
rect 611405 72457 611461 72473
rect 611547 72457 611603 72473
rect 611689 72457 611745 72473
rect 611831 72457 611887 72473
rect 611973 72457 612029 72473
rect 612115 72457 612171 72473
rect 610269 72417 610308 72457
rect 610308 72417 610325 72457
rect 610411 72417 610432 72457
rect 610432 72417 610467 72457
rect 610553 72417 610556 72457
rect 610556 72417 610609 72457
rect 610695 72417 610748 72457
rect 610748 72417 610751 72457
rect 610837 72417 610872 72457
rect 610872 72417 610893 72457
rect 610979 72417 610996 72457
rect 610996 72417 611035 72457
rect 611121 72417 611176 72457
rect 611176 72417 611177 72457
rect 611263 72417 611300 72457
rect 611300 72417 611319 72457
rect 611405 72417 611424 72457
rect 611424 72417 611461 72457
rect 611547 72417 611548 72457
rect 611548 72417 611603 72457
rect 611689 72417 611740 72457
rect 611740 72417 611745 72457
rect 611831 72417 611864 72457
rect 611864 72417 611887 72457
rect 611973 72417 611988 72457
rect 611988 72417 612029 72457
rect 612115 72417 612168 72457
rect 612168 72417 612171 72457
rect 610269 72277 610308 72331
rect 610308 72277 610325 72331
rect 610411 72277 610432 72331
rect 610432 72277 610467 72331
rect 610553 72277 610556 72331
rect 610556 72277 610609 72331
rect 610695 72277 610748 72331
rect 610748 72277 610751 72331
rect 610837 72277 610872 72331
rect 610872 72277 610893 72331
rect 610979 72277 610996 72331
rect 610996 72277 611035 72331
rect 611121 72277 611176 72331
rect 611176 72277 611177 72331
rect 611263 72277 611300 72331
rect 611300 72277 611319 72331
rect 611405 72277 611424 72331
rect 611424 72277 611461 72331
rect 611547 72277 611548 72331
rect 611548 72277 611603 72331
rect 611689 72277 611740 72331
rect 611740 72277 611745 72331
rect 611831 72277 611864 72331
rect 611864 72277 611887 72331
rect 611973 72277 611988 72331
rect 611988 72277 612029 72331
rect 612115 72277 612168 72331
rect 612168 72277 612171 72331
rect 610269 72275 610325 72277
rect 610411 72275 610467 72277
rect 610553 72275 610609 72277
rect 610695 72275 610751 72277
rect 610837 72275 610893 72277
rect 610979 72275 611035 72277
rect 611121 72275 611177 72277
rect 611263 72275 611319 72277
rect 611405 72275 611461 72277
rect 611547 72275 611603 72277
rect 611689 72275 611745 72277
rect 611831 72275 611887 72277
rect 611973 72275 612029 72277
rect 612115 72275 612171 72277
rect 610269 72153 610308 72189
rect 610308 72153 610325 72189
rect 610411 72153 610432 72189
rect 610432 72153 610467 72189
rect 610553 72153 610556 72189
rect 610556 72153 610609 72189
rect 610695 72153 610748 72189
rect 610748 72153 610751 72189
rect 610837 72153 610872 72189
rect 610872 72153 610893 72189
rect 610979 72153 610996 72189
rect 610996 72153 611035 72189
rect 611121 72153 611176 72189
rect 611176 72153 611177 72189
rect 611263 72153 611300 72189
rect 611300 72153 611319 72189
rect 611405 72153 611424 72189
rect 611424 72153 611461 72189
rect 611547 72153 611548 72189
rect 611548 72153 611603 72189
rect 611689 72153 611740 72189
rect 611740 72153 611745 72189
rect 611831 72153 611864 72189
rect 611864 72153 611887 72189
rect 611973 72153 611988 72189
rect 611988 72153 612029 72189
rect 612115 72153 612168 72189
rect 612168 72153 612171 72189
rect 610269 72133 610325 72153
rect 610411 72133 610467 72153
rect 610553 72133 610609 72153
rect 610695 72133 610751 72153
rect 610837 72133 610893 72153
rect 610979 72133 611035 72153
rect 611121 72133 611177 72153
rect 611263 72133 611319 72153
rect 611405 72133 611461 72153
rect 611547 72133 611603 72153
rect 611689 72133 611745 72153
rect 611831 72133 611887 72153
rect 611973 72133 612029 72153
rect 612115 72133 612171 72153
rect 612899 73979 612955 74035
rect 613041 73979 613097 74035
rect 613183 73979 613239 74035
rect 613325 73979 613381 74035
rect 613467 73979 613523 74035
rect 613609 73979 613665 74035
rect 613751 73979 613807 74035
rect 613893 73979 613949 74035
rect 614035 73979 614091 74035
rect 614177 73979 614233 74035
rect 614319 73979 614375 74035
rect 614461 73979 614517 74035
rect 614603 73979 614659 74035
rect 612899 73889 612938 73893
rect 612938 73889 612955 73893
rect 613041 73889 613062 73893
rect 613062 73889 613097 73893
rect 613183 73889 613186 73893
rect 613186 73889 613239 73893
rect 613325 73889 613378 73893
rect 613378 73889 613381 73893
rect 613467 73889 613502 73893
rect 613502 73889 613523 73893
rect 613609 73889 613626 73893
rect 613626 73889 613665 73893
rect 613751 73889 613806 73893
rect 613806 73889 613807 73893
rect 613893 73889 613930 73893
rect 613930 73889 613949 73893
rect 614035 73889 614054 73893
rect 614054 73889 614091 73893
rect 614177 73889 614178 73893
rect 614178 73889 614233 73893
rect 614319 73889 614370 73893
rect 614370 73889 614375 73893
rect 614461 73889 614494 73893
rect 614494 73889 614517 73893
rect 614603 73889 614618 73893
rect 614618 73889 614659 73893
rect 612899 73837 612955 73889
rect 613041 73837 613097 73889
rect 613183 73837 613239 73889
rect 613325 73837 613381 73889
rect 613467 73837 613523 73889
rect 613609 73837 613665 73889
rect 613751 73837 613807 73889
rect 613893 73837 613949 73889
rect 614035 73837 614091 73889
rect 614177 73837 614233 73889
rect 614319 73837 614375 73889
rect 614461 73837 614517 73889
rect 614603 73837 614659 73889
rect 612899 73697 612955 73751
rect 613041 73697 613097 73751
rect 613183 73697 613239 73751
rect 613325 73697 613381 73751
rect 613467 73697 613523 73751
rect 613609 73697 613665 73751
rect 613751 73697 613807 73751
rect 613893 73697 613949 73751
rect 614035 73697 614091 73751
rect 614177 73697 614233 73751
rect 614319 73697 614375 73751
rect 614461 73697 614517 73751
rect 614603 73697 614659 73751
rect 612899 73695 612938 73697
rect 612938 73695 612955 73697
rect 613041 73695 613062 73697
rect 613062 73695 613097 73697
rect 613183 73695 613186 73697
rect 613186 73695 613239 73697
rect 613325 73695 613378 73697
rect 613378 73695 613381 73697
rect 613467 73695 613502 73697
rect 613502 73695 613523 73697
rect 613609 73695 613626 73697
rect 613626 73695 613665 73697
rect 613751 73695 613806 73697
rect 613806 73695 613807 73697
rect 613893 73695 613930 73697
rect 613930 73695 613949 73697
rect 614035 73695 614054 73697
rect 614054 73695 614091 73697
rect 614177 73695 614178 73697
rect 614178 73695 614233 73697
rect 614319 73695 614370 73697
rect 614370 73695 614375 73697
rect 614461 73695 614494 73697
rect 614494 73695 614517 73697
rect 614603 73695 614618 73697
rect 614618 73695 614659 73697
rect 612899 73573 612955 73609
rect 613041 73573 613097 73609
rect 613183 73573 613239 73609
rect 613325 73573 613381 73609
rect 613467 73573 613523 73609
rect 613609 73573 613665 73609
rect 613751 73573 613807 73609
rect 613893 73573 613949 73609
rect 614035 73573 614091 73609
rect 614177 73573 614233 73609
rect 614319 73573 614375 73609
rect 614461 73573 614517 73609
rect 614603 73573 614659 73609
rect 612899 73553 612938 73573
rect 612938 73553 612955 73573
rect 613041 73553 613062 73573
rect 613062 73553 613097 73573
rect 613183 73553 613186 73573
rect 613186 73553 613239 73573
rect 613325 73553 613378 73573
rect 613378 73553 613381 73573
rect 613467 73553 613502 73573
rect 613502 73553 613523 73573
rect 613609 73553 613626 73573
rect 613626 73553 613665 73573
rect 613751 73553 613806 73573
rect 613806 73553 613807 73573
rect 613893 73553 613930 73573
rect 613930 73553 613949 73573
rect 614035 73553 614054 73573
rect 614054 73553 614091 73573
rect 614177 73553 614178 73573
rect 614178 73553 614233 73573
rect 614319 73553 614370 73573
rect 614370 73553 614375 73573
rect 614461 73553 614494 73573
rect 614494 73553 614517 73573
rect 614603 73553 614618 73573
rect 614618 73553 614659 73573
rect 612899 73449 612955 73467
rect 613041 73449 613097 73467
rect 613183 73449 613239 73467
rect 613325 73449 613381 73467
rect 613467 73449 613523 73467
rect 613609 73449 613665 73467
rect 613751 73449 613807 73467
rect 613893 73449 613949 73467
rect 614035 73449 614091 73467
rect 614177 73449 614233 73467
rect 614319 73449 614375 73467
rect 614461 73449 614517 73467
rect 614603 73449 614659 73467
rect 612899 73411 612938 73449
rect 612938 73411 612955 73449
rect 613041 73411 613062 73449
rect 613062 73411 613097 73449
rect 613183 73411 613186 73449
rect 613186 73411 613239 73449
rect 613325 73411 613378 73449
rect 613378 73411 613381 73449
rect 613467 73411 613502 73449
rect 613502 73411 613523 73449
rect 613609 73411 613626 73449
rect 613626 73411 613665 73449
rect 613751 73411 613806 73449
rect 613806 73411 613807 73449
rect 613893 73411 613930 73449
rect 613930 73411 613949 73449
rect 614035 73411 614054 73449
rect 614054 73411 614091 73449
rect 614177 73411 614178 73449
rect 614178 73411 614233 73449
rect 614319 73411 614370 73449
rect 614370 73411 614375 73449
rect 614461 73411 614494 73449
rect 614494 73411 614517 73449
rect 614603 73411 614618 73449
rect 614618 73411 614659 73449
rect 612899 73269 612938 73325
rect 612938 73269 612955 73325
rect 613041 73269 613062 73325
rect 613062 73269 613097 73325
rect 613183 73269 613186 73325
rect 613186 73269 613239 73325
rect 613325 73269 613378 73325
rect 613378 73269 613381 73325
rect 613467 73269 613502 73325
rect 613502 73269 613523 73325
rect 613609 73269 613626 73325
rect 613626 73269 613665 73325
rect 613751 73269 613806 73325
rect 613806 73269 613807 73325
rect 613893 73269 613930 73325
rect 613930 73269 613949 73325
rect 614035 73269 614054 73325
rect 614054 73269 614091 73325
rect 614177 73269 614178 73325
rect 614178 73269 614233 73325
rect 614319 73269 614370 73325
rect 614370 73269 614375 73325
rect 614461 73269 614494 73325
rect 614494 73269 614517 73325
rect 614603 73269 614618 73325
rect 614618 73269 614659 73325
rect 612899 73145 612938 73183
rect 612938 73145 612955 73183
rect 613041 73145 613062 73183
rect 613062 73145 613097 73183
rect 613183 73145 613186 73183
rect 613186 73145 613239 73183
rect 613325 73145 613378 73183
rect 613378 73145 613381 73183
rect 613467 73145 613502 73183
rect 613502 73145 613523 73183
rect 613609 73145 613626 73183
rect 613626 73145 613665 73183
rect 613751 73145 613806 73183
rect 613806 73145 613807 73183
rect 613893 73145 613930 73183
rect 613930 73145 613949 73183
rect 614035 73145 614054 73183
rect 614054 73145 614091 73183
rect 614177 73145 614178 73183
rect 614178 73145 614233 73183
rect 614319 73145 614370 73183
rect 614370 73145 614375 73183
rect 614461 73145 614494 73183
rect 614494 73145 614517 73183
rect 614603 73145 614618 73183
rect 614618 73145 614659 73183
rect 612899 73127 612955 73145
rect 613041 73127 613097 73145
rect 613183 73127 613239 73145
rect 613325 73127 613381 73145
rect 613467 73127 613523 73145
rect 613609 73127 613665 73145
rect 613751 73127 613807 73145
rect 613893 73127 613949 73145
rect 614035 73127 614091 73145
rect 614177 73127 614233 73145
rect 614319 73127 614375 73145
rect 614461 73127 614517 73145
rect 614603 73127 614659 73145
rect 612899 73021 612938 73041
rect 612938 73021 612955 73041
rect 613041 73021 613062 73041
rect 613062 73021 613097 73041
rect 613183 73021 613186 73041
rect 613186 73021 613239 73041
rect 613325 73021 613378 73041
rect 613378 73021 613381 73041
rect 613467 73021 613502 73041
rect 613502 73021 613523 73041
rect 613609 73021 613626 73041
rect 613626 73021 613665 73041
rect 613751 73021 613806 73041
rect 613806 73021 613807 73041
rect 613893 73021 613930 73041
rect 613930 73021 613949 73041
rect 614035 73021 614054 73041
rect 614054 73021 614091 73041
rect 614177 73021 614178 73041
rect 614178 73021 614233 73041
rect 614319 73021 614370 73041
rect 614370 73021 614375 73041
rect 614461 73021 614494 73041
rect 614494 73021 614517 73041
rect 614603 73021 614618 73041
rect 614618 73021 614659 73041
rect 612899 72985 612955 73021
rect 613041 72985 613097 73021
rect 613183 72985 613239 73021
rect 613325 72985 613381 73021
rect 613467 72985 613523 73021
rect 613609 72985 613665 73021
rect 613751 72985 613807 73021
rect 613893 72985 613949 73021
rect 614035 72985 614091 73021
rect 614177 72985 614233 73021
rect 614319 72985 614375 73021
rect 614461 72985 614517 73021
rect 614603 72985 614659 73021
rect 612899 72897 612938 72899
rect 612938 72897 612955 72899
rect 613041 72897 613062 72899
rect 613062 72897 613097 72899
rect 613183 72897 613186 72899
rect 613186 72897 613239 72899
rect 613325 72897 613378 72899
rect 613378 72897 613381 72899
rect 613467 72897 613502 72899
rect 613502 72897 613523 72899
rect 613609 72897 613626 72899
rect 613626 72897 613665 72899
rect 613751 72897 613806 72899
rect 613806 72897 613807 72899
rect 613893 72897 613930 72899
rect 613930 72897 613949 72899
rect 614035 72897 614054 72899
rect 614054 72897 614091 72899
rect 614177 72897 614178 72899
rect 614178 72897 614233 72899
rect 614319 72897 614370 72899
rect 614370 72897 614375 72899
rect 614461 72897 614494 72899
rect 614494 72897 614517 72899
rect 614603 72897 614618 72899
rect 614618 72897 614659 72899
rect 612899 72843 612955 72897
rect 613041 72843 613097 72897
rect 613183 72843 613239 72897
rect 613325 72843 613381 72897
rect 613467 72843 613523 72897
rect 613609 72843 613665 72897
rect 613751 72843 613807 72897
rect 613893 72843 613949 72897
rect 614035 72843 614091 72897
rect 614177 72843 614233 72897
rect 614319 72843 614375 72897
rect 614461 72843 614517 72897
rect 614603 72843 614659 72897
rect 612899 72705 612955 72757
rect 613041 72705 613097 72757
rect 613183 72705 613239 72757
rect 613325 72705 613381 72757
rect 613467 72705 613523 72757
rect 613609 72705 613665 72757
rect 613751 72705 613807 72757
rect 613893 72705 613949 72757
rect 614035 72705 614091 72757
rect 614177 72705 614233 72757
rect 614319 72705 614375 72757
rect 614461 72705 614517 72757
rect 614603 72705 614659 72757
rect 612899 72701 612938 72705
rect 612938 72701 612955 72705
rect 613041 72701 613062 72705
rect 613062 72701 613097 72705
rect 613183 72701 613186 72705
rect 613186 72701 613239 72705
rect 613325 72701 613378 72705
rect 613378 72701 613381 72705
rect 613467 72701 613502 72705
rect 613502 72701 613523 72705
rect 613609 72701 613626 72705
rect 613626 72701 613665 72705
rect 613751 72701 613806 72705
rect 613806 72701 613807 72705
rect 613893 72701 613930 72705
rect 613930 72701 613949 72705
rect 614035 72701 614054 72705
rect 614054 72701 614091 72705
rect 614177 72701 614178 72705
rect 614178 72701 614233 72705
rect 614319 72701 614370 72705
rect 614370 72701 614375 72705
rect 614461 72701 614494 72705
rect 614494 72701 614517 72705
rect 614603 72701 614618 72705
rect 614618 72701 614659 72705
rect 612899 72581 612955 72615
rect 613041 72581 613097 72615
rect 613183 72581 613239 72615
rect 613325 72581 613381 72615
rect 613467 72581 613523 72615
rect 613609 72581 613665 72615
rect 613751 72581 613807 72615
rect 613893 72581 613949 72615
rect 614035 72581 614091 72615
rect 614177 72581 614233 72615
rect 614319 72581 614375 72615
rect 614461 72581 614517 72615
rect 614603 72581 614659 72615
rect 612899 72559 612938 72581
rect 612938 72559 612955 72581
rect 613041 72559 613062 72581
rect 613062 72559 613097 72581
rect 613183 72559 613186 72581
rect 613186 72559 613239 72581
rect 613325 72559 613378 72581
rect 613378 72559 613381 72581
rect 613467 72559 613502 72581
rect 613502 72559 613523 72581
rect 613609 72559 613626 72581
rect 613626 72559 613665 72581
rect 613751 72559 613806 72581
rect 613806 72559 613807 72581
rect 613893 72559 613930 72581
rect 613930 72559 613949 72581
rect 614035 72559 614054 72581
rect 614054 72559 614091 72581
rect 614177 72559 614178 72581
rect 614178 72559 614233 72581
rect 614319 72559 614370 72581
rect 614370 72559 614375 72581
rect 614461 72559 614494 72581
rect 614494 72559 614517 72581
rect 614603 72559 614618 72581
rect 614618 72559 614659 72581
rect 612899 72457 612955 72473
rect 613041 72457 613097 72473
rect 613183 72457 613239 72473
rect 613325 72457 613381 72473
rect 613467 72457 613523 72473
rect 613609 72457 613665 72473
rect 613751 72457 613807 72473
rect 613893 72457 613949 72473
rect 614035 72457 614091 72473
rect 614177 72457 614233 72473
rect 614319 72457 614375 72473
rect 614461 72457 614517 72473
rect 614603 72457 614659 72473
rect 612899 72417 612938 72457
rect 612938 72417 612955 72457
rect 613041 72417 613062 72457
rect 613062 72417 613097 72457
rect 613183 72417 613186 72457
rect 613186 72417 613239 72457
rect 613325 72417 613378 72457
rect 613378 72417 613381 72457
rect 613467 72417 613502 72457
rect 613502 72417 613523 72457
rect 613609 72417 613626 72457
rect 613626 72417 613665 72457
rect 613751 72417 613806 72457
rect 613806 72417 613807 72457
rect 613893 72417 613930 72457
rect 613930 72417 613949 72457
rect 614035 72417 614054 72457
rect 614054 72417 614091 72457
rect 614177 72417 614178 72457
rect 614178 72417 614233 72457
rect 614319 72417 614370 72457
rect 614370 72417 614375 72457
rect 614461 72417 614494 72457
rect 614494 72417 614517 72457
rect 614603 72417 614618 72457
rect 614618 72417 614659 72457
rect 612899 72277 612938 72331
rect 612938 72277 612955 72331
rect 613041 72277 613062 72331
rect 613062 72277 613097 72331
rect 613183 72277 613186 72331
rect 613186 72277 613239 72331
rect 613325 72277 613378 72331
rect 613378 72277 613381 72331
rect 613467 72277 613502 72331
rect 613502 72277 613523 72331
rect 613609 72277 613626 72331
rect 613626 72277 613665 72331
rect 613751 72277 613806 72331
rect 613806 72277 613807 72331
rect 613893 72277 613930 72331
rect 613930 72277 613949 72331
rect 614035 72277 614054 72331
rect 614054 72277 614091 72331
rect 614177 72277 614178 72331
rect 614178 72277 614233 72331
rect 614319 72277 614370 72331
rect 614370 72277 614375 72331
rect 614461 72277 614494 72331
rect 614494 72277 614517 72331
rect 614603 72277 614618 72331
rect 614618 72277 614659 72331
rect 612899 72275 612955 72277
rect 613041 72275 613097 72277
rect 613183 72275 613239 72277
rect 613325 72275 613381 72277
rect 613467 72275 613523 72277
rect 613609 72275 613665 72277
rect 613751 72275 613807 72277
rect 613893 72275 613949 72277
rect 614035 72275 614091 72277
rect 614177 72275 614233 72277
rect 614319 72275 614375 72277
rect 614461 72275 614517 72277
rect 614603 72275 614659 72277
rect 612899 72153 612938 72189
rect 612938 72153 612955 72189
rect 613041 72153 613062 72189
rect 613062 72153 613097 72189
rect 613183 72153 613186 72189
rect 613186 72153 613239 72189
rect 613325 72153 613378 72189
rect 613378 72153 613381 72189
rect 613467 72153 613502 72189
rect 613502 72153 613523 72189
rect 613609 72153 613626 72189
rect 613626 72153 613665 72189
rect 613751 72153 613806 72189
rect 613806 72153 613807 72189
rect 613893 72153 613930 72189
rect 613930 72153 613949 72189
rect 614035 72153 614054 72189
rect 614054 72153 614091 72189
rect 614177 72153 614178 72189
rect 614178 72153 614233 72189
rect 614319 72153 614370 72189
rect 614370 72153 614375 72189
rect 614461 72153 614494 72189
rect 614494 72153 614517 72189
rect 614603 72153 614618 72189
rect 614618 72153 614659 72189
rect 612899 72133 612955 72153
rect 613041 72133 613097 72153
rect 613183 72133 613239 72153
rect 613325 72133 613381 72153
rect 613467 72133 613523 72153
rect 613609 72133 613665 72153
rect 613751 72133 613807 72153
rect 613893 72133 613949 72153
rect 614035 72133 614091 72153
rect 614177 72133 614233 72153
rect 614319 72133 614375 72153
rect 614461 72133 614517 72153
rect 614603 72133 614659 72153
<< metal4 >>
rect 379272 941675 380016 941720
rect 379272 941619 379341 941675
rect 379397 941619 379483 941675
rect 379539 941619 379625 941675
rect 379681 941619 379767 941675
rect 379823 941619 379909 941675
rect 379965 941619 380016 941675
rect 379272 941533 380016 941619
rect 379272 941477 379341 941533
rect 379397 941477 379483 941533
rect 379539 941477 379625 941533
rect 379681 941477 379767 941533
rect 379823 941477 379909 941533
rect 379965 941477 380016 941533
rect 379272 941391 380016 941477
rect 379272 941335 379341 941391
rect 379397 941335 379483 941391
rect 379539 941335 379625 941391
rect 379681 941335 379767 941391
rect 379823 941335 379909 941391
rect 379965 941335 380016 941391
rect 379272 941249 380016 941335
rect 379272 941193 379341 941249
rect 379397 941193 379483 941249
rect 379539 941193 379625 941249
rect 379681 941193 379767 941249
rect 379823 941193 379909 941249
rect 379965 941193 380016 941249
rect 379272 941107 380016 941193
rect 379272 941051 379341 941107
rect 379397 941051 379483 941107
rect 379539 941051 379625 941107
rect 379681 941051 379767 941107
rect 379823 941051 379909 941107
rect 379965 941051 380016 941107
rect 379272 940965 380016 941051
rect 379272 940909 379341 940965
rect 379397 940909 379483 940965
rect 379539 940909 379625 940965
rect 379681 940909 379767 940965
rect 379823 940909 379909 940965
rect 379965 940909 380016 940965
rect 379272 940823 380016 940909
rect 379272 940767 379341 940823
rect 379397 940767 379483 940823
rect 379539 940767 379625 940823
rect 379681 940767 379767 940823
rect 379823 940767 379909 940823
rect 379965 940767 380016 940823
rect 379272 940681 380016 940767
rect 379272 940625 379341 940681
rect 379397 940625 379483 940681
rect 379539 940625 379625 940681
rect 379681 940625 379767 940681
rect 379823 940625 379909 940681
rect 379965 940625 380016 940681
rect 379272 940539 380016 940625
rect 379272 940483 379341 940539
rect 379397 940483 379483 940539
rect 379539 940483 379625 940539
rect 379681 940483 379767 940539
rect 379823 940483 379909 940539
rect 379965 940483 380016 940539
rect 379272 940397 380016 940483
rect 379272 940341 379341 940397
rect 379397 940341 379483 940397
rect 379539 940341 379625 940397
rect 379681 940341 379767 940397
rect 379823 940341 379909 940397
rect 379965 940341 380016 940397
rect 379272 940255 380016 940341
rect 379272 940199 379341 940255
rect 379397 940199 379483 940255
rect 379539 940199 379625 940255
rect 379681 940199 379767 940255
rect 379823 940199 379909 940255
rect 379965 940199 380016 940255
rect 379272 940113 380016 940199
rect 379272 940057 379341 940113
rect 379397 940057 379483 940113
rect 379539 940057 379625 940113
rect 379681 940057 379767 940113
rect 379823 940057 379909 940113
rect 379965 940057 380016 940113
rect 379272 939971 380016 940057
rect 379272 939915 379341 939971
rect 379397 939915 379483 939971
rect 379539 939915 379625 939971
rect 379681 939915 379767 939971
rect 379823 939915 379909 939971
rect 379965 939915 380016 939971
rect 379272 939829 380016 939915
rect 379272 939773 379341 939829
rect 379397 939773 379483 939829
rect 379539 939773 379625 939829
rect 379681 939773 379767 939829
rect 379823 939773 379909 939829
rect 379965 939773 380016 939829
rect 379272 939720 380016 939773
rect 381752 941675 383802 941720
rect 381752 941619 381829 941675
rect 381885 941619 381971 941675
rect 382027 941619 382113 941675
rect 382169 941619 382255 941675
rect 382311 941619 382397 941675
rect 382453 941619 382539 941675
rect 382595 941619 382681 941675
rect 382737 941619 382823 941675
rect 382879 941619 382965 941675
rect 383021 941619 383107 941675
rect 383163 941619 383249 941675
rect 383305 941619 383391 941675
rect 383447 941619 383533 941675
rect 383589 941619 383675 941675
rect 383731 941619 383802 941675
rect 381752 941533 383802 941619
rect 381752 941477 381829 941533
rect 381885 941477 381971 941533
rect 382027 941477 382113 941533
rect 382169 941477 382255 941533
rect 382311 941477 382397 941533
rect 382453 941477 382539 941533
rect 382595 941477 382681 941533
rect 382737 941477 382823 941533
rect 382879 941477 382965 941533
rect 383021 941477 383107 941533
rect 383163 941477 383249 941533
rect 383305 941477 383391 941533
rect 383447 941477 383533 941533
rect 383589 941477 383675 941533
rect 383731 941477 383802 941533
rect 381752 941391 383802 941477
rect 381752 941335 381829 941391
rect 381885 941335 381971 941391
rect 382027 941335 382113 941391
rect 382169 941335 382255 941391
rect 382311 941335 382397 941391
rect 382453 941335 382539 941391
rect 382595 941335 382681 941391
rect 382737 941335 382823 941391
rect 382879 941335 382965 941391
rect 383021 941335 383107 941391
rect 383163 941335 383249 941391
rect 383305 941335 383391 941391
rect 383447 941335 383533 941391
rect 383589 941335 383675 941391
rect 383731 941335 383802 941391
rect 381752 941249 383802 941335
rect 381752 941193 381829 941249
rect 381885 941193 381971 941249
rect 382027 941193 382113 941249
rect 382169 941193 382255 941249
rect 382311 941193 382397 941249
rect 382453 941193 382539 941249
rect 382595 941193 382681 941249
rect 382737 941193 382823 941249
rect 382879 941193 382965 941249
rect 383021 941193 383107 941249
rect 383163 941193 383249 941249
rect 383305 941193 383391 941249
rect 383447 941193 383533 941249
rect 383589 941193 383675 941249
rect 383731 941193 383802 941249
rect 381752 941107 383802 941193
rect 381752 941051 381829 941107
rect 381885 941051 381971 941107
rect 382027 941051 382113 941107
rect 382169 941051 382255 941107
rect 382311 941051 382397 941107
rect 382453 941051 382539 941107
rect 382595 941051 382681 941107
rect 382737 941051 382823 941107
rect 382879 941051 382965 941107
rect 383021 941051 383107 941107
rect 383163 941051 383249 941107
rect 383305 941051 383391 941107
rect 383447 941051 383533 941107
rect 383589 941051 383675 941107
rect 383731 941051 383802 941107
rect 381752 940965 383802 941051
rect 381752 940909 381829 940965
rect 381885 940909 381971 940965
rect 382027 940909 382113 940965
rect 382169 940909 382255 940965
rect 382311 940909 382397 940965
rect 382453 940909 382539 940965
rect 382595 940909 382681 940965
rect 382737 940909 382823 940965
rect 382879 940909 382965 940965
rect 383021 940909 383107 940965
rect 383163 940909 383249 940965
rect 383305 940909 383391 940965
rect 383447 940909 383533 940965
rect 383589 940909 383675 940965
rect 383731 940909 383802 940965
rect 381752 940823 383802 940909
rect 381752 940767 381829 940823
rect 381885 940767 381971 940823
rect 382027 940767 382113 940823
rect 382169 940767 382255 940823
rect 382311 940767 382397 940823
rect 382453 940767 382539 940823
rect 382595 940767 382681 940823
rect 382737 940767 382823 940823
rect 382879 940767 382965 940823
rect 383021 940767 383107 940823
rect 383163 940767 383249 940823
rect 383305 940767 383391 940823
rect 383447 940767 383533 940823
rect 383589 940767 383675 940823
rect 383731 940767 383802 940823
rect 381752 940681 383802 940767
rect 381752 940625 381829 940681
rect 381885 940625 381971 940681
rect 382027 940625 382113 940681
rect 382169 940625 382255 940681
rect 382311 940625 382397 940681
rect 382453 940625 382539 940681
rect 382595 940625 382681 940681
rect 382737 940625 382823 940681
rect 382879 940625 382965 940681
rect 383021 940625 383107 940681
rect 383163 940625 383249 940681
rect 383305 940625 383391 940681
rect 383447 940625 383533 940681
rect 383589 940625 383675 940681
rect 383731 940625 383802 940681
rect 381752 940539 383802 940625
rect 381752 940483 381829 940539
rect 381885 940483 381971 940539
rect 382027 940483 382113 940539
rect 382169 940483 382255 940539
rect 382311 940483 382397 940539
rect 382453 940483 382539 940539
rect 382595 940483 382681 940539
rect 382737 940483 382823 940539
rect 382879 940483 382965 940539
rect 383021 940483 383107 940539
rect 383163 940483 383249 940539
rect 383305 940483 383391 940539
rect 383447 940483 383533 940539
rect 383589 940483 383675 940539
rect 383731 940483 383802 940539
rect 381752 940397 383802 940483
rect 381752 940341 381829 940397
rect 381885 940341 381971 940397
rect 382027 940341 382113 940397
rect 382169 940341 382255 940397
rect 382311 940341 382397 940397
rect 382453 940341 382539 940397
rect 382595 940341 382681 940397
rect 382737 940341 382823 940397
rect 382879 940341 382965 940397
rect 383021 940341 383107 940397
rect 383163 940341 383249 940397
rect 383305 940341 383391 940397
rect 383447 940341 383533 940397
rect 383589 940341 383675 940397
rect 383731 940341 383802 940397
rect 381752 940255 383802 940341
rect 381752 940199 381829 940255
rect 381885 940199 381971 940255
rect 382027 940199 382113 940255
rect 382169 940199 382255 940255
rect 382311 940199 382397 940255
rect 382453 940199 382539 940255
rect 382595 940199 382681 940255
rect 382737 940199 382823 940255
rect 382879 940199 382965 940255
rect 383021 940199 383107 940255
rect 383163 940199 383249 940255
rect 383305 940199 383391 940255
rect 383447 940199 383533 940255
rect 383589 940199 383675 940255
rect 383731 940199 383802 940255
rect 381752 940113 383802 940199
rect 381752 940057 381829 940113
rect 381885 940057 381971 940113
rect 382027 940057 382113 940113
rect 382169 940057 382255 940113
rect 382311 940057 382397 940113
rect 382453 940057 382539 940113
rect 382595 940057 382681 940113
rect 382737 940057 382823 940113
rect 382879 940057 382965 940113
rect 383021 940057 383107 940113
rect 383163 940057 383249 940113
rect 383305 940057 383391 940113
rect 383447 940057 383533 940113
rect 383589 940057 383675 940113
rect 383731 940057 383802 940113
rect 381752 939971 383802 940057
rect 381752 939915 381829 939971
rect 381885 939915 381971 939971
rect 382027 939915 382113 939971
rect 382169 939915 382255 939971
rect 382311 939915 382397 939971
rect 382453 939915 382539 939971
rect 382595 939915 382681 939971
rect 382737 939915 382823 939971
rect 382879 939915 382965 939971
rect 383021 939915 383107 939971
rect 383163 939915 383249 939971
rect 383305 939915 383391 939971
rect 383447 939915 383533 939971
rect 383589 939915 383675 939971
rect 383731 939915 383802 939971
rect 381752 939829 383802 939915
rect 381752 939773 381829 939829
rect 381885 939773 381971 939829
rect 382027 939773 382113 939829
rect 382169 939773 382255 939829
rect 382311 939773 382397 939829
rect 382453 939773 382539 939829
rect 382595 939773 382681 939829
rect 382737 939773 382823 939829
rect 382879 939773 382965 939829
rect 383021 939773 383107 939829
rect 383163 939773 383249 939829
rect 383305 939773 383391 939829
rect 383447 939773 383533 939829
rect 383589 939773 383675 939829
rect 383731 939773 383802 939829
rect 381752 939720 383802 939773
rect 384122 941675 386172 941720
rect 384122 941619 384199 941675
rect 384255 941619 384341 941675
rect 384397 941619 384483 941675
rect 384539 941619 384625 941675
rect 384681 941619 384767 941675
rect 384823 941619 384909 941675
rect 384965 941619 385051 941675
rect 385107 941619 385193 941675
rect 385249 941619 385335 941675
rect 385391 941619 385477 941675
rect 385533 941619 385619 941675
rect 385675 941619 385761 941675
rect 385817 941619 385903 941675
rect 385959 941619 386045 941675
rect 386101 941619 386172 941675
rect 384122 941533 386172 941619
rect 384122 941477 384199 941533
rect 384255 941477 384341 941533
rect 384397 941477 384483 941533
rect 384539 941477 384625 941533
rect 384681 941477 384767 941533
rect 384823 941477 384909 941533
rect 384965 941477 385051 941533
rect 385107 941477 385193 941533
rect 385249 941477 385335 941533
rect 385391 941477 385477 941533
rect 385533 941477 385619 941533
rect 385675 941477 385761 941533
rect 385817 941477 385903 941533
rect 385959 941477 386045 941533
rect 386101 941477 386172 941533
rect 384122 941391 386172 941477
rect 384122 941335 384199 941391
rect 384255 941335 384341 941391
rect 384397 941335 384483 941391
rect 384539 941335 384625 941391
rect 384681 941335 384767 941391
rect 384823 941335 384909 941391
rect 384965 941335 385051 941391
rect 385107 941335 385193 941391
rect 385249 941335 385335 941391
rect 385391 941335 385477 941391
rect 385533 941335 385619 941391
rect 385675 941335 385761 941391
rect 385817 941335 385903 941391
rect 385959 941335 386045 941391
rect 386101 941335 386172 941391
rect 384122 941249 386172 941335
rect 384122 941193 384199 941249
rect 384255 941193 384341 941249
rect 384397 941193 384483 941249
rect 384539 941193 384625 941249
rect 384681 941193 384767 941249
rect 384823 941193 384909 941249
rect 384965 941193 385051 941249
rect 385107 941193 385193 941249
rect 385249 941193 385335 941249
rect 385391 941193 385477 941249
rect 385533 941193 385619 941249
rect 385675 941193 385761 941249
rect 385817 941193 385903 941249
rect 385959 941193 386045 941249
rect 386101 941193 386172 941249
rect 384122 941107 386172 941193
rect 384122 941051 384199 941107
rect 384255 941051 384341 941107
rect 384397 941051 384483 941107
rect 384539 941051 384625 941107
rect 384681 941051 384767 941107
rect 384823 941051 384909 941107
rect 384965 941051 385051 941107
rect 385107 941051 385193 941107
rect 385249 941051 385335 941107
rect 385391 941051 385477 941107
rect 385533 941051 385619 941107
rect 385675 941051 385761 941107
rect 385817 941051 385903 941107
rect 385959 941051 386045 941107
rect 386101 941051 386172 941107
rect 384122 940965 386172 941051
rect 384122 940909 384199 940965
rect 384255 940909 384341 940965
rect 384397 940909 384483 940965
rect 384539 940909 384625 940965
rect 384681 940909 384767 940965
rect 384823 940909 384909 940965
rect 384965 940909 385051 940965
rect 385107 940909 385193 940965
rect 385249 940909 385335 940965
rect 385391 940909 385477 940965
rect 385533 940909 385619 940965
rect 385675 940909 385761 940965
rect 385817 940909 385903 940965
rect 385959 940909 386045 940965
rect 386101 940909 386172 940965
rect 384122 940823 386172 940909
rect 384122 940767 384199 940823
rect 384255 940767 384341 940823
rect 384397 940767 384483 940823
rect 384539 940767 384625 940823
rect 384681 940767 384767 940823
rect 384823 940767 384909 940823
rect 384965 940767 385051 940823
rect 385107 940767 385193 940823
rect 385249 940767 385335 940823
rect 385391 940767 385477 940823
rect 385533 940767 385619 940823
rect 385675 940767 385761 940823
rect 385817 940767 385903 940823
rect 385959 940767 386045 940823
rect 386101 940767 386172 940823
rect 384122 940681 386172 940767
rect 384122 940625 384199 940681
rect 384255 940625 384341 940681
rect 384397 940625 384483 940681
rect 384539 940625 384625 940681
rect 384681 940625 384767 940681
rect 384823 940625 384909 940681
rect 384965 940625 385051 940681
rect 385107 940625 385193 940681
rect 385249 940625 385335 940681
rect 385391 940625 385477 940681
rect 385533 940625 385619 940681
rect 385675 940625 385761 940681
rect 385817 940625 385903 940681
rect 385959 940625 386045 940681
rect 386101 940625 386172 940681
rect 384122 940539 386172 940625
rect 384122 940483 384199 940539
rect 384255 940483 384341 940539
rect 384397 940483 384483 940539
rect 384539 940483 384625 940539
rect 384681 940483 384767 940539
rect 384823 940483 384909 940539
rect 384965 940483 385051 940539
rect 385107 940483 385193 940539
rect 385249 940483 385335 940539
rect 385391 940483 385477 940539
rect 385533 940483 385619 940539
rect 385675 940483 385761 940539
rect 385817 940483 385903 940539
rect 385959 940483 386045 940539
rect 386101 940483 386172 940539
rect 384122 940397 386172 940483
rect 384122 940341 384199 940397
rect 384255 940341 384341 940397
rect 384397 940341 384483 940397
rect 384539 940341 384625 940397
rect 384681 940341 384767 940397
rect 384823 940341 384909 940397
rect 384965 940341 385051 940397
rect 385107 940341 385193 940397
rect 385249 940341 385335 940397
rect 385391 940341 385477 940397
rect 385533 940341 385619 940397
rect 385675 940341 385761 940397
rect 385817 940341 385903 940397
rect 385959 940341 386045 940397
rect 386101 940341 386172 940397
rect 384122 940255 386172 940341
rect 384122 940199 384199 940255
rect 384255 940199 384341 940255
rect 384397 940199 384483 940255
rect 384539 940199 384625 940255
rect 384681 940199 384767 940255
rect 384823 940199 384909 940255
rect 384965 940199 385051 940255
rect 385107 940199 385193 940255
rect 385249 940199 385335 940255
rect 385391 940199 385477 940255
rect 385533 940199 385619 940255
rect 385675 940199 385761 940255
rect 385817 940199 385903 940255
rect 385959 940199 386045 940255
rect 386101 940199 386172 940255
rect 384122 940113 386172 940199
rect 384122 940057 384199 940113
rect 384255 940057 384341 940113
rect 384397 940057 384483 940113
rect 384539 940057 384625 940113
rect 384681 940057 384767 940113
rect 384823 940057 384909 940113
rect 384965 940057 385051 940113
rect 385107 940057 385193 940113
rect 385249 940057 385335 940113
rect 385391 940057 385477 940113
rect 385533 940057 385619 940113
rect 385675 940057 385761 940113
rect 385817 940057 385903 940113
rect 385959 940057 386045 940113
rect 386101 940057 386172 940113
rect 384122 939971 386172 940057
rect 384122 939915 384199 939971
rect 384255 939915 384341 939971
rect 384397 939915 384483 939971
rect 384539 939915 384625 939971
rect 384681 939915 384767 939971
rect 384823 939915 384909 939971
rect 384965 939915 385051 939971
rect 385107 939915 385193 939971
rect 385249 939915 385335 939971
rect 385391 939915 385477 939971
rect 385533 939915 385619 939971
rect 385675 939915 385761 939971
rect 385817 939915 385903 939971
rect 385959 939915 386045 939971
rect 386101 939915 386172 939971
rect 384122 939829 386172 939915
rect 384122 939773 384199 939829
rect 384255 939773 384341 939829
rect 384397 939773 384483 939829
rect 384539 939773 384625 939829
rect 384681 939773 384767 939829
rect 384823 939773 384909 939829
rect 384965 939773 385051 939829
rect 385107 939773 385193 939829
rect 385249 939773 385335 939829
rect 385391 939773 385477 939829
rect 385533 939773 385619 939829
rect 385675 939773 385761 939829
rect 385817 939773 385903 939829
rect 385959 939773 386045 939829
rect 386101 939773 386172 939829
rect 384122 939720 386172 939773
rect 386828 941675 388878 941720
rect 386828 941619 386905 941675
rect 386961 941619 387047 941675
rect 387103 941619 387189 941675
rect 387245 941619 387331 941675
rect 387387 941619 387473 941675
rect 387529 941619 387615 941675
rect 387671 941619 387757 941675
rect 387813 941619 387899 941675
rect 387955 941619 388041 941675
rect 388097 941619 388183 941675
rect 388239 941619 388325 941675
rect 388381 941619 388467 941675
rect 388523 941619 388609 941675
rect 388665 941619 388751 941675
rect 388807 941619 388878 941675
rect 386828 941533 388878 941619
rect 386828 941477 386905 941533
rect 386961 941477 387047 941533
rect 387103 941477 387189 941533
rect 387245 941477 387331 941533
rect 387387 941477 387473 941533
rect 387529 941477 387615 941533
rect 387671 941477 387757 941533
rect 387813 941477 387899 941533
rect 387955 941477 388041 941533
rect 388097 941477 388183 941533
rect 388239 941477 388325 941533
rect 388381 941477 388467 941533
rect 388523 941477 388609 941533
rect 388665 941477 388751 941533
rect 388807 941477 388878 941533
rect 386828 941391 388878 941477
rect 386828 941335 386905 941391
rect 386961 941335 387047 941391
rect 387103 941335 387189 941391
rect 387245 941335 387331 941391
rect 387387 941335 387473 941391
rect 387529 941335 387615 941391
rect 387671 941335 387757 941391
rect 387813 941335 387899 941391
rect 387955 941335 388041 941391
rect 388097 941335 388183 941391
rect 388239 941335 388325 941391
rect 388381 941335 388467 941391
rect 388523 941335 388609 941391
rect 388665 941335 388751 941391
rect 388807 941335 388878 941391
rect 386828 941249 388878 941335
rect 386828 941193 386905 941249
rect 386961 941193 387047 941249
rect 387103 941193 387189 941249
rect 387245 941193 387331 941249
rect 387387 941193 387473 941249
rect 387529 941193 387615 941249
rect 387671 941193 387757 941249
rect 387813 941193 387899 941249
rect 387955 941193 388041 941249
rect 388097 941193 388183 941249
rect 388239 941193 388325 941249
rect 388381 941193 388467 941249
rect 388523 941193 388609 941249
rect 388665 941193 388751 941249
rect 388807 941193 388878 941249
rect 386828 941107 388878 941193
rect 386828 941051 386905 941107
rect 386961 941051 387047 941107
rect 387103 941051 387189 941107
rect 387245 941051 387331 941107
rect 387387 941051 387473 941107
rect 387529 941051 387615 941107
rect 387671 941051 387757 941107
rect 387813 941051 387899 941107
rect 387955 941051 388041 941107
rect 388097 941051 388183 941107
rect 388239 941051 388325 941107
rect 388381 941051 388467 941107
rect 388523 941051 388609 941107
rect 388665 941051 388751 941107
rect 388807 941051 388878 941107
rect 386828 940965 388878 941051
rect 386828 940909 386905 940965
rect 386961 940909 387047 940965
rect 387103 940909 387189 940965
rect 387245 940909 387331 940965
rect 387387 940909 387473 940965
rect 387529 940909 387615 940965
rect 387671 940909 387757 940965
rect 387813 940909 387899 940965
rect 387955 940909 388041 940965
rect 388097 940909 388183 940965
rect 388239 940909 388325 940965
rect 388381 940909 388467 940965
rect 388523 940909 388609 940965
rect 388665 940909 388751 940965
rect 388807 940909 388878 940965
rect 386828 940823 388878 940909
rect 386828 940767 386905 940823
rect 386961 940767 387047 940823
rect 387103 940767 387189 940823
rect 387245 940767 387331 940823
rect 387387 940767 387473 940823
rect 387529 940767 387615 940823
rect 387671 940767 387757 940823
rect 387813 940767 387899 940823
rect 387955 940767 388041 940823
rect 388097 940767 388183 940823
rect 388239 940767 388325 940823
rect 388381 940767 388467 940823
rect 388523 940767 388609 940823
rect 388665 940767 388751 940823
rect 388807 940767 388878 940823
rect 386828 940681 388878 940767
rect 386828 940625 386905 940681
rect 386961 940625 387047 940681
rect 387103 940625 387189 940681
rect 387245 940625 387331 940681
rect 387387 940625 387473 940681
rect 387529 940625 387615 940681
rect 387671 940625 387757 940681
rect 387813 940625 387899 940681
rect 387955 940625 388041 940681
rect 388097 940625 388183 940681
rect 388239 940625 388325 940681
rect 388381 940625 388467 940681
rect 388523 940625 388609 940681
rect 388665 940625 388751 940681
rect 388807 940625 388878 940681
rect 386828 940539 388878 940625
rect 386828 940483 386905 940539
rect 386961 940483 387047 940539
rect 387103 940483 387189 940539
rect 387245 940483 387331 940539
rect 387387 940483 387473 940539
rect 387529 940483 387615 940539
rect 387671 940483 387757 940539
rect 387813 940483 387899 940539
rect 387955 940483 388041 940539
rect 388097 940483 388183 940539
rect 388239 940483 388325 940539
rect 388381 940483 388467 940539
rect 388523 940483 388609 940539
rect 388665 940483 388751 940539
rect 388807 940483 388878 940539
rect 386828 940397 388878 940483
rect 386828 940341 386905 940397
rect 386961 940341 387047 940397
rect 387103 940341 387189 940397
rect 387245 940341 387331 940397
rect 387387 940341 387473 940397
rect 387529 940341 387615 940397
rect 387671 940341 387757 940397
rect 387813 940341 387899 940397
rect 387955 940341 388041 940397
rect 388097 940341 388183 940397
rect 388239 940341 388325 940397
rect 388381 940341 388467 940397
rect 388523 940341 388609 940397
rect 388665 940341 388751 940397
rect 388807 940341 388878 940397
rect 386828 940255 388878 940341
rect 386828 940199 386905 940255
rect 386961 940199 387047 940255
rect 387103 940199 387189 940255
rect 387245 940199 387331 940255
rect 387387 940199 387473 940255
rect 387529 940199 387615 940255
rect 387671 940199 387757 940255
rect 387813 940199 387899 940255
rect 387955 940199 388041 940255
rect 388097 940199 388183 940255
rect 388239 940199 388325 940255
rect 388381 940199 388467 940255
rect 388523 940199 388609 940255
rect 388665 940199 388751 940255
rect 388807 940199 388878 940255
rect 386828 940113 388878 940199
rect 386828 940057 386905 940113
rect 386961 940057 387047 940113
rect 387103 940057 387189 940113
rect 387245 940057 387331 940113
rect 387387 940057 387473 940113
rect 387529 940057 387615 940113
rect 387671 940057 387757 940113
rect 387813 940057 387899 940113
rect 387955 940057 388041 940113
rect 388097 940057 388183 940113
rect 388239 940057 388325 940113
rect 388381 940057 388467 940113
rect 388523 940057 388609 940113
rect 388665 940057 388751 940113
rect 388807 940057 388878 940113
rect 386828 939971 388878 940057
rect 386828 939915 386905 939971
rect 386961 939915 387047 939971
rect 387103 939915 387189 939971
rect 387245 939915 387331 939971
rect 387387 939915 387473 939971
rect 387529 939915 387615 939971
rect 387671 939915 387757 939971
rect 387813 939915 387899 939971
rect 387955 939915 388041 939971
rect 388097 939915 388183 939971
rect 388239 939915 388325 939971
rect 388381 939915 388467 939971
rect 388523 939915 388609 939971
rect 388665 939915 388751 939971
rect 388807 939915 388878 939971
rect 386828 939829 388878 939915
rect 386828 939773 386905 939829
rect 386961 939773 387047 939829
rect 387103 939773 387189 939829
rect 387245 939773 387331 939829
rect 387387 939773 387473 939829
rect 387529 939773 387615 939829
rect 387671 939773 387757 939829
rect 387813 939773 387899 939829
rect 387955 939773 388041 939829
rect 388097 939773 388183 939829
rect 388239 939773 388325 939829
rect 388381 939773 388467 939829
rect 388523 939773 388609 939829
rect 388665 939773 388751 939829
rect 388807 939773 388878 939829
rect 386828 939720 388878 939773
rect 389198 941675 391248 941720
rect 389198 941619 389275 941675
rect 389331 941619 389417 941675
rect 389473 941619 389559 941675
rect 389615 941619 389701 941675
rect 389757 941619 389843 941675
rect 389899 941619 389985 941675
rect 390041 941619 390127 941675
rect 390183 941619 390269 941675
rect 390325 941619 390411 941675
rect 390467 941619 390553 941675
rect 390609 941619 390695 941675
rect 390751 941619 390837 941675
rect 390893 941619 390979 941675
rect 391035 941619 391121 941675
rect 391177 941619 391248 941675
rect 389198 941533 391248 941619
rect 389198 941477 389275 941533
rect 389331 941477 389417 941533
rect 389473 941477 389559 941533
rect 389615 941477 389701 941533
rect 389757 941477 389843 941533
rect 389899 941477 389985 941533
rect 390041 941477 390127 941533
rect 390183 941477 390269 941533
rect 390325 941477 390411 941533
rect 390467 941477 390553 941533
rect 390609 941477 390695 941533
rect 390751 941477 390837 941533
rect 390893 941477 390979 941533
rect 391035 941477 391121 941533
rect 391177 941477 391248 941533
rect 389198 941391 391248 941477
rect 389198 941335 389275 941391
rect 389331 941335 389417 941391
rect 389473 941335 389559 941391
rect 389615 941335 389701 941391
rect 389757 941335 389843 941391
rect 389899 941335 389985 941391
rect 390041 941335 390127 941391
rect 390183 941335 390269 941391
rect 390325 941335 390411 941391
rect 390467 941335 390553 941391
rect 390609 941335 390695 941391
rect 390751 941335 390837 941391
rect 390893 941335 390979 941391
rect 391035 941335 391121 941391
rect 391177 941335 391248 941391
rect 389198 941249 391248 941335
rect 389198 941193 389275 941249
rect 389331 941193 389417 941249
rect 389473 941193 389559 941249
rect 389615 941193 389701 941249
rect 389757 941193 389843 941249
rect 389899 941193 389985 941249
rect 390041 941193 390127 941249
rect 390183 941193 390269 941249
rect 390325 941193 390411 941249
rect 390467 941193 390553 941249
rect 390609 941193 390695 941249
rect 390751 941193 390837 941249
rect 390893 941193 390979 941249
rect 391035 941193 391121 941249
rect 391177 941193 391248 941249
rect 389198 941107 391248 941193
rect 389198 941051 389275 941107
rect 389331 941051 389417 941107
rect 389473 941051 389559 941107
rect 389615 941051 389701 941107
rect 389757 941051 389843 941107
rect 389899 941051 389985 941107
rect 390041 941051 390127 941107
rect 390183 941051 390269 941107
rect 390325 941051 390411 941107
rect 390467 941051 390553 941107
rect 390609 941051 390695 941107
rect 390751 941051 390837 941107
rect 390893 941051 390979 941107
rect 391035 941051 391121 941107
rect 391177 941051 391248 941107
rect 389198 940965 391248 941051
rect 389198 940909 389275 940965
rect 389331 940909 389417 940965
rect 389473 940909 389559 940965
rect 389615 940909 389701 940965
rect 389757 940909 389843 940965
rect 389899 940909 389985 940965
rect 390041 940909 390127 940965
rect 390183 940909 390269 940965
rect 390325 940909 390411 940965
rect 390467 940909 390553 940965
rect 390609 940909 390695 940965
rect 390751 940909 390837 940965
rect 390893 940909 390979 940965
rect 391035 940909 391121 940965
rect 391177 940909 391248 940965
rect 389198 940823 391248 940909
rect 389198 940767 389275 940823
rect 389331 940767 389417 940823
rect 389473 940767 389559 940823
rect 389615 940767 389701 940823
rect 389757 940767 389843 940823
rect 389899 940767 389985 940823
rect 390041 940767 390127 940823
rect 390183 940767 390269 940823
rect 390325 940767 390411 940823
rect 390467 940767 390553 940823
rect 390609 940767 390695 940823
rect 390751 940767 390837 940823
rect 390893 940767 390979 940823
rect 391035 940767 391121 940823
rect 391177 940767 391248 940823
rect 389198 940681 391248 940767
rect 389198 940625 389275 940681
rect 389331 940625 389417 940681
rect 389473 940625 389559 940681
rect 389615 940625 389701 940681
rect 389757 940625 389843 940681
rect 389899 940625 389985 940681
rect 390041 940625 390127 940681
rect 390183 940625 390269 940681
rect 390325 940625 390411 940681
rect 390467 940625 390553 940681
rect 390609 940625 390695 940681
rect 390751 940625 390837 940681
rect 390893 940625 390979 940681
rect 391035 940625 391121 940681
rect 391177 940625 391248 940681
rect 389198 940539 391248 940625
rect 389198 940483 389275 940539
rect 389331 940483 389417 940539
rect 389473 940483 389559 940539
rect 389615 940483 389701 940539
rect 389757 940483 389843 940539
rect 389899 940483 389985 940539
rect 390041 940483 390127 940539
rect 390183 940483 390269 940539
rect 390325 940483 390411 940539
rect 390467 940483 390553 940539
rect 390609 940483 390695 940539
rect 390751 940483 390837 940539
rect 390893 940483 390979 940539
rect 391035 940483 391121 940539
rect 391177 940483 391248 940539
rect 389198 940397 391248 940483
rect 389198 940341 389275 940397
rect 389331 940341 389417 940397
rect 389473 940341 389559 940397
rect 389615 940341 389701 940397
rect 389757 940341 389843 940397
rect 389899 940341 389985 940397
rect 390041 940341 390127 940397
rect 390183 940341 390269 940397
rect 390325 940341 390411 940397
rect 390467 940341 390553 940397
rect 390609 940341 390695 940397
rect 390751 940341 390837 940397
rect 390893 940341 390979 940397
rect 391035 940341 391121 940397
rect 391177 940341 391248 940397
rect 389198 940255 391248 940341
rect 389198 940199 389275 940255
rect 389331 940199 389417 940255
rect 389473 940199 389559 940255
rect 389615 940199 389701 940255
rect 389757 940199 389843 940255
rect 389899 940199 389985 940255
rect 390041 940199 390127 940255
rect 390183 940199 390269 940255
rect 390325 940199 390411 940255
rect 390467 940199 390553 940255
rect 390609 940199 390695 940255
rect 390751 940199 390837 940255
rect 390893 940199 390979 940255
rect 391035 940199 391121 940255
rect 391177 940199 391248 940255
rect 389198 940113 391248 940199
rect 389198 940057 389275 940113
rect 389331 940057 389417 940113
rect 389473 940057 389559 940113
rect 389615 940057 389701 940113
rect 389757 940057 389843 940113
rect 389899 940057 389985 940113
rect 390041 940057 390127 940113
rect 390183 940057 390269 940113
rect 390325 940057 390411 940113
rect 390467 940057 390553 940113
rect 390609 940057 390695 940113
rect 390751 940057 390837 940113
rect 390893 940057 390979 940113
rect 391035 940057 391121 940113
rect 391177 940057 391248 940113
rect 389198 939971 391248 940057
rect 389198 939915 389275 939971
rect 389331 939915 389417 939971
rect 389473 939915 389559 939971
rect 389615 939915 389701 939971
rect 389757 939915 389843 939971
rect 389899 939915 389985 939971
rect 390041 939915 390127 939971
rect 390183 939915 390269 939971
rect 390325 939915 390411 939971
rect 390467 939915 390553 939971
rect 390609 939915 390695 939971
rect 390751 939915 390837 939971
rect 390893 939915 390979 939971
rect 391035 939915 391121 939971
rect 391177 939915 391248 939971
rect 389198 939829 391248 939915
rect 389198 939773 389275 939829
rect 389331 939773 389417 939829
rect 389473 939773 389559 939829
rect 389615 939773 389701 939829
rect 389757 939773 389843 939829
rect 389899 939773 389985 939829
rect 390041 939773 390127 939829
rect 390183 939773 390269 939829
rect 390325 939773 390411 939829
rect 390467 939773 390553 939829
rect 390609 939773 390695 939829
rect 390751 939773 390837 939829
rect 390893 939773 390979 939829
rect 391035 939773 391121 939829
rect 391177 939773 391248 939829
rect 389198 939720 391248 939773
rect 391828 941675 393728 941720
rect 391828 941619 391897 941675
rect 391953 941619 392039 941675
rect 392095 941619 392181 941675
rect 392237 941619 392323 941675
rect 392379 941619 392465 941675
rect 392521 941619 392607 941675
rect 392663 941619 392749 941675
rect 392805 941619 392891 941675
rect 392947 941619 393033 941675
rect 393089 941619 393175 941675
rect 393231 941619 393317 941675
rect 393373 941619 393459 941675
rect 393515 941619 393601 941675
rect 393657 941619 393728 941675
rect 391828 941533 393728 941619
rect 391828 941477 391897 941533
rect 391953 941477 392039 941533
rect 392095 941477 392181 941533
rect 392237 941477 392323 941533
rect 392379 941477 392465 941533
rect 392521 941477 392607 941533
rect 392663 941477 392749 941533
rect 392805 941477 392891 941533
rect 392947 941477 393033 941533
rect 393089 941477 393175 941533
rect 393231 941477 393317 941533
rect 393373 941477 393459 941533
rect 393515 941477 393601 941533
rect 393657 941477 393728 941533
rect 391828 941391 393728 941477
rect 391828 941335 391897 941391
rect 391953 941335 392039 941391
rect 392095 941335 392181 941391
rect 392237 941335 392323 941391
rect 392379 941335 392465 941391
rect 392521 941335 392607 941391
rect 392663 941335 392749 941391
rect 392805 941335 392891 941391
rect 392947 941335 393033 941391
rect 393089 941335 393175 941391
rect 393231 941335 393317 941391
rect 393373 941335 393459 941391
rect 393515 941335 393601 941391
rect 393657 941335 393728 941391
rect 391828 941249 393728 941335
rect 391828 941193 391897 941249
rect 391953 941193 392039 941249
rect 392095 941193 392181 941249
rect 392237 941193 392323 941249
rect 392379 941193 392465 941249
rect 392521 941193 392607 941249
rect 392663 941193 392749 941249
rect 392805 941193 392891 941249
rect 392947 941193 393033 941249
rect 393089 941193 393175 941249
rect 393231 941193 393317 941249
rect 393373 941193 393459 941249
rect 393515 941193 393601 941249
rect 393657 941193 393728 941249
rect 391828 941107 393728 941193
rect 391828 941051 391897 941107
rect 391953 941051 392039 941107
rect 392095 941051 392181 941107
rect 392237 941051 392323 941107
rect 392379 941051 392465 941107
rect 392521 941051 392607 941107
rect 392663 941051 392749 941107
rect 392805 941051 392891 941107
rect 392947 941051 393033 941107
rect 393089 941051 393175 941107
rect 393231 941051 393317 941107
rect 393373 941051 393459 941107
rect 393515 941051 393601 941107
rect 393657 941051 393728 941107
rect 391828 940965 393728 941051
rect 391828 940909 391897 940965
rect 391953 940909 392039 940965
rect 392095 940909 392181 940965
rect 392237 940909 392323 940965
rect 392379 940909 392465 940965
rect 392521 940909 392607 940965
rect 392663 940909 392749 940965
rect 392805 940909 392891 940965
rect 392947 940909 393033 940965
rect 393089 940909 393175 940965
rect 393231 940909 393317 940965
rect 393373 940909 393459 940965
rect 393515 940909 393601 940965
rect 393657 940909 393728 940965
rect 391828 940823 393728 940909
rect 391828 940767 391897 940823
rect 391953 940767 392039 940823
rect 392095 940767 392181 940823
rect 392237 940767 392323 940823
rect 392379 940767 392465 940823
rect 392521 940767 392607 940823
rect 392663 940767 392749 940823
rect 392805 940767 392891 940823
rect 392947 940767 393033 940823
rect 393089 940767 393175 940823
rect 393231 940767 393317 940823
rect 393373 940767 393459 940823
rect 393515 940767 393601 940823
rect 393657 940767 393728 940823
rect 391828 940681 393728 940767
rect 391828 940625 391897 940681
rect 391953 940625 392039 940681
rect 392095 940625 392181 940681
rect 392237 940625 392323 940681
rect 392379 940625 392465 940681
rect 392521 940625 392607 940681
rect 392663 940625 392749 940681
rect 392805 940625 392891 940681
rect 392947 940625 393033 940681
rect 393089 940625 393175 940681
rect 393231 940625 393317 940681
rect 393373 940625 393459 940681
rect 393515 940625 393601 940681
rect 393657 940625 393728 940681
rect 391828 940539 393728 940625
rect 391828 940483 391897 940539
rect 391953 940483 392039 940539
rect 392095 940483 392181 940539
rect 392237 940483 392323 940539
rect 392379 940483 392465 940539
rect 392521 940483 392607 940539
rect 392663 940483 392749 940539
rect 392805 940483 392891 940539
rect 392947 940483 393033 940539
rect 393089 940483 393175 940539
rect 393231 940483 393317 940539
rect 393373 940483 393459 940539
rect 393515 940483 393601 940539
rect 393657 940483 393728 940539
rect 391828 940397 393728 940483
rect 391828 940341 391897 940397
rect 391953 940341 392039 940397
rect 392095 940341 392181 940397
rect 392237 940341 392323 940397
rect 392379 940341 392465 940397
rect 392521 940341 392607 940397
rect 392663 940341 392749 940397
rect 392805 940341 392891 940397
rect 392947 940341 393033 940397
rect 393089 940341 393175 940397
rect 393231 940341 393317 940397
rect 393373 940341 393459 940397
rect 393515 940341 393601 940397
rect 393657 940341 393728 940397
rect 391828 940255 393728 940341
rect 391828 940199 391897 940255
rect 391953 940199 392039 940255
rect 392095 940199 392181 940255
rect 392237 940199 392323 940255
rect 392379 940199 392465 940255
rect 392521 940199 392607 940255
rect 392663 940199 392749 940255
rect 392805 940199 392891 940255
rect 392947 940199 393033 940255
rect 393089 940199 393175 940255
rect 393231 940199 393317 940255
rect 393373 940199 393459 940255
rect 393515 940199 393601 940255
rect 393657 940199 393728 940255
rect 391828 940113 393728 940199
rect 391828 940057 391897 940113
rect 391953 940057 392039 940113
rect 392095 940057 392181 940113
rect 392237 940057 392323 940113
rect 392379 940057 392465 940113
rect 392521 940057 392607 940113
rect 392663 940057 392749 940113
rect 392805 940057 392891 940113
rect 392947 940057 393033 940113
rect 393089 940057 393175 940113
rect 393231 940057 393317 940113
rect 393373 940057 393459 940113
rect 393515 940057 393601 940113
rect 393657 940057 393728 940113
rect 391828 939971 393728 940057
rect 391828 939915 391897 939971
rect 391953 939915 392039 939971
rect 392095 939915 392181 939971
rect 392237 939915 392323 939971
rect 392379 939915 392465 939971
rect 392521 939915 392607 939971
rect 392663 939915 392749 939971
rect 392805 939915 392891 939971
rect 392947 939915 393033 939971
rect 393089 939915 393175 939971
rect 393231 939915 393317 939971
rect 393373 939915 393459 939971
rect 393515 939915 393601 939971
rect 393657 939915 393728 939971
rect 391828 939829 393728 939915
rect 391828 939773 391897 939829
rect 391953 939773 392039 939829
rect 392095 939773 392181 939829
rect 392237 939773 392323 939829
rect 392379 939773 392465 939829
rect 392521 939773 392607 939829
rect 392663 939773 392749 939829
rect 392805 939773 392891 939829
rect 392947 939773 393033 939829
rect 393089 939773 393175 939829
rect 393231 939773 393317 939829
rect 393373 939773 393459 939829
rect 393515 939773 393601 939829
rect 393657 939773 393728 939829
rect 391828 939720 393728 939773
rect 599272 941675 601172 941720
rect 599272 941619 599341 941675
rect 599397 941619 599483 941675
rect 599539 941619 599625 941675
rect 599681 941619 599767 941675
rect 599823 941619 599909 941675
rect 599965 941619 600051 941675
rect 600107 941619 600193 941675
rect 600249 941619 600335 941675
rect 600391 941619 600477 941675
rect 600533 941619 600619 941675
rect 600675 941619 600761 941675
rect 600817 941619 600903 941675
rect 600959 941619 601045 941675
rect 601101 941619 601172 941675
rect 599272 941533 601172 941619
rect 599272 941477 599341 941533
rect 599397 941477 599483 941533
rect 599539 941477 599625 941533
rect 599681 941477 599767 941533
rect 599823 941477 599909 941533
rect 599965 941477 600051 941533
rect 600107 941477 600193 941533
rect 600249 941477 600335 941533
rect 600391 941477 600477 941533
rect 600533 941477 600619 941533
rect 600675 941477 600761 941533
rect 600817 941477 600903 941533
rect 600959 941477 601045 941533
rect 601101 941477 601172 941533
rect 599272 941391 601172 941477
rect 599272 941335 599341 941391
rect 599397 941335 599483 941391
rect 599539 941335 599625 941391
rect 599681 941335 599767 941391
rect 599823 941335 599909 941391
rect 599965 941335 600051 941391
rect 600107 941335 600193 941391
rect 600249 941335 600335 941391
rect 600391 941335 600477 941391
rect 600533 941335 600619 941391
rect 600675 941335 600761 941391
rect 600817 941335 600903 941391
rect 600959 941335 601045 941391
rect 601101 941335 601172 941391
rect 599272 941249 601172 941335
rect 599272 941193 599341 941249
rect 599397 941193 599483 941249
rect 599539 941193 599625 941249
rect 599681 941193 599767 941249
rect 599823 941193 599909 941249
rect 599965 941193 600051 941249
rect 600107 941193 600193 941249
rect 600249 941193 600335 941249
rect 600391 941193 600477 941249
rect 600533 941193 600619 941249
rect 600675 941193 600761 941249
rect 600817 941193 600903 941249
rect 600959 941193 601045 941249
rect 601101 941193 601172 941249
rect 599272 941107 601172 941193
rect 599272 941051 599341 941107
rect 599397 941051 599483 941107
rect 599539 941051 599625 941107
rect 599681 941051 599767 941107
rect 599823 941051 599909 941107
rect 599965 941051 600051 941107
rect 600107 941051 600193 941107
rect 600249 941051 600335 941107
rect 600391 941051 600477 941107
rect 600533 941051 600619 941107
rect 600675 941051 600761 941107
rect 600817 941051 600903 941107
rect 600959 941051 601045 941107
rect 601101 941051 601172 941107
rect 599272 940965 601172 941051
rect 599272 940909 599341 940965
rect 599397 940909 599483 940965
rect 599539 940909 599625 940965
rect 599681 940909 599767 940965
rect 599823 940909 599909 940965
rect 599965 940909 600051 940965
rect 600107 940909 600193 940965
rect 600249 940909 600335 940965
rect 600391 940909 600477 940965
rect 600533 940909 600619 940965
rect 600675 940909 600761 940965
rect 600817 940909 600903 940965
rect 600959 940909 601045 940965
rect 601101 940909 601172 940965
rect 599272 940823 601172 940909
rect 599272 940767 599341 940823
rect 599397 940767 599483 940823
rect 599539 940767 599625 940823
rect 599681 940767 599767 940823
rect 599823 940767 599909 940823
rect 599965 940767 600051 940823
rect 600107 940767 600193 940823
rect 600249 940767 600335 940823
rect 600391 940767 600477 940823
rect 600533 940767 600619 940823
rect 600675 940767 600761 940823
rect 600817 940767 600903 940823
rect 600959 940767 601045 940823
rect 601101 940767 601172 940823
rect 599272 940681 601172 940767
rect 599272 940625 599341 940681
rect 599397 940625 599483 940681
rect 599539 940625 599625 940681
rect 599681 940625 599767 940681
rect 599823 940625 599909 940681
rect 599965 940625 600051 940681
rect 600107 940625 600193 940681
rect 600249 940625 600335 940681
rect 600391 940625 600477 940681
rect 600533 940625 600619 940681
rect 600675 940625 600761 940681
rect 600817 940625 600903 940681
rect 600959 940625 601045 940681
rect 601101 940625 601172 940681
rect 599272 940539 601172 940625
rect 599272 940483 599341 940539
rect 599397 940483 599483 940539
rect 599539 940483 599625 940539
rect 599681 940483 599767 940539
rect 599823 940483 599909 940539
rect 599965 940483 600051 940539
rect 600107 940483 600193 940539
rect 600249 940483 600335 940539
rect 600391 940483 600477 940539
rect 600533 940483 600619 940539
rect 600675 940483 600761 940539
rect 600817 940483 600903 940539
rect 600959 940483 601045 940539
rect 601101 940483 601172 940539
rect 599272 940397 601172 940483
rect 599272 940341 599341 940397
rect 599397 940341 599483 940397
rect 599539 940341 599625 940397
rect 599681 940341 599767 940397
rect 599823 940341 599909 940397
rect 599965 940341 600051 940397
rect 600107 940341 600193 940397
rect 600249 940341 600335 940397
rect 600391 940341 600477 940397
rect 600533 940341 600619 940397
rect 600675 940341 600761 940397
rect 600817 940341 600903 940397
rect 600959 940341 601045 940397
rect 601101 940341 601172 940397
rect 599272 940255 601172 940341
rect 599272 940199 599341 940255
rect 599397 940199 599483 940255
rect 599539 940199 599625 940255
rect 599681 940199 599767 940255
rect 599823 940199 599909 940255
rect 599965 940199 600051 940255
rect 600107 940199 600193 940255
rect 600249 940199 600335 940255
rect 600391 940199 600477 940255
rect 600533 940199 600619 940255
rect 600675 940199 600761 940255
rect 600817 940199 600903 940255
rect 600959 940199 601045 940255
rect 601101 940199 601172 940255
rect 599272 940113 601172 940199
rect 599272 940057 599341 940113
rect 599397 940057 599483 940113
rect 599539 940057 599625 940113
rect 599681 940057 599767 940113
rect 599823 940057 599909 940113
rect 599965 940057 600051 940113
rect 600107 940057 600193 940113
rect 600249 940057 600335 940113
rect 600391 940057 600477 940113
rect 600533 940057 600619 940113
rect 600675 940057 600761 940113
rect 600817 940057 600903 940113
rect 600959 940057 601045 940113
rect 601101 940057 601172 940113
rect 599272 939971 601172 940057
rect 599272 939915 599341 939971
rect 599397 939915 599483 939971
rect 599539 939915 599625 939971
rect 599681 939915 599767 939971
rect 599823 939915 599909 939971
rect 599965 939915 600051 939971
rect 600107 939915 600193 939971
rect 600249 939915 600335 939971
rect 600391 939915 600477 939971
rect 600533 939915 600619 939971
rect 600675 939915 600761 939971
rect 600817 939915 600903 939971
rect 600959 939915 601045 939971
rect 601101 939915 601172 939971
rect 599272 939829 601172 939915
rect 599272 939773 599341 939829
rect 599397 939773 599483 939829
rect 599539 939773 599625 939829
rect 599681 939773 599767 939829
rect 599823 939773 599909 939829
rect 599965 939773 600051 939829
rect 600107 939773 600193 939829
rect 600249 939773 600335 939829
rect 600391 939773 600477 939829
rect 600533 939773 600619 939829
rect 600675 939773 600761 939829
rect 600817 939773 600903 939829
rect 600959 939773 601045 939829
rect 601101 939773 601172 939829
rect 599272 939720 601172 939773
rect 601752 941675 603802 941720
rect 601752 941619 601829 941675
rect 601885 941619 601971 941675
rect 602027 941619 602113 941675
rect 602169 941619 602255 941675
rect 602311 941619 602397 941675
rect 602453 941619 602539 941675
rect 602595 941619 602681 941675
rect 602737 941619 602823 941675
rect 602879 941619 602965 941675
rect 603021 941619 603107 941675
rect 603163 941619 603249 941675
rect 603305 941619 603391 941675
rect 603447 941619 603533 941675
rect 603589 941619 603675 941675
rect 603731 941619 603802 941675
rect 601752 941533 603802 941619
rect 601752 941477 601829 941533
rect 601885 941477 601971 941533
rect 602027 941477 602113 941533
rect 602169 941477 602255 941533
rect 602311 941477 602397 941533
rect 602453 941477 602539 941533
rect 602595 941477 602681 941533
rect 602737 941477 602823 941533
rect 602879 941477 602965 941533
rect 603021 941477 603107 941533
rect 603163 941477 603249 941533
rect 603305 941477 603391 941533
rect 603447 941477 603533 941533
rect 603589 941477 603675 941533
rect 603731 941477 603802 941533
rect 601752 941391 603802 941477
rect 601752 941335 601829 941391
rect 601885 941335 601971 941391
rect 602027 941335 602113 941391
rect 602169 941335 602255 941391
rect 602311 941335 602397 941391
rect 602453 941335 602539 941391
rect 602595 941335 602681 941391
rect 602737 941335 602823 941391
rect 602879 941335 602965 941391
rect 603021 941335 603107 941391
rect 603163 941335 603249 941391
rect 603305 941335 603391 941391
rect 603447 941335 603533 941391
rect 603589 941335 603675 941391
rect 603731 941335 603802 941391
rect 601752 941249 603802 941335
rect 601752 941193 601829 941249
rect 601885 941193 601971 941249
rect 602027 941193 602113 941249
rect 602169 941193 602255 941249
rect 602311 941193 602397 941249
rect 602453 941193 602539 941249
rect 602595 941193 602681 941249
rect 602737 941193 602823 941249
rect 602879 941193 602965 941249
rect 603021 941193 603107 941249
rect 603163 941193 603249 941249
rect 603305 941193 603391 941249
rect 603447 941193 603533 941249
rect 603589 941193 603675 941249
rect 603731 941193 603802 941249
rect 601752 941107 603802 941193
rect 601752 941051 601829 941107
rect 601885 941051 601971 941107
rect 602027 941051 602113 941107
rect 602169 941051 602255 941107
rect 602311 941051 602397 941107
rect 602453 941051 602539 941107
rect 602595 941051 602681 941107
rect 602737 941051 602823 941107
rect 602879 941051 602965 941107
rect 603021 941051 603107 941107
rect 603163 941051 603249 941107
rect 603305 941051 603391 941107
rect 603447 941051 603533 941107
rect 603589 941051 603675 941107
rect 603731 941051 603802 941107
rect 601752 940965 603802 941051
rect 601752 940909 601829 940965
rect 601885 940909 601971 940965
rect 602027 940909 602113 940965
rect 602169 940909 602255 940965
rect 602311 940909 602397 940965
rect 602453 940909 602539 940965
rect 602595 940909 602681 940965
rect 602737 940909 602823 940965
rect 602879 940909 602965 940965
rect 603021 940909 603107 940965
rect 603163 940909 603249 940965
rect 603305 940909 603391 940965
rect 603447 940909 603533 940965
rect 603589 940909 603675 940965
rect 603731 940909 603802 940965
rect 601752 940823 603802 940909
rect 601752 940767 601829 940823
rect 601885 940767 601971 940823
rect 602027 940767 602113 940823
rect 602169 940767 602255 940823
rect 602311 940767 602397 940823
rect 602453 940767 602539 940823
rect 602595 940767 602681 940823
rect 602737 940767 602823 940823
rect 602879 940767 602965 940823
rect 603021 940767 603107 940823
rect 603163 940767 603249 940823
rect 603305 940767 603391 940823
rect 603447 940767 603533 940823
rect 603589 940767 603675 940823
rect 603731 940767 603802 940823
rect 601752 940681 603802 940767
rect 601752 940625 601829 940681
rect 601885 940625 601971 940681
rect 602027 940625 602113 940681
rect 602169 940625 602255 940681
rect 602311 940625 602397 940681
rect 602453 940625 602539 940681
rect 602595 940625 602681 940681
rect 602737 940625 602823 940681
rect 602879 940625 602965 940681
rect 603021 940625 603107 940681
rect 603163 940625 603249 940681
rect 603305 940625 603391 940681
rect 603447 940625 603533 940681
rect 603589 940625 603675 940681
rect 603731 940625 603802 940681
rect 601752 940539 603802 940625
rect 601752 940483 601829 940539
rect 601885 940483 601971 940539
rect 602027 940483 602113 940539
rect 602169 940483 602255 940539
rect 602311 940483 602397 940539
rect 602453 940483 602539 940539
rect 602595 940483 602681 940539
rect 602737 940483 602823 940539
rect 602879 940483 602965 940539
rect 603021 940483 603107 940539
rect 603163 940483 603249 940539
rect 603305 940483 603391 940539
rect 603447 940483 603533 940539
rect 603589 940483 603675 940539
rect 603731 940483 603802 940539
rect 601752 940397 603802 940483
rect 601752 940341 601829 940397
rect 601885 940341 601971 940397
rect 602027 940341 602113 940397
rect 602169 940341 602255 940397
rect 602311 940341 602397 940397
rect 602453 940341 602539 940397
rect 602595 940341 602681 940397
rect 602737 940341 602823 940397
rect 602879 940341 602965 940397
rect 603021 940341 603107 940397
rect 603163 940341 603249 940397
rect 603305 940341 603391 940397
rect 603447 940341 603533 940397
rect 603589 940341 603675 940397
rect 603731 940341 603802 940397
rect 601752 940255 603802 940341
rect 601752 940199 601829 940255
rect 601885 940199 601971 940255
rect 602027 940199 602113 940255
rect 602169 940199 602255 940255
rect 602311 940199 602397 940255
rect 602453 940199 602539 940255
rect 602595 940199 602681 940255
rect 602737 940199 602823 940255
rect 602879 940199 602965 940255
rect 603021 940199 603107 940255
rect 603163 940199 603249 940255
rect 603305 940199 603391 940255
rect 603447 940199 603533 940255
rect 603589 940199 603675 940255
rect 603731 940199 603802 940255
rect 601752 940113 603802 940199
rect 601752 940057 601829 940113
rect 601885 940057 601971 940113
rect 602027 940057 602113 940113
rect 602169 940057 602255 940113
rect 602311 940057 602397 940113
rect 602453 940057 602539 940113
rect 602595 940057 602681 940113
rect 602737 940057 602823 940113
rect 602879 940057 602965 940113
rect 603021 940057 603107 940113
rect 603163 940057 603249 940113
rect 603305 940057 603391 940113
rect 603447 940057 603533 940113
rect 603589 940057 603675 940113
rect 603731 940057 603802 940113
rect 601752 939971 603802 940057
rect 601752 939915 601829 939971
rect 601885 939915 601971 939971
rect 602027 939915 602113 939971
rect 602169 939915 602255 939971
rect 602311 939915 602397 939971
rect 602453 939915 602539 939971
rect 602595 939915 602681 939971
rect 602737 939915 602823 939971
rect 602879 939915 602965 939971
rect 603021 939915 603107 939971
rect 603163 939915 603249 939971
rect 603305 939915 603391 939971
rect 603447 939915 603533 939971
rect 603589 939915 603675 939971
rect 603731 939915 603802 939971
rect 601752 939829 603802 939915
rect 601752 939773 601829 939829
rect 601885 939773 601971 939829
rect 602027 939773 602113 939829
rect 602169 939773 602255 939829
rect 602311 939773 602397 939829
rect 602453 939773 602539 939829
rect 602595 939773 602681 939829
rect 602737 939773 602823 939829
rect 602879 939773 602965 939829
rect 603021 939773 603107 939829
rect 603163 939773 603249 939829
rect 603305 939773 603391 939829
rect 603447 939773 603533 939829
rect 603589 939773 603675 939829
rect 603731 939773 603802 939829
rect 601752 939720 603802 939773
rect 605020 941675 606172 941720
rect 605020 941619 605051 941675
rect 605107 941619 605193 941675
rect 605249 941619 605335 941675
rect 605391 941619 605477 941675
rect 605533 941619 605619 941675
rect 605675 941619 605761 941675
rect 605817 941619 605903 941675
rect 605959 941619 606045 941675
rect 606101 941619 606172 941675
rect 605020 941533 606172 941619
rect 605020 941477 605051 941533
rect 605107 941477 605193 941533
rect 605249 941477 605335 941533
rect 605391 941477 605477 941533
rect 605533 941477 605619 941533
rect 605675 941477 605761 941533
rect 605817 941477 605903 941533
rect 605959 941477 606045 941533
rect 606101 941477 606172 941533
rect 605020 941391 606172 941477
rect 605020 941335 605051 941391
rect 605107 941335 605193 941391
rect 605249 941335 605335 941391
rect 605391 941335 605477 941391
rect 605533 941335 605619 941391
rect 605675 941335 605761 941391
rect 605817 941335 605903 941391
rect 605959 941335 606045 941391
rect 606101 941335 606172 941391
rect 605020 941249 606172 941335
rect 605020 941193 605051 941249
rect 605107 941193 605193 941249
rect 605249 941193 605335 941249
rect 605391 941193 605477 941249
rect 605533 941193 605619 941249
rect 605675 941193 605761 941249
rect 605817 941193 605903 941249
rect 605959 941193 606045 941249
rect 606101 941193 606172 941249
rect 605020 941107 606172 941193
rect 605020 941051 605051 941107
rect 605107 941051 605193 941107
rect 605249 941051 605335 941107
rect 605391 941051 605477 941107
rect 605533 941051 605619 941107
rect 605675 941051 605761 941107
rect 605817 941051 605903 941107
rect 605959 941051 606045 941107
rect 606101 941051 606172 941107
rect 605020 940965 606172 941051
rect 605020 940909 605051 940965
rect 605107 940909 605193 940965
rect 605249 940909 605335 940965
rect 605391 940909 605477 940965
rect 605533 940909 605619 940965
rect 605675 940909 605761 940965
rect 605817 940909 605903 940965
rect 605959 940909 606045 940965
rect 606101 940909 606172 940965
rect 605020 940823 606172 940909
rect 605020 940767 605051 940823
rect 605107 940767 605193 940823
rect 605249 940767 605335 940823
rect 605391 940767 605477 940823
rect 605533 940767 605619 940823
rect 605675 940767 605761 940823
rect 605817 940767 605903 940823
rect 605959 940767 606045 940823
rect 606101 940767 606172 940823
rect 605020 940681 606172 940767
rect 605020 940625 605051 940681
rect 605107 940625 605193 940681
rect 605249 940625 605335 940681
rect 605391 940625 605477 940681
rect 605533 940625 605619 940681
rect 605675 940625 605761 940681
rect 605817 940625 605903 940681
rect 605959 940625 606045 940681
rect 606101 940625 606172 940681
rect 605020 940539 606172 940625
rect 605020 940483 605051 940539
rect 605107 940483 605193 940539
rect 605249 940483 605335 940539
rect 605391 940483 605477 940539
rect 605533 940483 605619 940539
rect 605675 940483 605761 940539
rect 605817 940483 605903 940539
rect 605959 940483 606045 940539
rect 606101 940483 606172 940539
rect 605020 940397 606172 940483
rect 605020 940341 605051 940397
rect 605107 940341 605193 940397
rect 605249 940341 605335 940397
rect 605391 940341 605477 940397
rect 605533 940341 605619 940397
rect 605675 940341 605761 940397
rect 605817 940341 605903 940397
rect 605959 940341 606045 940397
rect 606101 940341 606172 940397
rect 605020 940255 606172 940341
rect 605020 940199 605051 940255
rect 605107 940199 605193 940255
rect 605249 940199 605335 940255
rect 605391 940199 605477 940255
rect 605533 940199 605619 940255
rect 605675 940199 605761 940255
rect 605817 940199 605903 940255
rect 605959 940199 606045 940255
rect 606101 940199 606172 940255
rect 605020 940113 606172 940199
rect 605020 940057 605051 940113
rect 605107 940057 605193 940113
rect 605249 940057 605335 940113
rect 605391 940057 605477 940113
rect 605533 940057 605619 940113
rect 605675 940057 605761 940113
rect 605817 940057 605903 940113
rect 605959 940057 606045 940113
rect 606101 940057 606172 940113
rect 605020 939971 606172 940057
rect 605020 939915 605051 939971
rect 605107 939915 605193 939971
rect 605249 939915 605335 939971
rect 605391 939915 605477 939971
rect 605533 939915 605619 939971
rect 605675 939915 605761 939971
rect 605817 939915 605903 939971
rect 605959 939915 606045 939971
rect 606101 939915 606172 939971
rect 605020 939829 606172 939915
rect 605020 939773 605051 939829
rect 605107 939773 605193 939829
rect 605249 939773 605335 939829
rect 605391 939773 605477 939829
rect 605533 939773 605619 939829
rect 605675 939773 605761 939829
rect 605817 939773 605903 939829
rect 605959 939773 606045 939829
rect 606101 939773 606172 939829
rect 605020 939720 606172 939773
rect 606828 941675 608878 941720
rect 606828 941619 606905 941675
rect 606961 941619 607047 941675
rect 607103 941619 607189 941675
rect 607245 941619 607331 941675
rect 607387 941619 607473 941675
rect 607529 941619 607615 941675
rect 607671 941619 607757 941675
rect 607813 941619 607899 941675
rect 607955 941619 608041 941675
rect 608097 941619 608183 941675
rect 608239 941619 608325 941675
rect 608381 941619 608467 941675
rect 608523 941619 608609 941675
rect 608665 941619 608751 941675
rect 608807 941619 608878 941675
rect 606828 941533 608878 941619
rect 606828 941477 606905 941533
rect 606961 941477 607047 941533
rect 607103 941477 607189 941533
rect 607245 941477 607331 941533
rect 607387 941477 607473 941533
rect 607529 941477 607615 941533
rect 607671 941477 607757 941533
rect 607813 941477 607899 941533
rect 607955 941477 608041 941533
rect 608097 941477 608183 941533
rect 608239 941477 608325 941533
rect 608381 941477 608467 941533
rect 608523 941477 608609 941533
rect 608665 941477 608751 941533
rect 608807 941477 608878 941533
rect 606828 941391 608878 941477
rect 606828 941335 606905 941391
rect 606961 941335 607047 941391
rect 607103 941335 607189 941391
rect 607245 941335 607331 941391
rect 607387 941335 607473 941391
rect 607529 941335 607615 941391
rect 607671 941335 607757 941391
rect 607813 941335 607899 941391
rect 607955 941335 608041 941391
rect 608097 941335 608183 941391
rect 608239 941335 608325 941391
rect 608381 941335 608467 941391
rect 608523 941335 608609 941391
rect 608665 941335 608751 941391
rect 608807 941335 608878 941391
rect 606828 941249 608878 941335
rect 606828 941193 606905 941249
rect 606961 941193 607047 941249
rect 607103 941193 607189 941249
rect 607245 941193 607331 941249
rect 607387 941193 607473 941249
rect 607529 941193 607615 941249
rect 607671 941193 607757 941249
rect 607813 941193 607899 941249
rect 607955 941193 608041 941249
rect 608097 941193 608183 941249
rect 608239 941193 608325 941249
rect 608381 941193 608467 941249
rect 608523 941193 608609 941249
rect 608665 941193 608751 941249
rect 608807 941193 608878 941249
rect 606828 941107 608878 941193
rect 606828 941051 606905 941107
rect 606961 941051 607047 941107
rect 607103 941051 607189 941107
rect 607245 941051 607331 941107
rect 607387 941051 607473 941107
rect 607529 941051 607615 941107
rect 607671 941051 607757 941107
rect 607813 941051 607899 941107
rect 607955 941051 608041 941107
rect 608097 941051 608183 941107
rect 608239 941051 608325 941107
rect 608381 941051 608467 941107
rect 608523 941051 608609 941107
rect 608665 941051 608751 941107
rect 608807 941051 608878 941107
rect 606828 940965 608878 941051
rect 606828 940909 606905 940965
rect 606961 940909 607047 940965
rect 607103 940909 607189 940965
rect 607245 940909 607331 940965
rect 607387 940909 607473 940965
rect 607529 940909 607615 940965
rect 607671 940909 607757 940965
rect 607813 940909 607899 940965
rect 607955 940909 608041 940965
rect 608097 940909 608183 940965
rect 608239 940909 608325 940965
rect 608381 940909 608467 940965
rect 608523 940909 608609 940965
rect 608665 940909 608751 940965
rect 608807 940909 608878 940965
rect 606828 940823 608878 940909
rect 606828 940767 606905 940823
rect 606961 940767 607047 940823
rect 607103 940767 607189 940823
rect 607245 940767 607331 940823
rect 607387 940767 607473 940823
rect 607529 940767 607615 940823
rect 607671 940767 607757 940823
rect 607813 940767 607899 940823
rect 607955 940767 608041 940823
rect 608097 940767 608183 940823
rect 608239 940767 608325 940823
rect 608381 940767 608467 940823
rect 608523 940767 608609 940823
rect 608665 940767 608751 940823
rect 608807 940767 608878 940823
rect 606828 940681 608878 940767
rect 606828 940625 606905 940681
rect 606961 940625 607047 940681
rect 607103 940625 607189 940681
rect 607245 940625 607331 940681
rect 607387 940625 607473 940681
rect 607529 940625 607615 940681
rect 607671 940625 607757 940681
rect 607813 940625 607899 940681
rect 607955 940625 608041 940681
rect 608097 940625 608183 940681
rect 608239 940625 608325 940681
rect 608381 940625 608467 940681
rect 608523 940625 608609 940681
rect 608665 940625 608751 940681
rect 608807 940625 608878 940681
rect 606828 940539 608878 940625
rect 606828 940483 606905 940539
rect 606961 940483 607047 940539
rect 607103 940483 607189 940539
rect 607245 940483 607331 940539
rect 607387 940483 607473 940539
rect 607529 940483 607615 940539
rect 607671 940483 607757 940539
rect 607813 940483 607899 940539
rect 607955 940483 608041 940539
rect 608097 940483 608183 940539
rect 608239 940483 608325 940539
rect 608381 940483 608467 940539
rect 608523 940483 608609 940539
rect 608665 940483 608751 940539
rect 608807 940483 608878 940539
rect 606828 940397 608878 940483
rect 606828 940341 606905 940397
rect 606961 940341 607047 940397
rect 607103 940341 607189 940397
rect 607245 940341 607331 940397
rect 607387 940341 607473 940397
rect 607529 940341 607615 940397
rect 607671 940341 607757 940397
rect 607813 940341 607899 940397
rect 607955 940341 608041 940397
rect 608097 940341 608183 940397
rect 608239 940341 608325 940397
rect 608381 940341 608467 940397
rect 608523 940341 608609 940397
rect 608665 940341 608751 940397
rect 608807 940341 608878 940397
rect 606828 940255 608878 940341
rect 606828 940199 606905 940255
rect 606961 940199 607047 940255
rect 607103 940199 607189 940255
rect 607245 940199 607331 940255
rect 607387 940199 607473 940255
rect 607529 940199 607615 940255
rect 607671 940199 607757 940255
rect 607813 940199 607899 940255
rect 607955 940199 608041 940255
rect 608097 940199 608183 940255
rect 608239 940199 608325 940255
rect 608381 940199 608467 940255
rect 608523 940199 608609 940255
rect 608665 940199 608751 940255
rect 608807 940199 608878 940255
rect 606828 940113 608878 940199
rect 606828 940057 606905 940113
rect 606961 940057 607047 940113
rect 607103 940057 607189 940113
rect 607245 940057 607331 940113
rect 607387 940057 607473 940113
rect 607529 940057 607615 940113
rect 607671 940057 607757 940113
rect 607813 940057 607899 940113
rect 607955 940057 608041 940113
rect 608097 940057 608183 940113
rect 608239 940057 608325 940113
rect 608381 940057 608467 940113
rect 608523 940057 608609 940113
rect 608665 940057 608751 940113
rect 608807 940057 608878 940113
rect 606828 939971 608878 940057
rect 606828 939915 606905 939971
rect 606961 939915 607047 939971
rect 607103 939915 607189 939971
rect 607245 939915 607331 939971
rect 607387 939915 607473 939971
rect 607529 939915 607615 939971
rect 607671 939915 607757 939971
rect 607813 939915 607899 939971
rect 607955 939915 608041 939971
rect 608097 939915 608183 939971
rect 608239 939915 608325 939971
rect 608381 939915 608467 939971
rect 608523 939915 608609 939971
rect 608665 939915 608751 939971
rect 608807 939915 608878 939971
rect 606828 939829 608878 939915
rect 606828 939773 606905 939829
rect 606961 939773 607047 939829
rect 607103 939773 607189 939829
rect 607245 939773 607331 939829
rect 607387 939773 607473 939829
rect 607529 939773 607615 939829
rect 607671 939773 607757 939829
rect 607813 939773 607899 939829
rect 607955 939773 608041 939829
rect 608097 939773 608183 939829
rect 608239 939773 608325 939829
rect 608381 939773 608467 939829
rect 608523 939773 608609 939829
rect 608665 939773 608751 939829
rect 608807 939773 608878 939829
rect 606828 939720 608878 939773
rect 609198 941675 611248 941720
rect 609198 941619 609275 941675
rect 609331 941619 609417 941675
rect 609473 941619 609559 941675
rect 609615 941619 609701 941675
rect 609757 941619 609843 941675
rect 609899 941619 609985 941675
rect 610041 941619 610127 941675
rect 610183 941619 610269 941675
rect 610325 941619 610411 941675
rect 610467 941619 610553 941675
rect 610609 941619 610695 941675
rect 610751 941619 610837 941675
rect 610893 941619 610979 941675
rect 611035 941619 611121 941675
rect 611177 941619 611248 941675
rect 609198 941533 611248 941619
rect 609198 941477 609275 941533
rect 609331 941477 609417 941533
rect 609473 941477 609559 941533
rect 609615 941477 609701 941533
rect 609757 941477 609843 941533
rect 609899 941477 609985 941533
rect 610041 941477 610127 941533
rect 610183 941477 610269 941533
rect 610325 941477 610411 941533
rect 610467 941477 610553 941533
rect 610609 941477 610695 941533
rect 610751 941477 610837 941533
rect 610893 941477 610979 941533
rect 611035 941477 611121 941533
rect 611177 941477 611248 941533
rect 609198 941391 611248 941477
rect 609198 941335 609275 941391
rect 609331 941335 609417 941391
rect 609473 941335 609559 941391
rect 609615 941335 609701 941391
rect 609757 941335 609843 941391
rect 609899 941335 609985 941391
rect 610041 941335 610127 941391
rect 610183 941335 610269 941391
rect 610325 941335 610411 941391
rect 610467 941335 610553 941391
rect 610609 941335 610695 941391
rect 610751 941335 610837 941391
rect 610893 941335 610979 941391
rect 611035 941335 611121 941391
rect 611177 941335 611248 941391
rect 609198 941249 611248 941335
rect 609198 941193 609275 941249
rect 609331 941193 609417 941249
rect 609473 941193 609559 941249
rect 609615 941193 609701 941249
rect 609757 941193 609843 941249
rect 609899 941193 609985 941249
rect 610041 941193 610127 941249
rect 610183 941193 610269 941249
rect 610325 941193 610411 941249
rect 610467 941193 610553 941249
rect 610609 941193 610695 941249
rect 610751 941193 610837 941249
rect 610893 941193 610979 941249
rect 611035 941193 611121 941249
rect 611177 941193 611248 941249
rect 609198 941107 611248 941193
rect 609198 941051 609275 941107
rect 609331 941051 609417 941107
rect 609473 941051 609559 941107
rect 609615 941051 609701 941107
rect 609757 941051 609843 941107
rect 609899 941051 609985 941107
rect 610041 941051 610127 941107
rect 610183 941051 610269 941107
rect 610325 941051 610411 941107
rect 610467 941051 610553 941107
rect 610609 941051 610695 941107
rect 610751 941051 610837 941107
rect 610893 941051 610979 941107
rect 611035 941051 611121 941107
rect 611177 941051 611248 941107
rect 609198 940965 611248 941051
rect 609198 940909 609275 940965
rect 609331 940909 609417 940965
rect 609473 940909 609559 940965
rect 609615 940909 609701 940965
rect 609757 940909 609843 940965
rect 609899 940909 609985 940965
rect 610041 940909 610127 940965
rect 610183 940909 610269 940965
rect 610325 940909 610411 940965
rect 610467 940909 610553 940965
rect 610609 940909 610695 940965
rect 610751 940909 610837 940965
rect 610893 940909 610979 940965
rect 611035 940909 611121 940965
rect 611177 940909 611248 940965
rect 609198 940823 611248 940909
rect 609198 940767 609275 940823
rect 609331 940767 609417 940823
rect 609473 940767 609559 940823
rect 609615 940767 609701 940823
rect 609757 940767 609843 940823
rect 609899 940767 609985 940823
rect 610041 940767 610127 940823
rect 610183 940767 610269 940823
rect 610325 940767 610411 940823
rect 610467 940767 610553 940823
rect 610609 940767 610695 940823
rect 610751 940767 610837 940823
rect 610893 940767 610979 940823
rect 611035 940767 611121 940823
rect 611177 940767 611248 940823
rect 609198 940681 611248 940767
rect 609198 940625 609275 940681
rect 609331 940625 609417 940681
rect 609473 940625 609559 940681
rect 609615 940625 609701 940681
rect 609757 940625 609843 940681
rect 609899 940625 609985 940681
rect 610041 940625 610127 940681
rect 610183 940625 610269 940681
rect 610325 940625 610411 940681
rect 610467 940625 610553 940681
rect 610609 940625 610695 940681
rect 610751 940625 610837 940681
rect 610893 940625 610979 940681
rect 611035 940625 611121 940681
rect 611177 940625 611248 940681
rect 609198 940539 611248 940625
rect 609198 940483 609275 940539
rect 609331 940483 609417 940539
rect 609473 940483 609559 940539
rect 609615 940483 609701 940539
rect 609757 940483 609843 940539
rect 609899 940483 609985 940539
rect 610041 940483 610127 940539
rect 610183 940483 610269 940539
rect 610325 940483 610411 940539
rect 610467 940483 610553 940539
rect 610609 940483 610695 940539
rect 610751 940483 610837 940539
rect 610893 940483 610979 940539
rect 611035 940483 611121 940539
rect 611177 940483 611248 940539
rect 609198 940397 611248 940483
rect 609198 940341 609275 940397
rect 609331 940341 609417 940397
rect 609473 940341 609559 940397
rect 609615 940341 609701 940397
rect 609757 940341 609843 940397
rect 609899 940341 609985 940397
rect 610041 940341 610127 940397
rect 610183 940341 610269 940397
rect 610325 940341 610411 940397
rect 610467 940341 610553 940397
rect 610609 940341 610695 940397
rect 610751 940341 610837 940397
rect 610893 940341 610979 940397
rect 611035 940341 611121 940397
rect 611177 940341 611248 940397
rect 609198 940255 611248 940341
rect 609198 940199 609275 940255
rect 609331 940199 609417 940255
rect 609473 940199 609559 940255
rect 609615 940199 609701 940255
rect 609757 940199 609843 940255
rect 609899 940199 609985 940255
rect 610041 940199 610127 940255
rect 610183 940199 610269 940255
rect 610325 940199 610411 940255
rect 610467 940199 610553 940255
rect 610609 940199 610695 940255
rect 610751 940199 610837 940255
rect 610893 940199 610979 940255
rect 611035 940199 611121 940255
rect 611177 940199 611248 940255
rect 609198 940113 611248 940199
rect 609198 940057 609275 940113
rect 609331 940057 609417 940113
rect 609473 940057 609559 940113
rect 609615 940057 609701 940113
rect 609757 940057 609843 940113
rect 609899 940057 609985 940113
rect 610041 940057 610127 940113
rect 610183 940057 610269 940113
rect 610325 940057 610411 940113
rect 610467 940057 610553 940113
rect 610609 940057 610695 940113
rect 610751 940057 610837 940113
rect 610893 940057 610979 940113
rect 611035 940057 611121 940113
rect 611177 940057 611248 940113
rect 609198 939971 611248 940057
rect 609198 939915 609275 939971
rect 609331 939915 609417 939971
rect 609473 939915 609559 939971
rect 609615 939915 609701 939971
rect 609757 939915 609843 939971
rect 609899 939915 609985 939971
rect 610041 939915 610127 939971
rect 610183 939915 610269 939971
rect 610325 939915 610411 939971
rect 610467 939915 610553 939971
rect 610609 939915 610695 939971
rect 610751 939915 610837 939971
rect 610893 939915 610979 939971
rect 611035 939915 611121 939971
rect 611177 939915 611248 939971
rect 609198 939829 611248 939915
rect 609198 939773 609275 939829
rect 609331 939773 609417 939829
rect 609473 939773 609559 939829
rect 609615 939773 609701 939829
rect 609757 939773 609843 939829
rect 609899 939773 609985 939829
rect 610041 939773 610127 939829
rect 610183 939773 610269 939829
rect 610325 939773 610411 939829
rect 610467 939773 610553 939829
rect 610609 939773 610695 939829
rect 610751 939773 610837 939829
rect 610893 939773 610979 939829
rect 611035 939773 611121 939829
rect 611177 939773 611248 939829
rect 609198 939720 611248 939773
rect 611828 941675 613728 941720
rect 611828 941619 611897 941675
rect 611953 941619 612039 941675
rect 612095 941619 612181 941675
rect 612237 941619 612323 941675
rect 612379 941619 612465 941675
rect 612521 941619 612607 941675
rect 612663 941619 612749 941675
rect 612805 941619 612891 941675
rect 612947 941619 613033 941675
rect 613089 941619 613175 941675
rect 613231 941619 613317 941675
rect 613373 941619 613459 941675
rect 613515 941619 613601 941675
rect 613657 941619 613728 941675
rect 611828 941533 613728 941619
rect 611828 941477 611897 941533
rect 611953 941477 612039 941533
rect 612095 941477 612181 941533
rect 612237 941477 612323 941533
rect 612379 941477 612465 941533
rect 612521 941477 612607 941533
rect 612663 941477 612749 941533
rect 612805 941477 612891 941533
rect 612947 941477 613033 941533
rect 613089 941477 613175 941533
rect 613231 941477 613317 941533
rect 613373 941477 613459 941533
rect 613515 941477 613601 941533
rect 613657 941477 613728 941533
rect 611828 941391 613728 941477
rect 611828 941335 611897 941391
rect 611953 941335 612039 941391
rect 612095 941335 612181 941391
rect 612237 941335 612323 941391
rect 612379 941335 612465 941391
rect 612521 941335 612607 941391
rect 612663 941335 612749 941391
rect 612805 941335 612891 941391
rect 612947 941335 613033 941391
rect 613089 941335 613175 941391
rect 613231 941335 613317 941391
rect 613373 941335 613459 941391
rect 613515 941335 613601 941391
rect 613657 941335 613728 941391
rect 611828 941249 613728 941335
rect 611828 941193 611897 941249
rect 611953 941193 612039 941249
rect 612095 941193 612181 941249
rect 612237 941193 612323 941249
rect 612379 941193 612465 941249
rect 612521 941193 612607 941249
rect 612663 941193 612749 941249
rect 612805 941193 612891 941249
rect 612947 941193 613033 941249
rect 613089 941193 613175 941249
rect 613231 941193 613317 941249
rect 613373 941193 613459 941249
rect 613515 941193 613601 941249
rect 613657 941193 613728 941249
rect 611828 941107 613728 941193
rect 611828 941051 611897 941107
rect 611953 941051 612039 941107
rect 612095 941051 612181 941107
rect 612237 941051 612323 941107
rect 612379 941051 612465 941107
rect 612521 941051 612607 941107
rect 612663 941051 612749 941107
rect 612805 941051 612891 941107
rect 612947 941051 613033 941107
rect 613089 941051 613175 941107
rect 613231 941051 613317 941107
rect 613373 941051 613459 941107
rect 613515 941051 613601 941107
rect 613657 941051 613728 941107
rect 611828 940965 613728 941051
rect 611828 940909 611897 940965
rect 611953 940909 612039 940965
rect 612095 940909 612181 940965
rect 612237 940909 612323 940965
rect 612379 940909 612465 940965
rect 612521 940909 612607 940965
rect 612663 940909 612749 940965
rect 612805 940909 612891 940965
rect 612947 940909 613033 940965
rect 613089 940909 613175 940965
rect 613231 940909 613317 940965
rect 613373 940909 613459 940965
rect 613515 940909 613601 940965
rect 613657 940909 613728 940965
rect 611828 940823 613728 940909
rect 611828 940767 611897 940823
rect 611953 940767 612039 940823
rect 612095 940767 612181 940823
rect 612237 940767 612323 940823
rect 612379 940767 612465 940823
rect 612521 940767 612607 940823
rect 612663 940767 612749 940823
rect 612805 940767 612891 940823
rect 612947 940767 613033 940823
rect 613089 940767 613175 940823
rect 613231 940767 613317 940823
rect 613373 940767 613459 940823
rect 613515 940767 613601 940823
rect 613657 940767 613728 940823
rect 611828 940681 613728 940767
rect 611828 940625 611897 940681
rect 611953 940625 612039 940681
rect 612095 940625 612181 940681
rect 612237 940625 612323 940681
rect 612379 940625 612465 940681
rect 612521 940625 612607 940681
rect 612663 940625 612749 940681
rect 612805 940625 612891 940681
rect 612947 940625 613033 940681
rect 613089 940625 613175 940681
rect 613231 940625 613317 940681
rect 613373 940625 613459 940681
rect 613515 940625 613601 940681
rect 613657 940625 613728 940681
rect 611828 940539 613728 940625
rect 611828 940483 611897 940539
rect 611953 940483 612039 940539
rect 612095 940483 612181 940539
rect 612237 940483 612323 940539
rect 612379 940483 612465 940539
rect 612521 940483 612607 940539
rect 612663 940483 612749 940539
rect 612805 940483 612891 940539
rect 612947 940483 613033 940539
rect 613089 940483 613175 940539
rect 613231 940483 613317 940539
rect 613373 940483 613459 940539
rect 613515 940483 613601 940539
rect 613657 940483 613728 940539
rect 611828 940397 613728 940483
rect 611828 940341 611897 940397
rect 611953 940341 612039 940397
rect 612095 940341 612181 940397
rect 612237 940341 612323 940397
rect 612379 940341 612465 940397
rect 612521 940341 612607 940397
rect 612663 940341 612749 940397
rect 612805 940341 612891 940397
rect 612947 940341 613033 940397
rect 613089 940341 613175 940397
rect 613231 940341 613317 940397
rect 613373 940341 613459 940397
rect 613515 940341 613601 940397
rect 613657 940341 613728 940397
rect 611828 940255 613728 940341
rect 611828 940199 611897 940255
rect 611953 940199 612039 940255
rect 612095 940199 612181 940255
rect 612237 940199 612323 940255
rect 612379 940199 612465 940255
rect 612521 940199 612607 940255
rect 612663 940199 612749 940255
rect 612805 940199 612891 940255
rect 612947 940199 613033 940255
rect 613089 940199 613175 940255
rect 613231 940199 613317 940255
rect 613373 940199 613459 940255
rect 613515 940199 613601 940255
rect 613657 940199 613728 940255
rect 611828 940113 613728 940199
rect 611828 940057 611897 940113
rect 611953 940057 612039 940113
rect 612095 940057 612181 940113
rect 612237 940057 612323 940113
rect 612379 940057 612465 940113
rect 612521 940057 612607 940113
rect 612663 940057 612749 940113
rect 612805 940057 612891 940113
rect 612947 940057 613033 940113
rect 613089 940057 613175 940113
rect 613231 940057 613317 940113
rect 613373 940057 613459 940113
rect 613515 940057 613601 940113
rect 613657 940057 613728 940113
rect 611828 939971 613728 940057
rect 611828 939915 611897 939971
rect 611953 939915 612039 939971
rect 612095 939915 612181 939971
rect 612237 939915 612323 939971
rect 612379 939915 612465 939971
rect 612521 939915 612607 939971
rect 612663 939915 612749 939971
rect 612805 939915 612891 939971
rect 612947 939915 613033 939971
rect 613089 939915 613175 939971
rect 613231 939915 613317 939971
rect 613373 939915 613459 939971
rect 613515 939915 613601 939971
rect 613657 939915 613728 939971
rect 611828 939829 613728 939915
rect 611828 939773 611897 939829
rect 611953 939773 612039 939829
rect 612095 939773 612181 939829
rect 612237 939773 612323 939829
rect 612379 939773 612465 939829
rect 612521 939773 612607 939829
rect 612663 939773 612749 939829
rect 612805 939773 612891 939829
rect 612947 939773 613033 939829
rect 613089 939773 613175 939829
rect 613231 939773 613317 939829
rect 613373 939773 613459 939829
rect 613515 939773 613601 939829
rect 613657 939773 613728 939829
rect 611828 939720 613728 939773
rect 655272 76035 656420 76088
rect 655272 75979 655343 76035
rect 655399 75979 655485 76035
rect 655541 75979 655627 76035
rect 655683 75979 655769 76035
rect 655825 75979 655911 76035
rect 655967 75979 656053 76035
rect 656109 75979 656195 76035
rect 656251 75979 656337 76035
rect 656393 75979 656420 76035
rect 655272 75893 656420 75979
rect 655272 75837 655343 75893
rect 655399 75837 655485 75893
rect 655541 75837 655627 75893
rect 655683 75837 655769 75893
rect 655825 75837 655911 75893
rect 655967 75837 656053 75893
rect 656109 75837 656195 75893
rect 656251 75837 656337 75893
rect 656393 75837 656420 75893
rect 655272 75751 656420 75837
rect 655272 75695 655343 75751
rect 655399 75695 655485 75751
rect 655541 75695 655627 75751
rect 655683 75695 655769 75751
rect 655825 75695 655911 75751
rect 655967 75695 656053 75751
rect 656109 75695 656195 75751
rect 656251 75695 656337 75751
rect 656393 75695 656420 75751
rect 655272 75609 656420 75695
rect 655272 75553 655343 75609
rect 655399 75553 655485 75609
rect 655541 75553 655627 75609
rect 655683 75553 655769 75609
rect 655825 75553 655911 75609
rect 655967 75553 656053 75609
rect 656109 75553 656195 75609
rect 656251 75553 656337 75609
rect 656393 75553 656420 75609
rect 655272 75467 656420 75553
rect 655272 75411 655343 75467
rect 655399 75411 655485 75467
rect 655541 75411 655627 75467
rect 655683 75411 655769 75467
rect 655825 75411 655911 75467
rect 655967 75411 656053 75467
rect 656109 75411 656195 75467
rect 656251 75411 656337 75467
rect 656393 75411 656420 75467
rect 655272 75325 656420 75411
rect 655272 75269 655343 75325
rect 655399 75269 655485 75325
rect 655541 75269 655627 75325
rect 655683 75269 655769 75325
rect 655825 75269 655911 75325
rect 655967 75269 656053 75325
rect 656109 75269 656195 75325
rect 656251 75269 656337 75325
rect 656393 75269 656420 75325
rect 655272 75183 656420 75269
rect 655272 75127 655343 75183
rect 655399 75127 655485 75183
rect 655541 75127 655627 75183
rect 655683 75127 655769 75183
rect 655825 75127 655911 75183
rect 655967 75127 656053 75183
rect 656109 75127 656195 75183
rect 656251 75127 656337 75183
rect 656393 75127 656420 75183
rect 655272 75041 656420 75127
rect 655272 74985 655343 75041
rect 655399 74985 655485 75041
rect 655541 74985 655627 75041
rect 655683 74985 655769 75041
rect 655825 74985 655911 75041
rect 655967 74985 656053 75041
rect 656109 74985 656195 75041
rect 656251 74985 656337 75041
rect 656393 74985 656420 75041
rect 655272 74899 656420 74985
rect 655272 74843 655343 74899
rect 655399 74843 655485 74899
rect 655541 74843 655627 74899
rect 655683 74843 655769 74899
rect 655825 74843 655911 74899
rect 655967 74843 656053 74899
rect 656109 74843 656195 74899
rect 656251 74843 656337 74899
rect 656393 74843 656420 74899
rect 655272 74757 656420 74843
rect 655272 74701 655343 74757
rect 655399 74701 655485 74757
rect 655541 74701 655627 74757
rect 655683 74701 655769 74757
rect 655825 74701 655911 74757
rect 655967 74701 656053 74757
rect 656109 74701 656195 74757
rect 656251 74701 656337 74757
rect 656393 74701 656420 74757
rect 655272 74615 656420 74701
rect 655272 74559 655343 74615
rect 655399 74559 655485 74615
rect 655541 74559 655627 74615
rect 655683 74559 655769 74615
rect 655825 74559 655911 74615
rect 655967 74559 656053 74615
rect 656109 74559 656195 74615
rect 656251 74559 656337 74615
rect 656393 74559 656420 74615
rect 655272 74488 656420 74559
rect 657752 76035 659802 76088
rect 657752 75979 657823 76035
rect 657879 75979 657965 76035
rect 658021 75979 658107 76035
rect 658163 75979 658249 76035
rect 658305 75979 658391 76035
rect 658447 75979 658533 76035
rect 658589 75979 658675 76035
rect 658731 75979 658817 76035
rect 658873 75979 658959 76035
rect 659015 75979 659101 76035
rect 659157 75979 659243 76035
rect 659299 75979 659385 76035
rect 659441 75979 659527 76035
rect 659583 75979 659669 76035
rect 659725 75979 659802 76035
rect 657752 75893 659802 75979
rect 657752 75837 657823 75893
rect 657879 75837 657965 75893
rect 658021 75837 658107 75893
rect 658163 75837 658249 75893
rect 658305 75837 658391 75893
rect 658447 75837 658533 75893
rect 658589 75837 658675 75893
rect 658731 75837 658817 75893
rect 658873 75837 658959 75893
rect 659015 75837 659101 75893
rect 659157 75837 659243 75893
rect 659299 75837 659385 75893
rect 659441 75837 659527 75893
rect 659583 75837 659669 75893
rect 659725 75837 659802 75893
rect 657752 75751 659802 75837
rect 657752 75695 657823 75751
rect 657879 75695 657965 75751
rect 658021 75695 658107 75751
rect 658163 75695 658249 75751
rect 658305 75695 658391 75751
rect 658447 75695 658533 75751
rect 658589 75695 658675 75751
rect 658731 75695 658817 75751
rect 658873 75695 658959 75751
rect 659015 75695 659101 75751
rect 659157 75695 659243 75751
rect 659299 75695 659385 75751
rect 659441 75695 659527 75751
rect 659583 75695 659669 75751
rect 659725 75695 659802 75751
rect 657752 75609 659802 75695
rect 657752 75553 657823 75609
rect 657879 75553 657965 75609
rect 658021 75553 658107 75609
rect 658163 75553 658249 75609
rect 658305 75553 658391 75609
rect 658447 75553 658533 75609
rect 658589 75553 658675 75609
rect 658731 75553 658817 75609
rect 658873 75553 658959 75609
rect 659015 75553 659101 75609
rect 659157 75553 659243 75609
rect 659299 75553 659385 75609
rect 659441 75553 659527 75609
rect 659583 75553 659669 75609
rect 659725 75553 659802 75609
rect 657752 75467 659802 75553
rect 657752 75411 657823 75467
rect 657879 75411 657965 75467
rect 658021 75411 658107 75467
rect 658163 75411 658249 75467
rect 658305 75411 658391 75467
rect 658447 75411 658533 75467
rect 658589 75411 658675 75467
rect 658731 75411 658817 75467
rect 658873 75411 658959 75467
rect 659015 75411 659101 75467
rect 659157 75411 659243 75467
rect 659299 75411 659385 75467
rect 659441 75411 659527 75467
rect 659583 75411 659669 75467
rect 659725 75411 659802 75467
rect 657752 75325 659802 75411
rect 657752 75269 657823 75325
rect 657879 75269 657965 75325
rect 658021 75269 658107 75325
rect 658163 75269 658249 75325
rect 658305 75269 658391 75325
rect 658447 75269 658533 75325
rect 658589 75269 658675 75325
rect 658731 75269 658817 75325
rect 658873 75269 658959 75325
rect 659015 75269 659101 75325
rect 659157 75269 659243 75325
rect 659299 75269 659385 75325
rect 659441 75269 659527 75325
rect 659583 75269 659669 75325
rect 659725 75269 659802 75325
rect 657752 75183 659802 75269
rect 657752 75127 657823 75183
rect 657879 75127 657965 75183
rect 658021 75127 658107 75183
rect 658163 75127 658249 75183
rect 658305 75127 658391 75183
rect 658447 75127 658533 75183
rect 658589 75127 658675 75183
rect 658731 75127 658817 75183
rect 658873 75127 658959 75183
rect 659015 75127 659101 75183
rect 659157 75127 659243 75183
rect 659299 75127 659385 75183
rect 659441 75127 659527 75183
rect 659583 75127 659669 75183
rect 659725 75127 659802 75183
rect 657752 75041 659802 75127
rect 657752 74985 657823 75041
rect 657879 74985 657965 75041
rect 658021 74985 658107 75041
rect 658163 74985 658249 75041
rect 658305 74985 658391 75041
rect 658447 74985 658533 75041
rect 658589 74985 658675 75041
rect 658731 74985 658817 75041
rect 658873 74985 658959 75041
rect 659015 74985 659101 75041
rect 659157 74985 659243 75041
rect 659299 74985 659385 75041
rect 659441 74985 659527 75041
rect 659583 74985 659669 75041
rect 659725 74985 659802 75041
rect 657752 74899 659802 74985
rect 657752 74843 657823 74899
rect 657879 74843 657965 74899
rect 658021 74843 658107 74899
rect 658163 74843 658249 74899
rect 658305 74843 658391 74899
rect 658447 74843 658533 74899
rect 658589 74843 658675 74899
rect 658731 74843 658817 74899
rect 658873 74843 658959 74899
rect 659015 74843 659101 74899
rect 659157 74843 659243 74899
rect 659299 74843 659385 74899
rect 659441 74843 659527 74899
rect 659583 74843 659669 74899
rect 659725 74843 659802 74899
rect 657752 74757 659802 74843
rect 657752 74701 657823 74757
rect 657879 74701 657965 74757
rect 658021 74701 658107 74757
rect 658163 74701 658249 74757
rect 658305 74701 658391 74757
rect 658447 74701 658533 74757
rect 658589 74701 658675 74757
rect 658731 74701 658817 74757
rect 658873 74701 658959 74757
rect 659015 74701 659101 74757
rect 659157 74701 659243 74757
rect 659299 74701 659385 74757
rect 659441 74701 659527 74757
rect 659583 74701 659669 74757
rect 659725 74701 659802 74757
rect 657752 74615 659802 74701
rect 657752 74559 657823 74615
rect 657879 74559 657965 74615
rect 658021 74559 658107 74615
rect 658163 74559 658249 74615
rect 658305 74559 658391 74615
rect 658447 74559 658533 74615
rect 658589 74559 658675 74615
rect 658731 74559 658817 74615
rect 658873 74559 658959 74615
rect 659015 74559 659101 74615
rect 659157 74559 659243 74615
rect 659299 74559 659385 74615
rect 659441 74559 659527 74615
rect 659583 74559 659669 74615
rect 659725 74559 659802 74615
rect 657752 74488 659802 74559
rect 660122 76035 662172 76088
rect 660122 75979 660193 76035
rect 660249 75979 660335 76035
rect 660391 75979 660477 76035
rect 660533 75979 660619 76035
rect 660675 75979 660761 76035
rect 660817 75979 660903 76035
rect 660959 75979 661045 76035
rect 661101 75979 661187 76035
rect 661243 75979 661329 76035
rect 661385 75979 661471 76035
rect 661527 75979 661613 76035
rect 661669 75979 661755 76035
rect 661811 75979 661897 76035
rect 661953 75979 662039 76035
rect 662095 75979 662172 76035
rect 660122 75893 662172 75979
rect 660122 75837 660193 75893
rect 660249 75837 660335 75893
rect 660391 75837 660477 75893
rect 660533 75837 660619 75893
rect 660675 75837 660761 75893
rect 660817 75837 660903 75893
rect 660959 75837 661045 75893
rect 661101 75837 661187 75893
rect 661243 75837 661329 75893
rect 661385 75837 661471 75893
rect 661527 75837 661613 75893
rect 661669 75837 661755 75893
rect 661811 75837 661897 75893
rect 661953 75837 662039 75893
rect 662095 75837 662172 75893
rect 660122 75751 662172 75837
rect 660122 75695 660193 75751
rect 660249 75695 660335 75751
rect 660391 75695 660477 75751
rect 660533 75695 660619 75751
rect 660675 75695 660761 75751
rect 660817 75695 660903 75751
rect 660959 75695 661045 75751
rect 661101 75695 661187 75751
rect 661243 75695 661329 75751
rect 661385 75695 661471 75751
rect 661527 75695 661613 75751
rect 661669 75695 661755 75751
rect 661811 75695 661897 75751
rect 661953 75695 662039 75751
rect 662095 75695 662172 75751
rect 660122 75609 662172 75695
rect 660122 75553 660193 75609
rect 660249 75553 660335 75609
rect 660391 75553 660477 75609
rect 660533 75553 660619 75609
rect 660675 75553 660761 75609
rect 660817 75553 660903 75609
rect 660959 75553 661045 75609
rect 661101 75553 661187 75609
rect 661243 75553 661329 75609
rect 661385 75553 661471 75609
rect 661527 75553 661613 75609
rect 661669 75553 661755 75609
rect 661811 75553 661897 75609
rect 661953 75553 662039 75609
rect 662095 75553 662172 75609
rect 660122 75467 662172 75553
rect 660122 75411 660193 75467
rect 660249 75411 660335 75467
rect 660391 75411 660477 75467
rect 660533 75411 660619 75467
rect 660675 75411 660761 75467
rect 660817 75411 660903 75467
rect 660959 75411 661045 75467
rect 661101 75411 661187 75467
rect 661243 75411 661329 75467
rect 661385 75411 661471 75467
rect 661527 75411 661613 75467
rect 661669 75411 661755 75467
rect 661811 75411 661897 75467
rect 661953 75411 662039 75467
rect 662095 75411 662172 75467
rect 660122 75325 662172 75411
rect 660122 75269 660193 75325
rect 660249 75269 660335 75325
rect 660391 75269 660477 75325
rect 660533 75269 660619 75325
rect 660675 75269 660761 75325
rect 660817 75269 660903 75325
rect 660959 75269 661045 75325
rect 661101 75269 661187 75325
rect 661243 75269 661329 75325
rect 661385 75269 661471 75325
rect 661527 75269 661613 75325
rect 661669 75269 661755 75325
rect 661811 75269 661897 75325
rect 661953 75269 662039 75325
rect 662095 75269 662172 75325
rect 660122 75183 662172 75269
rect 660122 75127 660193 75183
rect 660249 75127 660335 75183
rect 660391 75127 660477 75183
rect 660533 75127 660619 75183
rect 660675 75127 660761 75183
rect 660817 75127 660903 75183
rect 660959 75127 661045 75183
rect 661101 75127 661187 75183
rect 661243 75127 661329 75183
rect 661385 75127 661471 75183
rect 661527 75127 661613 75183
rect 661669 75127 661755 75183
rect 661811 75127 661897 75183
rect 661953 75127 662039 75183
rect 662095 75127 662172 75183
rect 660122 75041 662172 75127
rect 660122 74985 660193 75041
rect 660249 74985 660335 75041
rect 660391 74985 660477 75041
rect 660533 74985 660619 75041
rect 660675 74985 660761 75041
rect 660817 74985 660903 75041
rect 660959 74985 661045 75041
rect 661101 74985 661187 75041
rect 661243 74985 661329 75041
rect 661385 74985 661471 75041
rect 661527 74985 661613 75041
rect 661669 74985 661755 75041
rect 661811 74985 661897 75041
rect 661953 74985 662039 75041
rect 662095 74985 662172 75041
rect 660122 74899 662172 74985
rect 660122 74843 660193 74899
rect 660249 74843 660335 74899
rect 660391 74843 660477 74899
rect 660533 74843 660619 74899
rect 660675 74843 660761 74899
rect 660817 74843 660903 74899
rect 660959 74843 661045 74899
rect 661101 74843 661187 74899
rect 661243 74843 661329 74899
rect 661385 74843 661471 74899
rect 661527 74843 661613 74899
rect 661669 74843 661755 74899
rect 661811 74843 661897 74899
rect 661953 74843 662039 74899
rect 662095 74843 662172 74899
rect 660122 74757 662172 74843
rect 660122 74701 660193 74757
rect 660249 74701 660335 74757
rect 660391 74701 660477 74757
rect 660533 74701 660619 74757
rect 660675 74701 660761 74757
rect 660817 74701 660903 74757
rect 660959 74701 661045 74757
rect 661101 74701 661187 74757
rect 661243 74701 661329 74757
rect 661385 74701 661471 74757
rect 661527 74701 661613 74757
rect 661669 74701 661755 74757
rect 661811 74701 661897 74757
rect 661953 74701 662039 74757
rect 662095 74701 662172 74757
rect 660122 74615 662172 74701
rect 660122 74559 660193 74615
rect 660249 74559 660335 74615
rect 660391 74559 660477 74615
rect 660533 74559 660619 74615
rect 660675 74559 660761 74615
rect 660817 74559 660903 74615
rect 660959 74559 661045 74615
rect 661101 74559 661187 74615
rect 661243 74559 661329 74615
rect 661385 74559 661471 74615
rect 661527 74559 661613 74615
rect 661669 74559 661755 74615
rect 661811 74559 661897 74615
rect 661953 74559 662039 74615
rect 662095 74559 662172 74615
rect 660122 74488 662172 74559
rect 662828 76035 664878 76088
rect 662828 75979 662899 76035
rect 662955 75979 663041 76035
rect 663097 75979 663183 76035
rect 663239 75979 663325 76035
rect 663381 75979 663467 76035
rect 663523 75979 663609 76035
rect 663665 75979 663751 76035
rect 663807 75979 663893 76035
rect 663949 75979 664035 76035
rect 664091 75979 664177 76035
rect 664233 75979 664319 76035
rect 664375 75979 664461 76035
rect 664517 75979 664603 76035
rect 664659 75979 664745 76035
rect 664801 75979 664878 76035
rect 662828 75893 664878 75979
rect 662828 75837 662899 75893
rect 662955 75837 663041 75893
rect 663097 75837 663183 75893
rect 663239 75837 663325 75893
rect 663381 75837 663467 75893
rect 663523 75837 663609 75893
rect 663665 75837 663751 75893
rect 663807 75837 663893 75893
rect 663949 75837 664035 75893
rect 664091 75837 664177 75893
rect 664233 75837 664319 75893
rect 664375 75837 664461 75893
rect 664517 75837 664603 75893
rect 664659 75837 664745 75893
rect 664801 75837 664878 75893
rect 662828 75751 664878 75837
rect 662828 75695 662899 75751
rect 662955 75695 663041 75751
rect 663097 75695 663183 75751
rect 663239 75695 663325 75751
rect 663381 75695 663467 75751
rect 663523 75695 663609 75751
rect 663665 75695 663751 75751
rect 663807 75695 663893 75751
rect 663949 75695 664035 75751
rect 664091 75695 664177 75751
rect 664233 75695 664319 75751
rect 664375 75695 664461 75751
rect 664517 75695 664603 75751
rect 664659 75695 664745 75751
rect 664801 75695 664878 75751
rect 662828 75609 664878 75695
rect 662828 75553 662899 75609
rect 662955 75553 663041 75609
rect 663097 75553 663183 75609
rect 663239 75553 663325 75609
rect 663381 75553 663467 75609
rect 663523 75553 663609 75609
rect 663665 75553 663751 75609
rect 663807 75553 663893 75609
rect 663949 75553 664035 75609
rect 664091 75553 664177 75609
rect 664233 75553 664319 75609
rect 664375 75553 664461 75609
rect 664517 75553 664603 75609
rect 664659 75553 664745 75609
rect 664801 75553 664878 75609
rect 662828 75467 664878 75553
rect 662828 75411 662899 75467
rect 662955 75411 663041 75467
rect 663097 75411 663183 75467
rect 663239 75411 663325 75467
rect 663381 75411 663467 75467
rect 663523 75411 663609 75467
rect 663665 75411 663751 75467
rect 663807 75411 663893 75467
rect 663949 75411 664035 75467
rect 664091 75411 664177 75467
rect 664233 75411 664319 75467
rect 664375 75411 664461 75467
rect 664517 75411 664603 75467
rect 664659 75411 664745 75467
rect 664801 75411 664878 75467
rect 662828 75325 664878 75411
rect 662828 75269 662899 75325
rect 662955 75269 663041 75325
rect 663097 75269 663183 75325
rect 663239 75269 663325 75325
rect 663381 75269 663467 75325
rect 663523 75269 663609 75325
rect 663665 75269 663751 75325
rect 663807 75269 663893 75325
rect 663949 75269 664035 75325
rect 664091 75269 664177 75325
rect 664233 75269 664319 75325
rect 664375 75269 664461 75325
rect 664517 75269 664603 75325
rect 664659 75269 664745 75325
rect 664801 75269 664878 75325
rect 662828 75183 664878 75269
rect 662828 75127 662899 75183
rect 662955 75127 663041 75183
rect 663097 75127 663183 75183
rect 663239 75127 663325 75183
rect 663381 75127 663467 75183
rect 663523 75127 663609 75183
rect 663665 75127 663751 75183
rect 663807 75127 663893 75183
rect 663949 75127 664035 75183
rect 664091 75127 664177 75183
rect 664233 75127 664319 75183
rect 664375 75127 664461 75183
rect 664517 75127 664603 75183
rect 664659 75127 664745 75183
rect 664801 75127 664878 75183
rect 662828 75041 664878 75127
rect 662828 74985 662899 75041
rect 662955 74985 663041 75041
rect 663097 74985 663183 75041
rect 663239 74985 663325 75041
rect 663381 74985 663467 75041
rect 663523 74985 663609 75041
rect 663665 74985 663751 75041
rect 663807 74985 663893 75041
rect 663949 74985 664035 75041
rect 664091 74985 664177 75041
rect 664233 74985 664319 75041
rect 664375 74985 664461 75041
rect 664517 74985 664603 75041
rect 664659 74985 664745 75041
rect 664801 74985 664878 75041
rect 662828 74899 664878 74985
rect 662828 74843 662899 74899
rect 662955 74843 663041 74899
rect 663097 74843 663183 74899
rect 663239 74843 663325 74899
rect 663381 74843 663467 74899
rect 663523 74843 663609 74899
rect 663665 74843 663751 74899
rect 663807 74843 663893 74899
rect 663949 74843 664035 74899
rect 664091 74843 664177 74899
rect 664233 74843 664319 74899
rect 664375 74843 664461 74899
rect 664517 74843 664603 74899
rect 664659 74843 664745 74899
rect 664801 74843 664878 74899
rect 662828 74757 664878 74843
rect 662828 74701 662899 74757
rect 662955 74701 663041 74757
rect 663097 74701 663183 74757
rect 663239 74701 663325 74757
rect 663381 74701 663467 74757
rect 663523 74701 663609 74757
rect 663665 74701 663751 74757
rect 663807 74701 663893 74757
rect 663949 74701 664035 74757
rect 664091 74701 664177 74757
rect 664233 74701 664319 74757
rect 664375 74701 664461 74757
rect 664517 74701 664603 74757
rect 664659 74701 664745 74757
rect 664801 74701 664878 74757
rect 662828 74615 664878 74701
rect 662828 74559 662899 74615
rect 662955 74559 663041 74615
rect 663097 74559 663183 74615
rect 663239 74559 663325 74615
rect 663381 74559 663467 74615
rect 663523 74559 663609 74615
rect 663665 74559 663751 74615
rect 663807 74559 663893 74615
rect 663949 74559 664035 74615
rect 664091 74559 664177 74615
rect 664233 74559 664319 74615
rect 664375 74559 664461 74615
rect 664517 74559 664603 74615
rect 664659 74559 664745 74615
rect 664801 74559 664878 74615
rect 662828 74488 664878 74559
rect 665198 76035 667248 76088
rect 665198 75979 665269 76035
rect 665325 75979 665411 76035
rect 665467 75979 665553 76035
rect 665609 75979 665695 76035
rect 665751 75979 665837 76035
rect 665893 75979 665979 76035
rect 666035 75979 666121 76035
rect 666177 75979 666263 76035
rect 666319 75979 666405 76035
rect 666461 75979 666547 76035
rect 666603 75979 666689 76035
rect 666745 75979 666831 76035
rect 666887 75979 666973 76035
rect 667029 75979 667115 76035
rect 667171 75979 667248 76035
rect 665198 75893 667248 75979
rect 665198 75837 665269 75893
rect 665325 75837 665411 75893
rect 665467 75837 665553 75893
rect 665609 75837 665695 75893
rect 665751 75837 665837 75893
rect 665893 75837 665979 75893
rect 666035 75837 666121 75893
rect 666177 75837 666263 75893
rect 666319 75837 666405 75893
rect 666461 75837 666547 75893
rect 666603 75837 666689 75893
rect 666745 75837 666831 75893
rect 666887 75837 666973 75893
rect 667029 75837 667115 75893
rect 667171 75837 667248 75893
rect 665198 75751 667248 75837
rect 665198 75695 665269 75751
rect 665325 75695 665411 75751
rect 665467 75695 665553 75751
rect 665609 75695 665695 75751
rect 665751 75695 665837 75751
rect 665893 75695 665979 75751
rect 666035 75695 666121 75751
rect 666177 75695 666263 75751
rect 666319 75695 666405 75751
rect 666461 75695 666547 75751
rect 666603 75695 666689 75751
rect 666745 75695 666831 75751
rect 666887 75695 666973 75751
rect 667029 75695 667115 75751
rect 667171 75695 667248 75751
rect 665198 75609 667248 75695
rect 665198 75553 665269 75609
rect 665325 75553 665411 75609
rect 665467 75553 665553 75609
rect 665609 75553 665695 75609
rect 665751 75553 665837 75609
rect 665893 75553 665979 75609
rect 666035 75553 666121 75609
rect 666177 75553 666263 75609
rect 666319 75553 666405 75609
rect 666461 75553 666547 75609
rect 666603 75553 666689 75609
rect 666745 75553 666831 75609
rect 666887 75553 666973 75609
rect 667029 75553 667115 75609
rect 667171 75553 667248 75609
rect 665198 75467 667248 75553
rect 665198 75411 665269 75467
rect 665325 75411 665411 75467
rect 665467 75411 665553 75467
rect 665609 75411 665695 75467
rect 665751 75411 665837 75467
rect 665893 75411 665979 75467
rect 666035 75411 666121 75467
rect 666177 75411 666263 75467
rect 666319 75411 666405 75467
rect 666461 75411 666547 75467
rect 666603 75411 666689 75467
rect 666745 75411 666831 75467
rect 666887 75411 666973 75467
rect 667029 75411 667115 75467
rect 667171 75411 667248 75467
rect 665198 75325 667248 75411
rect 665198 75269 665269 75325
rect 665325 75269 665411 75325
rect 665467 75269 665553 75325
rect 665609 75269 665695 75325
rect 665751 75269 665837 75325
rect 665893 75269 665979 75325
rect 666035 75269 666121 75325
rect 666177 75269 666263 75325
rect 666319 75269 666405 75325
rect 666461 75269 666547 75325
rect 666603 75269 666689 75325
rect 666745 75269 666831 75325
rect 666887 75269 666973 75325
rect 667029 75269 667115 75325
rect 667171 75269 667248 75325
rect 665198 75183 667248 75269
rect 665198 75127 665269 75183
rect 665325 75127 665411 75183
rect 665467 75127 665553 75183
rect 665609 75127 665695 75183
rect 665751 75127 665837 75183
rect 665893 75127 665979 75183
rect 666035 75127 666121 75183
rect 666177 75127 666263 75183
rect 666319 75127 666405 75183
rect 666461 75127 666547 75183
rect 666603 75127 666689 75183
rect 666745 75127 666831 75183
rect 666887 75127 666973 75183
rect 667029 75127 667115 75183
rect 667171 75127 667248 75183
rect 665198 75041 667248 75127
rect 665198 74985 665269 75041
rect 665325 74985 665411 75041
rect 665467 74985 665553 75041
rect 665609 74985 665695 75041
rect 665751 74985 665837 75041
rect 665893 74985 665979 75041
rect 666035 74985 666121 75041
rect 666177 74985 666263 75041
rect 666319 74985 666405 75041
rect 666461 74985 666547 75041
rect 666603 74985 666689 75041
rect 666745 74985 666831 75041
rect 666887 74985 666973 75041
rect 667029 74985 667115 75041
rect 667171 74985 667248 75041
rect 665198 74899 667248 74985
rect 665198 74843 665269 74899
rect 665325 74843 665411 74899
rect 665467 74843 665553 74899
rect 665609 74843 665695 74899
rect 665751 74843 665837 74899
rect 665893 74843 665979 74899
rect 666035 74843 666121 74899
rect 666177 74843 666263 74899
rect 666319 74843 666405 74899
rect 666461 74843 666547 74899
rect 666603 74843 666689 74899
rect 666745 74843 666831 74899
rect 666887 74843 666973 74899
rect 667029 74843 667115 74899
rect 667171 74843 667248 74899
rect 665198 74757 667248 74843
rect 665198 74701 665269 74757
rect 665325 74701 665411 74757
rect 665467 74701 665553 74757
rect 665609 74701 665695 74757
rect 665751 74701 665837 74757
rect 665893 74701 665979 74757
rect 666035 74701 666121 74757
rect 666177 74701 666263 74757
rect 666319 74701 666405 74757
rect 666461 74701 666547 74757
rect 666603 74701 666689 74757
rect 666745 74701 666831 74757
rect 666887 74701 666973 74757
rect 667029 74701 667115 74757
rect 667171 74701 667248 74757
rect 665198 74615 667248 74701
rect 665198 74559 665269 74615
rect 665325 74559 665411 74615
rect 665467 74559 665553 74615
rect 665609 74559 665695 74615
rect 665751 74559 665837 74615
rect 665893 74559 665979 74615
rect 666035 74559 666121 74615
rect 666177 74559 666263 74615
rect 666319 74559 666405 74615
rect 666461 74559 666547 74615
rect 666603 74559 666689 74615
rect 666745 74559 666831 74615
rect 666887 74559 666973 74615
rect 667029 74559 667115 74615
rect 667171 74559 667248 74615
rect 665198 74488 667248 74559
rect 667828 76035 669728 76088
rect 667828 75979 667899 76035
rect 667955 75979 668041 76035
rect 668097 75979 668183 76035
rect 668239 75979 668325 76035
rect 668381 75979 668467 76035
rect 668523 75979 668609 76035
rect 668665 75979 668751 76035
rect 668807 75979 668893 76035
rect 668949 75979 669035 76035
rect 669091 75979 669177 76035
rect 669233 75979 669319 76035
rect 669375 75979 669461 76035
rect 669517 75979 669603 76035
rect 669659 75979 669728 76035
rect 667828 75893 669728 75979
rect 667828 75837 667899 75893
rect 667955 75837 668041 75893
rect 668097 75837 668183 75893
rect 668239 75837 668325 75893
rect 668381 75837 668467 75893
rect 668523 75837 668609 75893
rect 668665 75837 668751 75893
rect 668807 75837 668893 75893
rect 668949 75837 669035 75893
rect 669091 75837 669177 75893
rect 669233 75837 669319 75893
rect 669375 75837 669461 75893
rect 669517 75837 669603 75893
rect 669659 75837 669728 75893
rect 667828 75751 669728 75837
rect 667828 75695 667899 75751
rect 667955 75695 668041 75751
rect 668097 75695 668183 75751
rect 668239 75695 668325 75751
rect 668381 75695 668467 75751
rect 668523 75695 668609 75751
rect 668665 75695 668751 75751
rect 668807 75695 668893 75751
rect 668949 75695 669035 75751
rect 669091 75695 669177 75751
rect 669233 75695 669319 75751
rect 669375 75695 669461 75751
rect 669517 75695 669603 75751
rect 669659 75695 669728 75751
rect 667828 75609 669728 75695
rect 667828 75553 667899 75609
rect 667955 75553 668041 75609
rect 668097 75553 668183 75609
rect 668239 75553 668325 75609
rect 668381 75553 668467 75609
rect 668523 75553 668609 75609
rect 668665 75553 668751 75609
rect 668807 75553 668893 75609
rect 668949 75553 669035 75609
rect 669091 75553 669177 75609
rect 669233 75553 669319 75609
rect 669375 75553 669461 75609
rect 669517 75553 669603 75609
rect 669659 75553 669728 75609
rect 667828 75467 669728 75553
rect 667828 75411 667899 75467
rect 667955 75411 668041 75467
rect 668097 75411 668183 75467
rect 668239 75411 668325 75467
rect 668381 75411 668467 75467
rect 668523 75411 668609 75467
rect 668665 75411 668751 75467
rect 668807 75411 668893 75467
rect 668949 75411 669035 75467
rect 669091 75411 669177 75467
rect 669233 75411 669319 75467
rect 669375 75411 669461 75467
rect 669517 75411 669603 75467
rect 669659 75411 669728 75467
rect 667828 75325 669728 75411
rect 667828 75269 667899 75325
rect 667955 75269 668041 75325
rect 668097 75269 668183 75325
rect 668239 75269 668325 75325
rect 668381 75269 668467 75325
rect 668523 75269 668609 75325
rect 668665 75269 668751 75325
rect 668807 75269 668893 75325
rect 668949 75269 669035 75325
rect 669091 75269 669177 75325
rect 669233 75269 669319 75325
rect 669375 75269 669461 75325
rect 669517 75269 669603 75325
rect 669659 75269 669728 75325
rect 667828 75183 669728 75269
rect 667828 75127 667899 75183
rect 667955 75127 668041 75183
rect 668097 75127 668183 75183
rect 668239 75127 668325 75183
rect 668381 75127 668467 75183
rect 668523 75127 668609 75183
rect 668665 75127 668751 75183
rect 668807 75127 668893 75183
rect 668949 75127 669035 75183
rect 669091 75127 669177 75183
rect 669233 75127 669319 75183
rect 669375 75127 669461 75183
rect 669517 75127 669603 75183
rect 669659 75127 669728 75183
rect 667828 75041 669728 75127
rect 667828 74985 667899 75041
rect 667955 74985 668041 75041
rect 668097 74985 668183 75041
rect 668239 74985 668325 75041
rect 668381 74985 668467 75041
rect 668523 74985 668609 75041
rect 668665 74985 668751 75041
rect 668807 74985 668893 75041
rect 668949 74985 669035 75041
rect 669091 74985 669177 75041
rect 669233 74985 669319 75041
rect 669375 74985 669461 75041
rect 669517 74985 669603 75041
rect 669659 74985 669728 75041
rect 667828 74899 669728 74985
rect 667828 74843 667899 74899
rect 667955 74843 668041 74899
rect 668097 74843 668183 74899
rect 668239 74843 668325 74899
rect 668381 74843 668467 74899
rect 668523 74843 668609 74899
rect 668665 74843 668751 74899
rect 668807 74843 668893 74899
rect 668949 74843 669035 74899
rect 669091 74843 669177 74899
rect 669233 74843 669319 74899
rect 669375 74843 669461 74899
rect 669517 74843 669603 74899
rect 669659 74843 669728 74899
rect 667828 74757 669728 74843
rect 667828 74701 667899 74757
rect 667955 74701 668041 74757
rect 668097 74701 668183 74757
rect 668239 74701 668325 74757
rect 668381 74701 668467 74757
rect 668523 74701 668609 74757
rect 668665 74701 668751 74757
rect 668807 74701 668893 74757
rect 668949 74701 669035 74757
rect 669091 74701 669177 74757
rect 669233 74701 669319 74757
rect 669375 74701 669461 74757
rect 669517 74701 669603 74757
rect 669659 74701 669728 74757
rect 667828 74615 669728 74701
rect 667828 74559 667899 74615
rect 667955 74559 668041 74615
rect 668097 74559 668183 74615
rect 668239 74559 668325 74615
rect 668381 74559 668467 74615
rect 668523 74559 668609 74615
rect 668665 74559 668751 74615
rect 668807 74559 668893 74615
rect 668949 74559 669035 74615
rect 669091 74559 669177 74615
rect 669233 74559 669319 74615
rect 669375 74559 669461 74615
rect 669517 74559 669603 74615
rect 669659 74559 669728 74615
rect 667828 74488 669728 74559
rect 105272 74035 107172 74088
rect 105272 73979 105343 74035
rect 105399 73979 105485 74035
rect 105541 73979 105627 74035
rect 105683 73979 105769 74035
rect 105825 73979 105911 74035
rect 105967 73979 106053 74035
rect 106109 73979 106195 74035
rect 106251 73979 106337 74035
rect 106393 73979 106479 74035
rect 106535 73979 106621 74035
rect 106677 73979 106763 74035
rect 106819 73979 106905 74035
rect 106961 73979 107047 74035
rect 107103 73979 107172 74035
rect 105272 73893 107172 73979
rect 105272 73837 105343 73893
rect 105399 73837 105485 73893
rect 105541 73837 105627 73893
rect 105683 73837 105769 73893
rect 105825 73837 105911 73893
rect 105967 73837 106053 73893
rect 106109 73837 106195 73893
rect 106251 73837 106337 73893
rect 106393 73837 106479 73893
rect 106535 73837 106621 73893
rect 106677 73837 106763 73893
rect 106819 73837 106905 73893
rect 106961 73837 107047 73893
rect 107103 73837 107172 73893
rect 105272 73751 107172 73837
rect 105272 73695 105343 73751
rect 105399 73695 105485 73751
rect 105541 73695 105627 73751
rect 105683 73695 105769 73751
rect 105825 73695 105911 73751
rect 105967 73695 106053 73751
rect 106109 73695 106195 73751
rect 106251 73695 106337 73751
rect 106393 73695 106479 73751
rect 106535 73695 106621 73751
rect 106677 73695 106763 73751
rect 106819 73695 106905 73751
rect 106961 73695 107047 73751
rect 107103 73695 107172 73751
rect 105272 73609 107172 73695
rect 105272 73553 105343 73609
rect 105399 73553 105485 73609
rect 105541 73553 105627 73609
rect 105683 73553 105769 73609
rect 105825 73553 105911 73609
rect 105967 73553 106053 73609
rect 106109 73553 106195 73609
rect 106251 73553 106337 73609
rect 106393 73553 106479 73609
rect 106535 73553 106621 73609
rect 106677 73553 106763 73609
rect 106819 73553 106905 73609
rect 106961 73553 107047 73609
rect 107103 73553 107172 73609
rect 105272 73467 107172 73553
rect 105272 73411 105343 73467
rect 105399 73411 105485 73467
rect 105541 73411 105627 73467
rect 105683 73411 105769 73467
rect 105825 73411 105911 73467
rect 105967 73411 106053 73467
rect 106109 73411 106195 73467
rect 106251 73411 106337 73467
rect 106393 73411 106479 73467
rect 106535 73411 106621 73467
rect 106677 73411 106763 73467
rect 106819 73411 106905 73467
rect 106961 73411 107047 73467
rect 107103 73411 107172 73467
rect 105272 73325 107172 73411
rect 105272 73269 105343 73325
rect 105399 73269 105485 73325
rect 105541 73269 105627 73325
rect 105683 73269 105769 73325
rect 105825 73269 105911 73325
rect 105967 73269 106053 73325
rect 106109 73269 106195 73325
rect 106251 73269 106337 73325
rect 106393 73269 106479 73325
rect 106535 73269 106621 73325
rect 106677 73269 106763 73325
rect 106819 73269 106905 73325
rect 106961 73269 107047 73325
rect 107103 73269 107172 73325
rect 105272 73183 107172 73269
rect 105272 73127 105343 73183
rect 105399 73127 105485 73183
rect 105541 73127 105627 73183
rect 105683 73127 105769 73183
rect 105825 73127 105911 73183
rect 105967 73127 106053 73183
rect 106109 73127 106195 73183
rect 106251 73127 106337 73183
rect 106393 73127 106479 73183
rect 106535 73127 106621 73183
rect 106677 73127 106763 73183
rect 106819 73127 106905 73183
rect 106961 73127 107047 73183
rect 107103 73127 107172 73183
rect 105272 73041 107172 73127
rect 105272 72985 105343 73041
rect 105399 72985 105485 73041
rect 105541 72985 105627 73041
rect 105683 72985 105769 73041
rect 105825 72985 105911 73041
rect 105967 72985 106053 73041
rect 106109 72985 106195 73041
rect 106251 72985 106337 73041
rect 106393 72985 106479 73041
rect 106535 72985 106621 73041
rect 106677 72985 106763 73041
rect 106819 72985 106905 73041
rect 106961 72985 107047 73041
rect 107103 72985 107172 73041
rect 105272 72899 107172 72985
rect 105272 72843 105343 72899
rect 105399 72843 105485 72899
rect 105541 72843 105627 72899
rect 105683 72843 105769 72899
rect 105825 72843 105911 72899
rect 105967 72843 106053 72899
rect 106109 72843 106195 72899
rect 106251 72843 106337 72899
rect 106393 72843 106479 72899
rect 106535 72843 106621 72899
rect 106677 72843 106763 72899
rect 106819 72843 106905 72899
rect 106961 72843 107047 72899
rect 107103 72843 107172 72899
rect 105272 72757 107172 72843
rect 105272 72701 105343 72757
rect 105399 72701 105485 72757
rect 105541 72701 105627 72757
rect 105683 72701 105769 72757
rect 105825 72701 105911 72757
rect 105967 72701 106053 72757
rect 106109 72701 106195 72757
rect 106251 72701 106337 72757
rect 106393 72701 106479 72757
rect 106535 72701 106621 72757
rect 106677 72701 106763 72757
rect 106819 72701 106905 72757
rect 106961 72701 107047 72757
rect 107103 72701 107172 72757
rect 105272 72615 107172 72701
rect 105272 72559 105343 72615
rect 105399 72559 105485 72615
rect 105541 72559 105627 72615
rect 105683 72559 105769 72615
rect 105825 72559 105911 72615
rect 105967 72559 106053 72615
rect 106109 72559 106195 72615
rect 106251 72559 106337 72615
rect 106393 72559 106479 72615
rect 106535 72559 106621 72615
rect 106677 72559 106763 72615
rect 106819 72559 106905 72615
rect 106961 72559 107047 72615
rect 107103 72559 107172 72615
rect 105272 72473 107172 72559
rect 105272 72417 105343 72473
rect 105399 72417 105485 72473
rect 105541 72417 105627 72473
rect 105683 72417 105769 72473
rect 105825 72417 105911 72473
rect 105967 72417 106053 72473
rect 106109 72417 106195 72473
rect 106251 72417 106337 72473
rect 106393 72417 106479 72473
rect 106535 72417 106621 72473
rect 106677 72417 106763 72473
rect 106819 72417 106905 72473
rect 106961 72417 107047 72473
rect 107103 72417 107172 72473
rect 105272 72331 107172 72417
rect 105272 72275 105343 72331
rect 105399 72275 105485 72331
rect 105541 72275 105627 72331
rect 105683 72275 105769 72331
rect 105825 72275 105911 72331
rect 105967 72275 106053 72331
rect 106109 72275 106195 72331
rect 106251 72275 106337 72331
rect 106393 72275 106479 72331
rect 106535 72275 106621 72331
rect 106677 72275 106763 72331
rect 106819 72275 106905 72331
rect 106961 72275 107047 72331
rect 107103 72275 107172 72331
rect 105272 72189 107172 72275
rect 105272 72133 105343 72189
rect 105399 72133 105485 72189
rect 105541 72133 105627 72189
rect 105683 72133 105769 72189
rect 105825 72133 105911 72189
rect 105967 72133 106053 72189
rect 106109 72133 106195 72189
rect 106251 72133 106337 72189
rect 106393 72133 106479 72189
rect 106535 72133 106621 72189
rect 106677 72133 106763 72189
rect 106819 72133 106905 72189
rect 106961 72133 107047 72189
rect 107103 72133 107172 72189
rect 105272 72088 107172 72133
rect 108948 74035 109802 74088
rect 108948 73979 108995 74035
rect 109051 73979 109137 74035
rect 109193 73979 109279 74035
rect 109335 73979 109421 74035
rect 109477 73979 109563 74035
rect 109619 73979 109705 74035
rect 109761 73979 109802 74035
rect 108948 73893 109802 73979
rect 108948 73837 108995 73893
rect 109051 73837 109137 73893
rect 109193 73837 109279 73893
rect 109335 73837 109421 73893
rect 109477 73837 109563 73893
rect 109619 73837 109705 73893
rect 109761 73837 109802 73893
rect 108948 73751 109802 73837
rect 108948 73695 108995 73751
rect 109051 73695 109137 73751
rect 109193 73695 109279 73751
rect 109335 73695 109421 73751
rect 109477 73695 109563 73751
rect 109619 73695 109705 73751
rect 109761 73695 109802 73751
rect 108948 73609 109802 73695
rect 108948 73553 108995 73609
rect 109051 73553 109137 73609
rect 109193 73553 109279 73609
rect 109335 73553 109421 73609
rect 109477 73553 109563 73609
rect 109619 73553 109705 73609
rect 109761 73553 109802 73609
rect 108948 73467 109802 73553
rect 108948 73411 108995 73467
rect 109051 73411 109137 73467
rect 109193 73411 109279 73467
rect 109335 73411 109421 73467
rect 109477 73411 109563 73467
rect 109619 73411 109705 73467
rect 109761 73411 109802 73467
rect 108948 73325 109802 73411
rect 108948 73269 108995 73325
rect 109051 73269 109137 73325
rect 109193 73269 109279 73325
rect 109335 73269 109421 73325
rect 109477 73269 109563 73325
rect 109619 73269 109705 73325
rect 109761 73269 109802 73325
rect 108948 73183 109802 73269
rect 108948 73127 108995 73183
rect 109051 73127 109137 73183
rect 109193 73127 109279 73183
rect 109335 73127 109421 73183
rect 109477 73127 109563 73183
rect 109619 73127 109705 73183
rect 109761 73127 109802 73183
rect 108948 73041 109802 73127
rect 108948 72985 108995 73041
rect 109051 72985 109137 73041
rect 109193 72985 109279 73041
rect 109335 72985 109421 73041
rect 109477 72985 109563 73041
rect 109619 72985 109705 73041
rect 109761 72985 109802 73041
rect 108948 72899 109802 72985
rect 108948 72843 108995 72899
rect 109051 72843 109137 72899
rect 109193 72843 109279 72899
rect 109335 72843 109421 72899
rect 109477 72843 109563 72899
rect 109619 72843 109705 72899
rect 109761 72843 109802 72899
rect 108948 72757 109802 72843
rect 108948 72701 108995 72757
rect 109051 72701 109137 72757
rect 109193 72701 109279 72757
rect 109335 72701 109421 72757
rect 109477 72701 109563 72757
rect 109619 72701 109705 72757
rect 109761 72701 109802 72757
rect 108948 72615 109802 72701
rect 108948 72559 108995 72615
rect 109051 72559 109137 72615
rect 109193 72559 109279 72615
rect 109335 72559 109421 72615
rect 109477 72559 109563 72615
rect 109619 72559 109705 72615
rect 109761 72559 109802 72615
rect 108948 72473 109802 72559
rect 108948 72417 108995 72473
rect 109051 72417 109137 72473
rect 109193 72417 109279 72473
rect 109335 72417 109421 72473
rect 109477 72417 109563 72473
rect 109619 72417 109705 72473
rect 109761 72417 109802 72473
rect 108948 72331 109802 72417
rect 108948 72275 108995 72331
rect 109051 72275 109137 72331
rect 109193 72275 109279 72331
rect 109335 72275 109421 72331
rect 109477 72275 109563 72331
rect 109619 72275 109705 72331
rect 109761 72275 109802 72331
rect 108948 72189 109802 72275
rect 108948 72133 108995 72189
rect 109051 72133 109137 72189
rect 109193 72133 109279 72189
rect 109335 72133 109421 72189
rect 109477 72133 109563 72189
rect 109619 72133 109705 72189
rect 109761 72133 109802 72189
rect 108948 72088 109802 72133
rect 110122 74035 112172 74088
rect 110122 73979 110193 74035
rect 110249 73979 110335 74035
rect 110391 73979 110477 74035
rect 110533 73979 110619 74035
rect 110675 73979 110761 74035
rect 110817 73979 110903 74035
rect 110959 73979 111045 74035
rect 111101 73979 111187 74035
rect 111243 73979 111329 74035
rect 111385 73979 111471 74035
rect 111527 73979 111613 74035
rect 111669 73979 111755 74035
rect 111811 73979 111897 74035
rect 111953 73979 112039 74035
rect 112095 73979 112172 74035
rect 110122 73893 112172 73979
rect 110122 73837 110193 73893
rect 110249 73837 110335 73893
rect 110391 73837 110477 73893
rect 110533 73837 110619 73893
rect 110675 73837 110761 73893
rect 110817 73837 110903 73893
rect 110959 73837 111045 73893
rect 111101 73837 111187 73893
rect 111243 73837 111329 73893
rect 111385 73837 111471 73893
rect 111527 73837 111613 73893
rect 111669 73837 111755 73893
rect 111811 73837 111897 73893
rect 111953 73837 112039 73893
rect 112095 73837 112172 73893
rect 110122 73751 112172 73837
rect 110122 73695 110193 73751
rect 110249 73695 110335 73751
rect 110391 73695 110477 73751
rect 110533 73695 110619 73751
rect 110675 73695 110761 73751
rect 110817 73695 110903 73751
rect 110959 73695 111045 73751
rect 111101 73695 111187 73751
rect 111243 73695 111329 73751
rect 111385 73695 111471 73751
rect 111527 73695 111613 73751
rect 111669 73695 111755 73751
rect 111811 73695 111897 73751
rect 111953 73695 112039 73751
rect 112095 73695 112172 73751
rect 110122 73609 112172 73695
rect 110122 73553 110193 73609
rect 110249 73553 110335 73609
rect 110391 73553 110477 73609
rect 110533 73553 110619 73609
rect 110675 73553 110761 73609
rect 110817 73553 110903 73609
rect 110959 73553 111045 73609
rect 111101 73553 111187 73609
rect 111243 73553 111329 73609
rect 111385 73553 111471 73609
rect 111527 73553 111613 73609
rect 111669 73553 111755 73609
rect 111811 73553 111897 73609
rect 111953 73553 112039 73609
rect 112095 73553 112172 73609
rect 110122 73467 112172 73553
rect 110122 73411 110193 73467
rect 110249 73411 110335 73467
rect 110391 73411 110477 73467
rect 110533 73411 110619 73467
rect 110675 73411 110761 73467
rect 110817 73411 110903 73467
rect 110959 73411 111045 73467
rect 111101 73411 111187 73467
rect 111243 73411 111329 73467
rect 111385 73411 111471 73467
rect 111527 73411 111613 73467
rect 111669 73411 111755 73467
rect 111811 73411 111897 73467
rect 111953 73411 112039 73467
rect 112095 73411 112172 73467
rect 110122 73325 112172 73411
rect 110122 73269 110193 73325
rect 110249 73269 110335 73325
rect 110391 73269 110477 73325
rect 110533 73269 110619 73325
rect 110675 73269 110761 73325
rect 110817 73269 110903 73325
rect 110959 73269 111045 73325
rect 111101 73269 111187 73325
rect 111243 73269 111329 73325
rect 111385 73269 111471 73325
rect 111527 73269 111613 73325
rect 111669 73269 111755 73325
rect 111811 73269 111897 73325
rect 111953 73269 112039 73325
rect 112095 73269 112172 73325
rect 110122 73183 112172 73269
rect 110122 73127 110193 73183
rect 110249 73127 110335 73183
rect 110391 73127 110477 73183
rect 110533 73127 110619 73183
rect 110675 73127 110761 73183
rect 110817 73127 110903 73183
rect 110959 73127 111045 73183
rect 111101 73127 111187 73183
rect 111243 73127 111329 73183
rect 111385 73127 111471 73183
rect 111527 73127 111613 73183
rect 111669 73127 111755 73183
rect 111811 73127 111897 73183
rect 111953 73127 112039 73183
rect 112095 73127 112172 73183
rect 110122 73041 112172 73127
rect 110122 72985 110193 73041
rect 110249 72985 110335 73041
rect 110391 72985 110477 73041
rect 110533 72985 110619 73041
rect 110675 72985 110761 73041
rect 110817 72985 110903 73041
rect 110959 72985 111045 73041
rect 111101 72985 111187 73041
rect 111243 72985 111329 73041
rect 111385 72985 111471 73041
rect 111527 72985 111613 73041
rect 111669 72985 111755 73041
rect 111811 72985 111897 73041
rect 111953 72985 112039 73041
rect 112095 72985 112172 73041
rect 110122 72899 112172 72985
rect 110122 72843 110193 72899
rect 110249 72843 110335 72899
rect 110391 72843 110477 72899
rect 110533 72843 110619 72899
rect 110675 72843 110761 72899
rect 110817 72843 110903 72899
rect 110959 72843 111045 72899
rect 111101 72843 111187 72899
rect 111243 72843 111329 72899
rect 111385 72843 111471 72899
rect 111527 72843 111613 72899
rect 111669 72843 111755 72899
rect 111811 72843 111897 72899
rect 111953 72843 112039 72899
rect 112095 72843 112172 72899
rect 110122 72757 112172 72843
rect 110122 72701 110193 72757
rect 110249 72701 110335 72757
rect 110391 72701 110477 72757
rect 110533 72701 110619 72757
rect 110675 72701 110761 72757
rect 110817 72701 110903 72757
rect 110959 72701 111045 72757
rect 111101 72701 111187 72757
rect 111243 72701 111329 72757
rect 111385 72701 111471 72757
rect 111527 72701 111613 72757
rect 111669 72701 111755 72757
rect 111811 72701 111897 72757
rect 111953 72701 112039 72757
rect 112095 72701 112172 72757
rect 110122 72615 112172 72701
rect 110122 72559 110193 72615
rect 110249 72559 110335 72615
rect 110391 72559 110477 72615
rect 110533 72559 110619 72615
rect 110675 72559 110761 72615
rect 110817 72559 110903 72615
rect 110959 72559 111045 72615
rect 111101 72559 111187 72615
rect 111243 72559 111329 72615
rect 111385 72559 111471 72615
rect 111527 72559 111613 72615
rect 111669 72559 111755 72615
rect 111811 72559 111897 72615
rect 111953 72559 112039 72615
rect 112095 72559 112172 72615
rect 110122 72473 112172 72559
rect 110122 72417 110193 72473
rect 110249 72417 110335 72473
rect 110391 72417 110477 72473
rect 110533 72417 110619 72473
rect 110675 72417 110761 72473
rect 110817 72417 110903 72473
rect 110959 72417 111045 72473
rect 111101 72417 111187 72473
rect 111243 72417 111329 72473
rect 111385 72417 111471 72473
rect 111527 72417 111613 72473
rect 111669 72417 111755 72473
rect 111811 72417 111897 72473
rect 111953 72417 112039 72473
rect 112095 72417 112172 72473
rect 110122 72331 112172 72417
rect 110122 72275 110193 72331
rect 110249 72275 110335 72331
rect 110391 72275 110477 72331
rect 110533 72275 110619 72331
rect 110675 72275 110761 72331
rect 110817 72275 110903 72331
rect 110959 72275 111045 72331
rect 111101 72275 111187 72331
rect 111243 72275 111329 72331
rect 111385 72275 111471 72331
rect 111527 72275 111613 72331
rect 111669 72275 111755 72331
rect 111811 72275 111897 72331
rect 111953 72275 112039 72331
rect 112095 72275 112172 72331
rect 110122 72189 112172 72275
rect 110122 72133 110193 72189
rect 110249 72133 110335 72189
rect 110391 72133 110477 72189
rect 110533 72133 110619 72189
rect 110675 72133 110761 72189
rect 110817 72133 110903 72189
rect 110959 72133 111045 72189
rect 111101 72133 111187 72189
rect 111243 72133 111329 72189
rect 111385 72133 111471 72189
rect 111527 72133 111613 72189
rect 111669 72133 111755 72189
rect 111811 72133 111897 72189
rect 111953 72133 112039 72189
rect 112095 72133 112172 72189
rect 110122 72088 112172 72133
rect 112828 74035 114878 74088
rect 112828 73979 113325 74035
rect 113381 73979 113467 74035
rect 113523 73979 113609 74035
rect 113665 73979 113751 74035
rect 113807 73979 113893 74035
rect 113949 73979 114035 74035
rect 114091 73979 114177 74035
rect 114233 73979 114319 74035
rect 114375 73979 114461 74035
rect 114517 73979 114603 74035
rect 114659 73979 114745 74035
rect 114801 73979 114878 74035
rect 112828 73893 114878 73979
rect 112828 73837 113325 73893
rect 113381 73837 113467 73893
rect 113523 73837 113609 73893
rect 113665 73837 113751 73893
rect 113807 73837 113893 73893
rect 113949 73837 114035 73893
rect 114091 73837 114177 73893
rect 114233 73837 114319 73893
rect 114375 73837 114461 73893
rect 114517 73837 114603 73893
rect 114659 73837 114745 73893
rect 114801 73837 114878 73893
rect 112828 73751 114878 73837
rect 112828 73695 113325 73751
rect 113381 73695 113467 73751
rect 113523 73695 113609 73751
rect 113665 73695 113751 73751
rect 113807 73695 113893 73751
rect 113949 73695 114035 73751
rect 114091 73695 114177 73751
rect 114233 73695 114319 73751
rect 114375 73695 114461 73751
rect 114517 73695 114603 73751
rect 114659 73695 114745 73751
rect 114801 73695 114878 73751
rect 112828 73609 114878 73695
rect 112828 73553 113325 73609
rect 113381 73553 113467 73609
rect 113523 73553 113609 73609
rect 113665 73553 113751 73609
rect 113807 73553 113893 73609
rect 113949 73553 114035 73609
rect 114091 73553 114177 73609
rect 114233 73553 114319 73609
rect 114375 73553 114461 73609
rect 114517 73553 114603 73609
rect 114659 73553 114745 73609
rect 114801 73553 114878 73609
rect 112828 73467 114878 73553
rect 112828 73411 113325 73467
rect 113381 73411 113467 73467
rect 113523 73411 113609 73467
rect 113665 73411 113751 73467
rect 113807 73411 113893 73467
rect 113949 73411 114035 73467
rect 114091 73411 114177 73467
rect 114233 73411 114319 73467
rect 114375 73411 114461 73467
rect 114517 73411 114603 73467
rect 114659 73411 114745 73467
rect 114801 73411 114878 73467
rect 112828 73325 114878 73411
rect 112828 73269 113325 73325
rect 113381 73269 113467 73325
rect 113523 73269 113609 73325
rect 113665 73269 113751 73325
rect 113807 73269 113893 73325
rect 113949 73269 114035 73325
rect 114091 73269 114177 73325
rect 114233 73269 114319 73325
rect 114375 73269 114461 73325
rect 114517 73269 114603 73325
rect 114659 73269 114745 73325
rect 114801 73269 114878 73325
rect 112828 73183 114878 73269
rect 112828 73127 113325 73183
rect 113381 73127 113467 73183
rect 113523 73127 113609 73183
rect 113665 73127 113751 73183
rect 113807 73127 113893 73183
rect 113949 73127 114035 73183
rect 114091 73127 114177 73183
rect 114233 73127 114319 73183
rect 114375 73127 114461 73183
rect 114517 73127 114603 73183
rect 114659 73127 114745 73183
rect 114801 73127 114878 73183
rect 112828 73041 114878 73127
rect 112828 72985 113325 73041
rect 113381 72985 113467 73041
rect 113523 72985 113609 73041
rect 113665 72985 113751 73041
rect 113807 72985 113893 73041
rect 113949 72985 114035 73041
rect 114091 72985 114177 73041
rect 114233 72985 114319 73041
rect 114375 72985 114461 73041
rect 114517 72985 114603 73041
rect 114659 72985 114745 73041
rect 114801 72985 114878 73041
rect 112828 72899 114878 72985
rect 112828 72843 113325 72899
rect 113381 72843 113467 72899
rect 113523 72843 113609 72899
rect 113665 72843 113751 72899
rect 113807 72843 113893 72899
rect 113949 72843 114035 72899
rect 114091 72843 114177 72899
rect 114233 72843 114319 72899
rect 114375 72843 114461 72899
rect 114517 72843 114603 72899
rect 114659 72843 114745 72899
rect 114801 72843 114878 72899
rect 112828 72757 114878 72843
rect 112828 72701 113325 72757
rect 113381 72701 113467 72757
rect 113523 72701 113609 72757
rect 113665 72701 113751 72757
rect 113807 72701 113893 72757
rect 113949 72701 114035 72757
rect 114091 72701 114177 72757
rect 114233 72701 114319 72757
rect 114375 72701 114461 72757
rect 114517 72701 114603 72757
rect 114659 72701 114745 72757
rect 114801 72701 114878 72757
rect 112828 72615 114878 72701
rect 112828 72559 113325 72615
rect 113381 72559 113467 72615
rect 113523 72559 113609 72615
rect 113665 72559 113751 72615
rect 113807 72559 113893 72615
rect 113949 72559 114035 72615
rect 114091 72559 114177 72615
rect 114233 72559 114319 72615
rect 114375 72559 114461 72615
rect 114517 72559 114603 72615
rect 114659 72559 114745 72615
rect 114801 72559 114878 72615
rect 112828 72473 114878 72559
rect 112828 72417 113325 72473
rect 113381 72417 113467 72473
rect 113523 72417 113609 72473
rect 113665 72417 113751 72473
rect 113807 72417 113893 72473
rect 113949 72417 114035 72473
rect 114091 72417 114177 72473
rect 114233 72417 114319 72473
rect 114375 72417 114461 72473
rect 114517 72417 114603 72473
rect 114659 72417 114745 72473
rect 114801 72417 114878 72473
rect 112828 72331 114878 72417
rect 112828 72275 113325 72331
rect 113381 72275 113467 72331
rect 113523 72275 113609 72331
rect 113665 72275 113751 72331
rect 113807 72275 113893 72331
rect 113949 72275 114035 72331
rect 114091 72275 114177 72331
rect 114233 72275 114319 72331
rect 114375 72275 114461 72331
rect 114517 72275 114603 72331
rect 114659 72275 114745 72331
rect 114801 72275 114878 72331
rect 112828 72189 114878 72275
rect 112828 72133 113325 72189
rect 113381 72133 113467 72189
rect 113523 72133 113609 72189
rect 113665 72133 113751 72189
rect 113807 72133 113893 72189
rect 113949 72133 114035 72189
rect 114091 72133 114177 72189
rect 114233 72133 114319 72189
rect 114375 72133 114461 72189
rect 114517 72133 114603 72189
rect 114659 72133 114745 72189
rect 114801 72133 114878 72189
rect 112828 72088 114878 72133
rect 115198 74035 117248 74088
rect 115198 73979 115269 74035
rect 115325 73979 115411 74035
rect 115467 73979 115553 74035
rect 115609 73979 115695 74035
rect 115751 73979 115837 74035
rect 115893 73979 115979 74035
rect 116035 73979 116121 74035
rect 116177 73979 116263 74035
rect 116319 73979 116405 74035
rect 116461 73979 116547 74035
rect 116603 73979 116689 74035
rect 116745 73979 116831 74035
rect 116887 73979 116973 74035
rect 117029 73979 117115 74035
rect 117171 73979 117248 74035
rect 115198 73893 117248 73979
rect 115198 73837 115269 73893
rect 115325 73837 115411 73893
rect 115467 73837 115553 73893
rect 115609 73837 115695 73893
rect 115751 73837 115837 73893
rect 115893 73837 115979 73893
rect 116035 73837 116121 73893
rect 116177 73837 116263 73893
rect 116319 73837 116405 73893
rect 116461 73837 116547 73893
rect 116603 73837 116689 73893
rect 116745 73837 116831 73893
rect 116887 73837 116973 73893
rect 117029 73837 117115 73893
rect 117171 73837 117248 73893
rect 115198 73751 117248 73837
rect 115198 73695 115269 73751
rect 115325 73695 115411 73751
rect 115467 73695 115553 73751
rect 115609 73695 115695 73751
rect 115751 73695 115837 73751
rect 115893 73695 115979 73751
rect 116035 73695 116121 73751
rect 116177 73695 116263 73751
rect 116319 73695 116405 73751
rect 116461 73695 116547 73751
rect 116603 73695 116689 73751
rect 116745 73695 116831 73751
rect 116887 73695 116973 73751
rect 117029 73695 117115 73751
rect 117171 73695 117248 73751
rect 115198 73609 117248 73695
rect 115198 73553 115269 73609
rect 115325 73553 115411 73609
rect 115467 73553 115553 73609
rect 115609 73553 115695 73609
rect 115751 73553 115837 73609
rect 115893 73553 115979 73609
rect 116035 73553 116121 73609
rect 116177 73553 116263 73609
rect 116319 73553 116405 73609
rect 116461 73553 116547 73609
rect 116603 73553 116689 73609
rect 116745 73553 116831 73609
rect 116887 73553 116973 73609
rect 117029 73553 117115 73609
rect 117171 73553 117248 73609
rect 115198 73467 117248 73553
rect 115198 73411 115269 73467
rect 115325 73411 115411 73467
rect 115467 73411 115553 73467
rect 115609 73411 115695 73467
rect 115751 73411 115837 73467
rect 115893 73411 115979 73467
rect 116035 73411 116121 73467
rect 116177 73411 116263 73467
rect 116319 73411 116405 73467
rect 116461 73411 116547 73467
rect 116603 73411 116689 73467
rect 116745 73411 116831 73467
rect 116887 73411 116973 73467
rect 117029 73411 117115 73467
rect 117171 73411 117248 73467
rect 115198 73325 117248 73411
rect 115198 73269 115269 73325
rect 115325 73269 115411 73325
rect 115467 73269 115553 73325
rect 115609 73269 115695 73325
rect 115751 73269 115837 73325
rect 115893 73269 115979 73325
rect 116035 73269 116121 73325
rect 116177 73269 116263 73325
rect 116319 73269 116405 73325
rect 116461 73269 116547 73325
rect 116603 73269 116689 73325
rect 116745 73269 116831 73325
rect 116887 73269 116973 73325
rect 117029 73269 117115 73325
rect 117171 73269 117248 73325
rect 115198 73183 117248 73269
rect 115198 73127 115269 73183
rect 115325 73127 115411 73183
rect 115467 73127 115553 73183
rect 115609 73127 115695 73183
rect 115751 73127 115837 73183
rect 115893 73127 115979 73183
rect 116035 73127 116121 73183
rect 116177 73127 116263 73183
rect 116319 73127 116405 73183
rect 116461 73127 116547 73183
rect 116603 73127 116689 73183
rect 116745 73127 116831 73183
rect 116887 73127 116973 73183
rect 117029 73127 117115 73183
rect 117171 73127 117248 73183
rect 115198 73041 117248 73127
rect 115198 72985 115269 73041
rect 115325 72985 115411 73041
rect 115467 72985 115553 73041
rect 115609 72985 115695 73041
rect 115751 72985 115837 73041
rect 115893 72985 115979 73041
rect 116035 72985 116121 73041
rect 116177 72985 116263 73041
rect 116319 72985 116405 73041
rect 116461 72985 116547 73041
rect 116603 72985 116689 73041
rect 116745 72985 116831 73041
rect 116887 72985 116973 73041
rect 117029 72985 117115 73041
rect 117171 72985 117248 73041
rect 115198 72899 117248 72985
rect 115198 72843 115269 72899
rect 115325 72843 115411 72899
rect 115467 72843 115553 72899
rect 115609 72843 115695 72899
rect 115751 72843 115837 72899
rect 115893 72843 115979 72899
rect 116035 72843 116121 72899
rect 116177 72843 116263 72899
rect 116319 72843 116405 72899
rect 116461 72843 116547 72899
rect 116603 72843 116689 72899
rect 116745 72843 116831 72899
rect 116887 72843 116973 72899
rect 117029 72843 117115 72899
rect 117171 72843 117248 72899
rect 115198 72757 117248 72843
rect 115198 72701 115269 72757
rect 115325 72701 115411 72757
rect 115467 72701 115553 72757
rect 115609 72701 115695 72757
rect 115751 72701 115837 72757
rect 115893 72701 115979 72757
rect 116035 72701 116121 72757
rect 116177 72701 116263 72757
rect 116319 72701 116405 72757
rect 116461 72701 116547 72757
rect 116603 72701 116689 72757
rect 116745 72701 116831 72757
rect 116887 72701 116973 72757
rect 117029 72701 117115 72757
rect 117171 72701 117248 72757
rect 115198 72615 117248 72701
rect 115198 72559 115269 72615
rect 115325 72559 115411 72615
rect 115467 72559 115553 72615
rect 115609 72559 115695 72615
rect 115751 72559 115837 72615
rect 115893 72559 115979 72615
rect 116035 72559 116121 72615
rect 116177 72559 116263 72615
rect 116319 72559 116405 72615
rect 116461 72559 116547 72615
rect 116603 72559 116689 72615
rect 116745 72559 116831 72615
rect 116887 72559 116973 72615
rect 117029 72559 117115 72615
rect 117171 72559 117248 72615
rect 115198 72473 117248 72559
rect 115198 72417 115269 72473
rect 115325 72417 115411 72473
rect 115467 72417 115553 72473
rect 115609 72417 115695 72473
rect 115751 72417 115837 72473
rect 115893 72417 115979 72473
rect 116035 72417 116121 72473
rect 116177 72417 116263 72473
rect 116319 72417 116405 72473
rect 116461 72417 116547 72473
rect 116603 72417 116689 72473
rect 116745 72417 116831 72473
rect 116887 72417 116973 72473
rect 117029 72417 117115 72473
rect 117171 72417 117248 72473
rect 115198 72331 117248 72417
rect 115198 72275 115269 72331
rect 115325 72275 115411 72331
rect 115467 72275 115553 72331
rect 115609 72275 115695 72331
rect 115751 72275 115837 72331
rect 115893 72275 115979 72331
rect 116035 72275 116121 72331
rect 116177 72275 116263 72331
rect 116319 72275 116405 72331
rect 116461 72275 116547 72331
rect 116603 72275 116689 72331
rect 116745 72275 116831 72331
rect 116887 72275 116973 72331
rect 117029 72275 117115 72331
rect 117171 72275 117248 72331
rect 115198 72189 117248 72275
rect 115198 72133 115269 72189
rect 115325 72133 115411 72189
rect 115467 72133 115553 72189
rect 115609 72133 115695 72189
rect 115751 72133 115837 72189
rect 115893 72133 115979 72189
rect 116035 72133 116121 72189
rect 116177 72133 116263 72189
rect 116319 72133 116405 72189
rect 116461 72133 116547 72189
rect 116603 72133 116689 72189
rect 116745 72133 116831 72189
rect 116887 72133 116973 72189
rect 117029 72133 117115 72189
rect 117171 72133 117248 72189
rect 115198 72088 117248 72133
rect 117828 74035 119728 74088
rect 117828 73979 117899 74035
rect 117955 73979 118041 74035
rect 118097 73979 118183 74035
rect 118239 73979 118325 74035
rect 118381 73979 118467 74035
rect 118523 73979 118609 74035
rect 118665 73979 118751 74035
rect 118807 73979 118893 74035
rect 118949 73979 119035 74035
rect 119091 73979 119177 74035
rect 119233 73979 119319 74035
rect 119375 73979 119461 74035
rect 119517 73979 119603 74035
rect 119659 73979 119728 74035
rect 117828 73893 119728 73979
rect 117828 73837 117899 73893
rect 117955 73837 118041 73893
rect 118097 73837 118183 73893
rect 118239 73837 118325 73893
rect 118381 73837 118467 73893
rect 118523 73837 118609 73893
rect 118665 73837 118751 73893
rect 118807 73837 118893 73893
rect 118949 73837 119035 73893
rect 119091 73837 119177 73893
rect 119233 73837 119319 73893
rect 119375 73837 119461 73893
rect 119517 73837 119603 73893
rect 119659 73837 119728 73893
rect 117828 73751 119728 73837
rect 117828 73695 117899 73751
rect 117955 73695 118041 73751
rect 118097 73695 118183 73751
rect 118239 73695 118325 73751
rect 118381 73695 118467 73751
rect 118523 73695 118609 73751
rect 118665 73695 118751 73751
rect 118807 73695 118893 73751
rect 118949 73695 119035 73751
rect 119091 73695 119177 73751
rect 119233 73695 119319 73751
rect 119375 73695 119461 73751
rect 119517 73695 119603 73751
rect 119659 73695 119728 73751
rect 117828 73609 119728 73695
rect 117828 73553 117899 73609
rect 117955 73553 118041 73609
rect 118097 73553 118183 73609
rect 118239 73553 118325 73609
rect 118381 73553 118467 73609
rect 118523 73553 118609 73609
rect 118665 73553 118751 73609
rect 118807 73553 118893 73609
rect 118949 73553 119035 73609
rect 119091 73553 119177 73609
rect 119233 73553 119319 73609
rect 119375 73553 119461 73609
rect 119517 73553 119603 73609
rect 119659 73553 119728 73609
rect 117828 73467 119728 73553
rect 117828 73411 117899 73467
rect 117955 73411 118041 73467
rect 118097 73411 118183 73467
rect 118239 73411 118325 73467
rect 118381 73411 118467 73467
rect 118523 73411 118609 73467
rect 118665 73411 118751 73467
rect 118807 73411 118893 73467
rect 118949 73411 119035 73467
rect 119091 73411 119177 73467
rect 119233 73411 119319 73467
rect 119375 73411 119461 73467
rect 119517 73411 119603 73467
rect 119659 73411 119728 73467
rect 117828 73325 119728 73411
rect 117828 73269 117899 73325
rect 117955 73269 118041 73325
rect 118097 73269 118183 73325
rect 118239 73269 118325 73325
rect 118381 73269 118467 73325
rect 118523 73269 118609 73325
rect 118665 73269 118751 73325
rect 118807 73269 118893 73325
rect 118949 73269 119035 73325
rect 119091 73269 119177 73325
rect 119233 73269 119319 73325
rect 119375 73269 119461 73325
rect 119517 73269 119603 73325
rect 119659 73269 119728 73325
rect 117828 73183 119728 73269
rect 117828 73127 117899 73183
rect 117955 73127 118041 73183
rect 118097 73127 118183 73183
rect 118239 73127 118325 73183
rect 118381 73127 118467 73183
rect 118523 73127 118609 73183
rect 118665 73127 118751 73183
rect 118807 73127 118893 73183
rect 118949 73127 119035 73183
rect 119091 73127 119177 73183
rect 119233 73127 119319 73183
rect 119375 73127 119461 73183
rect 119517 73127 119603 73183
rect 119659 73127 119728 73183
rect 117828 73041 119728 73127
rect 117828 72985 117899 73041
rect 117955 72985 118041 73041
rect 118097 72985 118183 73041
rect 118239 72985 118325 73041
rect 118381 72985 118467 73041
rect 118523 72985 118609 73041
rect 118665 72985 118751 73041
rect 118807 72985 118893 73041
rect 118949 72985 119035 73041
rect 119091 72985 119177 73041
rect 119233 72985 119319 73041
rect 119375 72985 119461 73041
rect 119517 72985 119603 73041
rect 119659 72985 119728 73041
rect 117828 72899 119728 72985
rect 117828 72843 117899 72899
rect 117955 72843 118041 72899
rect 118097 72843 118183 72899
rect 118239 72843 118325 72899
rect 118381 72843 118467 72899
rect 118523 72843 118609 72899
rect 118665 72843 118751 72899
rect 118807 72843 118893 72899
rect 118949 72843 119035 72899
rect 119091 72843 119177 72899
rect 119233 72843 119319 72899
rect 119375 72843 119461 72899
rect 119517 72843 119603 72899
rect 119659 72843 119728 72899
rect 117828 72757 119728 72843
rect 117828 72701 117899 72757
rect 117955 72701 118041 72757
rect 118097 72701 118183 72757
rect 118239 72701 118325 72757
rect 118381 72701 118467 72757
rect 118523 72701 118609 72757
rect 118665 72701 118751 72757
rect 118807 72701 118893 72757
rect 118949 72701 119035 72757
rect 119091 72701 119177 72757
rect 119233 72701 119319 72757
rect 119375 72701 119461 72757
rect 119517 72701 119603 72757
rect 119659 72701 119728 72757
rect 117828 72615 119728 72701
rect 117828 72559 117899 72615
rect 117955 72559 118041 72615
rect 118097 72559 118183 72615
rect 118239 72559 118325 72615
rect 118381 72559 118467 72615
rect 118523 72559 118609 72615
rect 118665 72559 118751 72615
rect 118807 72559 118893 72615
rect 118949 72559 119035 72615
rect 119091 72559 119177 72615
rect 119233 72559 119319 72615
rect 119375 72559 119461 72615
rect 119517 72559 119603 72615
rect 119659 72559 119728 72615
rect 117828 72473 119728 72559
rect 117828 72417 117899 72473
rect 117955 72417 118041 72473
rect 118097 72417 118183 72473
rect 118239 72417 118325 72473
rect 118381 72417 118467 72473
rect 118523 72417 118609 72473
rect 118665 72417 118751 72473
rect 118807 72417 118893 72473
rect 118949 72417 119035 72473
rect 119091 72417 119177 72473
rect 119233 72417 119319 72473
rect 119375 72417 119461 72473
rect 119517 72417 119603 72473
rect 119659 72417 119728 72473
rect 117828 72331 119728 72417
rect 117828 72275 117899 72331
rect 117955 72275 118041 72331
rect 118097 72275 118183 72331
rect 118239 72275 118325 72331
rect 118381 72275 118467 72331
rect 118523 72275 118609 72331
rect 118665 72275 118751 72331
rect 118807 72275 118893 72331
rect 118949 72275 119035 72331
rect 119091 72275 119177 72331
rect 119233 72275 119319 72331
rect 119375 72275 119461 72331
rect 119517 72275 119603 72331
rect 119659 72275 119728 72331
rect 117828 72189 119728 72275
rect 117828 72133 117899 72189
rect 117955 72133 118041 72189
rect 118097 72133 118183 72189
rect 118239 72133 118325 72189
rect 118381 72133 118467 72189
rect 118523 72133 118609 72189
rect 118665 72133 118751 72189
rect 118807 72133 118893 72189
rect 118949 72133 119035 72189
rect 119091 72133 119177 72189
rect 119233 72133 119319 72189
rect 119375 72133 119461 72189
rect 119517 72133 119603 72189
rect 119659 72133 119728 72189
rect 117828 72088 119728 72133
rect 270272 74035 272172 74088
rect 270272 73979 270343 74035
rect 270399 73979 270485 74035
rect 270541 73979 270627 74035
rect 270683 73979 270769 74035
rect 270825 73979 270911 74035
rect 270967 73979 271053 74035
rect 271109 73979 271195 74035
rect 271251 73979 271337 74035
rect 271393 73979 271479 74035
rect 271535 73979 271621 74035
rect 271677 73979 271763 74035
rect 271819 73979 271905 74035
rect 271961 73979 272047 74035
rect 272103 73979 272172 74035
rect 270272 73893 272172 73979
rect 270272 73837 270343 73893
rect 270399 73837 270485 73893
rect 270541 73837 270627 73893
rect 270683 73837 270769 73893
rect 270825 73837 270911 73893
rect 270967 73837 271053 73893
rect 271109 73837 271195 73893
rect 271251 73837 271337 73893
rect 271393 73837 271479 73893
rect 271535 73837 271621 73893
rect 271677 73837 271763 73893
rect 271819 73837 271905 73893
rect 271961 73837 272047 73893
rect 272103 73837 272172 73893
rect 270272 73751 272172 73837
rect 270272 73695 270343 73751
rect 270399 73695 270485 73751
rect 270541 73695 270627 73751
rect 270683 73695 270769 73751
rect 270825 73695 270911 73751
rect 270967 73695 271053 73751
rect 271109 73695 271195 73751
rect 271251 73695 271337 73751
rect 271393 73695 271479 73751
rect 271535 73695 271621 73751
rect 271677 73695 271763 73751
rect 271819 73695 271905 73751
rect 271961 73695 272047 73751
rect 272103 73695 272172 73751
rect 270272 73609 272172 73695
rect 270272 73553 270343 73609
rect 270399 73553 270485 73609
rect 270541 73553 270627 73609
rect 270683 73553 270769 73609
rect 270825 73553 270911 73609
rect 270967 73553 271053 73609
rect 271109 73553 271195 73609
rect 271251 73553 271337 73609
rect 271393 73553 271479 73609
rect 271535 73553 271621 73609
rect 271677 73553 271763 73609
rect 271819 73553 271905 73609
rect 271961 73553 272047 73609
rect 272103 73553 272172 73609
rect 270272 73467 272172 73553
rect 270272 73411 270343 73467
rect 270399 73411 270485 73467
rect 270541 73411 270627 73467
rect 270683 73411 270769 73467
rect 270825 73411 270911 73467
rect 270967 73411 271053 73467
rect 271109 73411 271195 73467
rect 271251 73411 271337 73467
rect 271393 73411 271479 73467
rect 271535 73411 271621 73467
rect 271677 73411 271763 73467
rect 271819 73411 271905 73467
rect 271961 73411 272047 73467
rect 272103 73411 272172 73467
rect 270272 73325 272172 73411
rect 270272 73269 270343 73325
rect 270399 73269 270485 73325
rect 270541 73269 270627 73325
rect 270683 73269 270769 73325
rect 270825 73269 270911 73325
rect 270967 73269 271053 73325
rect 271109 73269 271195 73325
rect 271251 73269 271337 73325
rect 271393 73269 271479 73325
rect 271535 73269 271621 73325
rect 271677 73269 271763 73325
rect 271819 73269 271905 73325
rect 271961 73269 272047 73325
rect 272103 73269 272172 73325
rect 270272 73183 272172 73269
rect 270272 73127 270343 73183
rect 270399 73127 270485 73183
rect 270541 73127 270627 73183
rect 270683 73127 270769 73183
rect 270825 73127 270911 73183
rect 270967 73127 271053 73183
rect 271109 73127 271195 73183
rect 271251 73127 271337 73183
rect 271393 73127 271479 73183
rect 271535 73127 271621 73183
rect 271677 73127 271763 73183
rect 271819 73127 271905 73183
rect 271961 73127 272047 73183
rect 272103 73127 272172 73183
rect 270272 73041 272172 73127
rect 270272 72985 270343 73041
rect 270399 72985 270485 73041
rect 270541 72985 270627 73041
rect 270683 72985 270769 73041
rect 270825 72985 270911 73041
rect 270967 72985 271053 73041
rect 271109 72985 271195 73041
rect 271251 72985 271337 73041
rect 271393 72985 271479 73041
rect 271535 72985 271621 73041
rect 271677 72985 271763 73041
rect 271819 72985 271905 73041
rect 271961 72985 272047 73041
rect 272103 72985 272172 73041
rect 270272 72899 272172 72985
rect 270272 72843 270343 72899
rect 270399 72843 270485 72899
rect 270541 72843 270627 72899
rect 270683 72843 270769 72899
rect 270825 72843 270911 72899
rect 270967 72843 271053 72899
rect 271109 72843 271195 72899
rect 271251 72843 271337 72899
rect 271393 72843 271479 72899
rect 271535 72843 271621 72899
rect 271677 72843 271763 72899
rect 271819 72843 271905 72899
rect 271961 72843 272047 72899
rect 272103 72843 272172 72899
rect 270272 72757 272172 72843
rect 270272 72701 270343 72757
rect 270399 72701 270485 72757
rect 270541 72701 270627 72757
rect 270683 72701 270769 72757
rect 270825 72701 270911 72757
rect 270967 72701 271053 72757
rect 271109 72701 271195 72757
rect 271251 72701 271337 72757
rect 271393 72701 271479 72757
rect 271535 72701 271621 72757
rect 271677 72701 271763 72757
rect 271819 72701 271905 72757
rect 271961 72701 272047 72757
rect 272103 72701 272172 72757
rect 270272 72615 272172 72701
rect 270272 72559 270343 72615
rect 270399 72559 270485 72615
rect 270541 72559 270627 72615
rect 270683 72559 270769 72615
rect 270825 72559 270911 72615
rect 270967 72559 271053 72615
rect 271109 72559 271195 72615
rect 271251 72559 271337 72615
rect 271393 72559 271479 72615
rect 271535 72559 271621 72615
rect 271677 72559 271763 72615
rect 271819 72559 271905 72615
rect 271961 72559 272047 72615
rect 272103 72559 272172 72615
rect 270272 72473 272172 72559
rect 270272 72417 270343 72473
rect 270399 72417 270485 72473
rect 270541 72417 270627 72473
rect 270683 72417 270769 72473
rect 270825 72417 270911 72473
rect 270967 72417 271053 72473
rect 271109 72417 271195 72473
rect 271251 72417 271337 72473
rect 271393 72417 271479 72473
rect 271535 72417 271621 72473
rect 271677 72417 271763 72473
rect 271819 72417 271905 72473
rect 271961 72417 272047 72473
rect 272103 72417 272172 72473
rect 270272 72331 272172 72417
rect 270272 72275 270343 72331
rect 270399 72275 270485 72331
rect 270541 72275 270627 72331
rect 270683 72275 270769 72331
rect 270825 72275 270911 72331
rect 270967 72275 271053 72331
rect 271109 72275 271195 72331
rect 271251 72275 271337 72331
rect 271393 72275 271479 72331
rect 271535 72275 271621 72331
rect 271677 72275 271763 72331
rect 271819 72275 271905 72331
rect 271961 72275 272047 72331
rect 272103 72275 272172 72331
rect 270272 72189 272172 72275
rect 270272 72133 270343 72189
rect 270399 72133 270485 72189
rect 270541 72133 270627 72189
rect 270683 72133 270769 72189
rect 270825 72133 270911 72189
rect 270967 72133 271053 72189
rect 271109 72133 271195 72189
rect 271251 72133 271337 72189
rect 271393 72133 271479 72189
rect 271535 72133 271621 72189
rect 271677 72133 271763 72189
rect 271819 72133 271905 72189
rect 271961 72133 272047 72189
rect 272103 72133 272172 72189
rect 270272 72088 272172 72133
rect 272752 74035 274802 74088
rect 272752 73979 272823 74035
rect 272879 73979 272965 74035
rect 273021 73979 273107 74035
rect 273163 73979 273249 74035
rect 273305 73979 273391 74035
rect 273447 73979 273533 74035
rect 273589 73979 273675 74035
rect 273731 73979 273817 74035
rect 273873 73979 273959 74035
rect 274015 73979 274101 74035
rect 274157 73979 274243 74035
rect 274299 73979 274385 74035
rect 274441 73979 274527 74035
rect 274583 73979 274669 74035
rect 274725 73979 274802 74035
rect 272752 73893 274802 73979
rect 272752 73837 272823 73893
rect 272879 73837 272965 73893
rect 273021 73837 273107 73893
rect 273163 73837 273249 73893
rect 273305 73837 273391 73893
rect 273447 73837 273533 73893
rect 273589 73837 273675 73893
rect 273731 73837 273817 73893
rect 273873 73837 273959 73893
rect 274015 73837 274101 73893
rect 274157 73837 274243 73893
rect 274299 73837 274385 73893
rect 274441 73837 274527 73893
rect 274583 73837 274669 73893
rect 274725 73837 274802 73893
rect 272752 73751 274802 73837
rect 272752 73695 272823 73751
rect 272879 73695 272965 73751
rect 273021 73695 273107 73751
rect 273163 73695 273249 73751
rect 273305 73695 273391 73751
rect 273447 73695 273533 73751
rect 273589 73695 273675 73751
rect 273731 73695 273817 73751
rect 273873 73695 273959 73751
rect 274015 73695 274101 73751
rect 274157 73695 274243 73751
rect 274299 73695 274385 73751
rect 274441 73695 274527 73751
rect 274583 73695 274669 73751
rect 274725 73695 274802 73751
rect 272752 73609 274802 73695
rect 272752 73553 272823 73609
rect 272879 73553 272965 73609
rect 273021 73553 273107 73609
rect 273163 73553 273249 73609
rect 273305 73553 273391 73609
rect 273447 73553 273533 73609
rect 273589 73553 273675 73609
rect 273731 73553 273817 73609
rect 273873 73553 273959 73609
rect 274015 73553 274101 73609
rect 274157 73553 274243 73609
rect 274299 73553 274385 73609
rect 274441 73553 274527 73609
rect 274583 73553 274669 73609
rect 274725 73553 274802 73609
rect 272752 73467 274802 73553
rect 272752 73411 272823 73467
rect 272879 73411 272965 73467
rect 273021 73411 273107 73467
rect 273163 73411 273249 73467
rect 273305 73411 273391 73467
rect 273447 73411 273533 73467
rect 273589 73411 273675 73467
rect 273731 73411 273817 73467
rect 273873 73411 273959 73467
rect 274015 73411 274101 73467
rect 274157 73411 274243 73467
rect 274299 73411 274385 73467
rect 274441 73411 274527 73467
rect 274583 73411 274669 73467
rect 274725 73411 274802 73467
rect 272752 73325 274802 73411
rect 272752 73269 272823 73325
rect 272879 73269 272965 73325
rect 273021 73269 273107 73325
rect 273163 73269 273249 73325
rect 273305 73269 273391 73325
rect 273447 73269 273533 73325
rect 273589 73269 273675 73325
rect 273731 73269 273817 73325
rect 273873 73269 273959 73325
rect 274015 73269 274101 73325
rect 274157 73269 274243 73325
rect 274299 73269 274385 73325
rect 274441 73269 274527 73325
rect 274583 73269 274669 73325
rect 274725 73269 274802 73325
rect 272752 73183 274802 73269
rect 272752 73127 272823 73183
rect 272879 73127 272965 73183
rect 273021 73127 273107 73183
rect 273163 73127 273249 73183
rect 273305 73127 273391 73183
rect 273447 73127 273533 73183
rect 273589 73127 273675 73183
rect 273731 73127 273817 73183
rect 273873 73127 273959 73183
rect 274015 73127 274101 73183
rect 274157 73127 274243 73183
rect 274299 73127 274385 73183
rect 274441 73127 274527 73183
rect 274583 73127 274669 73183
rect 274725 73127 274802 73183
rect 272752 73041 274802 73127
rect 272752 72985 272823 73041
rect 272879 72985 272965 73041
rect 273021 72985 273107 73041
rect 273163 72985 273249 73041
rect 273305 72985 273391 73041
rect 273447 72985 273533 73041
rect 273589 72985 273675 73041
rect 273731 72985 273817 73041
rect 273873 72985 273959 73041
rect 274015 72985 274101 73041
rect 274157 72985 274243 73041
rect 274299 72985 274385 73041
rect 274441 72985 274527 73041
rect 274583 72985 274669 73041
rect 274725 72985 274802 73041
rect 272752 72899 274802 72985
rect 272752 72843 272823 72899
rect 272879 72843 272965 72899
rect 273021 72843 273107 72899
rect 273163 72843 273249 72899
rect 273305 72843 273391 72899
rect 273447 72843 273533 72899
rect 273589 72843 273675 72899
rect 273731 72843 273817 72899
rect 273873 72843 273959 72899
rect 274015 72843 274101 72899
rect 274157 72843 274243 72899
rect 274299 72843 274385 72899
rect 274441 72843 274527 72899
rect 274583 72843 274669 72899
rect 274725 72843 274802 72899
rect 272752 72757 274802 72843
rect 272752 72701 272823 72757
rect 272879 72701 272965 72757
rect 273021 72701 273107 72757
rect 273163 72701 273249 72757
rect 273305 72701 273391 72757
rect 273447 72701 273533 72757
rect 273589 72701 273675 72757
rect 273731 72701 273817 72757
rect 273873 72701 273959 72757
rect 274015 72701 274101 72757
rect 274157 72701 274243 72757
rect 274299 72701 274385 72757
rect 274441 72701 274527 72757
rect 274583 72701 274669 72757
rect 274725 72701 274802 72757
rect 272752 72615 274802 72701
rect 272752 72559 272823 72615
rect 272879 72559 272965 72615
rect 273021 72559 273107 72615
rect 273163 72559 273249 72615
rect 273305 72559 273391 72615
rect 273447 72559 273533 72615
rect 273589 72559 273675 72615
rect 273731 72559 273817 72615
rect 273873 72559 273959 72615
rect 274015 72559 274101 72615
rect 274157 72559 274243 72615
rect 274299 72559 274385 72615
rect 274441 72559 274527 72615
rect 274583 72559 274669 72615
rect 274725 72559 274802 72615
rect 272752 72473 274802 72559
rect 272752 72417 272823 72473
rect 272879 72417 272965 72473
rect 273021 72417 273107 72473
rect 273163 72417 273249 72473
rect 273305 72417 273391 72473
rect 273447 72417 273533 72473
rect 273589 72417 273675 72473
rect 273731 72417 273817 72473
rect 273873 72417 273959 72473
rect 274015 72417 274101 72473
rect 274157 72417 274243 72473
rect 274299 72417 274385 72473
rect 274441 72417 274527 72473
rect 274583 72417 274669 72473
rect 274725 72417 274802 72473
rect 272752 72331 274802 72417
rect 272752 72275 272823 72331
rect 272879 72275 272965 72331
rect 273021 72275 273107 72331
rect 273163 72275 273249 72331
rect 273305 72275 273391 72331
rect 273447 72275 273533 72331
rect 273589 72275 273675 72331
rect 273731 72275 273817 72331
rect 273873 72275 273959 72331
rect 274015 72275 274101 72331
rect 274157 72275 274243 72331
rect 274299 72275 274385 72331
rect 274441 72275 274527 72331
rect 274583 72275 274669 72331
rect 274725 72275 274802 72331
rect 272752 72189 274802 72275
rect 272752 72133 272823 72189
rect 272879 72133 272965 72189
rect 273021 72133 273107 72189
rect 273163 72133 273249 72189
rect 273305 72133 273391 72189
rect 273447 72133 273533 72189
rect 273589 72133 273675 72189
rect 273731 72133 273817 72189
rect 273873 72133 273959 72189
rect 274015 72133 274101 72189
rect 274157 72133 274243 72189
rect 274299 72133 274385 72189
rect 274441 72133 274527 72189
rect 274583 72133 274669 72189
rect 274725 72133 274802 72189
rect 272752 72088 274802 72133
rect 275122 74035 277172 74088
rect 275122 73979 275193 74035
rect 275249 73979 275335 74035
rect 275391 73979 275477 74035
rect 275533 73979 275619 74035
rect 275675 73979 275761 74035
rect 275817 73979 275903 74035
rect 275959 73979 276045 74035
rect 276101 73979 276187 74035
rect 276243 73979 276329 74035
rect 276385 73979 276471 74035
rect 276527 73979 276613 74035
rect 276669 73979 276755 74035
rect 276811 73979 276897 74035
rect 276953 73979 277039 74035
rect 277095 73979 277172 74035
rect 275122 73893 277172 73979
rect 275122 73837 275193 73893
rect 275249 73837 275335 73893
rect 275391 73837 275477 73893
rect 275533 73837 275619 73893
rect 275675 73837 275761 73893
rect 275817 73837 275903 73893
rect 275959 73837 276045 73893
rect 276101 73837 276187 73893
rect 276243 73837 276329 73893
rect 276385 73837 276471 73893
rect 276527 73837 276613 73893
rect 276669 73837 276755 73893
rect 276811 73837 276897 73893
rect 276953 73837 277039 73893
rect 277095 73837 277172 73893
rect 275122 73751 277172 73837
rect 275122 73695 275193 73751
rect 275249 73695 275335 73751
rect 275391 73695 275477 73751
rect 275533 73695 275619 73751
rect 275675 73695 275761 73751
rect 275817 73695 275903 73751
rect 275959 73695 276045 73751
rect 276101 73695 276187 73751
rect 276243 73695 276329 73751
rect 276385 73695 276471 73751
rect 276527 73695 276613 73751
rect 276669 73695 276755 73751
rect 276811 73695 276897 73751
rect 276953 73695 277039 73751
rect 277095 73695 277172 73751
rect 275122 73609 277172 73695
rect 275122 73553 275193 73609
rect 275249 73553 275335 73609
rect 275391 73553 275477 73609
rect 275533 73553 275619 73609
rect 275675 73553 275761 73609
rect 275817 73553 275903 73609
rect 275959 73553 276045 73609
rect 276101 73553 276187 73609
rect 276243 73553 276329 73609
rect 276385 73553 276471 73609
rect 276527 73553 276613 73609
rect 276669 73553 276755 73609
rect 276811 73553 276897 73609
rect 276953 73553 277039 73609
rect 277095 73553 277172 73609
rect 275122 73467 277172 73553
rect 275122 73411 275193 73467
rect 275249 73411 275335 73467
rect 275391 73411 275477 73467
rect 275533 73411 275619 73467
rect 275675 73411 275761 73467
rect 275817 73411 275903 73467
rect 275959 73411 276045 73467
rect 276101 73411 276187 73467
rect 276243 73411 276329 73467
rect 276385 73411 276471 73467
rect 276527 73411 276613 73467
rect 276669 73411 276755 73467
rect 276811 73411 276897 73467
rect 276953 73411 277039 73467
rect 277095 73411 277172 73467
rect 275122 73325 277172 73411
rect 275122 73269 275193 73325
rect 275249 73269 275335 73325
rect 275391 73269 275477 73325
rect 275533 73269 275619 73325
rect 275675 73269 275761 73325
rect 275817 73269 275903 73325
rect 275959 73269 276045 73325
rect 276101 73269 276187 73325
rect 276243 73269 276329 73325
rect 276385 73269 276471 73325
rect 276527 73269 276613 73325
rect 276669 73269 276755 73325
rect 276811 73269 276897 73325
rect 276953 73269 277039 73325
rect 277095 73269 277172 73325
rect 275122 73183 277172 73269
rect 275122 73127 275193 73183
rect 275249 73127 275335 73183
rect 275391 73127 275477 73183
rect 275533 73127 275619 73183
rect 275675 73127 275761 73183
rect 275817 73127 275903 73183
rect 275959 73127 276045 73183
rect 276101 73127 276187 73183
rect 276243 73127 276329 73183
rect 276385 73127 276471 73183
rect 276527 73127 276613 73183
rect 276669 73127 276755 73183
rect 276811 73127 276897 73183
rect 276953 73127 277039 73183
rect 277095 73127 277172 73183
rect 275122 73041 277172 73127
rect 275122 72985 275193 73041
rect 275249 72985 275335 73041
rect 275391 72985 275477 73041
rect 275533 72985 275619 73041
rect 275675 72985 275761 73041
rect 275817 72985 275903 73041
rect 275959 72985 276045 73041
rect 276101 72985 276187 73041
rect 276243 72985 276329 73041
rect 276385 72985 276471 73041
rect 276527 72985 276613 73041
rect 276669 72985 276755 73041
rect 276811 72985 276897 73041
rect 276953 72985 277039 73041
rect 277095 72985 277172 73041
rect 275122 72899 277172 72985
rect 275122 72843 275193 72899
rect 275249 72843 275335 72899
rect 275391 72843 275477 72899
rect 275533 72843 275619 72899
rect 275675 72843 275761 72899
rect 275817 72843 275903 72899
rect 275959 72843 276045 72899
rect 276101 72843 276187 72899
rect 276243 72843 276329 72899
rect 276385 72843 276471 72899
rect 276527 72843 276613 72899
rect 276669 72843 276755 72899
rect 276811 72843 276897 72899
rect 276953 72843 277039 72899
rect 277095 72843 277172 72899
rect 275122 72757 277172 72843
rect 275122 72701 275193 72757
rect 275249 72701 275335 72757
rect 275391 72701 275477 72757
rect 275533 72701 275619 72757
rect 275675 72701 275761 72757
rect 275817 72701 275903 72757
rect 275959 72701 276045 72757
rect 276101 72701 276187 72757
rect 276243 72701 276329 72757
rect 276385 72701 276471 72757
rect 276527 72701 276613 72757
rect 276669 72701 276755 72757
rect 276811 72701 276897 72757
rect 276953 72701 277039 72757
rect 277095 72701 277172 72757
rect 275122 72615 277172 72701
rect 275122 72559 275193 72615
rect 275249 72559 275335 72615
rect 275391 72559 275477 72615
rect 275533 72559 275619 72615
rect 275675 72559 275761 72615
rect 275817 72559 275903 72615
rect 275959 72559 276045 72615
rect 276101 72559 276187 72615
rect 276243 72559 276329 72615
rect 276385 72559 276471 72615
rect 276527 72559 276613 72615
rect 276669 72559 276755 72615
rect 276811 72559 276897 72615
rect 276953 72559 277039 72615
rect 277095 72559 277172 72615
rect 275122 72473 277172 72559
rect 275122 72417 275193 72473
rect 275249 72417 275335 72473
rect 275391 72417 275477 72473
rect 275533 72417 275619 72473
rect 275675 72417 275761 72473
rect 275817 72417 275903 72473
rect 275959 72417 276045 72473
rect 276101 72417 276187 72473
rect 276243 72417 276329 72473
rect 276385 72417 276471 72473
rect 276527 72417 276613 72473
rect 276669 72417 276755 72473
rect 276811 72417 276897 72473
rect 276953 72417 277039 72473
rect 277095 72417 277172 72473
rect 275122 72331 277172 72417
rect 275122 72275 275193 72331
rect 275249 72275 275335 72331
rect 275391 72275 275477 72331
rect 275533 72275 275619 72331
rect 275675 72275 275761 72331
rect 275817 72275 275903 72331
rect 275959 72275 276045 72331
rect 276101 72275 276187 72331
rect 276243 72275 276329 72331
rect 276385 72275 276471 72331
rect 276527 72275 276613 72331
rect 276669 72275 276755 72331
rect 276811 72275 276897 72331
rect 276953 72275 277039 72331
rect 277095 72275 277172 72331
rect 275122 72189 277172 72275
rect 275122 72133 275193 72189
rect 275249 72133 275335 72189
rect 275391 72133 275477 72189
rect 275533 72133 275619 72189
rect 275675 72133 275761 72189
rect 275817 72133 275903 72189
rect 275959 72133 276045 72189
rect 276101 72133 276187 72189
rect 276243 72133 276329 72189
rect 276385 72133 276471 72189
rect 276527 72133 276613 72189
rect 276669 72133 276755 72189
rect 276811 72133 276897 72189
rect 276953 72133 277039 72189
rect 277095 72133 277172 72189
rect 275122 72088 277172 72133
rect 277828 74035 279878 74088
rect 277828 73979 277899 74035
rect 277955 73979 278041 74035
rect 278097 73979 278183 74035
rect 278239 73979 278325 74035
rect 278381 73979 278467 74035
rect 278523 73979 278609 74035
rect 278665 73979 278751 74035
rect 278807 73979 278893 74035
rect 278949 73979 279035 74035
rect 279091 73979 279177 74035
rect 279233 73979 279319 74035
rect 279375 73979 279461 74035
rect 279517 73979 279603 74035
rect 279659 73979 279745 74035
rect 279801 73979 279878 74035
rect 277828 73893 279878 73979
rect 277828 73837 277899 73893
rect 277955 73837 278041 73893
rect 278097 73837 278183 73893
rect 278239 73837 278325 73893
rect 278381 73837 278467 73893
rect 278523 73837 278609 73893
rect 278665 73837 278751 73893
rect 278807 73837 278893 73893
rect 278949 73837 279035 73893
rect 279091 73837 279177 73893
rect 279233 73837 279319 73893
rect 279375 73837 279461 73893
rect 279517 73837 279603 73893
rect 279659 73837 279745 73893
rect 279801 73837 279878 73893
rect 277828 73751 279878 73837
rect 277828 73695 277899 73751
rect 277955 73695 278041 73751
rect 278097 73695 278183 73751
rect 278239 73695 278325 73751
rect 278381 73695 278467 73751
rect 278523 73695 278609 73751
rect 278665 73695 278751 73751
rect 278807 73695 278893 73751
rect 278949 73695 279035 73751
rect 279091 73695 279177 73751
rect 279233 73695 279319 73751
rect 279375 73695 279461 73751
rect 279517 73695 279603 73751
rect 279659 73695 279745 73751
rect 279801 73695 279878 73751
rect 277828 73609 279878 73695
rect 277828 73553 277899 73609
rect 277955 73553 278041 73609
rect 278097 73553 278183 73609
rect 278239 73553 278325 73609
rect 278381 73553 278467 73609
rect 278523 73553 278609 73609
rect 278665 73553 278751 73609
rect 278807 73553 278893 73609
rect 278949 73553 279035 73609
rect 279091 73553 279177 73609
rect 279233 73553 279319 73609
rect 279375 73553 279461 73609
rect 279517 73553 279603 73609
rect 279659 73553 279745 73609
rect 279801 73553 279878 73609
rect 277828 73467 279878 73553
rect 277828 73411 277899 73467
rect 277955 73411 278041 73467
rect 278097 73411 278183 73467
rect 278239 73411 278325 73467
rect 278381 73411 278467 73467
rect 278523 73411 278609 73467
rect 278665 73411 278751 73467
rect 278807 73411 278893 73467
rect 278949 73411 279035 73467
rect 279091 73411 279177 73467
rect 279233 73411 279319 73467
rect 279375 73411 279461 73467
rect 279517 73411 279603 73467
rect 279659 73411 279745 73467
rect 279801 73411 279878 73467
rect 277828 73325 279878 73411
rect 277828 73269 277899 73325
rect 277955 73269 278041 73325
rect 278097 73269 278183 73325
rect 278239 73269 278325 73325
rect 278381 73269 278467 73325
rect 278523 73269 278609 73325
rect 278665 73269 278751 73325
rect 278807 73269 278893 73325
rect 278949 73269 279035 73325
rect 279091 73269 279177 73325
rect 279233 73269 279319 73325
rect 279375 73269 279461 73325
rect 279517 73269 279603 73325
rect 279659 73269 279745 73325
rect 279801 73269 279878 73325
rect 277828 73183 279878 73269
rect 277828 73127 277899 73183
rect 277955 73127 278041 73183
rect 278097 73127 278183 73183
rect 278239 73127 278325 73183
rect 278381 73127 278467 73183
rect 278523 73127 278609 73183
rect 278665 73127 278751 73183
rect 278807 73127 278893 73183
rect 278949 73127 279035 73183
rect 279091 73127 279177 73183
rect 279233 73127 279319 73183
rect 279375 73127 279461 73183
rect 279517 73127 279603 73183
rect 279659 73127 279745 73183
rect 279801 73127 279878 73183
rect 277828 73041 279878 73127
rect 277828 72985 277899 73041
rect 277955 72985 278041 73041
rect 278097 72985 278183 73041
rect 278239 72985 278325 73041
rect 278381 72985 278467 73041
rect 278523 72985 278609 73041
rect 278665 72985 278751 73041
rect 278807 72985 278893 73041
rect 278949 72985 279035 73041
rect 279091 72985 279177 73041
rect 279233 72985 279319 73041
rect 279375 72985 279461 73041
rect 279517 72985 279603 73041
rect 279659 72985 279745 73041
rect 279801 72985 279878 73041
rect 277828 72899 279878 72985
rect 277828 72843 277899 72899
rect 277955 72843 278041 72899
rect 278097 72843 278183 72899
rect 278239 72843 278325 72899
rect 278381 72843 278467 72899
rect 278523 72843 278609 72899
rect 278665 72843 278751 72899
rect 278807 72843 278893 72899
rect 278949 72843 279035 72899
rect 279091 72843 279177 72899
rect 279233 72843 279319 72899
rect 279375 72843 279461 72899
rect 279517 72843 279603 72899
rect 279659 72843 279745 72899
rect 279801 72843 279878 72899
rect 277828 72757 279878 72843
rect 277828 72701 277899 72757
rect 277955 72701 278041 72757
rect 278097 72701 278183 72757
rect 278239 72701 278325 72757
rect 278381 72701 278467 72757
rect 278523 72701 278609 72757
rect 278665 72701 278751 72757
rect 278807 72701 278893 72757
rect 278949 72701 279035 72757
rect 279091 72701 279177 72757
rect 279233 72701 279319 72757
rect 279375 72701 279461 72757
rect 279517 72701 279603 72757
rect 279659 72701 279745 72757
rect 279801 72701 279878 72757
rect 277828 72615 279878 72701
rect 277828 72559 277899 72615
rect 277955 72559 278041 72615
rect 278097 72559 278183 72615
rect 278239 72559 278325 72615
rect 278381 72559 278467 72615
rect 278523 72559 278609 72615
rect 278665 72559 278751 72615
rect 278807 72559 278893 72615
rect 278949 72559 279035 72615
rect 279091 72559 279177 72615
rect 279233 72559 279319 72615
rect 279375 72559 279461 72615
rect 279517 72559 279603 72615
rect 279659 72559 279745 72615
rect 279801 72559 279878 72615
rect 277828 72473 279878 72559
rect 277828 72417 277899 72473
rect 277955 72417 278041 72473
rect 278097 72417 278183 72473
rect 278239 72417 278325 72473
rect 278381 72417 278467 72473
rect 278523 72417 278609 72473
rect 278665 72417 278751 72473
rect 278807 72417 278893 72473
rect 278949 72417 279035 72473
rect 279091 72417 279177 72473
rect 279233 72417 279319 72473
rect 279375 72417 279461 72473
rect 279517 72417 279603 72473
rect 279659 72417 279745 72473
rect 279801 72417 279878 72473
rect 277828 72331 279878 72417
rect 277828 72275 277899 72331
rect 277955 72275 278041 72331
rect 278097 72275 278183 72331
rect 278239 72275 278325 72331
rect 278381 72275 278467 72331
rect 278523 72275 278609 72331
rect 278665 72275 278751 72331
rect 278807 72275 278893 72331
rect 278949 72275 279035 72331
rect 279091 72275 279177 72331
rect 279233 72275 279319 72331
rect 279375 72275 279461 72331
rect 279517 72275 279603 72331
rect 279659 72275 279745 72331
rect 279801 72275 279878 72331
rect 277828 72189 279878 72275
rect 277828 72133 277899 72189
rect 277955 72133 278041 72189
rect 278097 72133 278183 72189
rect 278239 72133 278325 72189
rect 278381 72133 278467 72189
rect 278523 72133 278609 72189
rect 278665 72133 278751 72189
rect 278807 72133 278893 72189
rect 278949 72133 279035 72189
rect 279091 72133 279177 72189
rect 279233 72133 279319 72189
rect 279375 72133 279461 72189
rect 279517 72133 279603 72189
rect 279659 72133 279745 72189
rect 279801 72133 279878 72189
rect 277828 72088 279878 72133
rect 280198 74035 282248 74088
rect 280198 73979 280269 74035
rect 280325 73979 280411 74035
rect 280467 73979 280553 74035
rect 280609 73979 280695 74035
rect 280751 73979 280837 74035
rect 280893 73979 280979 74035
rect 281035 73979 281121 74035
rect 281177 73979 281263 74035
rect 281319 73979 281405 74035
rect 281461 73979 281547 74035
rect 281603 73979 281689 74035
rect 281745 73979 281831 74035
rect 281887 73979 281973 74035
rect 282029 73979 282115 74035
rect 282171 73979 282248 74035
rect 280198 73893 282248 73979
rect 280198 73837 280269 73893
rect 280325 73837 280411 73893
rect 280467 73837 280553 73893
rect 280609 73837 280695 73893
rect 280751 73837 280837 73893
rect 280893 73837 280979 73893
rect 281035 73837 281121 73893
rect 281177 73837 281263 73893
rect 281319 73837 281405 73893
rect 281461 73837 281547 73893
rect 281603 73837 281689 73893
rect 281745 73837 281831 73893
rect 281887 73837 281973 73893
rect 282029 73837 282115 73893
rect 282171 73837 282248 73893
rect 280198 73751 282248 73837
rect 280198 73695 280269 73751
rect 280325 73695 280411 73751
rect 280467 73695 280553 73751
rect 280609 73695 280695 73751
rect 280751 73695 280837 73751
rect 280893 73695 280979 73751
rect 281035 73695 281121 73751
rect 281177 73695 281263 73751
rect 281319 73695 281405 73751
rect 281461 73695 281547 73751
rect 281603 73695 281689 73751
rect 281745 73695 281831 73751
rect 281887 73695 281973 73751
rect 282029 73695 282115 73751
rect 282171 73695 282248 73751
rect 280198 73609 282248 73695
rect 280198 73553 280269 73609
rect 280325 73553 280411 73609
rect 280467 73553 280553 73609
rect 280609 73553 280695 73609
rect 280751 73553 280837 73609
rect 280893 73553 280979 73609
rect 281035 73553 281121 73609
rect 281177 73553 281263 73609
rect 281319 73553 281405 73609
rect 281461 73553 281547 73609
rect 281603 73553 281689 73609
rect 281745 73553 281831 73609
rect 281887 73553 281973 73609
rect 282029 73553 282115 73609
rect 282171 73553 282248 73609
rect 280198 73467 282248 73553
rect 280198 73411 280269 73467
rect 280325 73411 280411 73467
rect 280467 73411 280553 73467
rect 280609 73411 280695 73467
rect 280751 73411 280837 73467
rect 280893 73411 280979 73467
rect 281035 73411 281121 73467
rect 281177 73411 281263 73467
rect 281319 73411 281405 73467
rect 281461 73411 281547 73467
rect 281603 73411 281689 73467
rect 281745 73411 281831 73467
rect 281887 73411 281973 73467
rect 282029 73411 282115 73467
rect 282171 73411 282248 73467
rect 280198 73325 282248 73411
rect 280198 73269 280269 73325
rect 280325 73269 280411 73325
rect 280467 73269 280553 73325
rect 280609 73269 280695 73325
rect 280751 73269 280837 73325
rect 280893 73269 280979 73325
rect 281035 73269 281121 73325
rect 281177 73269 281263 73325
rect 281319 73269 281405 73325
rect 281461 73269 281547 73325
rect 281603 73269 281689 73325
rect 281745 73269 281831 73325
rect 281887 73269 281973 73325
rect 282029 73269 282115 73325
rect 282171 73269 282248 73325
rect 280198 73183 282248 73269
rect 280198 73127 280269 73183
rect 280325 73127 280411 73183
rect 280467 73127 280553 73183
rect 280609 73127 280695 73183
rect 280751 73127 280837 73183
rect 280893 73127 280979 73183
rect 281035 73127 281121 73183
rect 281177 73127 281263 73183
rect 281319 73127 281405 73183
rect 281461 73127 281547 73183
rect 281603 73127 281689 73183
rect 281745 73127 281831 73183
rect 281887 73127 281973 73183
rect 282029 73127 282115 73183
rect 282171 73127 282248 73183
rect 280198 73041 282248 73127
rect 280198 72985 280269 73041
rect 280325 72985 280411 73041
rect 280467 72985 280553 73041
rect 280609 72985 280695 73041
rect 280751 72985 280837 73041
rect 280893 72985 280979 73041
rect 281035 72985 281121 73041
rect 281177 72985 281263 73041
rect 281319 72985 281405 73041
rect 281461 72985 281547 73041
rect 281603 72985 281689 73041
rect 281745 72985 281831 73041
rect 281887 72985 281973 73041
rect 282029 72985 282115 73041
rect 282171 72985 282248 73041
rect 280198 72899 282248 72985
rect 280198 72843 280269 72899
rect 280325 72843 280411 72899
rect 280467 72843 280553 72899
rect 280609 72843 280695 72899
rect 280751 72843 280837 72899
rect 280893 72843 280979 72899
rect 281035 72843 281121 72899
rect 281177 72843 281263 72899
rect 281319 72843 281405 72899
rect 281461 72843 281547 72899
rect 281603 72843 281689 72899
rect 281745 72843 281831 72899
rect 281887 72843 281973 72899
rect 282029 72843 282115 72899
rect 282171 72843 282248 72899
rect 280198 72757 282248 72843
rect 280198 72701 280269 72757
rect 280325 72701 280411 72757
rect 280467 72701 280553 72757
rect 280609 72701 280695 72757
rect 280751 72701 280837 72757
rect 280893 72701 280979 72757
rect 281035 72701 281121 72757
rect 281177 72701 281263 72757
rect 281319 72701 281405 72757
rect 281461 72701 281547 72757
rect 281603 72701 281689 72757
rect 281745 72701 281831 72757
rect 281887 72701 281973 72757
rect 282029 72701 282115 72757
rect 282171 72701 282248 72757
rect 280198 72615 282248 72701
rect 280198 72559 280269 72615
rect 280325 72559 280411 72615
rect 280467 72559 280553 72615
rect 280609 72559 280695 72615
rect 280751 72559 280837 72615
rect 280893 72559 280979 72615
rect 281035 72559 281121 72615
rect 281177 72559 281263 72615
rect 281319 72559 281405 72615
rect 281461 72559 281547 72615
rect 281603 72559 281689 72615
rect 281745 72559 281831 72615
rect 281887 72559 281973 72615
rect 282029 72559 282115 72615
rect 282171 72559 282248 72615
rect 280198 72473 282248 72559
rect 280198 72417 280269 72473
rect 280325 72417 280411 72473
rect 280467 72417 280553 72473
rect 280609 72417 280695 72473
rect 280751 72417 280837 72473
rect 280893 72417 280979 72473
rect 281035 72417 281121 72473
rect 281177 72417 281263 72473
rect 281319 72417 281405 72473
rect 281461 72417 281547 72473
rect 281603 72417 281689 72473
rect 281745 72417 281831 72473
rect 281887 72417 281973 72473
rect 282029 72417 282115 72473
rect 282171 72417 282248 72473
rect 280198 72331 282248 72417
rect 280198 72275 280269 72331
rect 280325 72275 280411 72331
rect 280467 72275 280553 72331
rect 280609 72275 280695 72331
rect 280751 72275 280837 72331
rect 280893 72275 280979 72331
rect 281035 72275 281121 72331
rect 281177 72275 281263 72331
rect 281319 72275 281405 72331
rect 281461 72275 281547 72331
rect 281603 72275 281689 72331
rect 281745 72275 281831 72331
rect 281887 72275 281973 72331
rect 282029 72275 282115 72331
rect 282171 72275 282248 72331
rect 280198 72189 282248 72275
rect 280198 72133 280269 72189
rect 280325 72133 280411 72189
rect 280467 72133 280553 72189
rect 280609 72133 280695 72189
rect 280751 72133 280837 72189
rect 280893 72133 280979 72189
rect 281035 72133 281121 72189
rect 281177 72133 281263 72189
rect 281319 72133 281405 72189
rect 281461 72133 281547 72189
rect 281603 72133 281689 72189
rect 281745 72133 281831 72189
rect 281887 72133 281973 72189
rect 282029 72133 282115 72189
rect 282171 72133 282248 72189
rect 280198 72088 282248 72133
rect 282828 74035 284016 74088
rect 282828 73979 282899 74035
rect 282955 73979 283041 74035
rect 283097 73979 283183 74035
rect 283239 73979 283325 74035
rect 283381 73979 283467 74035
rect 283523 73979 283609 74035
rect 283665 73979 283751 74035
rect 283807 73979 283893 74035
rect 283949 73979 284016 74035
rect 282828 73893 284016 73979
rect 282828 73837 282899 73893
rect 282955 73837 283041 73893
rect 283097 73837 283183 73893
rect 283239 73837 283325 73893
rect 283381 73837 283467 73893
rect 283523 73837 283609 73893
rect 283665 73837 283751 73893
rect 283807 73837 283893 73893
rect 283949 73837 284016 73893
rect 282828 73751 284016 73837
rect 282828 73695 282899 73751
rect 282955 73695 283041 73751
rect 283097 73695 283183 73751
rect 283239 73695 283325 73751
rect 283381 73695 283467 73751
rect 283523 73695 283609 73751
rect 283665 73695 283751 73751
rect 283807 73695 283893 73751
rect 283949 73695 284016 73751
rect 282828 73609 284016 73695
rect 282828 73553 282899 73609
rect 282955 73553 283041 73609
rect 283097 73553 283183 73609
rect 283239 73553 283325 73609
rect 283381 73553 283467 73609
rect 283523 73553 283609 73609
rect 283665 73553 283751 73609
rect 283807 73553 283893 73609
rect 283949 73553 284016 73609
rect 282828 73467 284016 73553
rect 282828 73411 282899 73467
rect 282955 73411 283041 73467
rect 283097 73411 283183 73467
rect 283239 73411 283325 73467
rect 283381 73411 283467 73467
rect 283523 73411 283609 73467
rect 283665 73411 283751 73467
rect 283807 73411 283893 73467
rect 283949 73411 284016 73467
rect 282828 73325 284016 73411
rect 282828 73269 282899 73325
rect 282955 73269 283041 73325
rect 283097 73269 283183 73325
rect 283239 73269 283325 73325
rect 283381 73269 283467 73325
rect 283523 73269 283609 73325
rect 283665 73269 283751 73325
rect 283807 73269 283893 73325
rect 283949 73269 284016 73325
rect 282828 73183 284016 73269
rect 282828 73127 282899 73183
rect 282955 73127 283041 73183
rect 283097 73127 283183 73183
rect 283239 73127 283325 73183
rect 283381 73127 283467 73183
rect 283523 73127 283609 73183
rect 283665 73127 283751 73183
rect 283807 73127 283893 73183
rect 283949 73127 284016 73183
rect 282828 73041 284016 73127
rect 282828 72985 282899 73041
rect 282955 72985 283041 73041
rect 283097 72985 283183 73041
rect 283239 72985 283325 73041
rect 283381 72985 283467 73041
rect 283523 72985 283609 73041
rect 283665 72985 283751 73041
rect 283807 72985 283893 73041
rect 283949 72985 284016 73041
rect 282828 72899 284016 72985
rect 282828 72843 282899 72899
rect 282955 72843 283041 72899
rect 283097 72843 283183 72899
rect 283239 72843 283325 72899
rect 283381 72843 283467 72899
rect 283523 72843 283609 72899
rect 283665 72843 283751 72899
rect 283807 72843 283893 72899
rect 283949 72843 284016 72899
rect 282828 72757 284016 72843
rect 282828 72701 282899 72757
rect 282955 72701 283041 72757
rect 283097 72701 283183 72757
rect 283239 72701 283325 72757
rect 283381 72701 283467 72757
rect 283523 72701 283609 72757
rect 283665 72701 283751 72757
rect 283807 72701 283893 72757
rect 283949 72701 284016 72757
rect 282828 72615 284016 72701
rect 282828 72559 282899 72615
rect 282955 72559 283041 72615
rect 283097 72559 283183 72615
rect 283239 72559 283325 72615
rect 283381 72559 283467 72615
rect 283523 72559 283609 72615
rect 283665 72559 283751 72615
rect 283807 72559 283893 72615
rect 283949 72559 284016 72615
rect 282828 72473 284016 72559
rect 282828 72417 282899 72473
rect 282955 72417 283041 72473
rect 283097 72417 283183 72473
rect 283239 72417 283325 72473
rect 283381 72417 283467 72473
rect 283523 72417 283609 72473
rect 283665 72417 283751 72473
rect 283807 72417 283893 72473
rect 283949 72417 284016 72473
rect 282828 72331 284016 72417
rect 282828 72275 282899 72331
rect 282955 72275 283041 72331
rect 283097 72275 283183 72331
rect 283239 72275 283325 72331
rect 283381 72275 283467 72331
rect 283523 72275 283609 72331
rect 283665 72275 283751 72331
rect 283807 72275 283893 72331
rect 283949 72275 284016 72331
rect 282828 72189 284016 72275
rect 282828 72133 282899 72189
rect 282955 72133 283041 72189
rect 283097 72133 283183 72189
rect 283239 72133 283325 72189
rect 283381 72133 283467 72189
rect 283523 72133 283609 72189
rect 283665 72133 283751 72189
rect 283807 72133 283893 72189
rect 283949 72133 284016 72189
rect 282828 72088 284016 72133
rect 600272 74035 602172 74088
rect 600272 73979 600343 74035
rect 600399 73979 600485 74035
rect 600541 73979 600627 74035
rect 600683 73979 600769 74035
rect 600825 73979 600911 74035
rect 600967 73979 601053 74035
rect 601109 73979 601195 74035
rect 601251 73979 601337 74035
rect 601393 73979 601479 74035
rect 601535 73979 601621 74035
rect 601677 73979 601763 74035
rect 601819 73979 601905 74035
rect 601961 73979 602047 74035
rect 602103 73979 602172 74035
rect 600272 73893 602172 73979
rect 600272 73837 600343 73893
rect 600399 73837 600485 73893
rect 600541 73837 600627 73893
rect 600683 73837 600769 73893
rect 600825 73837 600911 73893
rect 600967 73837 601053 73893
rect 601109 73837 601195 73893
rect 601251 73837 601337 73893
rect 601393 73837 601479 73893
rect 601535 73837 601621 73893
rect 601677 73837 601763 73893
rect 601819 73837 601905 73893
rect 601961 73837 602047 73893
rect 602103 73837 602172 73893
rect 600272 73751 602172 73837
rect 600272 73695 600343 73751
rect 600399 73695 600485 73751
rect 600541 73695 600627 73751
rect 600683 73695 600769 73751
rect 600825 73695 600911 73751
rect 600967 73695 601053 73751
rect 601109 73695 601195 73751
rect 601251 73695 601337 73751
rect 601393 73695 601479 73751
rect 601535 73695 601621 73751
rect 601677 73695 601763 73751
rect 601819 73695 601905 73751
rect 601961 73695 602047 73751
rect 602103 73695 602172 73751
rect 600272 73609 602172 73695
rect 600272 73553 600343 73609
rect 600399 73553 600485 73609
rect 600541 73553 600627 73609
rect 600683 73553 600769 73609
rect 600825 73553 600911 73609
rect 600967 73553 601053 73609
rect 601109 73553 601195 73609
rect 601251 73553 601337 73609
rect 601393 73553 601479 73609
rect 601535 73553 601621 73609
rect 601677 73553 601763 73609
rect 601819 73553 601905 73609
rect 601961 73553 602047 73609
rect 602103 73553 602172 73609
rect 600272 73467 602172 73553
rect 600272 73411 600343 73467
rect 600399 73411 600485 73467
rect 600541 73411 600627 73467
rect 600683 73411 600769 73467
rect 600825 73411 600911 73467
rect 600967 73411 601053 73467
rect 601109 73411 601195 73467
rect 601251 73411 601337 73467
rect 601393 73411 601479 73467
rect 601535 73411 601621 73467
rect 601677 73411 601763 73467
rect 601819 73411 601905 73467
rect 601961 73411 602047 73467
rect 602103 73411 602172 73467
rect 600272 73325 602172 73411
rect 600272 73269 600343 73325
rect 600399 73269 600485 73325
rect 600541 73269 600627 73325
rect 600683 73269 600769 73325
rect 600825 73269 600911 73325
rect 600967 73269 601053 73325
rect 601109 73269 601195 73325
rect 601251 73269 601337 73325
rect 601393 73269 601479 73325
rect 601535 73269 601621 73325
rect 601677 73269 601763 73325
rect 601819 73269 601905 73325
rect 601961 73269 602047 73325
rect 602103 73269 602172 73325
rect 600272 73183 602172 73269
rect 600272 73127 600343 73183
rect 600399 73127 600485 73183
rect 600541 73127 600627 73183
rect 600683 73127 600769 73183
rect 600825 73127 600911 73183
rect 600967 73127 601053 73183
rect 601109 73127 601195 73183
rect 601251 73127 601337 73183
rect 601393 73127 601479 73183
rect 601535 73127 601621 73183
rect 601677 73127 601763 73183
rect 601819 73127 601905 73183
rect 601961 73127 602047 73183
rect 602103 73127 602172 73183
rect 600272 73041 602172 73127
rect 600272 72985 600343 73041
rect 600399 72985 600485 73041
rect 600541 72985 600627 73041
rect 600683 72985 600769 73041
rect 600825 72985 600911 73041
rect 600967 72985 601053 73041
rect 601109 72985 601195 73041
rect 601251 72985 601337 73041
rect 601393 72985 601479 73041
rect 601535 72985 601621 73041
rect 601677 72985 601763 73041
rect 601819 72985 601905 73041
rect 601961 72985 602047 73041
rect 602103 72985 602172 73041
rect 600272 72899 602172 72985
rect 600272 72843 600343 72899
rect 600399 72843 600485 72899
rect 600541 72843 600627 72899
rect 600683 72843 600769 72899
rect 600825 72843 600911 72899
rect 600967 72843 601053 72899
rect 601109 72843 601195 72899
rect 601251 72843 601337 72899
rect 601393 72843 601479 72899
rect 601535 72843 601621 72899
rect 601677 72843 601763 72899
rect 601819 72843 601905 72899
rect 601961 72843 602047 72899
rect 602103 72843 602172 72899
rect 600272 72757 602172 72843
rect 600272 72701 600343 72757
rect 600399 72701 600485 72757
rect 600541 72701 600627 72757
rect 600683 72701 600769 72757
rect 600825 72701 600911 72757
rect 600967 72701 601053 72757
rect 601109 72701 601195 72757
rect 601251 72701 601337 72757
rect 601393 72701 601479 72757
rect 601535 72701 601621 72757
rect 601677 72701 601763 72757
rect 601819 72701 601905 72757
rect 601961 72701 602047 72757
rect 602103 72701 602172 72757
rect 600272 72615 602172 72701
rect 600272 72559 600343 72615
rect 600399 72559 600485 72615
rect 600541 72559 600627 72615
rect 600683 72559 600769 72615
rect 600825 72559 600911 72615
rect 600967 72559 601053 72615
rect 601109 72559 601195 72615
rect 601251 72559 601337 72615
rect 601393 72559 601479 72615
rect 601535 72559 601621 72615
rect 601677 72559 601763 72615
rect 601819 72559 601905 72615
rect 601961 72559 602047 72615
rect 602103 72559 602172 72615
rect 600272 72473 602172 72559
rect 600272 72417 600343 72473
rect 600399 72417 600485 72473
rect 600541 72417 600627 72473
rect 600683 72417 600769 72473
rect 600825 72417 600911 72473
rect 600967 72417 601053 72473
rect 601109 72417 601195 72473
rect 601251 72417 601337 72473
rect 601393 72417 601479 72473
rect 601535 72417 601621 72473
rect 601677 72417 601763 72473
rect 601819 72417 601905 72473
rect 601961 72417 602047 72473
rect 602103 72417 602172 72473
rect 600272 72331 602172 72417
rect 600272 72275 600343 72331
rect 600399 72275 600485 72331
rect 600541 72275 600627 72331
rect 600683 72275 600769 72331
rect 600825 72275 600911 72331
rect 600967 72275 601053 72331
rect 601109 72275 601195 72331
rect 601251 72275 601337 72331
rect 601393 72275 601479 72331
rect 601535 72275 601621 72331
rect 601677 72275 601763 72331
rect 601819 72275 601905 72331
rect 601961 72275 602047 72331
rect 602103 72275 602172 72331
rect 600272 72189 602172 72275
rect 600272 72133 600343 72189
rect 600399 72133 600485 72189
rect 600541 72133 600627 72189
rect 600683 72133 600769 72189
rect 600825 72133 600911 72189
rect 600967 72133 601053 72189
rect 601109 72133 601195 72189
rect 601251 72133 601337 72189
rect 601393 72133 601479 72189
rect 601535 72133 601621 72189
rect 601677 72133 601763 72189
rect 601819 72133 601905 72189
rect 601961 72133 602047 72189
rect 602103 72133 602172 72189
rect 600272 72088 602172 72133
rect 602752 74035 604040 74088
rect 602752 73979 602823 74035
rect 602879 73979 602965 74035
rect 603021 73979 603107 74035
rect 603163 73979 603249 74035
rect 603305 73979 603391 74035
rect 603447 73979 603533 74035
rect 603589 73979 603675 74035
rect 603731 73979 603817 74035
rect 603873 73979 603959 74035
rect 604015 73979 604040 74035
rect 602752 73893 604040 73979
rect 602752 73837 602823 73893
rect 602879 73837 602965 73893
rect 603021 73837 603107 73893
rect 603163 73837 603249 73893
rect 603305 73837 603391 73893
rect 603447 73837 603533 73893
rect 603589 73837 603675 73893
rect 603731 73837 603817 73893
rect 603873 73837 603959 73893
rect 604015 73837 604040 73893
rect 602752 73751 604040 73837
rect 602752 73695 602823 73751
rect 602879 73695 602965 73751
rect 603021 73695 603107 73751
rect 603163 73695 603249 73751
rect 603305 73695 603391 73751
rect 603447 73695 603533 73751
rect 603589 73695 603675 73751
rect 603731 73695 603817 73751
rect 603873 73695 603959 73751
rect 604015 73695 604040 73751
rect 602752 73609 604040 73695
rect 602752 73553 602823 73609
rect 602879 73553 602965 73609
rect 603021 73553 603107 73609
rect 603163 73553 603249 73609
rect 603305 73553 603391 73609
rect 603447 73553 603533 73609
rect 603589 73553 603675 73609
rect 603731 73553 603817 73609
rect 603873 73553 603959 73609
rect 604015 73553 604040 73609
rect 602752 73467 604040 73553
rect 602752 73411 602823 73467
rect 602879 73411 602965 73467
rect 603021 73411 603107 73467
rect 603163 73411 603249 73467
rect 603305 73411 603391 73467
rect 603447 73411 603533 73467
rect 603589 73411 603675 73467
rect 603731 73411 603817 73467
rect 603873 73411 603959 73467
rect 604015 73411 604040 73467
rect 602752 73325 604040 73411
rect 602752 73269 602823 73325
rect 602879 73269 602965 73325
rect 603021 73269 603107 73325
rect 603163 73269 603249 73325
rect 603305 73269 603391 73325
rect 603447 73269 603533 73325
rect 603589 73269 603675 73325
rect 603731 73269 603817 73325
rect 603873 73269 603959 73325
rect 604015 73269 604040 73325
rect 602752 73183 604040 73269
rect 602752 73127 602823 73183
rect 602879 73127 602965 73183
rect 603021 73127 603107 73183
rect 603163 73127 603249 73183
rect 603305 73127 603391 73183
rect 603447 73127 603533 73183
rect 603589 73127 603675 73183
rect 603731 73127 603817 73183
rect 603873 73127 603959 73183
rect 604015 73127 604040 73183
rect 602752 73041 604040 73127
rect 602752 72985 602823 73041
rect 602879 72985 602965 73041
rect 603021 72985 603107 73041
rect 603163 72985 603249 73041
rect 603305 72985 603391 73041
rect 603447 72985 603533 73041
rect 603589 72985 603675 73041
rect 603731 72985 603817 73041
rect 603873 72985 603959 73041
rect 604015 72985 604040 73041
rect 602752 72899 604040 72985
rect 602752 72843 602823 72899
rect 602879 72843 602965 72899
rect 603021 72843 603107 72899
rect 603163 72843 603249 72899
rect 603305 72843 603391 72899
rect 603447 72843 603533 72899
rect 603589 72843 603675 72899
rect 603731 72843 603817 72899
rect 603873 72843 603959 72899
rect 604015 72843 604040 72899
rect 602752 72757 604040 72843
rect 602752 72701 602823 72757
rect 602879 72701 602965 72757
rect 603021 72701 603107 72757
rect 603163 72701 603249 72757
rect 603305 72701 603391 72757
rect 603447 72701 603533 72757
rect 603589 72701 603675 72757
rect 603731 72701 603817 72757
rect 603873 72701 603959 72757
rect 604015 72701 604040 72757
rect 602752 72615 604040 72701
rect 602752 72559 602823 72615
rect 602879 72559 602965 72615
rect 603021 72559 603107 72615
rect 603163 72559 603249 72615
rect 603305 72559 603391 72615
rect 603447 72559 603533 72615
rect 603589 72559 603675 72615
rect 603731 72559 603817 72615
rect 603873 72559 603959 72615
rect 604015 72559 604040 72615
rect 602752 72473 604040 72559
rect 602752 72417 602823 72473
rect 602879 72417 602965 72473
rect 603021 72417 603107 72473
rect 603163 72417 603249 72473
rect 603305 72417 603391 72473
rect 603447 72417 603533 72473
rect 603589 72417 603675 72473
rect 603731 72417 603817 72473
rect 603873 72417 603959 72473
rect 604015 72417 604040 72473
rect 602752 72331 604040 72417
rect 602752 72275 602823 72331
rect 602879 72275 602965 72331
rect 603021 72275 603107 72331
rect 603163 72275 603249 72331
rect 603305 72275 603391 72331
rect 603447 72275 603533 72331
rect 603589 72275 603675 72331
rect 603731 72275 603817 72331
rect 603873 72275 603959 72331
rect 604015 72275 604040 72331
rect 602752 72189 604040 72275
rect 602752 72133 602823 72189
rect 602879 72133 602965 72189
rect 603021 72133 603107 72189
rect 603163 72133 603249 72189
rect 603305 72133 603391 72189
rect 603447 72133 603533 72189
rect 603589 72133 603675 72189
rect 603731 72133 603817 72189
rect 603873 72133 603959 72189
rect 604015 72133 604040 72189
rect 602752 72088 604040 72133
rect 605122 74035 607172 74088
rect 605122 73979 605193 74035
rect 605249 73979 605335 74035
rect 605391 73979 605477 74035
rect 605533 73979 605619 74035
rect 605675 73979 605761 74035
rect 605817 73979 605903 74035
rect 605959 73979 606045 74035
rect 606101 73979 606187 74035
rect 606243 73979 606329 74035
rect 606385 73979 606471 74035
rect 606527 73979 606613 74035
rect 606669 73979 606755 74035
rect 606811 73979 606897 74035
rect 606953 73979 607039 74035
rect 607095 73979 607172 74035
rect 605122 73893 607172 73979
rect 605122 73837 605193 73893
rect 605249 73837 605335 73893
rect 605391 73837 605477 73893
rect 605533 73837 605619 73893
rect 605675 73837 605761 73893
rect 605817 73837 605903 73893
rect 605959 73837 606045 73893
rect 606101 73837 606187 73893
rect 606243 73837 606329 73893
rect 606385 73837 606471 73893
rect 606527 73837 606613 73893
rect 606669 73837 606755 73893
rect 606811 73837 606897 73893
rect 606953 73837 607039 73893
rect 607095 73837 607172 73893
rect 605122 73751 607172 73837
rect 605122 73695 605193 73751
rect 605249 73695 605335 73751
rect 605391 73695 605477 73751
rect 605533 73695 605619 73751
rect 605675 73695 605761 73751
rect 605817 73695 605903 73751
rect 605959 73695 606045 73751
rect 606101 73695 606187 73751
rect 606243 73695 606329 73751
rect 606385 73695 606471 73751
rect 606527 73695 606613 73751
rect 606669 73695 606755 73751
rect 606811 73695 606897 73751
rect 606953 73695 607039 73751
rect 607095 73695 607172 73751
rect 605122 73609 607172 73695
rect 605122 73553 605193 73609
rect 605249 73553 605335 73609
rect 605391 73553 605477 73609
rect 605533 73553 605619 73609
rect 605675 73553 605761 73609
rect 605817 73553 605903 73609
rect 605959 73553 606045 73609
rect 606101 73553 606187 73609
rect 606243 73553 606329 73609
rect 606385 73553 606471 73609
rect 606527 73553 606613 73609
rect 606669 73553 606755 73609
rect 606811 73553 606897 73609
rect 606953 73553 607039 73609
rect 607095 73553 607172 73609
rect 605122 73467 607172 73553
rect 605122 73411 605193 73467
rect 605249 73411 605335 73467
rect 605391 73411 605477 73467
rect 605533 73411 605619 73467
rect 605675 73411 605761 73467
rect 605817 73411 605903 73467
rect 605959 73411 606045 73467
rect 606101 73411 606187 73467
rect 606243 73411 606329 73467
rect 606385 73411 606471 73467
rect 606527 73411 606613 73467
rect 606669 73411 606755 73467
rect 606811 73411 606897 73467
rect 606953 73411 607039 73467
rect 607095 73411 607172 73467
rect 605122 73325 607172 73411
rect 605122 73269 605193 73325
rect 605249 73269 605335 73325
rect 605391 73269 605477 73325
rect 605533 73269 605619 73325
rect 605675 73269 605761 73325
rect 605817 73269 605903 73325
rect 605959 73269 606045 73325
rect 606101 73269 606187 73325
rect 606243 73269 606329 73325
rect 606385 73269 606471 73325
rect 606527 73269 606613 73325
rect 606669 73269 606755 73325
rect 606811 73269 606897 73325
rect 606953 73269 607039 73325
rect 607095 73269 607172 73325
rect 605122 73183 607172 73269
rect 605122 73127 605193 73183
rect 605249 73127 605335 73183
rect 605391 73127 605477 73183
rect 605533 73127 605619 73183
rect 605675 73127 605761 73183
rect 605817 73127 605903 73183
rect 605959 73127 606045 73183
rect 606101 73127 606187 73183
rect 606243 73127 606329 73183
rect 606385 73127 606471 73183
rect 606527 73127 606613 73183
rect 606669 73127 606755 73183
rect 606811 73127 606897 73183
rect 606953 73127 607039 73183
rect 607095 73127 607172 73183
rect 605122 73041 607172 73127
rect 605122 72985 605193 73041
rect 605249 72985 605335 73041
rect 605391 72985 605477 73041
rect 605533 72985 605619 73041
rect 605675 72985 605761 73041
rect 605817 72985 605903 73041
rect 605959 72985 606045 73041
rect 606101 72985 606187 73041
rect 606243 72985 606329 73041
rect 606385 72985 606471 73041
rect 606527 72985 606613 73041
rect 606669 72985 606755 73041
rect 606811 72985 606897 73041
rect 606953 72985 607039 73041
rect 607095 72985 607172 73041
rect 605122 72899 607172 72985
rect 605122 72843 605193 72899
rect 605249 72843 605335 72899
rect 605391 72843 605477 72899
rect 605533 72843 605619 72899
rect 605675 72843 605761 72899
rect 605817 72843 605903 72899
rect 605959 72843 606045 72899
rect 606101 72843 606187 72899
rect 606243 72843 606329 72899
rect 606385 72843 606471 72899
rect 606527 72843 606613 72899
rect 606669 72843 606755 72899
rect 606811 72843 606897 72899
rect 606953 72843 607039 72899
rect 607095 72843 607172 72899
rect 605122 72757 607172 72843
rect 605122 72701 605193 72757
rect 605249 72701 605335 72757
rect 605391 72701 605477 72757
rect 605533 72701 605619 72757
rect 605675 72701 605761 72757
rect 605817 72701 605903 72757
rect 605959 72701 606045 72757
rect 606101 72701 606187 72757
rect 606243 72701 606329 72757
rect 606385 72701 606471 72757
rect 606527 72701 606613 72757
rect 606669 72701 606755 72757
rect 606811 72701 606897 72757
rect 606953 72701 607039 72757
rect 607095 72701 607172 72757
rect 605122 72615 607172 72701
rect 605122 72559 605193 72615
rect 605249 72559 605335 72615
rect 605391 72559 605477 72615
rect 605533 72559 605619 72615
rect 605675 72559 605761 72615
rect 605817 72559 605903 72615
rect 605959 72559 606045 72615
rect 606101 72559 606187 72615
rect 606243 72559 606329 72615
rect 606385 72559 606471 72615
rect 606527 72559 606613 72615
rect 606669 72559 606755 72615
rect 606811 72559 606897 72615
rect 606953 72559 607039 72615
rect 607095 72559 607172 72615
rect 605122 72473 607172 72559
rect 605122 72417 605193 72473
rect 605249 72417 605335 72473
rect 605391 72417 605477 72473
rect 605533 72417 605619 72473
rect 605675 72417 605761 72473
rect 605817 72417 605903 72473
rect 605959 72417 606045 72473
rect 606101 72417 606187 72473
rect 606243 72417 606329 72473
rect 606385 72417 606471 72473
rect 606527 72417 606613 72473
rect 606669 72417 606755 72473
rect 606811 72417 606897 72473
rect 606953 72417 607039 72473
rect 607095 72417 607172 72473
rect 605122 72331 607172 72417
rect 605122 72275 605193 72331
rect 605249 72275 605335 72331
rect 605391 72275 605477 72331
rect 605533 72275 605619 72331
rect 605675 72275 605761 72331
rect 605817 72275 605903 72331
rect 605959 72275 606045 72331
rect 606101 72275 606187 72331
rect 606243 72275 606329 72331
rect 606385 72275 606471 72331
rect 606527 72275 606613 72331
rect 606669 72275 606755 72331
rect 606811 72275 606897 72331
rect 606953 72275 607039 72331
rect 607095 72275 607172 72331
rect 605122 72189 607172 72275
rect 605122 72133 605193 72189
rect 605249 72133 605335 72189
rect 605391 72133 605477 72189
rect 605533 72133 605619 72189
rect 605675 72133 605761 72189
rect 605817 72133 605903 72189
rect 605959 72133 606045 72189
rect 606101 72133 606187 72189
rect 606243 72133 606329 72189
rect 606385 72133 606471 72189
rect 606527 72133 606613 72189
rect 606669 72133 606755 72189
rect 606811 72133 606897 72189
rect 606953 72133 607039 72189
rect 607095 72133 607172 72189
rect 605122 72088 607172 72133
rect 607828 74035 609878 74088
rect 607828 73979 607899 74035
rect 607955 73979 608041 74035
rect 608097 73979 608183 74035
rect 608239 73979 608325 74035
rect 608381 73979 608467 74035
rect 608523 73979 608609 74035
rect 608665 73979 608751 74035
rect 608807 73979 608893 74035
rect 608949 73979 609035 74035
rect 609091 73979 609177 74035
rect 609233 73979 609319 74035
rect 609375 73979 609461 74035
rect 609517 73979 609603 74035
rect 609659 73979 609745 74035
rect 609801 73979 609878 74035
rect 607828 73893 609878 73979
rect 607828 73837 607899 73893
rect 607955 73837 608041 73893
rect 608097 73837 608183 73893
rect 608239 73837 608325 73893
rect 608381 73837 608467 73893
rect 608523 73837 608609 73893
rect 608665 73837 608751 73893
rect 608807 73837 608893 73893
rect 608949 73837 609035 73893
rect 609091 73837 609177 73893
rect 609233 73837 609319 73893
rect 609375 73837 609461 73893
rect 609517 73837 609603 73893
rect 609659 73837 609745 73893
rect 609801 73837 609878 73893
rect 607828 73751 609878 73837
rect 607828 73695 607899 73751
rect 607955 73695 608041 73751
rect 608097 73695 608183 73751
rect 608239 73695 608325 73751
rect 608381 73695 608467 73751
rect 608523 73695 608609 73751
rect 608665 73695 608751 73751
rect 608807 73695 608893 73751
rect 608949 73695 609035 73751
rect 609091 73695 609177 73751
rect 609233 73695 609319 73751
rect 609375 73695 609461 73751
rect 609517 73695 609603 73751
rect 609659 73695 609745 73751
rect 609801 73695 609878 73751
rect 607828 73609 609878 73695
rect 607828 73553 607899 73609
rect 607955 73553 608041 73609
rect 608097 73553 608183 73609
rect 608239 73553 608325 73609
rect 608381 73553 608467 73609
rect 608523 73553 608609 73609
rect 608665 73553 608751 73609
rect 608807 73553 608893 73609
rect 608949 73553 609035 73609
rect 609091 73553 609177 73609
rect 609233 73553 609319 73609
rect 609375 73553 609461 73609
rect 609517 73553 609603 73609
rect 609659 73553 609745 73609
rect 609801 73553 609878 73609
rect 607828 73467 609878 73553
rect 607828 73411 607899 73467
rect 607955 73411 608041 73467
rect 608097 73411 608183 73467
rect 608239 73411 608325 73467
rect 608381 73411 608467 73467
rect 608523 73411 608609 73467
rect 608665 73411 608751 73467
rect 608807 73411 608893 73467
rect 608949 73411 609035 73467
rect 609091 73411 609177 73467
rect 609233 73411 609319 73467
rect 609375 73411 609461 73467
rect 609517 73411 609603 73467
rect 609659 73411 609745 73467
rect 609801 73411 609878 73467
rect 607828 73325 609878 73411
rect 607828 73269 607899 73325
rect 607955 73269 608041 73325
rect 608097 73269 608183 73325
rect 608239 73269 608325 73325
rect 608381 73269 608467 73325
rect 608523 73269 608609 73325
rect 608665 73269 608751 73325
rect 608807 73269 608893 73325
rect 608949 73269 609035 73325
rect 609091 73269 609177 73325
rect 609233 73269 609319 73325
rect 609375 73269 609461 73325
rect 609517 73269 609603 73325
rect 609659 73269 609745 73325
rect 609801 73269 609878 73325
rect 607828 73183 609878 73269
rect 607828 73127 607899 73183
rect 607955 73127 608041 73183
rect 608097 73127 608183 73183
rect 608239 73127 608325 73183
rect 608381 73127 608467 73183
rect 608523 73127 608609 73183
rect 608665 73127 608751 73183
rect 608807 73127 608893 73183
rect 608949 73127 609035 73183
rect 609091 73127 609177 73183
rect 609233 73127 609319 73183
rect 609375 73127 609461 73183
rect 609517 73127 609603 73183
rect 609659 73127 609745 73183
rect 609801 73127 609878 73183
rect 607828 73041 609878 73127
rect 607828 72985 607899 73041
rect 607955 72985 608041 73041
rect 608097 72985 608183 73041
rect 608239 72985 608325 73041
rect 608381 72985 608467 73041
rect 608523 72985 608609 73041
rect 608665 72985 608751 73041
rect 608807 72985 608893 73041
rect 608949 72985 609035 73041
rect 609091 72985 609177 73041
rect 609233 72985 609319 73041
rect 609375 72985 609461 73041
rect 609517 72985 609603 73041
rect 609659 72985 609745 73041
rect 609801 72985 609878 73041
rect 607828 72899 609878 72985
rect 607828 72843 607899 72899
rect 607955 72843 608041 72899
rect 608097 72843 608183 72899
rect 608239 72843 608325 72899
rect 608381 72843 608467 72899
rect 608523 72843 608609 72899
rect 608665 72843 608751 72899
rect 608807 72843 608893 72899
rect 608949 72843 609035 72899
rect 609091 72843 609177 72899
rect 609233 72843 609319 72899
rect 609375 72843 609461 72899
rect 609517 72843 609603 72899
rect 609659 72843 609745 72899
rect 609801 72843 609878 72899
rect 607828 72757 609878 72843
rect 607828 72701 607899 72757
rect 607955 72701 608041 72757
rect 608097 72701 608183 72757
rect 608239 72701 608325 72757
rect 608381 72701 608467 72757
rect 608523 72701 608609 72757
rect 608665 72701 608751 72757
rect 608807 72701 608893 72757
rect 608949 72701 609035 72757
rect 609091 72701 609177 72757
rect 609233 72701 609319 72757
rect 609375 72701 609461 72757
rect 609517 72701 609603 72757
rect 609659 72701 609745 72757
rect 609801 72701 609878 72757
rect 607828 72615 609878 72701
rect 607828 72559 607899 72615
rect 607955 72559 608041 72615
rect 608097 72559 608183 72615
rect 608239 72559 608325 72615
rect 608381 72559 608467 72615
rect 608523 72559 608609 72615
rect 608665 72559 608751 72615
rect 608807 72559 608893 72615
rect 608949 72559 609035 72615
rect 609091 72559 609177 72615
rect 609233 72559 609319 72615
rect 609375 72559 609461 72615
rect 609517 72559 609603 72615
rect 609659 72559 609745 72615
rect 609801 72559 609878 72615
rect 607828 72473 609878 72559
rect 607828 72417 607899 72473
rect 607955 72417 608041 72473
rect 608097 72417 608183 72473
rect 608239 72417 608325 72473
rect 608381 72417 608467 72473
rect 608523 72417 608609 72473
rect 608665 72417 608751 72473
rect 608807 72417 608893 72473
rect 608949 72417 609035 72473
rect 609091 72417 609177 72473
rect 609233 72417 609319 72473
rect 609375 72417 609461 72473
rect 609517 72417 609603 72473
rect 609659 72417 609745 72473
rect 609801 72417 609878 72473
rect 607828 72331 609878 72417
rect 607828 72275 607899 72331
rect 607955 72275 608041 72331
rect 608097 72275 608183 72331
rect 608239 72275 608325 72331
rect 608381 72275 608467 72331
rect 608523 72275 608609 72331
rect 608665 72275 608751 72331
rect 608807 72275 608893 72331
rect 608949 72275 609035 72331
rect 609091 72275 609177 72331
rect 609233 72275 609319 72331
rect 609375 72275 609461 72331
rect 609517 72275 609603 72331
rect 609659 72275 609745 72331
rect 609801 72275 609878 72331
rect 607828 72189 609878 72275
rect 607828 72133 607899 72189
rect 607955 72133 608041 72189
rect 608097 72133 608183 72189
rect 608239 72133 608325 72189
rect 608381 72133 608467 72189
rect 608523 72133 608609 72189
rect 608665 72133 608751 72189
rect 608807 72133 608893 72189
rect 608949 72133 609035 72189
rect 609091 72133 609177 72189
rect 609233 72133 609319 72189
rect 609375 72133 609461 72189
rect 609517 72133 609603 72189
rect 609659 72133 609745 72189
rect 609801 72133 609878 72189
rect 607828 72088 609878 72133
rect 610198 74035 612248 74088
rect 610198 73979 610269 74035
rect 610325 73979 610411 74035
rect 610467 73979 610553 74035
rect 610609 73979 610695 74035
rect 610751 73979 610837 74035
rect 610893 73979 610979 74035
rect 611035 73979 611121 74035
rect 611177 73979 611263 74035
rect 611319 73979 611405 74035
rect 611461 73979 611547 74035
rect 611603 73979 611689 74035
rect 611745 73979 611831 74035
rect 611887 73979 611973 74035
rect 612029 73979 612115 74035
rect 612171 73979 612248 74035
rect 610198 73893 612248 73979
rect 610198 73837 610269 73893
rect 610325 73837 610411 73893
rect 610467 73837 610553 73893
rect 610609 73837 610695 73893
rect 610751 73837 610837 73893
rect 610893 73837 610979 73893
rect 611035 73837 611121 73893
rect 611177 73837 611263 73893
rect 611319 73837 611405 73893
rect 611461 73837 611547 73893
rect 611603 73837 611689 73893
rect 611745 73837 611831 73893
rect 611887 73837 611973 73893
rect 612029 73837 612115 73893
rect 612171 73837 612248 73893
rect 610198 73751 612248 73837
rect 610198 73695 610269 73751
rect 610325 73695 610411 73751
rect 610467 73695 610553 73751
rect 610609 73695 610695 73751
rect 610751 73695 610837 73751
rect 610893 73695 610979 73751
rect 611035 73695 611121 73751
rect 611177 73695 611263 73751
rect 611319 73695 611405 73751
rect 611461 73695 611547 73751
rect 611603 73695 611689 73751
rect 611745 73695 611831 73751
rect 611887 73695 611973 73751
rect 612029 73695 612115 73751
rect 612171 73695 612248 73751
rect 610198 73609 612248 73695
rect 610198 73553 610269 73609
rect 610325 73553 610411 73609
rect 610467 73553 610553 73609
rect 610609 73553 610695 73609
rect 610751 73553 610837 73609
rect 610893 73553 610979 73609
rect 611035 73553 611121 73609
rect 611177 73553 611263 73609
rect 611319 73553 611405 73609
rect 611461 73553 611547 73609
rect 611603 73553 611689 73609
rect 611745 73553 611831 73609
rect 611887 73553 611973 73609
rect 612029 73553 612115 73609
rect 612171 73553 612248 73609
rect 610198 73467 612248 73553
rect 610198 73411 610269 73467
rect 610325 73411 610411 73467
rect 610467 73411 610553 73467
rect 610609 73411 610695 73467
rect 610751 73411 610837 73467
rect 610893 73411 610979 73467
rect 611035 73411 611121 73467
rect 611177 73411 611263 73467
rect 611319 73411 611405 73467
rect 611461 73411 611547 73467
rect 611603 73411 611689 73467
rect 611745 73411 611831 73467
rect 611887 73411 611973 73467
rect 612029 73411 612115 73467
rect 612171 73411 612248 73467
rect 610198 73325 612248 73411
rect 610198 73269 610269 73325
rect 610325 73269 610411 73325
rect 610467 73269 610553 73325
rect 610609 73269 610695 73325
rect 610751 73269 610837 73325
rect 610893 73269 610979 73325
rect 611035 73269 611121 73325
rect 611177 73269 611263 73325
rect 611319 73269 611405 73325
rect 611461 73269 611547 73325
rect 611603 73269 611689 73325
rect 611745 73269 611831 73325
rect 611887 73269 611973 73325
rect 612029 73269 612115 73325
rect 612171 73269 612248 73325
rect 610198 73183 612248 73269
rect 610198 73127 610269 73183
rect 610325 73127 610411 73183
rect 610467 73127 610553 73183
rect 610609 73127 610695 73183
rect 610751 73127 610837 73183
rect 610893 73127 610979 73183
rect 611035 73127 611121 73183
rect 611177 73127 611263 73183
rect 611319 73127 611405 73183
rect 611461 73127 611547 73183
rect 611603 73127 611689 73183
rect 611745 73127 611831 73183
rect 611887 73127 611973 73183
rect 612029 73127 612115 73183
rect 612171 73127 612248 73183
rect 610198 73041 612248 73127
rect 610198 72985 610269 73041
rect 610325 72985 610411 73041
rect 610467 72985 610553 73041
rect 610609 72985 610695 73041
rect 610751 72985 610837 73041
rect 610893 72985 610979 73041
rect 611035 72985 611121 73041
rect 611177 72985 611263 73041
rect 611319 72985 611405 73041
rect 611461 72985 611547 73041
rect 611603 72985 611689 73041
rect 611745 72985 611831 73041
rect 611887 72985 611973 73041
rect 612029 72985 612115 73041
rect 612171 72985 612248 73041
rect 610198 72899 612248 72985
rect 610198 72843 610269 72899
rect 610325 72843 610411 72899
rect 610467 72843 610553 72899
rect 610609 72843 610695 72899
rect 610751 72843 610837 72899
rect 610893 72843 610979 72899
rect 611035 72843 611121 72899
rect 611177 72843 611263 72899
rect 611319 72843 611405 72899
rect 611461 72843 611547 72899
rect 611603 72843 611689 72899
rect 611745 72843 611831 72899
rect 611887 72843 611973 72899
rect 612029 72843 612115 72899
rect 612171 72843 612248 72899
rect 610198 72757 612248 72843
rect 610198 72701 610269 72757
rect 610325 72701 610411 72757
rect 610467 72701 610553 72757
rect 610609 72701 610695 72757
rect 610751 72701 610837 72757
rect 610893 72701 610979 72757
rect 611035 72701 611121 72757
rect 611177 72701 611263 72757
rect 611319 72701 611405 72757
rect 611461 72701 611547 72757
rect 611603 72701 611689 72757
rect 611745 72701 611831 72757
rect 611887 72701 611973 72757
rect 612029 72701 612115 72757
rect 612171 72701 612248 72757
rect 610198 72615 612248 72701
rect 610198 72559 610269 72615
rect 610325 72559 610411 72615
rect 610467 72559 610553 72615
rect 610609 72559 610695 72615
rect 610751 72559 610837 72615
rect 610893 72559 610979 72615
rect 611035 72559 611121 72615
rect 611177 72559 611263 72615
rect 611319 72559 611405 72615
rect 611461 72559 611547 72615
rect 611603 72559 611689 72615
rect 611745 72559 611831 72615
rect 611887 72559 611973 72615
rect 612029 72559 612115 72615
rect 612171 72559 612248 72615
rect 610198 72473 612248 72559
rect 610198 72417 610269 72473
rect 610325 72417 610411 72473
rect 610467 72417 610553 72473
rect 610609 72417 610695 72473
rect 610751 72417 610837 72473
rect 610893 72417 610979 72473
rect 611035 72417 611121 72473
rect 611177 72417 611263 72473
rect 611319 72417 611405 72473
rect 611461 72417 611547 72473
rect 611603 72417 611689 72473
rect 611745 72417 611831 72473
rect 611887 72417 611973 72473
rect 612029 72417 612115 72473
rect 612171 72417 612248 72473
rect 610198 72331 612248 72417
rect 610198 72275 610269 72331
rect 610325 72275 610411 72331
rect 610467 72275 610553 72331
rect 610609 72275 610695 72331
rect 610751 72275 610837 72331
rect 610893 72275 610979 72331
rect 611035 72275 611121 72331
rect 611177 72275 611263 72331
rect 611319 72275 611405 72331
rect 611461 72275 611547 72331
rect 611603 72275 611689 72331
rect 611745 72275 611831 72331
rect 611887 72275 611973 72331
rect 612029 72275 612115 72331
rect 612171 72275 612248 72331
rect 610198 72189 612248 72275
rect 610198 72133 610269 72189
rect 610325 72133 610411 72189
rect 610467 72133 610553 72189
rect 610609 72133 610695 72189
rect 610751 72133 610837 72189
rect 610893 72133 610979 72189
rect 611035 72133 611121 72189
rect 611177 72133 611263 72189
rect 611319 72133 611405 72189
rect 611461 72133 611547 72189
rect 611603 72133 611689 72189
rect 611745 72133 611831 72189
rect 611887 72133 611973 72189
rect 612029 72133 612115 72189
rect 612171 72133 612248 72189
rect 610198 72088 612248 72133
rect 612828 74035 614728 74088
rect 612828 73979 612899 74035
rect 612955 73979 613041 74035
rect 613097 73979 613183 74035
rect 613239 73979 613325 74035
rect 613381 73979 613467 74035
rect 613523 73979 613609 74035
rect 613665 73979 613751 74035
rect 613807 73979 613893 74035
rect 613949 73979 614035 74035
rect 614091 73979 614177 74035
rect 614233 73979 614319 74035
rect 614375 73979 614461 74035
rect 614517 73979 614603 74035
rect 614659 73979 614728 74035
rect 612828 73893 614728 73979
rect 612828 73837 612899 73893
rect 612955 73837 613041 73893
rect 613097 73837 613183 73893
rect 613239 73837 613325 73893
rect 613381 73837 613467 73893
rect 613523 73837 613609 73893
rect 613665 73837 613751 73893
rect 613807 73837 613893 73893
rect 613949 73837 614035 73893
rect 614091 73837 614177 73893
rect 614233 73837 614319 73893
rect 614375 73837 614461 73893
rect 614517 73837 614603 73893
rect 614659 73837 614728 73893
rect 612828 73751 614728 73837
rect 612828 73695 612899 73751
rect 612955 73695 613041 73751
rect 613097 73695 613183 73751
rect 613239 73695 613325 73751
rect 613381 73695 613467 73751
rect 613523 73695 613609 73751
rect 613665 73695 613751 73751
rect 613807 73695 613893 73751
rect 613949 73695 614035 73751
rect 614091 73695 614177 73751
rect 614233 73695 614319 73751
rect 614375 73695 614461 73751
rect 614517 73695 614603 73751
rect 614659 73695 614728 73751
rect 612828 73609 614728 73695
rect 612828 73553 612899 73609
rect 612955 73553 613041 73609
rect 613097 73553 613183 73609
rect 613239 73553 613325 73609
rect 613381 73553 613467 73609
rect 613523 73553 613609 73609
rect 613665 73553 613751 73609
rect 613807 73553 613893 73609
rect 613949 73553 614035 73609
rect 614091 73553 614177 73609
rect 614233 73553 614319 73609
rect 614375 73553 614461 73609
rect 614517 73553 614603 73609
rect 614659 73553 614728 73609
rect 612828 73467 614728 73553
rect 612828 73411 612899 73467
rect 612955 73411 613041 73467
rect 613097 73411 613183 73467
rect 613239 73411 613325 73467
rect 613381 73411 613467 73467
rect 613523 73411 613609 73467
rect 613665 73411 613751 73467
rect 613807 73411 613893 73467
rect 613949 73411 614035 73467
rect 614091 73411 614177 73467
rect 614233 73411 614319 73467
rect 614375 73411 614461 73467
rect 614517 73411 614603 73467
rect 614659 73411 614728 73467
rect 612828 73325 614728 73411
rect 612828 73269 612899 73325
rect 612955 73269 613041 73325
rect 613097 73269 613183 73325
rect 613239 73269 613325 73325
rect 613381 73269 613467 73325
rect 613523 73269 613609 73325
rect 613665 73269 613751 73325
rect 613807 73269 613893 73325
rect 613949 73269 614035 73325
rect 614091 73269 614177 73325
rect 614233 73269 614319 73325
rect 614375 73269 614461 73325
rect 614517 73269 614603 73325
rect 614659 73269 614728 73325
rect 612828 73183 614728 73269
rect 612828 73127 612899 73183
rect 612955 73127 613041 73183
rect 613097 73127 613183 73183
rect 613239 73127 613325 73183
rect 613381 73127 613467 73183
rect 613523 73127 613609 73183
rect 613665 73127 613751 73183
rect 613807 73127 613893 73183
rect 613949 73127 614035 73183
rect 614091 73127 614177 73183
rect 614233 73127 614319 73183
rect 614375 73127 614461 73183
rect 614517 73127 614603 73183
rect 614659 73127 614728 73183
rect 612828 73041 614728 73127
rect 612828 72985 612899 73041
rect 612955 72985 613041 73041
rect 613097 72985 613183 73041
rect 613239 72985 613325 73041
rect 613381 72985 613467 73041
rect 613523 72985 613609 73041
rect 613665 72985 613751 73041
rect 613807 72985 613893 73041
rect 613949 72985 614035 73041
rect 614091 72985 614177 73041
rect 614233 72985 614319 73041
rect 614375 72985 614461 73041
rect 614517 72985 614603 73041
rect 614659 72985 614728 73041
rect 612828 72899 614728 72985
rect 612828 72843 612899 72899
rect 612955 72843 613041 72899
rect 613097 72843 613183 72899
rect 613239 72843 613325 72899
rect 613381 72843 613467 72899
rect 613523 72843 613609 72899
rect 613665 72843 613751 72899
rect 613807 72843 613893 72899
rect 613949 72843 614035 72899
rect 614091 72843 614177 72899
rect 614233 72843 614319 72899
rect 614375 72843 614461 72899
rect 614517 72843 614603 72899
rect 614659 72843 614728 72899
rect 612828 72757 614728 72843
rect 612828 72701 612899 72757
rect 612955 72701 613041 72757
rect 613097 72701 613183 72757
rect 613239 72701 613325 72757
rect 613381 72701 613467 72757
rect 613523 72701 613609 72757
rect 613665 72701 613751 72757
rect 613807 72701 613893 72757
rect 613949 72701 614035 72757
rect 614091 72701 614177 72757
rect 614233 72701 614319 72757
rect 614375 72701 614461 72757
rect 614517 72701 614603 72757
rect 614659 72701 614728 72757
rect 612828 72615 614728 72701
rect 612828 72559 612899 72615
rect 612955 72559 613041 72615
rect 613097 72559 613183 72615
rect 613239 72559 613325 72615
rect 613381 72559 613467 72615
rect 613523 72559 613609 72615
rect 613665 72559 613751 72615
rect 613807 72559 613893 72615
rect 613949 72559 614035 72615
rect 614091 72559 614177 72615
rect 614233 72559 614319 72615
rect 614375 72559 614461 72615
rect 614517 72559 614603 72615
rect 614659 72559 614728 72615
rect 612828 72473 614728 72559
rect 612828 72417 612899 72473
rect 612955 72417 613041 72473
rect 613097 72417 613183 72473
rect 613239 72417 613325 72473
rect 613381 72417 613467 72473
rect 613523 72417 613609 72473
rect 613665 72417 613751 72473
rect 613807 72417 613893 72473
rect 613949 72417 614035 72473
rect 614091 72417 614177 72473
rect 614233 72417 614319 72473
rect 614375 72417 614461 72473
rect 614517 72417 614603 72473
rect 614659 72417 614728 72473
rect 612828 72331 614728 72417
rect 612828 72275 612899 72331
rect 612955 72275 613041 72331
rect 613097 72275 613183 72331
rect 613239 72275 613325 72331
rect 613381 72275 613467 72331
rect 613523 72275 613609 72331
rect 613665 72275 613751 72331
rect 613807 72275 613893 72331
rect 613949 72275 614035 72331
rect 614091 72275 614177 72331
rect 614233 72275 614319 72331
rect 614375 72275 614461 72331
rect 614517 72275 614603 72331
rect 614659 72275 614728 72331
rect 612828 72189 614728 72275
rect 612828 72133 612899 72189
rect 612955 72133 613041 72189
rect 613097 72133 613183 72189
rect 613239 72133 613325 72189
rect 613381 72133 613467 72189
rect 613523 72133 613609 72189
rect 613665 72133 613751 72189
rect 613807 72133 613893 72189
rect 613949 72133 614035 72189
rect 614091 72133 614177 72189
rect 614233 72133 614319 72189
rect 614375 72133 614461 72189
rect 614517 72133 614603 72189
rect 614659 72133 614728 72189
rect 612828 72088 614728 72133
<< via4 >>
rect 379341 941619 379397 941675
rect 379483 941619 379539 941675
rect 379625 941619 379681 941675
rect 379767 941619 379823 941675
rect 379909 941619 379965 941675
rect 379341 941477 379397 941533
rect 379483 941477 379539 941533
rect 379625 941477 379681 941533
rect 379767 941477 379823 941533
rect 379909 941477 379965 941533
rect 379341 941335 379397 941391
rect 379483 941335 379539 941391
rect 379625 941335 379681 941391
rect 379767 941335 379823 941391
rect 379909 941335 379965 941391
rect 379341 941193 379397 941249
rect 379483 941193 379539 941249
rect 379625 941193 379681 941249
rect 379767 941193 379823 941249
rect 379909 941193 379965 941249
rect 379341 941051 379397 941107
rect 379483 941051 379539 941107
rect 379625 941051 379681 941107
rect 379767 941051 379823 941107
rect 379909 941051 379965 941107
rect 379341 940909 379397 940965
rect 379483 940909 379539 940965
rect 379625 940909 379681 940965
rect 379767 940909 379823 940965
rect 379909 940909 379965 940965
rect 379341 940767 379397 940823
rect 379483 940767 379539 940823
rect 379625 940767 379681 940823
rect 379767 940767 379823 940823
rect 379909 940767 379965 940823
rect 379341 940625 379397 940681
rect 379483 940625 379539 940681
rect 379625 940625 379681 940681
rect 379767 940625 379823 940681
rect 379909 940625 379965 940681
rect 379341 940483 379397 940539
rect 379483 940483 379539 940539
rect 379625 940483 379681 940539
rect 379767 940483 379823 940539
rect 379909 940483 379965 940539
rect 379341 940341 379397 940397
rect 379483 940341 379539 940397
rect 379625 940341 379681 940397
rect 379767 940341 379823 940397
rect 379909 940341 379965 940397
rect 379341 940199 379397 940255
rect 379483 940199 379539 940255
rect 379625 940199 379681 940255
rect 379767 940199 379823 940255
rect 379909 940199 379965 940255
rect 379341 940057 379397 940113
rect 379483 940057 379539 940113
rect 379625 940057 379681 940113
rect 379767 940057 379823 940113
rect 379909 940057 379965 940113
rect 379341 939915 379397 939971
rect 379483 939915 379539 939971
rect 379625 939915 379681 939971
rect 379767 939915 379823 939971
rect 379909 939915 379965 939971
rect 379341 939773 379397 939829
rect 379483 939773 379539 939829
rect 379625 939773 379681 939829
rect 379767 939773 379823 939829
rect 379909 939773 379965 939829
rect 381829 941619 381885 941675
rect 381971 941619 382027 941675
rect 382113 941619 382169 941675
rect 382255 941619 382311 941675
rect 382397 941619 382453 941675
rect 382539 941619 382595 941675
rect 382681 941619 382737 941675
rect 382823 941619 382879 941675
rect 382965 941619 383021 941675
rect 383107 941619 383163 941675
rect 383249 941619 383305 941675
rect 383391 941619 383447 941675
rect 383533 941619 383589 941675
rect 383675 941619 383731 941675
rect 381829 941477 381885 941533
rect 381971 941477 382027 941533
rect 382113 941477 382169 941533
rect 382255 941477 382311 941533
rect 382397 941477 382453 941533
rect 382539 941477 382595 941533
rect 382681 941477 382737 941533
rect 382823 941477 382879 941533
rect 382965 941477 383021 941533
rect 383107 941477 383163 941533
rect 383249 941477 383305 941533
rect 383391 941477 383447 941533
rect 383533 941477 383589 941533
rect 383675 941477 383731 941533
rect 381829 941335 381885 941391
rect 381971 941335 382027 941391
rect 382113 941335 382169 941391
rect 382255 941335 382311 941391
rect 382397 941335 382453 941391
rect 382539 941335 382595 941391
rect 382681 941335 382737 941391
rect 382823 941335 382879 941391
rect 382965 941335 383021 941391
rect 383107 941335 383163 941391
rect 383249 941335 383305 941391
rect 383391 941335 383447 941391
rect 383533 941335 383589 941391
rect 383675 941335 383731 941391
rect 381829 941193 381885 941249
rect 381971 941193 382027 941249
rect 382113 941193 382169 941249
rect 382255 941193 382311 941249
rect 382397 941193 382453 941249
rect 382539 941193 382595 941249
rect 382681 941193 382737 941249
rect 382823 941193 382879 941249
rect 382965 941193 383021 941249
rect 383107 941193 383163 941249
rect 383249 941193 383305 941249
rect 383391 941193 383447 941249
rect 383533 941193 383589 941249
rect 383675 941193 383731 941249
rect 381829 941051 381885 941107
rect 381971 941051 382027 941107
rect 382113 941051 382169 941107
rect 382255 941051 382311 941107
rect 382397 941051 382453 941107
rect 382539 941051 382595 941107
rect 382681 941051 382737 941107
rect 382823 941051 382879 941107
rect 382965 941051 383021 941107
rect 383107 941051 383163 941107
rect 383249 941051 383305 941107
rect 383391 941051 383447 941107
rect 383533 941051 383589 941107
rect 383675 941051 383731 941107
rect 381829 940909 381885 940965
rect 381971 940909 382027 940965
rect 382113 940909 382169 940965
rect 382255 940909 382311 940965
rect 382397 940909 382453 940965
rect 382539 940909 382595 940965
rect 382681 940909 382737 940965
rect 382823 940909 382879 940965
rect 382965 940909 383021 940965
rect 383107 940909 383163 940965
rect 383249 940909 383305 940965
rect 383391 940909 383447 940965
rect 383533 940909 383589 940965
rect 383675 940909 383731 940965
rect 381829 940767 381885 940823
rect 381971 940767 382027 940823
rect 382113 940767 382169 940823
rect 382255 940767 382311 940823
rect 382397 940767 382453 940823
rect 382539 940767 382595 940823
rect 382681 940767 382737 940823
rect 382823 940767 382879 940823
rect 382965 940767 383021 940823
rect 383107 940767 383163 940823
rect 383249 940767 383305 940823
rect 383391 940767 383447 940823
rect 383533 940767 383589 940823
rect 383675 940767 383731 940823
rect 381829 940625 381885 940681
rect 381971 940625 382027 940681
rect 382113 940625 382169 940681
rect 382255 940625 382311 940681
rect 382397 940625 382453 940681
rect 382539 940625 382595 940681
rect 382681 940625 382737 940681
rect 382823 940625 382879 940681
rect 382965 940625 383021 940681
rect 383107 940625 383163 940681
rect 383249 940625 383305 940681
rect 383391 940625 383447 940681
rect 383533 940625 383589 940681
rect 383675 940625 383731 940681
rect 381829 940483 381885 940539
rect 381971 940483 382027 940539
rect 382113 940483 382169 940539
rect 382255 940483 382311 940539
rect 382397 940483 382453 940539
rect 382539 940483 382595 940539
rect 382681 940483 382737 940539
rect 382823 940483 382879 940539
rect 382965 940483 383021 940539
rect 383107 940483 383163 940539
rect 383249 940483 383305 940539
rect 383391 940483 383447 940539
rect 383533 940483 383589 940539
rect 383675 940483 383731 940539
rect 381829 940341 381885 940397
rect 381971 940341 382027 940397
rect 382113 940341 382169 940397
rect 382255 940341 382311 940397
rect 382397 940341 382453 940397
rect 382539 940341 382595 940397
rect 382681 940341 382737 940397
rect 382823 940341 382879 940397
rect 382965 940341 383021 940397
rect 383107 940341 383163 940397
rect 383249 940341 383305 940397
rect 383391 940341 383447 940397
rect 383533 940341 383589 940397
rect 383675 940341 383731 940397
rect 381829 940199 381885 940255
rect 381971 940199 382027 940255
rect 382113 940199 382169 940255
rect 382255 940199 382311 940255
rect 382397 940199 382453 940255
rect 382539 940199 382595 940255
rect 382681 940199 382737 940255
rect 382823 940199 382879 940255
rect 382965 940199 383021 940255
rect 383107 940199 383163 940255
rect 383249 940199 383305 940255
rect 383391 940199 383447 940255
rect 383533 940199 383589 940255
rect 383675 940199 383731 940255
rect 381829 940057 381885 940113
rect 381971 940057 382027 940113
rect 382113 940057 382169 940113
rect 382255 940057 382311 940113
rect 382397 940057 382453 940113
rect 382539 940057 382595 940113
rect 382681 940057 382737 940113
rect 382823 940057 382879 940113
rect 382965 940057 383021 940113
rect 383107 940057 383163 940113
rect 383249 940057 383305 940113
rect 383391 940057 383447 940113
rect 383533 940057 383589 940113
rect 383675 940057 383731 940113
rect 381829 939915 381885 939971
rect 381971 939915 382027 939971
rect 382113 939915 382169 939971
rect 382255 939915 382311 939971
rect 382397 939915 382453 939971
rect 382539 939915 382595 939971
rect 382681 939915 382737 939971
rect 382823 939915 382879 939971
rect 382965 939915 383021 939971
rect 383107 939915 383163 939971
rect 383249 939915 383305 939971
rect 383391 939915 383447 939971
rect 383533 939915 383589 939971
rect 383675 939915 383731 939971
rect 381829 939773 381885 939829
rect 381971 939773 382027 939829
rect 382113 939773 382169 939829
rect 382255 939773 382311 939829
rect 382397 939773 382453 939829
rect 382539 939773 382595 939829
rect 382681 939773 382737 939829
rect 382823 939773 382879 939829
rect 382965 939773 383021 939829
rect 383107 939773 383163 939829
rect 383249 939773 383305 939829
rect 383391 939773 383447 939829
rect 383533 939773 383589 939829
rect 383675 939773 383731 939829
rect 384199 941619 384255 941675
rect 384341 941619 384397 941675
rect 384483 941619 384539 941675
rect 385335 941619 385391 941675
rect 385477 941619 385533 941675
rect 385619 941619 385675 941675
rect 385761 941619 385817 941675
rect 385903 941619 385959 941675
rect 386045 941619 386101 941675
rect 384199 941477 384255 941533
rect 384341 941477 384397 941533
rect 384483 941477 384539 941533
rect 385335 941477 385391 941533
rect 385477 941477 385533 941533
rect 385619 941477 385675 941533
rect 385761 941477 385817 941533
rect 385903 941477 385959 941533
rect 386045 941477 386101 941533
rect 384199 941335 384255 941391
rect 384341 941335 384397 941391
rect 384483 941335 384539 941391
rect 385335 941335 385391 941391
rect 385477 941335 385533 941391
rect 385619 941335 385675 941391
rect 385761 941335 385817 941391
rect 385903 941335 385959 941391
rect 386045 941335 386101 941391
rect 384199 941193 384255 941249
rect 384341 941193 384397 941249
rect 384483 941193 384539 941249
rect 385335 941193 385391 941249
rect 385477 941193 385533 941249
rect 385619 941193 385675 941249
rect 385761 941193 385817 941249
rect 385903 941193 385959 941249
rect 386045 941193 386101 941249
rect 384199 941051 384255 941107
rect 384341 941051 384397 941107
rect 384483 941051 384539 941107
rect 385335 941051 385391 941107
rect 385477 941051 385533 941107
rect 385619 941051 385675 941107
rect 385761 941051 385817 941107
rect 385903 941051 385959 941107
rect 386045 941051 386101 941107
rect 384199 940909 384255 940965
rect 384341 940909 384397 940965
rect 384483 940909 384539 940965
rect 385335 940909 385391 940965
rect 385477 940909 385533 940965
rect 385619 940909 385675 940965
rect 385761 940909 385817 940965
rect 385903 940909 385959 940965
rect 386045 940909 386101 940965
rect 384199 940767 384255 940823
rect 384341 940767 384397 940823
rect 384483 940767 384539 940823
rect 385335 940767 385391 940823
rect 385477 940767 385533 940823
rect 385619 940767 385675 940823
rect 385761 940767 385817 940823
rect 385903 940767 385959 940823
rect 386045 940767 386101 940823
rect 384199 940625 384255 940681
rect 384341 940625 384397 940681
rect 384483 940625 384539 940681
rect 385335 940625 385391 940681
rect 385477 940625 385533 940681
rect 385619 940625 385675 940681
rect 385761 940625 385817 940681
rect 385903 940625 385959 940681
rect 386045 940625 386101 940681
rect 384199 940483 384255 940539
rect 384341 940483 384397 940539
rect 384483 940483 384539 940539
rect 385335 940483 385391 940539
rect 385477 940483 385533 940539
rect 385619 940483 385675 940539
rect 385761 940483 385817 940539
rect 385903 940483 385959 940539
rect 386045 940483 386101 940539
rect 384199 940341 384255 940397
rect 384341 940341 384397 940397
rect 384483 940341 384539 940397
rect 385335 940341 385391 940397
rect 385477 940341 385533 940397
rect 385619 940341 385675 940397
rect 385761 940341 385817 940397
rect 385903 940341 385959 940397
rect 386045 940341 386101 940397
rect 384199 940199 384255 940255
rect 384341 940199 384397 940255
rect 384483 940199 384539 940255
rect 385335 940199 385391 940255
rect 385477 940199 385533 940255
rect 385619 940199 385675 940255
rect 385761 940199 385817 940255
rect 385903 940199 385959 940255
rect 386045 940199 386101 940255
rect 384199 940057 384255 940113
rect 384341 940057 384397 940113
rect 384483 940057 384539 940113
rect 385335 940057 385391 940113
rect 385477 940057 385533 940113
rect 385619 940057 385675 940113
rect 385761 940057 385817 940113
rect 385903 940057 385959 940113
rect 386045 940057 386101 940113
rect 384199 939915 384255 939971
rect 384341 939915 384397 939971
rect 384483 939915 384539 939971
rect 385335 939915 385391 939971
rect 385477 939915 385533 939971
rect 385619 939915 385675 939971
rect 385761 939915 385817 939971
rect 385903 939915 385959 939971
rect 386045 939915 386101 939971
rect 384199 939773 384255 939829
rect 384341 939773 384397 939829
rect 384483 939773 384539 939829
rect 385335 939773 385391 939829
rect 385477 939773 385533 939829
rect 385619 939773 385675 939829
rect 385761 939773 385817 939829
rect 385903 939773 385959 939829
rect 386045 939773 386101 939829
rect 386905 941619 386961 941675
rect 387047 941619 387103 941675
rect 387189 941619 387245 941675
rect 387331 941619 387387 941675
rect 387473 941619 387529 941675
rect 387615 941619 387671 941675
rect 387757 941619 387813 941675
rect 387899 941619 387955 941675
rect 388041 941619 388097 941675
rect 388183 941619 388239 941675
rect 388325 941619 388381 941675
rect 388467 941619 388523 941675
rect 388609 941619 388665 941675
rect 388751 941619 388807 941675
rect 386905 941477 386961 941533
rect 387047 941477 387103 941533
rect 387189 941477 387245 941533
rect 387331 941477 387387 941533
rect 387473 941477 387529 941533
rect 387615 941477 387671 941533
rect 387757 941477 387813 941533
rect 387899 941477 387955 941533
rect 388041 941477 388097 941533
rect 388183 941477 388239 941533
rect 388325 941477 388381 941533
rect 388467 941477 388523 941533
rect 388609 941477 388665 941533
rect 388751 941477 388807 941533
rect 386905 941335 386961 941391
rect 387047 941335 387103 941391
rect 387189 941335 387245 941391
rect 387331 941335 387387 941391
rect 387473 941335 387529 941391
rect 387615 941335 387671 941391
rect 387757 941335 387813 941391
rect 387899 941335 387955 941391
rect 388041 941335 388097 941391
rect 388183 941335 388239 941391
rect 388325 941335 388381 941391
rect 388467 941335 388523 941391
rect 388609 941335 388665 941391
rect 388751 941335 388807 941391
rect 386905 941193 386961 941249
rect 387047 941193 387103 941249
rect 387189 941193 387245 941249
rect 387331 941193 387387 941249
rect 387473 941193 387529 941249
rect 387615 941193 387671 941249
rect 387757 941193 387813 941249
rect 387899 941193 387955 941249
rect 388041 941193 388097 941249
rect 388183 941193 388239 941249
rect 388325 941193 388381 941249
rect 388467 941193 388523 941249
rect 388609 941193 388665 941249
rect 388751 941193 388807 941249
rect 386905 941051 386961 941107
rect 387047 941051 387103 941107
rect 387189 941051 387245 941107
rect 387331 941051 387387 941107
rect 387473 941051 387529 941107
rect 387615 941051 387671 941107
rect 387757 941051 387813 941107
rect 387899 941051 387955 941107
rect 388041 941051 388097 941107
rect 388183 941051 388239 941107
rect 388325 941051 388381 941107
rect 388467 941051 388523 941107
rect 388609 941051 388665 941107
rect 388751 941051 388807 941107
rect 386905 940909 386961 940965
rect 387047 940909 387103 940965
rect 387189 940909 387245 940965
rect 387331 940909 387387 940965
rect 387473 940909 387529 940965
rect 387615 940909 387671 940965
rect 387757 940909 387813 940965
rect 387899 940909 387955 940965
rect 388041 940909 388097 940965
rect 388183 940909 388239 940965
rect 388325 940909 388381 940965
rect 388467 940909 388523 940965
rect 388609 940909 388665 940965
rect 388751 940909 388807 940965
rect 386905 940767 386961 940823
rect 387047 940767 387103 940823
rect 387189 940767 387245 940823
rect 387331 940767 387387 940823
rect 387473 940767 387529 940823
rect 387615 940767 387671 940823
rect 387757 940767 387813 940823
rect 387899 940767 387955 940823
rect 388041 940767 388097 940823
rect 388183 940767 388239 940823
rect 388325 940767 388381 940823
rect 388467 940767 388523 940823
rect 388609 940767 388665 940823
rect 388751 940767 388807 940823
rect 386905 940625 386961 940681
rect 387047 940625 387103 940681
rect 387189 940625 387245 940681
rect 387331 940625 387387 940681
rect 387473 940625 387529 940681
rect 387615 940625 387671 940681
rect 387757 940625 387813 940681
rect 387899 940625 387955 940681
rect 388041 940625 388097 940681
rect 388183 940625 388239 940681
rect 388325 940625 388381 940681
rect 388467 940625 388523 940681
rect 388609 940625 388665 940681
rect 388751 940625 388807 940681
rect 386905 940483 386961 940539
rect 387047 940483 387103 940539
rect 387189 940483 387245 940539
rect 387331 940483 387387 940539
rect 387473 940483 387529 940539
rect 387615 940483 387671 940539
rect 387757 940483 387813 940539
rect 387899 940483 387955 940539
rect 388041 940483 388097 940539
rect 388183 940483 388239 940539
rect 388325 940483 388381 940539
rect 388467 940483 388523 940539
rect 388609 940483 388665 940539
rect 388751 940483 388807 940539
rect 386905 940341 386961 940397
rect 387047 940341 387103 940397
rect 387189 940341 387245 940397
rect 387331 940341 387387 940397
rect 387473 940341 387529 940397
rect 387615 940341 387671 940397
rect 387757 940341 387813 940397
rect 387899 940341 387955 940397
rect 388041 940341 388097 940397
rect 388183 940341 388239 940397
rect 388325 940341 388381 940397
rect 388467 940341 388523 940397
rect 388609 940341 388665 940397
rect 388751 940341 388807 940397
rect 386905 940199 386961 940255
rect 387047 940199 387103 940255
rect 387189 940199 387245 940255
rect 387331 940199 387387 940255
rect 387473 940199 387529 940255
rect 387615 940199 387671 940255
rect 387757 940199 387813 940255
rect 387899 940199 387955 940255
rect 388041 940199 388097 940255
rect 388183 940199 388239 940255
rect 388325 940199 388381 940255
rect 388467 940199 388523 940255
rect 388609 940199 388665 940255
rect 388751 940199 388807 940255
rect 386905 940057 386961 940113
rect 387047 940057 387103 940113
rect 387189 940057 387245 940113
rect 387331 940057 387387 940113
rect 387473 940057 387529 940113
rect 387615 940057 387671 940113
rect 387757 940057 387813 940113
rect 387899 940057 387955 940113
rect 388041 940057 388097 940113
rect 388183 940057 388239 940113
rect 388325 940057 388381 940113
rect 388467 940057 388523 940113
rect 388609 940057 388665 940113
rect 388751 940057 388807 940113
rect 386905 939915 386961 939971
rect 387047 939915 387103 939971
rect 387189 939915 387245 939971
rect 387331 939915 387387 939971
rect 387473 939915 387529 939971
rect 387615 939915 387671 939971
rect 387757 939915 387813 939971
rect 387899 939915 387955 939971
rect 388041 939915 388097 939971
rect 388183 939915 388239 939971
rect 388325 939915 388381 939971
rect 388467 939915 388523 939971
rect 388609 939915 388665 939971
rect 388751 939915 388807 939971
rect 386905 939773 386961 939829
rect 387047 939773 387103 939829
rect 387189 939773 387245 939829
rect 387331 939773 387387 939829
rect 387473 939773 387529 939829
rect 387615 939773 387671 939829
rect 387757 939773 387813 939829
rect 387899 939773 387955 939829
rect 388041 939773 388097 939829
rect 388183 939773 388239 939829
rect 388325 939773 388381 939829
rect 388467 939773 388523 939829
rect 388609 939773 388665 939829
rect 388751 939773 388807 939829
rect 389275 941619 389331 941675
rect 389417 941619 389473 941675
rect 389559 941619 389615 941675
rect 389701 941619 389757 941675
rect 389843 941619 389899 941675
rect 389985 941619 390041 941675
rect 390127 941619 390183 941675
rect 390269 941619 390325 941675
rect 390411 941619 390467 941675
rect 390553 941619 390609 941675
rect 390695 941619 390751 941675
rect 390837 941619 390893 941675
rect 390979 941619 391035 941675
rect 391121 941619 391177 941675
rect 389275 941477 389331 941533
rect 389417 941477 389473 941533
rect 389559 941477 389615 941533
rect 389701 941477 389757 941533
rect 389843 941477 389899 941533
rect 389985 941477 390041 941533
rect 390127 941477 390183 941533
rect 390269 941477 390325 941533
rect 390411 941477 390467 941533
rect 390553 941477 390609 941533
rect 390695 941477 390751 941533
rect 390837 941477 390893 941533
rect 390979 941477 391035 941533
rect 391121 941477 391177 941533
rect 389275 941335 389331 941391
rect 389417 941335 389473 941391
rect 389559 941335 389615 941391
rect 389701 941335 389757 941391
rect 389843 941335 389899 941391
rect 389985 941335 390041 941391
rect 390127 941335 390183 941391
rect 390269 941335 390325 941391
rect 390411 941335 390467 941391
rect 390553 941335 390609 941391
rect 390695 941335 390751 941391
rect 390837 941335 390893 941391
rect 390979 941335 391035 941391
rect 391121 941335 391177 941391
rect 389275 941193 389331 941249
rect 389417 941193 389473 941249
rect 389559 941193 389615 941249
rect 389701 941193 389757 941249
rect 389843 941193 389899 941249
rect 389985 941193 390041 941249
rect 390127 941193 390183 941249
rect 390269 941193 390325 941249
rect 390411 941193 390467 941249
rect 390553 941193 390609 941249
rect 390695 941193 390751 941249
rect 390837 941193 390893 941249
rect 390979 941193 391035 941249
rect 391121 941193 391177 941249
rect 389275 941051 389331 941107
rect 389417 941051 389473 941107
rect 389559 941051 389615 941107
rect 389701 941051 389757 941107
rect 389843 941051 389899 941107
rect 389985 941051 390041 941107
rect 390127 941051 390183 941107
rect 390269 941051 390325 941107
rect 390411 941051 390467 941107
rect 390553 941051 390609 941107
rect 390695 941051 390751 941107
rect 390837 941051 390893 941107
rect 390979 941051 391035 941107
rect 391121 941051 391177 941107
rect 389275 940909 389331 940965
rect 389417 940909 389473 940965
rect 389559 940909 389615 940965
rect 389701 940909 389757 940965
rect 389843 940909 389899 940965
rect 389985 940909 390041 940965
rect 390127 940909 390183 940965
rect 390269 940909 390325 940965
rect 390411 940909 390467 940965
rect 390553 940909 390609 940965
rect 390695 940909 390751 940965
rect 390837 940909 390893 940965
rect 390979 940909 391035 940965
rect 391121 940909 391177 940965
rect 389275 940767 389331 940823
rect 389417 940767 389473 940823
rect 389559 940767 389615 940823
rect 389701 940767 389757 940823
rect 389843 940767 389899 940823
rect 389985 940767 390041 940823
rect 390127 940767 390183 940823
rect 390269 940767 390325 940823
rect 390411 940767 390467 940823
rect 390553 940767 390609 940823
rect 390695 940767 390751 940823
rect 390837 940767 390893 940823
rect 390979 940767 391035 940823
rect 391121 940767 391177 940823
rect 389275 940625 389331 940681
rect 389417 940625 389473 940681
rect 389559 940625 389615 940681
rect 389701 940625 389757 940681
rect 389843 940625 389899 940681
rect 389985 940625 390041 940681
rect 390127 940625 390183 940681
rect 390269 940625 390325 940681
rect 390411 940625 390467 940681
rect 390553 940625 390609 940681
rect 390695 940625 390751 940681
rect 390837 940625 390893 940681
rect 390979 940625 391035 940681
rect 391121 940625 391177 940681
rect 389275 940483 389331 940539
rect 389417 940483 389473 940539
rect 389559 940483 389615 940539
rect 389701 940483 389757 940539
rect 389843 940483 389899 940539
rect 389985 940483 390041 940539
rect 390127 940483 390183 940539
rect 390269 940483 390325 940539
rect 390411 940483 390467 940539
rect 390553 940483 390609 940539
rect 390695 940483 390751 940539
rect 390837 940483 390893 940539
rect 390979 940483 391035 940539
rect 391121 940483 391177 940539
rect 389275 940341 389331 940397
rect 389417 940341 389473 940397
rect 389559 940341 389615 940397
rect 389701 940341 389757 940397
rect 389843 940341 389899 940397
rect 389985 940341 390041 940397
rect 390127 940341 390183 940397
rect 390269 940341 390325 940397
rect 390411 940341 390467 940397
rect 390553 940341 390609 940397
rect 390695 940341 390751 940397
rect 390837 940341 390893 940397
rect 390979 940341 391035 940397
rect 391121 940341 391177 940397
rect 389275 940199 389331 940255
rect 389417 940199 389473 940255
rect 389559 940199 389615 940255
rect 389701 940199 389757 940255
rect 389843 940199 389899 940255
rect 389985 940199 390041 940255
rect 390127 940199 390183 940255
rect 390269 940199 390325 940255
rect 390411 940199 390467 940255
rect 390553 940199 390609 940255
rect 390695 940199 390751 940255
rect 390837 940199 390893 940255
rect 390979 940199 391035 940255
rect 391121 940199 391177 940255
rect 389275 940057 389331 940113
rect 389417 940057 389473 940113
rect 389559 940057 389615 940113
rect 389701 940057 389757 940113
rect 389843 940057 389899 940113
rect 389985 940057 390041 940113
rect 390127 940057 390183 940113
rect 390269 940057 390325 940113
rect 390411 940057 390467 940113
rect 390553 940057 390609 940113
rect 390695 940057 390751 940113
rect 390837 940057 390893 940113
rect 390979 940057 391035 940113
rect 391121 940057 391177 940113
rect 389275 939915 389331 939971
rect 389417 939915 389473 939971
rect 389559 939915 389615 939971
rect 389701 939915 389757 939971
rect 389843 939915 389899 939971
rect 389985 939915 390041 939971
rect 390127 939915 390183 939971
rect 390269 939915 390325 939971
rect 390411 939915 390467 939971
rect 390553 939915 390609 939971
rect 390695 939915 390751 939971
rect 390837 939915 390893 939971
rect 390979 939915 391035 939971
rect 391121 939915 391177 939971
rect 389275 939773 389331 939829
rect 389417 939773 389473 939829
rect 389559 939773 389615 939829
rect 389701 939773 389757 939829
rect 389843 939773 389899 939829
rect 389985 939773 390041 939829
rect 390127 939773 390183 939829
rect 390269 939773 390325 939829
rect 390411 939773 390467 939829
rect 390553 939773 390609 939829
rect 390695 939773 390751 939829
rect 390837 939773 390893 939829
rect 390979 939773 391035 939829
rect 391121 939773 391177 939829
rect 391897 941619 391953 941675
rect 392039 941619 392095 941675
rect 392181 941619 392237 941675
rect 392323 941619 392379 941675
rect 392465 941619 392521 941675
rect 392607 941619 392663 941675
rect 392749 941619 392805 941675
rect 392891 941619 392947 941675
rect 393033 941619 393089 941675
rect 393175 941619 393231 941675
rect 393317 941619 393373 941675
rect 393459 941619 393515 941675
rect 393601 941619 393657 941675
rect 391897 941477 391953 941533
rect 392039 941477 392095 941533
rect 392181 941477 392237 941533
rect 392323 941477 392379 941533
rect 392465 941477 392521 941533
rect 392607 941477 392663 941533
rect 392749 941477 392805 941533
rect 392891 941477 392947 941533
rect 393033 941477 393089 941533
rect 393175 941477 393231 941533
rect 393317 941477 393373 941533
rect 393459 941477 393515 941533
rect 393601 941477 393657 941533
rect 391897 941335 391953 941391
rect 392039 941335 392095 941391
rect 392181 941335 392237 941391
rect 392323 941335 392379 941391
rect 392465 941335 392521 941391
rect 392607 941335 392663 941391
rect 392749 941335 392805 941391
rect 392891 941335 392947 941391
rect 393033 941335 393089 941391
rect 393175 941335 393231 941391
rect 393317 941335 393373 941391
rect 393459 941335 393515 941391
rect 393601 941335 393657 941391
rect 391897 941193 391953 941249
rect 392039 941193 392095 941249
rect 392181 941193 392237 941249
rect 392323 941193 392379 941249
rect 392465 941193 392521 941249
rect 392607 941193 392663 941249
rect 392749 941193 392805 941249
rect 392891 941193 392947 941249
rect 393033 941193 393089 941249
rect 393175 941193 393231 941249
rect 393317 941193 393373 941249
rect 393459 941193 393515 941249
rect 393601 941193 393657 941249
rect 391897 941051 391953 941107
rect 392039 941051 392095 941107
rect 392181 941051 392237 941107
rect 392323 941051 392379 941107
rect 392465 941051 392521 941107
rect 392607 941051 392663 941107
rect 392749 941051 392805 941107
rect 392891 941051 392947 941107
rect 393033 941051 393089 941107
rect 393175 941051 393231 941107
rect 393317 941051 393373 941107
rect 393459 941051 393515 941107
rect 393601 941051 393657 941107
rect 391897 940909 391953 940965
rect 392039 940909 392095 940965
rect 392181 940909 392237 940965
rect 392323 940909 392379 940965
rect 392465 940909 392521 940965
rect 392607 940909 392663 940965
rect 392749 940909 392805 940965
rect 392891 940909 392947 940965
rect 393033 940909 393089 940965
rect 393175 940909 393231 940965
rect 393317 940909 393373 940965
rect 393459 940909 393515 940965
rect 393601 940909 393657 940965
rect 391897 940767 391953 940823
rect 392039 940767 392095 940823
rect 392181 940767 392237 940823
rect 392323 940767 392379 940823
rect 392465 940767 392521 940823
rect 392607 940767 392663 940823
rect 392749 940767 392805 940823
rect 392891 940767 392947 940823
rect 393033 940767 393089 940823
rect 393175 940767 393231 940823
rect 393317 940767 393373 940823
rect 393459 940767 393515 940823
rect 393601 940767 393657 940823
rect 391897 940625 391953 940681
rect 392039 940625 392095 940681
rect 392181 940625 392237 940681
rect 392323 940625 392379 940681
rect 392465 940625 392521 940681
rect 392607 940625 392663 940681
rect 392749 940625 392805 940681
rect 392891 940625 392947 940681
rect 393033 940625 393089 940681
rect 393175 940625 393231 940681
rect 393317 940625 393373 940681
rect 393459 940625 393515 940681
rect 393601 940625 393657 940681
rect 391897 940483 391953 940539
rect 392039 940483 392095 940539
rect 392181 940483 392237 940539
rect 392323 940483 392379 940539
rect 392465 940483 392521 940539
rect 392607 940483 392663 940539
rect 392749 940483 392805 940539
rect 392891 940483 392947 940539
rect 393033 940483 393089 940539
rect 393175 940483 393231 940539
rect 393317 940483 393373 940539
rect 393459 940483 393515 940539
rect 393601 940483 393657 940539
rect 391897 940341 391953 940397
rect 392039 940341 392095 940397
rect 392181 940341 392237 940397
rect 392323 940341 392379 940397
rect 392465 940341 392521 940397
rect 392607 940341 392663 940397
rect 392749 940341 392805 940397
rect 392891 940341 392947 940397
rect 393033 940341 393089 940397
rect 393175 940341 393231 940397
rect 393317 940341 393373 940397
rect 393459 940341 393515 940397
rect 393601 940341 393657 940397
rect 391897 940199 391953 940255
rect 392039 940199 392095 940255
rect 392181 940199 392237 940255
rect 392323 940199 392379 940255
rect 392465 940199 392521 940255
rect 392607 940199 392663 940255
rect 392749 940199 392805 940255
rect 392891 940199 392947 940255
rect 393033 940199 393089 940255
rect 393175 940199 393231 940255
rect 393317 940199 393373 940255
rect 393459 940199 393515 940255
rect 393601 940199 393657 940255
rect 391897 940057 391953 940113
rect 392039 940057 392095 940113
rect 392181 940057 392237 940113
rect 392323 940057 392379 940113
rect 392465 940057 392521 940113
rect 392607 940057 392663 940113
rect 392749 940057 392805 940113
rect 392891 940057 392947 940113
rect 393033 940057 393089 940113
rect 393175 940057 393231 940113
rect 393317 940057 393373 940113
rect 393459 940057 393515 940113
rect 393601 940057 393657 940113
rect 391897 939915 391953 939971
rect 392039 939915 392095 939971
rect 392181 939915 392237 939971
rect 392323 939915 392379 939971
rect 392465 939915 392521 939971
rect 392607 939915 392663 939971
rect 392749 939915 392805 939971
rect 392891 939915 392947 939971
rect 393033 939915 393089 939971
rect 393175 939915 393231 939971
rect 393317 939915 393373 939971
rect 393459 939915 393515 939971
rect 393601 939915 393657 939971
rect 391897 939773 391953 939829
rect 392039 939773 392095 939829
rect 392181 939773 392237 939829
rect 392323 939773 392379 939829
rect 392465 939773 392521 939829
rect 392607 939773 392663 939829
rect 392749 939773 392805 939829
rect 392891 939773 392947 939829
rect 393033 939773 393089 939829
rect 393175 939773 393231 939829
rect 393317 939773 393373 939829
rect 393459 939773 393515 939829
rect 393601 939773 393657 939829
rect 599341 941619 599397 941675
rect 599483 941619 599539 941675
rect 599625 941619 599681 941675
rect 599767 941619 599823 941675
rect 599909 941619 599965 941675
rect 600051 941619 600107 941675
rect 600193 941619 600249 941675
rect 600335 941619 600391 941675
rect 600477 941619 600533 941675
rect 600619 941619 600675 941675
rect 600761 941619 600817 941675
rect 600903 941619 600959 941675
rect 601045 941619 601101 941675
rect 599341 941477 599397 941533
rect 599483 941477 599539 941533
rect 599625 941477 599681 941533
rect 599767 941477 599823 941533
rect 599909 941477 599965 941533
rect 600051 941477 600107 941533
rect 600193 941477 600249 941533
rect 600335 941477 600391 941533
rect 600477 941477 600533 941533
rect 600619 941477 600675 941533
rect 600761 941477 600817 941533
rect 600903 941477 600959 941533
rect 601045 941477 601101 941533
rect 599341 941335 599397 941391
rect 599483 941335 599539 941391
rect 599625 941335 599681 941391
rect 599767 941335 599823 941391
rect 599909 941335 599965 941391
rect 600051 941335 600107 941391
rect 600193 941335 600249 941391
rect 600335 941335 600391 941391
rect 600477 941335 600533 941391
rect 600619 941335 600675 941391
rect 600761 941335 600817 941391
rect 600903 941335 600959 941391
rect 601045 941335 601101 941391
rect 599341 941193 599397 941249
rect 599483 941193 599539 941249
rect 599625 941193 599681 941249
rect 599767 941193 599823 941249
rect 599909 941193 599965 941249
rect 600051 941193 600107 941249
rect 600193 941193 600249 941249
rect 600335 941193 600391 941249
rect 600477 941193 600533 941249
rect 600619 941193 600675 941249
rect 600761 941193 600817 941249
rect 600903 941193 600959 941249
rect 601045 941193 601101 941249
rect 599341 941051 599397 941107
rect 599483 941051 599539 941107
rect 599625 941051 599681 941107
rect 599767 941051 599823 941107
rect 599909 941051 599965 941107
rect 600051 941051 600107 941107
rect 600193 941051 600249 941107
rect 600335 941051 600391 941107
rect 600477 941051 600533 941107
rect 600619 941051 600675 941107
rect 600761 941051 600817 941107
rect 600903 941051 600959 941107
rect 601045 941051 601101 941107
rect 599341 940909 599397 940965
rect 599483 940909 599539 940965
rect 599625 940909 599681 940965
rect 599767 940909 599823 940965
rect 599909 940909 599965 940965
rect 600051 940909 600107 940965
rect 600193 940909 600249 940965
rect 600335 940909 600391 940965
rect 600477 940909 600533 940965
rect 600619 940909 600675 940965
rect 600761 940909 600817 940965
rect 600903 940909 600959 940965
rect 601045 940909 601101 940965
rect 599341 940767 599397 940823
rect 599483 940767 599539 940823
rect 599625 940767 599681 940823
rect 599767 940767 599823 940823
rect 599909 940767 599965 940823
rect 600051 940767 600107 940823
rect 600193 940767 600249 940823
rect 600335 940767 600391 940823
rect 600477 940767 600533 940823
rect 600619 940767 600675 940823
rect 600761 940767 600817 940823
rect 600903 940767 600959 940823
rect 601045 940767 601101 940823
rect 599341 940625 599397 940681
rect 599483 940625 599539 940681
rect 599625 940625 599681 940681
rect 599767 940625 599823 940681
rect 599909 940625 599965 940681
rect 600051 940625 600107 940681
rect 600193 940625 600249 940681
rect 600335 940625 600391 940681
rect 600477 940625 600533 940681
rect 600619 940625 600675 940681
rect 600761 940625 600817 940681
rect 600903 940625 600959 940681
rect 601045 940625 601101 940681
rect 599341 940483 599397 940539
rect 599483 940483 599539 940539
rect 599625 940483 599681 940539
rect 599767 940483 599823 940539
rect 599909 940483 599965 940539
rect 600051 940483 600107 940539
rect 600193 940483 600249 940539
rect 600335 940483 600391 940539
rect 600477 940483 600533 940539
rect 600619 940483 600675 940539
rect 600761 940483 600817 940539
rect 600903 940483 600959 940539
rect 601045 940483 601101 940539
rect 599341 940341 599397 940397
rect 599483 940341 599539 940397
rect 599625 940341 599681 940397
rect 599767 940341 599823 940397
rect 599909 940341 599965 940397
rect 600051 940341 600107 940397
rect 600193 940341 600249 940397
rect 600335 940341 600391 940397
rect 600477 940341 600533 940397
rect 600619 940341 600675 940397
rect 600761 940341 600817 940397
rect 600903 940341 600959 940397
rect 601045 940341 601101 940397
rect 599341 940199 599397 940255
rect 599483 940199 599539 940255
rect 599625 940199 599681 940255
rect 599767 940199 599823 940255
rect 599909 940199 599965 940255
rect 600051 940199 600107 940255
rect 600193 940199 600249 940255
rect 600335 940199 600391 940255
rect 600477 940199 600533 940255
rect 600619 940199 600675 940255
rect 600761 940199 600817 940255
rect 600903 940199 600959 940255
rect 601045 940199 601101 940255
rect 599341 940057 599397 940113
rect 599483 940057 599539 940113
rect 599625 940057 599681 940113
rect 599767 940057 599823 940113
rect 599909 940057 599965 940113
rect 600051 940057 600107 940113
rect 600193 940057 600249 940113
rect 600335 940057 600391 940113
rect 600477 940057 600533 940113
rect 600619 940057 600675 940113
rect 600761 940057 600817 940113
rect 600903 940057 600959 940113
rect 601045 940057 601101 940113
rect 599341 939915 599397 939971
rect 599483 939915 599539 939971
rect 599625 939915 599681 939971
rect 599767 939915 599823 939971
rect 599909 939915 599965 939971
rect 600051 939915 600107 939971
rect 600193 939915 600249 939971
rect 600335 939915 600391 939971
rect 600477 939915 600533 939971
rect 600619 939915 600675 939971
rect 600761 939915 600817 939971
rect 600903 939915 600959 939971
rect 601045 939915 601101 939971
rect 599341 939773 599397 939829
rect 599483 939773 599539 939829
rect 599625 939773 599681 939829
rect 599767 939773 599823 939829
rect 599909 939773 599965 939829
rect 600051 939773 600107 939829
rect 600193 939773 600249 939829
rect 600335 939773 600391 939829
rect 600477 939773 600533 939829
rect 600619 939773 600675 939829
rect 600761 939773 600817 939829
rect 600903 939773 600959 939829
rect 601045 939773 601101 939829
rect 601829 941619 601885 941675
rect 601971 941619 602027 941675
rect 602113 941619 602169 941675
rect 602255 941619 602311 941675
rect 602397 941619 602453 941675
rect 602539 941619 602595 941675
rect 602681 941619 602737 941675
rect 602823 941619 602879 941675
rect 602965 941619 603021 941675
rect 603107 941619 603163 941675
rect 603249 941619 603305 941675
rect 603391 941619 603447 941675
rect 603533 941619 603589 941675
rect 603675 941619 603731 941675
rect 601829 941477 601885 941533
rect 601971 941477 602027 941533
rect 602113 941477 602169 941533
rect 602255 941477 602311 941533
rect 602397 941477 602453 941533
rect 602539 941477 602595 941533
rect 602681 941477 602737 941533
rect 602823 941477 602879 941533
rect 602965 941477 603021 941533
rect 603107 941477 603163 941533
rect 603249 941477 603305 941533
rect 603391 941477 603447 941533
rect 603533 941477 603589 941533
rect 603675 941477 603731 941533
rect 601829 941335 601885 941391
rect 601971 941335 602027 941391
rect 602113 941335 602169 941391
rect 602255 941335 602311 941391
rect 602397 941335 602453 941391
rect 602539 941335 602595 941391
rect 602681 941335 602737 941391
rect 602823 941335 602879 941391
rect 602965 941335 603021 941391
rect 603107 941335 603163 941391
rect 603249 941335 603305 941391
rect 603391 941335 603447 941391
rect 603533 941335 603589 941391
rect 603675 941335 603731 941391
rect 601829 941193 601885 941249
rect 601971 941193 602027 941249
rect 602113 941193 602169 941249
rect 602255 941193 602311 941249
rect 602397 941193 602453 941249
rect 602539 941193 602595 941249
rect 602681 941193 602737 941249
rect 602823 941193 602879 941249
rect 602965 941193 603021 941249
rect 603107 941193 603163 941249
rect 603249 941193 603305 941249
rect 603391 941193 603447 941249
rect 603533 941193 603589 941249
rect 603675 941193 603731 941249
rect 601829 941051 601885 941107
rect 601971 941051 602027 941107
rect 602113 941051 602169 941107
rect 602255 941051 602311 941107
rect 602397 941051 602453 941107
rect 602539 941051 602595 941107
rect 602681 941051 602737 941107
rect 602823 941051 602879 941107
rect 602965 941051 603021 941107
rect 603107 941051 603163 941107
rect 603249 941051 603305 941107
rect 603391 941051 603447 941107
rect 603533 941051 603589 941107
rect 603675 941051 603731 941107
rect 601829 940909 601885 940965
rect 601971 940909 602027 940965
rect 602113 940909 602169 940965
rect 602255 940909 602311 940965
rect 602397 940909 602453 940965
rect 602539 940909 602595 940965
rect 602681 940909 602737 940965
rect 602823 940909 602879 940965
rect 602965 940909 603021 940965
rect 603107 940909 603163 940965
rect 603249 940909 603305 940965
rect 603391 940909 603447 940965
rect 603533 940909 603589 940965
rect 603675 940909 603731 940965
rect 601829 940767 601885 940823
rect 601971 940767 602027 940823
rect 602113 940767 602169 940823
rect 602255 940767 602311 940823
rect 602397 940767 602453 940823
rect 602539 940767 602595 940823
rect 602681 940767 602737 940823
rect 602823 940767 602879 940823
rect 602965 940767 603021 940823
rect 603107 940767 603163 940823
rect 603249 940767 603305 940823
rect 603391 940767 603447 940823
rect 603533 940767 603589 940823
rect 603675 940767 603731 940823
rect 601829 940625 601885 940681
rect 601971 940625 602027 940681
rect 602113 940625 602169 940681
rect 602255 940625 602311 940681
rect 602397 940625 602453 940681
rect 602539 940625 602595 940681
rect 602681 940625 602737 940681
rect 602823 940625 602879 940681
rect 602965 940625 603021 940681
rect 603107 940625 603163 940681
rect 603249 940625 603305 940681
rect 603391 940625 603447 940681
rect 603533 940625 603589 940681
rect 603675 940625 603731 940681
rect 601829 940483 601885 940539
rect 601971 940483 602027 940539
rect 602113 940483 602169 940539
rect 602255 940483 602311 940539
rect 602397 940483 602453 940539
rect 602539 940483 602595 940539
rect 602681 940483 602737 940539
rect 602823 940483 602879 940539
rect 602965 940483 603021 940539
rect 603107 940483 603163 940539
rect 603249 940483 603305 940539
rect 603391 940483 603447 940539
rect 603533 940483 603589 940539
rect 603675 940483 603731 940539
rect 601829 940341 601885 940397
rect 601971 940341 602027 940397
rect 602113 940341 602169 940397
rect 602255 940341 602311 940397
rect 602397 940341 602453 940397
rect 602539 940341 602595 940397
rect 602681 940341 602737 940397
rect 602823 940341 602879 940397
rect 602965 940341 603021 940397
rect 603107 940341 603163 940397
rect 603249 940341 603305 940397
rect 603391 940341 603447 940397
rect 603533 940341 603589 940397
rect 603675 940341 603731 940397
rect 601829 940199 601885 940255
rect 601971 940199 602027 940255
rect 602113 940199 602169 940255
rect 602255 940199 602311 940255
rect 602397 940199 602453 940255
rect 602539 940199 602595 940255
rect 602681 940199 602737 940255
rect 602823 940199 602879 940255
rect 602965 940199 603021 940255
rect 603107 940199 603163 940255
rect 603249 940199 603305 940255
rect 603391 940199 603447 940255
rect 603533 940199 603589 940255
rect 603675 940199 603731 940255
rect 601829 940057 601885 940113
rect 601971 940057 602027 940113
rect 602113 940057 602169 940113
rect 602255 940057 602311 940113
rect 602397 940057 602453 940113
rect 602539 940057 602595 940113
rect 602681 940057 602737 940113
rect 602823 940057 602879 940113
rect 602965 940057 603021 940113
rect 603107 940057 603163 940113
rect 603249 940057 603305 940113
rect 603391 940057 603447 940113
rect 603533 940057 603589 940113
rect 603675 940057 603731 940113
rect 601829 939915 601885 939971
rect 601971 939915 602027 939971
rect 602113 939915 602169 939971
rect 602255 939915 602311 939971
rect 602397 939915 602453 939971
rect 602539 939915 602595 939971
rect 602681 939915 602737 939971
rect 602823 939915 602879 939971
rect 602965 939915 603021 939971
rect 603107 939915 603163 939971
rect 603249 939915 603305 939971
rect 603391 939915 603447 939971
rect 603533 939915 603589 939971
rect 603675 939915 603731 939971
rect 601829 939773 601885 939829
rect 601971 939773 602027 939829
rect 602113 939773 602169 939829
rect 602255 939773 602311 939829
rect 602397 939773 602453 939829
rect 602539 939773 602595 939829
rect 602681 939773 602737 939829
rect 602823 939773 602879 939829
rect 602965 939773 603021 939829
rect 603107 939773 603163 939829
rect 603249 939773 603305 939829
rect 603391 939773 603447 939829
rect 603533 939773 603589 939829
rect 603675 939773 603731 939829
rect 605051 941619 605107 941675
rect 605193 941619 605249 941675
rect 605335 941619 605391 941675
rect 605477 941619 605533 941675
rect 605619 941619 605675 941675
rect 605761 941619 605817 941675
rect 605903 941619 605959 941675
rect 606045 941619 606101 941675
rect 605051 941477 605107 941533
rect 605193 941477 605249 941533
rect 605335 941477 605391 941533
rect 605477 941477 605533 941533
rect 605619 941477 605675 941533
rect 605761 941477 605817 941533
rect 605903 941477 605959 941533
rect 606045 941477 606101 941533
rect 605051 941335 605107 941391
rect 605193 941335 605249 941391
rect 605335 941335 605391 941391
rect 605477 941335 605533 941391
rect 605619 941335 605675 941391
rect 605761 941335 605817 941391
rect 605903 941335 605959 941391
rect 606045 941335 606101 941391
rect 605051 941193 605107 941249
rect 605193 941193 605249 941249
rect 605335 941193 605391 941249
rect 605477 941193 605533 941249
rect 605619 941193 605675 941249
rect 605761 941193 605817 941249
rect 605903 941193 605959 941249
rect 606045 941193 606101 941249
rect 605051 941051 605107 941107
rect 605193 941051 605249 941107
rect 605335 941051 605391 941107
rect 605477 941051 605533 941107
rect 605619 941051 605675 941107
rect 605761 941051 605817 941107
rect 605903 941051 605959 941107
rect 606045 941051 606101 941107
rect 605051 940909 605107 940965
rect 605193 940909 605249 940965
rect 605335 940909 605391 940965
rect 605477 940909 605533 940965
rect 605619 940909 605675 940965
rect 605761 940909 605817 940965
rect 605903 940909 605959 940965
rect 606045 940909 606101 940965
rect 605051 940767 605107 940823
rect 605193 940767 605249 940823
rect 605335 940767 605391 940823
rect 605477 940767 605533 940823
rect 605619 940767 605675 940823
rect 605761 940767 605817 940823
rect 605903 940767 605959 940823
rect 606045 940767 606101 940823
rect 605051 940625 605107 940681
rect 605193 940625 605249 940681
rect 605335 940625 605391 940681
rect 605477 940625 605533 940681
rect 605619 940625 605675 940681
rect 605761 940625 605817 940681
rect 605903 940625 605959 940681
rect 606045 940625 606101 940681
rect 605051 940483 605107 940539
rect 605193 940483 605249 940539
rect 605335 940483 605391 940539
rect 605477 940483 605533 940539
rect 605619 940483 605675 940539
rect 605761 940483 605817 940539
rect 605903 940483 605959 940539
rect 606045 940483 606101 940539
rect 605051 940341 605107 940397
rect 605193 940341 605249 940397
rect 605335 940341 605391 940397
rect 605477 940341 605533 940397
rect 605619 940341 605675 940397
rect 605761 940341 605817 940397
rect 605903 940341 605959 940397
rect 606045 940341 606101 940397
rect 605051 940199 605107 940255
rect 605193 940199 605249 940255
rect 605335 940199 605391 940255
rect 605477 940199 605533 940255
rect 605619 940199 605675 940255
rect 605761 940199 605817 940255
rect 605903 940199 605959 940255
rect 606045 940199 606101 940255
rect 605051 940057 605107 940113
rect 605193 940057 605249 940113
rect 605335 940057 605391 940113
rect 605477 940057 605533 940113
rect 605619 940057 605675 940113
rect 605761 940057 605817 940113
rect 605903 940057 605959 940113
rect 606045 940057 606101 940113
rect 605051 939915 605107 939971
rect 605193 939915 605249 939971
rect 605335 939915 605391 939971
rect 605477 939915 605533 939971
rect 605619 939915 605675 939971
rect 605761 939915 605817 939971
rect 605903 939915 605959 939971
rect 606045 939915 606101 939971
rect 605051 939773 605107 939829
rect 605193 939773 605249 939829
rect 605335 939773 605391 939829
rect 605477 939773 605533 939829
rect 605619 939773 605675 939829
rect 605761 939773 605817 939829
rect 605903 939773 605959 939829
rect 606045 939773 606101 939829
rect 606905 941619 606961 941675
rect 607047 941619 607103 941675
rect 607189 941619 607245 941675
rect 607331 941619 607387 941675
rect 607473 941619 607529 941675
rect 607615 941619 607671 941675
rect 607757 941619 607813 941675
rect 607899 941619 607955 941675
rect 608041 941619 608097 941675
rect 608183 941619 608239 941675
rect 608325 941619 608381 941675
rect 608467 941619 608523 941675
rect 606905 941477 606961 941533
rect 607047 941477 607103 941533
rect 607189 941477 607245 941533
rect 607331 941477 607387 941533
rect 607473 941477 607529 941533
rect 607615 941477 607671 941533
rect 607757 941477 607813 941533
rect 607899 941477 607955 941533
rect 608041 941477 608097 941533
rect 608183 941477 608239 941533
rect 608325 941477 608381 941533
rect 608467 941477 608523 941533
rect 606905 941335 606961 941391
rect 607047 941335 607103 941391
rect 607189 941335 607245 941391
rect 607331 941335 607387 941391
rect 607473 941335 607529 941391
rect 607615 941335 607671 941391
rect 607757 941335 607813 941391
rect 607899 941335 607955 941391
rect 608041 941335 608097 941391
rect 608183 941335 608239 941391
rect 608325 941335 608381 941391
rect 608467 941335 608523 941391
rect 606905 941193 606961 941249
rect 607047 941193 607103 941249
rect 607189 941193 607245 941249
rect 607331 941193 607387 941249
rect 607473 941193 607529 941249
rect 607615 941193 607671 941249
rect 607757 941193 607813 941249
rect 607899 941193 607955 941249
rect 608041 941193 608097 941249
rect 608183 941193 608239 941249
rect 608325 941193 608381 941249
rect 608467 941193 608523 941249
rect 606905 941051 606961 941107
rect 607047 941051 607103 941107
rect 607189 941051 607245 941107
rect 607331 941051 607387 941107
rect 607473 941051 607529 941107
rect 607615 941051 607671 941107
rect 607757 941051 607813 941107
rect 607899 941051 607955 941107
rect 608041 941051 608097 941107
rect 608183 941051 608239 941107
rect 608325 941051 608381 941107
rect 608467 941051 608523 941107
rect 606905 940909 606961 940965
rect 607047 940909 607103 940965
rect 607189 940909 607245 940965
rect 607331 940909 607387 940965
rect 607473 940909 607529 940965
rect 607615 940909 607671 940965
rect 607757 940909 607813 940965
rect 607899 940909 607955 940965
rect 608041 940909 608097 940965
rect 608183 940909 608239 940965
rect 608325 940909 608381 940965
rect 608467 940909 608523 940965
rect 606905 940767 606961 940823
rect 607047 940767 607103 940823
rect 607189 940767 607245 940823
rect 607331 940767 607387 940823
rect 607473 940767 607529 940823
rect 607615 940767 607671 940823
rect 607757 940767 607813 940823
rect 607899 940767 607955 940823
rect 608041 940767 608097 940823
rect 608183 940767 608239 940823
rect 608325 940767 608381 940823
rect 608467 940767 608523 940823
rect 606905 940625 606961 940681
rect 607047 940625 607103 940681
rect 607189 940625 607245 940681
rect 607331 940625 607387 940681
rect 607473 940625 607529 940681
rect 607615 940625 607671 940681
rect 607757 940625 607813 940681
rect 607899 940625 607955 940681
rect 608041 940625 608097 940681
rect 608183 940625 608239 940681
rect 608325 940625 608381 940681
rect 608467 940625 608523 940681
rect 606905 940483 606961 940539
rect 607047 940483 607103 940539
rect 607189 940483 607245 940539
rect 607331 940483 607387 940539
rect 607473 940483 607529 940539
rect 607615 940483 607671 940539
rect 607757 940483 607813 940539
rect 607899 940483 607955 940539
rect 608041 940483 608097 940539
rect 608183 940483 608239 940539
rect 608325 940483 608381 940539
rect 608467 940483 608523 940539
rect 606905 940341 606961 940397
rect 607047 940341 607103 940397
rect 607189 940341 607245 940397
rect 607331 940341 607387 940397
rect 607473 940341 607529 940397
rect 607615 940341 607671 940397
rect 607757 940341 607813 940397
rect 607899 940341 607955 940397
rect 608041 940341 608097 940397
rect 608183 940341 608239 940397
rect 608325 940341 608381 940397
rect 608467 940341 608523 940397
rect 606905 940199 606961 940255
rect 607047 940199 607103 940255
rect 607189 940199 607245 940255
rect 607331 940199 607387 940255
rect 607473 940199 607529 940255
rect 607615 940199 607671 940255
rect 607757 940199 607813 940255
rect 607899 940199 607955 940255
rect 608041 940199 608097 940255
rect 608183 940199 608239 940255
rect 608325 940199 608381 940255
rect 608467 940199 608523 940255
rect 606905 940057 606961 940113
rect 607047 940057 607103 940113
rect 607189 940057 607245 940113
rect 607331 940057 607387 940113
rect 607473 940057 607529 940113
rect 607615 940057 607671 940113
rect 607757 940057 607813 940113
rect 607899 940057 607955 940113
rect 608041 940057 608097 940113
rect 608183 940057 608239 940113
rect 608325 940057 608381 940113
rect 608467 940057 608523 940113
rect 606905 939915 606961 939971
rect 607047 939915 607103 939971
rect 607189 939915 607245 939971
rect 607331 939915 607387 939971
rect 607473 939915 607529 939971
rect 607615 939915 607671 939971
rect 607757 939915 607813 939971
rect 607899 939915 607955 939971
rect 608041 939915 608097 939971
rect 608183 939915 608239 939971
rect 608325 939915 608381 939971
rect 608467 939915 608523 939971
rect 606905 939773 606961 939829
rect 607047 939773 607103 939829
rect 607189 939773 607245 939829
rect 607331 939773 607387 939829
rect 607473 939773 607529 939829
rect 607615 939773 607671 939829
rect 607757 939773 607813 939829
rect 607899 939773 607955 939829
rect 608041 939773 608097 939829
rect 608183 939773 608239 939829
rect 608325 939773 608381 939829
rect 608467 939773 608523 939829
rect 609275 941619 609331 941675
rect 609417 941619 609473 941675
rect 609559 941619 609615 941675
rect 609701 941619 609757 941675
rect 609843 941619 609899 941675
rect 609985 941619 610041 941675
rect 610127 941619 610183 941675
rect 610269 941619 610325 941675
rect 610411 941619 610467 941675
rect 610553 941619 610609 941675
rect 610695 941619 610751 941675
rect 610837 941619 610893 941675
rect 610979 941619 611035 941675
rect 611121 941619 611177 941675
rect 609275 941477 609331 941533
rect 609417 941477 609473 941533
rect 609559 941477 609615 941533
rect 609701 941477 609757 941533
rect 609843 941477 609899 941533
rect 609985 941477 610041 941533
rect 610127 941477 610183 941533
rect 610269 941477 610325 941533
rect 610411 941477 610467 941533
rect 610553 941477 610609 941533
rect 610695 941477 610751 941533
rect 610837 941477 610893 941533
rect 610979 941477 611035 941533
rect 611121 941477 611177 941533
rect 609275 941335 609331 941391
rect 609417 941335 609473 941391
rect 609559 941335 609615 941391
rect 609701 941335 609757 941391
rect 609843 941335 609899 941391
rect 609985 941335 610041 941391
rect 610127 941335 610183 941391
rect 610269 941335 610325 941391
rect 610411 941335 610467 941391
rect 610553 941335 610609 941391
rect 610695 941335 610751 941391
rect 610837 941335 610893 941391
rect 610979 941335 611035 941391
rect 611121 941335 611177 941391
rect 609275 941193 609331 941249
rect 609417 941193 609473 941249
rect 609559 941193 609615 941249
rect 609701 941193 609757 941249
rect 609843 941193 609899 941249
rect 609985 941193 610041 941249
rect 610127 941193 610183 941249
rect 610269 941193 610325 941249
rect 610411 941193 610467 941249
rect 610553 941193 610609 941249
rect 610695 941193 610751 941249
rect 610837 941193 610893 941249
rect 610979 941193 611035 941249
rect 611121 941193 611177 941249
rect 609275 941051 609331 941107
rect 609417 941051 609473 941107
rect 609559 941051 609615 941107
rect 609701 941051 609757 941107
rect 609843 941051 609899 941107
rect 609985 941051 610041 941107
rect 610127 941051 610183 941107
rect 610269 941051 610325 941107
rect 610411 941051 610467 941107
rect 610553 941051 610609 941107
rect 610695 941051 610751 941107
rect 610837 941051 610893 941107
rect 610979 941051 611035 941107
rect 611121 941051 611177 941107
rect 609275 940909 609331 940965
rect 609417 940909 609473 940965
rect 609559 940909 609615 940965
rect 609701 940909 609757 940965
rect 609843 940909 609899 940965
rect 609985 940909 610041 940965
rect 610127 940909 610183 940965
rect 610269 940909 610325 940965
rect 610411 940909 610467 940965
rect 610553 940909 610609 940965
rect 610695 940909 610751 940965
rect 610837 940909 610893 940965
rect 610979 940909 611035 940965
rect 611121 940909 611177 940965
rect 609275 940767 609331 940823
rect 609417 940767 609473 940823
rect 609559 940767 609615 940823
rect 609701 940767 609757 940823
rect 609843 940767 609899 940823
rect 609985 940767 610041 940823
rect 610127 940767 610183 940823
rect 610269 940767 610325 940823
rect 610411 940767 610467 940823
rect 610553 940767 610609 940823
rect 610695 940767 610751 940823
rect 610837 940767 610893 940823
rect 610979 940767 611035 940823
rect 611121 940767 611177 940823
rect 609275 940625 609331 940681
rect 609417 940625 609473 940681
rect 609559 940625 609615 940681
rect 609701 940625 609757 940681
rect 609843 940625 609899 940681
rect 609985 940625 610041 940681
rect 610127 940625 610183 940681
rect 610269 940625 610325 940681
rect 610411 940625 610467 940681
rect 610553 940625 610609 940681
rect 610695 940625 610751 940681
rect 610837 940625 610893 940681
rect 610979 940625 611035 940681
rect 611121 940625 611177 940681
rect 609275 940483 609331 940539
rect 609417 940483 609473 940539
rect 609559 940483 609615 940539
rect 609701 940483 609757 940539
rect 609843 940483 609899 940539
rect 609985 940483 610041 940539
rect 610127 940483 610183 940539
rect 610269 940483 610325 940539
rect 610411 940483 610467 940539
rect 610553 940483 610609 940539
rect 610695 940483 610751 940539
rect 610837 940483 610893 940539
rect 610979 940483 611035 940539
rect 611121 940483 611177 940539
rect 609275 940341 609331 940397
rect 609417 940341 609473 940397
rect 609559 940341 609615 940397
rect 609701 940341 609757 940397
rect 609843 940341 609899 940397
rect 609985 940341 610041 940397
rect 610127 940341 610183 940397
rect 610269 940341 610325 940397
rect 610411 940341 610467 940397
rect 610553 940341 610609 940397
rect 610695 940341 610751 940397
rect 610837 940341 610893 940397
rect 610979 940341 611035 940397
rect 611121 940341 611177 940397
rect 609275 940199 609331 940255
rect 609417 940199 609473 940255
rect 609559 940199 609615 940255
rect 609701 940199 609757 940255
rect 609843 940199 609899 940255
rect 609985 940199 610041 940255
rect 610127 940199 610183 940255
rect 610269 940199 610325 940255
rect 610411 940199 610467 940255
rect 610553 940199 610609 940255
rect 610695 940199 610751 940255
rect 610837 940199 610893 940255
rect 610979 940199 611035 940255
rect 611121 940199 611177 940255
rect 609275 940057 609331 940113
rect 609417 940057 609473 940113
rect 609559 940057 609615 940113
rect 609701 940057 609757 940113
rect 609843 940057 609899 940113
rect 609985 940057 610041 940113
rect 610127 940057 610183 940113
rect 610269 940057 610325 940113
rect 610411 940057 610467 940113
rect 610553 940057 610609 940113
rect 610695 940057 610751 940113
rect 610837 940057 610893 940113
rect 610979 940057 611035 940113
rect 611121 940057 611177 940113
rect 609275 939915 609331 939971
rect 609417 939915 609473 939971
rect 609559 939915 609615 939971
rect 609701 939915 609757 939971
rect 609843 939915 609899 939971
rect 609985 939915 610041 939971
rect 610127 939915 610183 939971
rect 610269 939915 610325 939971
rect 610411 939915 610467 939971
rect 610553 939915 610609 939971
rect 610695 939915 610751 939971
rect 610837 939915 610893 939971
rect 610979 939915 611035 939971
rect 611121 939915 611177 939971
rect 609275 939773 609331 939829
rect 609417 939773 609473 939829
rect 609559 939773 609615 939829
rect 609701 939773 609757 939829
rect 609843 939773 609899 939829
rect 609985 939773 610041 939829
rect 610127 939773 610183 939829
rect 610269 939773 610325 939829
rect 610411 939773 610467 939829
rect 610553 939773 610609 939829
rect 610695 939773 610751 939829
rect 610837 939773 610893 939829
rect 610979 939773 611035 939829
rect 611121 939773 611177 939829
rect 611897 941619 611953 941675
rect 612039 941619 612095 941675
rect 612181 941619 612237 941675
rect 612323 941619 612379 941675
rect 612465 941619 612521 941675
rect 612607 941619 612663 941675
rect 612749 941619 612805 941675
rect 612891 941619 612947 941675
rect 613033 941619 613089 941675
rect 613175 941619 613231 941675
rect 613317 941619 613373 941675
rect 613459 941619 613515 941675
rect 613601 941619 613657 941675
rect 611897 941477 611953 941533
rect 612039 941477 612095 941533
rect 612181 941477 612237 941533
rect 612323 941477 612379 941533
rect 612465 941477 612521 941533
rect 612607 941477 612663 941533
rect 612749 941477 612805 941533
rect 612891 941477 612947 941533
rect 613033 941477 613089 941533
rect 613175 941477 613231 941533
rect 613317 941477 613373 941533
rect 613459 941477 613515 941533
rect 613601 941477 613657 941533
rect 611897 941335 611953 941391
rect 612039 941335 612095 941391
rect 612181 941335 612237 941391
rect 612323 941335 612379 941391
rect 612465 941335 612521 941391
rect 612607 941335 612663 941391
rect 612749 941335 612805 941391
rect 612891 941335 612947 941391
rect 613033 941335 613089 941391
rect 613175 941335 613231 941391
rect 613317 941335 613373 941391
rect 613459 941335 613515 941391
rect 613601 941335 613657 941391
rect 611897 941193 611953 941249
rect 612039 941193 612095 941249
rect 612181 941193 612237 941249
rect 612323 941193 612379 941249
rect 612465 941193 612521 941249
rect 612607 941193 612663 941249
rect 612749 941193 612805 941249
rect 612891 941193 612947 941249
rect 613033 941193 613089 941249
rect 613175 941193 613231 941249
rect 613317 941193 613373 941249
rect 613459 941193 613515 941249
rect 613601 941193 613657 941249
rect 611897 941051 611953 941107
rect 612039 941051 612095 941107
rect 612181 941051 612237 941107
rect 612323 941051 612379 941107
rect 612465 941051 612521 941107
rect 612607 941051 612663 941107
rect 612749 941051 612805 941107
rect 612891 941051 612947 941107
rect 613033 941051 613089 941107
rect 613175 941051 613231 941107
rect 613317 941051 613373 941107
rect 613459 941051 613515 941107
rect 613601 941051 613657 941107
rect 611897 940909 611953 940965
rect 612039 940909 612095 940965
rect 612181 940909 612237 940965
rect 612323 940909 612379 940965
rect 612465 940909 612521 940965
rect 612607 940909 612663 940965
rect 612749 940909 612805 940965
rect 612891 940909 612947 940965
rect 613033 940909 613089 940965
rect 613175 940909 613231 940965
rect 613317 940909 613373 940965
rect 613459 940909 613515 940965
rect 613601 940909 613657 940965
rect 611897 940767 611953 940823
rect 612039 940767 612095 940823
rect 612181 940767 612237 940823
rect 612323 940767 612379 940823
rect 612465 940767 612521 940823
rect 612607 940767 612663 940823
rect 612749 940767 612805 940823
rect 612891 940767 612947 940823
rect 613033 940767 613089 940823
rect 613175 940767 613231 940823
rect 613317 940767 613373 940823
rect 613459 940767 613515 940823
rect 613601 940767 613657 940823
rect 611897 940625 611953 940681
rect 612039 940625 612095 940681
rect 612181 940625 612237 940681
rect 612323 940625 612379 940681
rect 612465 940625 612521 940681
rect 612607 940625 612663 940681
rect 612749 940625 612805 940681
rect 612891 940625 612947 940681
rect 613033 940625 613089 940681
rect 613175 940625 613231 940681
rect 613317 940625 613373 940681
rect 613459 940625 613515 940681
rect 613601 940625 613657 940681
rect 611897 940483 611953 940539
rect 612039 940483 612095 940539
rect 612181 940483 612237 940539
rect 612323 940483 612379 940539
rect 612465 940483 612521 940539
rect 612607 940483 612663 940539
rect 612749 940483 612805 940539
rect 612891 940483 612947 940539
rect 613033 940483 613089 940539
rect 613175 940483 613231 940539
rect 613317 940483 613373 940539
rect 613459 940483 613515 940539
rect 613601 940483 613657 940539
rect 611897 940341 611953 940397
rect 612039 940341 612095 940397
rect 612181 940341 612237 940397
rect 612323 940341 612379 940397
rect 612465 940341 612521 940397
rect 612607 940341 612663 940397
rect 612749 940341 612805 940397
rect 612891 940341 612947 940397
rect 613033 940341 613089 940397
rect 613175 940341 613231 940397
rect 613317 940341 613373 940397
rect 613459 940341 613515 940397
rect 613601 940341 613657 940397
rect 611897 940199 611953 940255
rect 612039 940199 612095 940255
rect 612181 940199 612237 940255
rect 612323 940199 612379 940255
rect 612465 940199 612521 940255
rect 612607 940199 612663 940255
rect 612749 940199 612805 940255
rect 612891 940199 612947 940255
rect 613033 940199 613089 940255
rect 613175 940199 613231 940255
rect 613317 940199 613373 940255
rect 613459 940199 613515 940255
rect 613601 940199 613657 940255
rect 611897 940057 611953 940113
rect 612039 940057 612095 940113
rect 612181 940057 612237 940113
rect 612323 940057 612379 940113
rect 612465 940057 612521 940113
rect 612607 940057 612663 940113
rect 612749 940057 612805 940113
rect 612891 940057 612947 940113
rect 613033 940057 613089 940113
rect 613175 940057 613231 940113
rect 613317 940057 613373 940113
rect 613459 940057 613515 940113
rect 613601 940057 613657 940113
rect 611897 939915 611953 939971
rect 612039 939915 612095 939971
rect 612181 939915 612237 939971
rect 612323 939915 612379 939971
rect 612465 939915 612521 939971
rect 612607 939915 612663 939971
rect 612749 939915 612805 939971
rect 612891 939915 612947 939971
rect 613033 939915 613089 939971
rect 613175 939915 613231 939971
rect 613317 939915 613373 939971
rect 613459 939915 613515 939971
rect 613601 939915 613657 939971
rect 611897 939773 611953 939829
rect 612039 939773 612095 939829
rect 612181 939773 612237 939829
rect 612323 939773 612379 939829
rect 612465 939773 612521 939829
rect 612607 939773 612663 939829
rect 612749 939773 612805 939829
rect 612891 939773 612947 939829
rect 613033 939773 613089 939829
rect 613175 939773 613231 939829
rect 613317 939773 613373 939829
rect 613459 939773 613515 939829
rect 613601 939773 613657 939829
rect 655343 75979 655399 76035
rect 655485 75979 655541 76035
rect 655627 75979 655683 76035
rect 655769 75979 655825 76035
rect 655911 75979 655967 76035
rect 656053 75979 656109 76035
rect 656195 75979 656251 76035
rect 656337 75979 656393 76035
rect 655343 75837 655399 75893
rect 655485 75837 655541 75893
rect 655627 75837 655683 75893
rect 655769 75837 655825 75893
rect 655911 75837 655967 75893
rect 656053 75837 656109 75893
rect 656195 75837 656251 75893
rect 656337 75837 656393 75893
rect 655343 75695 655399 75751
rect 655485 75695 655541 75751
rect 655627 75695 655683 75751
rect 655769 75695 655825 75751
rect 655911 75695 655967 75751
rect 656053 75695 656109 75751
rect 656195 75695 656251 75751
rect 656337 75695 656393 75751
rect 655343 75553 655399 75609
rect 655485 75553 655541 75609
rect 655627 75553 655683 75609
rect 655769 75553 655825 75609
rect 655911 75553 655967 75609
rect 656053 75553 656109 75609
rect 656195 75553 656251 75609
rect 656337 75553 656393 75609
rect 655343 75411 655399 75467
rect 655485 75411 655541 75467
rect 655627 75411 655683 75467
rect 655769 75411 655825 75467
rect 655911 75411 655967 75467
rect 656053 75411 656109 75467
rect 656195 75411 656251 75467
rect 656337 75411 656393 75467
rect 655343 75269 655399 75325
rect 655485 75269 655541 75325
rect 655627 75269 655683 75325
rect 655769 75269 655825 75325
rect 655911 75269 655967 75325
rect 656053 75269 656109 75325
rect 656195 75269 656251 75325
rect 656337 75269 656393 75325
rect 655343 75127 655399 75183
rect 655485 75127 655541 75183
rect 655627 75127 655683 75183
rect 655769 75127 655825 75183
rect 655911 75127 655967 75183
rect 656053 75127 656109 75183
rect 656195 75127 656251 75183
rect 656337 75127 656393 75183
rect 655343 74985 655399 75041
rect 655485 74985 655541 75041
rect 655627 74985 655683 75041
rect 655769 74985 655825 75041
rect 655911 74985 655967 75041
rect 656053 74985 656109 75041
rect 656195 74985 656251 75041
rect 656337 74985 656393 75041
rect 655343 74843 655399 74899
rect 655485 74843 655541 74899
rect 655627 74843 655683 74899
rect 655769 74843 655825 74899
rect 655911 74843 655967 74899
rect 656053 74843 656109 74899
rect 656195 74843 656251 74899
rect 656337 74843 656393 74899
rect 655343 74701 655399 74757
rect 655485 74701 655541 74757
rect 655627 74701 655683 74757
rect 655769 74701 655825 74757
rect 655911 74701 655967 74757
rect 656053 74701 656109 74757
rect 656195 74701 656251 74757
rect 656337 74701 656393 74757
rect 655343 74559 655399 74615
rect 655485 74559 655541 74615
rect 655627 74559 655683 74615
rect 655769 74559 655825 74615
rect 655911 74559 655967 74615
rect 656053 74559 656109 74615
rect 656195 74559 656251 74615
rect 656337 74559 656393 74615
rect 657823 75979 657879 76035
rect 657965 75979 658021 76035
rect 658107 75979 658163 76035
rect 658249 75979 658305 76035
rect 658391 75979 658447 76035
rect 658533 75979 658589 76035
rect 658675 75979 658731 76035
rect 658817 75979 658873 76035
rect 658959 75979 659015 76035
rect 659101 75979 659157 76035
rect 659243 75979 659299 76035
rect 659385 75979 659441 76035
rect 659527 75979 659583 76035
rect 659669 75979 659725 76035
rect 657823 75837 657879 75893
rect 657965 75837 658021 75893
rect 658107 75837 658163 75893
rect 658249 75837 658305 75893
rect 658391 75837 658447 75893
rect 658533 75837 658589 75893
rect 658675 75837 658731 75893
rect 658817 75837 658873 75893
rect 658959 75837 659015 75893
rect 659101 75837 659157 75893
rect 659243 75837 659299 75893
rect 659385 75837 659441 75893
rect 659527 75837 659583 75893
rect 659669 75837 659725 75893
rect 657823 75695 657879 75751
rect 657965 75695 658021 75751
rect 658107 75695 658163 75751
rect 658249 75695 658305 75751
rect 658391 75695 658447 75751
rect 658533 75695 658589 75751
rect 658675 75695 658731 75751
rect 658817 75695 658873 75751
rect 658959 75695 659015 75751
rect 659101 75695 659157 75751
rect 659243 75695 659299 75751
rect 659385 75695 659441 75751
rect 659527 75695 659583 75751
rect 659669 75695 659725 75751
rect 657823 75553 657879 75609
rect 657965 75553 658021 75609
rect 658107 75553 658163 75609
rect 658249 75553 658305 75609
rect 658391 75553 658447 75609
rect 658533 75553 658589 75609
rect 658675 75553 658731 75609
rect 658817 75553 658873 75609
rect 658959 75553 659015 75609
rect 659101 75553 659157 75609
rect 659243 75553 659299 75609
rect 659385 75553 659441 75609
rect 659527 75553 659583 75609
rect 659669 75553 659725 75609
rect 657823 75411 657879 75467
rect 657965 75411 658021 75467
rect 658107 75411 658163 75467
rect 658249 75411 658305 75467
rect 658391 75411 658447 75467
rect 658533 75411 658589 75467
rect 658675 75411 658731 75467
rect 658817 75411 658873 75467
rect 658959 75411 659015 75467
rect 659101 75411 659157 75467
rect 659243 75411 659299 75467
rect 659385 75411 659441 75467
rect 659527 75411 659583 75467
rect 659669 75411 659725 75467
rect 657823 75269 657879 75325
rect 657965 75269 658021 75325
rect 658107 75269 658163 75325
rect 658249 75269 658305 75325
rect 658391 75269 658447 75325
rect 658533 75269 658589 75325
rect 658675 75269 658731 75325
rect 658817 75269 658873 75325
rect 658959 75269 659015 75325
rect 659101 75269 659157 75325
rect 659243 75269 659299 75325
rect 659385 75269 659441 75325
rect 659527 75269 659583 75325
rect 659669 75269 659725 75325
rect 657823 75127 657879 75183
rect 657965 75127 658021 75183
rect 658107 75127 658163 75183
rect 658249 75127 658305 75183
rect 658391 75127 658447 75183
rect 658533 75127 658589 75183
rect 658675 75127 658731 75183
rect 658817 75127 658873 75183
rect 658959 75127 659015 75183
rect 659101 75127 659157 75183
rect 659243 75127 659299 75183
rect 659385 75127 659441 75183
rect 659527 75127 659583 75183
rect 659669 75127 659725 75183
rect 657823 74985 657879 75041
rect 657965 74985 658021 75041
rect 658107 74985 658163 75041
rect 658249 74985 658305 75041
rect 658391 74985 658447 75041
rect 658533 74985 658589 75041
rect 658675 74985 658731 75041
rect 658817 74985 658873 75041
rect 658959 74985 659015 75041
rect 659101 74985 659157 75041
rect 659243 74985 659299 75041
rect 659385 74985 659441 75041
rect 659527 74985 659583 75041
rect 659669 74985 659725 75041
rect 657823 74843 657879 74899
rect 657965 74843 658021 74899
rect 658107 74843 658163 74899
rect 658249 74843 658305 74899
rect 658391 74843 658447 74899
rect 658533 74843 658589 74899
rect 658675 74843 658731 74899
rect 658817 74843 658873 74899
rect 658959 74843 659015 74899
rect 659101 74843 659157 74899
rect 659243 74843 659299 74899
rect 659385 74843 659441 74899
rect 659527 74843 659583 74899
rect 659669 74843 659725 74899
rect 657823 74701 657879 74757
rect 657965 74701 658021 74757
rect 658107 74701 658163 74757
rect 658249 74701 658305 74757
rect 658391 74701 658447 74757
rect 658533 74701 658589 74757
rect 658675 74701 658731 74757
rect 658817 74701 658873 74757
rect 658959 74701 659015 74757
rect 659101 74701 659157 74757
rect 659243 74701 659299 74757
rect 659385 74701 659441 74757
rect 659527 74701 659583 74757
rect 659669 74701 659725 74757
rect 657823 74559 657879 74615
rect 657965 74559 658021 74615
rect 658107 74559 658163 74615
rect 658249 74559 658305 74615
rect 658391 74559 658447 74615
rect 658533 74559 658589 74615
rect 658675 74559 658731 74615
rect 658817 74559 658873 74615
rect 658959 74559 659015 74615
rect 659101 74559 659157 74615
rect 659243 74559 659299 74615
rect 659385 74559 659441 74615
rect 659527 74559 659583 74615
rect 659669 74559 659725 74615
rect 660193 75979 660249 76035
rect 660335 75979 660391 76035
rect 660477 75979 660533 76035
rect 660619 75979 660675 76035
rect 660761 75979 660817 76035
rect 660903 75979 660959 76035
rect 661045 75979 661101 76035
rect 661187 75979 661243 76035
rect 661329 75979 661385 76035
rect 661471 75979 661527 76035
rect 661613 75979 661669 76035
rect 661755 75979 661811 76035
rect 661897 75979 661953 76035
rect 662039 75979 662095 76035
rect 660193 75837 660249 75893
rect 660335 75837 660391 75893
rect 660477 75837 660533 75893
rect 660619 75837 660675 75893
rect 660761 75837 660817 75893
rect 660903 75837 660959 75893
rect 661045 75837 661101 75893
rect 661187 75837 661243 75893
rect 661329 75837 661385 75893
rect 661471 75837 661527 75893
rect 661613 75837 661669 75893
rect 661755 75837 661811 75893
rect 661897 75837 661953 75893
rect 662039 75837 662095 75893
rect 660193 75695 660249 75751
rect 660335 75695 660391 75751
rect 660477 75695 660533 75751
rect 660619 75695 660675 75751
rect 660761 75695 660817 75751
rect 660903 75695 660959 75751
rect 661045 75695 661101 75751
rect 661187 75695 661243 75751
rect 661329 75695 661385 75751
rect 661471 75695 661527 75751
rect 661613 75695 661669 75751
rect 661755 75695 661811 75751
rect 661897 75695 661953 75751
rect 662039 75695 662095 75751
rect 660193 75553 660249 75609
rect 660335 75553 660391 75609
rect 660477 75553 660533 75609
rect 660619 75553 660675 75609
rect 660761 75553 660817 75609
rect 660903 75553 660959 75609
rect 661045 75553 661101 75609
rect 661187 75553 661243 75609
rect 661329 75553 661385 75609
rect 661471 75553 661527 75609
rect 661613 75553 661669 75609
rect 661755 75553 661811 75609
rect 661897 75553 661953 75609
rect 662039 75553 662095 75609
rect 660193 75411 660249 75467
rect 660335 75411 660391 75467
rect 660477 75411 660533 75467
rect 660619 75411 660675 75467
rect 660761 75411 660817 75467
rect 660903 75411 660959 75467
rect 661045 75411 661101 75467
rect 661187 75411 661243 75467
rect 661329 75411 661385 75467
rect 661471 75411 661527 75467
rect 661613 75411 661669 75467
rect 661755 75411 661811 75467
rect 661897 75411 661953 75467
rect 662039 75411 662095 75467
rect 660193 75269 660249 75325
rect 660335 75269 660391 75325
rect 660477 75269 660533 75325
rect 660619 75269 660675 75325
rect 660761 75269 660817 75325
rect 660903 75269 660959 75325
rect 661045 75269 661101 75325
rect 661187 75269 661243 75325
rect 661329 75269 661385 75325
rect 661471 75269 661527 75325
rect 661613 75269 661669 75325
rect 661755 75269 661811 75325
rect 661897 75269 661953 75325
rect 662039 75269 662095 75325
rect 660193 75127 660249 75183
rect 660335 75127 660391 75183
rect 660477 75127 660533 75183
rect 660619 75127 660675 75183
rect 660761 75127 660817 75183
rect 660903 75127 660959 75183
rect 661045 75127 661101 75183
rect 661187 75127 661243 75183
rect 661329 75127 661385 75183
rect 661471 75127 661527 75183
rect 661613 75127 661669 75183
rect 661755 75127 661811 75183
rect 661897 75127 661953 75183
rect 662039 75127 662095 75183
rect 660193 74985 660249 75041
rect 660335 74985 660391 75041
rect 660477 74985 660533 75041
rect 660619 74985 660675 75041
rect 660761 74985 660817 75041
rect 660903 74985 660959 75041
rect 661045 74985 661101 75041
rect 661187 74985 661243 75041
rect 661329 74985 661385 75041
rect 661471 74985 661527 75041
rect 661613 74985 661669 75041
rect 661755 74985 661811 75041
rect 661897 74985 661953 75041
rect 662039 74985 662095 75041
rect 660193 74843 660249 74899
rect 660335 74843 660391 74899
rect 660477 74843 660533 74899
rect 660619 74843 660675 74899
rect 660761 74843 660817 74899
rect 660903 74843 660959 74899
rect 661045 74843 661101 74899
rect 661187 74843 661243 74899
rect 661329 74843 661385 74899
rect 661471 74843 661527 74899
rect 661613 74843 661669 74899
rect 661755 74843 661811 74899
rect 661897 74843 661953 74899
rect 662039 74843 662095 74899
rect 660193 74701 660249 74757
rect 660335 74701 660391 74757
rect 660477 74701 660533 74757
rect 660619 74701 660675 74757
rect 660761 74701 660817 74757
rect 660903 74701 660959 74757
rect 661045 74701 661101 74757
rect 661187 74701 661243 74757
rect 661329 74701 661385 74757
rect 661471 74701 661527 74757
rect 661613 74701 661669 74757
rect 661755 74701 661811 74757
rect 661897 74701 661953 74757
rect 662039 74701 662095 74757
rect 660193 74559 660249 74615
rect 660335 74559 660391 74615
rect 660477 74559 660533 74615
rect 660619 74559 660675 74615
rect 660761 74559 660817 74615
rect 660903 74559 660959 74615
rect 661045 74559 661101 74615
rect 661187 74559 661243 74615
rect 661329 74559 661385 74615
rect 661471 74559 661527 74615
rect 661613 74559 661669 74615
rect 661755 74559 661811 74615
rect 661897 74559 661953 74615
rect 662039 74559 662095 74615
rect 662899 75979 662955 76035
rect 663041 75979 663097 76035
rect 663183 75979 663239 76035
rect 663325 75979 663381 76035
rect 663467 75979 663523 76035
rect 663609 75979 663665 76035
rect 663751 75979 663807 76035
rect 663893 75979 663949 76035
rect 664035 75979 664091 76035
rect 664177 75979 664233 76035
rect 664319 75979 664375 76035
rect 664461 75979 664517 76035
rect 664603 75979 664659 76035
rect 664745 75979 664801 76035
rect 662899 75837 662955 75893
rect 663041 75837 663097 75893
rect 663183 75837 663239 75893
rect 663325 75837 663381 75893
rect 663467 75837 663523 75893
rect 663609 75837 663665 75893
rect 663751 75837 663807 75893
rect 663893 75837 663949 75893
rect 664035 75837 664091 75893
rect 664177 75837 664233 75893
rect 664319 75837 664375 75893
rect 664461 75837 664517 75893
rect 664603 75837 664659 75893
rect 664745 75837 664801 75893
rect 662899 75695 662955 75751
rect 663041 75695 663097 75751
rect 663183 75695 663239 75751
rect 663325 75695 663381 75751
rect 663467 75695 663523 75751
rect 663609 75695 663665 75751
rect 663751 75695 663807 75751
rect 663893 75695 663949 75751
rect 664035 75695 664091 75751
rect 664177 75695 664233 75751
rect 664319 75695 664375 75751
rect 664461 75695 664517 75751
rect 664603 75695 664659 75751
rect 664745 75695 664801 75751
rect 662899 75553 662955 75609
rect 663041 75553 663097 75609
rect 663183 75553 663239 75609
rect 663325 75553 663381 75609
rect 663467 75553 663523 75609
rect 663609 75553 663665 75609
rect 663751 75553 663807 75609
rect 663893 75553 663949 75609
rect 664035 75553 664091 75609
rect 664177 75553 664233 75609
rect 664319 75553 664375 75609
rect 664461 75553 664517 75609
rect 664603 75553 664659 75609
rect 664745 75553 664801 75609
rect 662899 75411 662955 75467
rect 663041 75411 663097 75467
rect 663183 75411 663239 75467
rect 663325 75411 663381 75467
rect 663467 75411 663523 75467
rect 663609 75411 663665 75467
rect 663751 75411 663807 75467
rect 663893 75411 663949 75467
rect 664035 75411 664091 75467
rect 664177 75411 664233 75467
rect 664319 75411 664375 75467
rect 664461 75411 664517 75467
rect 664603 75411 664659 75467
rect 664745 75411 664801 75467
rect 662899 75269 662955 75325
rect 663041 75269 663097 75325
rect 663183 75269 663239 75325
rect 663325 75269 663381 75325
rect 663467 75269 663523 75325
rect 663609 75269 663665 75325
rect 663751 75269 663807 75325
rect 663893 75269 663949 75325
rect 664035 75269 664091 75325
rect 664177 75269 664233 75325
rect 664319 75269 664375 75325
rect 664461 75269 664517 75325
rect 664603 75269 664659 75325
rect 664745 75269 664801 75325
rect 662899 75127 662955 75183
rect 663041 75127 663097 75183
rect 663183 75127 663239 75183
rect 663325 75127 663381 75183
rect 663467 75127 663523 75183
rect 663609 75127 663665 75183
rect 663751 75127 663807 75183
rect 663893 75127 663949 75183
rect 664035 75127 664091 75183
rect 664177 75127 664233 75183
rect 664319 75127 664375 75183
rect 664461 75127 664517 75183
rect 664603 75127 664659 75183
rect 664745 75127 664801 75183
rect 662899 74985 662955 75041
rect 663041 74985 663097 75041
rect 663183 74985 663239 75041
rect 663325 74985 663381 75041
rect 663467 74985 663523 75041
rect 663609 74985 663665 75041
rect 663751 74985 663807 75041
rect 663893 74985 663949 75041
rect 664035 74985 664091 75041
rect 664177 74985 664233 75041
rect 664319 74985 664375 75041
rect 664461 74985 664517 75041
rect 664603 74985 664659 75041
rect 664745 74985 664801 75041
rect 662899 74843 662955 74899
rect 663041 74843 663097 74899
rect 663183 74843 663239 74899
rect 663325 74843 663381 74899
rect 663467 74843 663523 74899
rect 663609 74843 663665 74899
rect 663751 74843 663807 74899
rect 663893 74843 663949 74899
rect 664035 74843 664091 74899
rect 664177 74843 664233 74899
rect 664319 74843 664375 74899
rect 664461 74843 664517 74899
rect 664603 74843 664659 74899
rect 664745 74843 664801 74899
rect 662899 74701 662955 74757
rect 663041 74701 663097 74757
rect 663183 74701 663239 74757
rect 663325 74701 663381 74757
rect 663467 74701 663523 74757
rect 663609 74701 663665 74757
rect 663751 74701 663807 74757
rect 663893 74701 663949 74757
rect 664035 74701 664091 74757
rect 664177 74701 664233 74757
rect 664319 74701 664375 74757
rect 664461 74701 664517 74757
rect 664603 74701 664659 74757
rect 664745 74701 664801 74757
rect 662899 74559 662955 74615
rect 663041 74559 663097 74615
rect 663183 74559 663239 74615
rect 663325 74559 663381 74615
rect 663467 74559 663523 74615
rect 663609 74559 663665 74615
rect 663751 74559 663807 74615
rect 663893 74559 663949 74615
rect 664035 74559 664091 74615
rect 664177 74559 664233 74615
rect 664319 74559 664375 74615
rect 664461 74559 664517 74615
rect 664603 74559 664659 74615
rect 664745 74559 664801 74615
rect 665269 75979 665325 76035
rect 665411 75979 665467 76035
rect 665553 75979 665609 76035
rect 665695 75979 665751 76035
rect 665837 75979 665893 76035
rect 665979 75979 666035 76035
rect 666121 75979 666177 76035
rect 666263 75979 666319 76035
rect 666405 75979 666461 76035
rect 666547 75979 666603 76035
rect 666689 75979 666745 76035
rect 666831 75979 666887 76035
rect 666973 75979 667029 76035
rect 667115 75979 667171 76035
rect 665269 75837 665325 75893
rect 665411 75837 665467 75893
rect 665553 75837 665609 75893
rect 665695 75837 665751 75893
rect 665837 75837 665893 75893
rect 665979 75837 666035 75893
rect 666121 75837 666177 75893
rect 666263 75837 666319 75893
rect 666405 75837 666461 75893
rect 666547 75837 666603 75893
rect 666689 75837 666745 75893
rect 666831 75837 666887 75893
rect 666973 75837 667029 75893
rect 667115 75837 667171 75893
rect 665269 75695 665325 75751
rect 665411 75695 665467 75751
rect 665553 75695 665609 75751
rect 665695 75695 665751 75751
rect 665837 75695 665893 75751
rect 665979 75695 666035 75751
rect 666121 75695 666177 75751
rect 666263 75695 666319 75751
rect 666405 75695 666461 75751
rect 666547 75695 666603 75751
rect 666689 75695 666745 75751
rect 666831 75695 666887 75751
rect 666973 75695 667029 75751
rect 667115 75695 667171 75751
rect 665269 75553 665325 75609
rect 665411 75553 665467 75609
rect 665553 75553 665609 75609
rect 665695 75553 665751 75609
rect 665837 75553 665893 75609
rect 665979 75553 666035 75609
rect 666121 75553 666177 75609
rect 666263 75553 666319 75609
rect 666405 75553 666461 75609
rect 666547 75553 666603 75609
rect 666689 75553 666745 75609
rect 666831 75553 666887 75609
rect 666973 75553 667029 75609
rect 667115 75553 667171 75609
rect 665269 75411 665325 75467
rect 665411 75411 665467 75467
rect 665553 75411 665609 75467
rect 665695 75411 665751 75467
rect 665837 75411 665893 75467
rect 665979 75411 666035 75467
rect 666121 75411 666177 75467
rect 666263 75411 666319 75467
rect 666405 75411 666461 75467
rect 666547 75411 666603 75467
rect 666689 75411 666745 75467
rect 666831 75411 666887 75467
rect 666973 75411 667029 75467
rect 667115 75411 667171 75467
rect 665269 75269 665325 75325
rect 665411 75269 665467 75325
rect 665553 75269 665609 75325
rect 665695 75269 665751 75325
rect 665837 75269 665893 75325
rect 665979 75269 666035 75325
rect 666121 75269 666177 75325
rect 666263 75269 666319 75325
rect 666405 75269 666461 75325
rect 666547 75269 666603 75325
rect 666689 75269 666745 75325
rect 666831 75269 666887 75325
rect 666973 75269 667029 75325
rect 667115 75269 667171 75325
rect 665269 75127 665325 75183
rect 665411 75127 665467 75183
rect 665553 75127 665609 75183
rect 665695 75127 665751 75183
rect 665837 75127 665893 75183
rect 665979 75127 666035 75183
rect 666121 75127 666177 75183
rect 666263 75127 666319 75183
rect 666405 75127 666461 75183
rect 666547 75127 666603 75183
rect 666689 75127 666745 75183
rect 666831 75127 666887 75183
rect 666973 75127 667029 75183
rect 667115 75127 667171 75183
rect 665269 74985 665325 75041
rect 665411 74985 665467 75041
rect 665553 74985 665609 75041
rect 665695 74985 665751 75041
rect 665837 74985 665893 75041
rect 665979 74985 666035 75041
rect 666121 74985 666177 75041
rect 666263 74985 666319 75041
rect 666405 74985 666461 75041
rect 666547 74985 666603 75041
rect 666689 74985 666745 75041
rect 666831 74985 666887 75041
rect 666973 74985 667029 75041
rect 667115 74985 667171 75041
rect 665269 74843 665325 74899
rect 665411 74843 665467 74899
rect 665553 74843 665609 74899
rect 665695 74843 665751 74899
rect 665837 74843 665893 74899
rect 665979 74843 666035 74899
rect 666121 74843 666177 74899
rect 666263 74843 666319 74899
rect 666405 74843 666461 74899
rect 666547 74843 666603 74899
rect 666689 74843 666745 74899
rect 666831 74843 666887 74899
rect 666973 74843 667029 74899
rect 667115 74843 667171 74899
rect 665269 74701 665325 74757
rect 665411 74701 665467 74757
rect 665553 74701 665609 74757
rect 665695 74701 665751 74757
rect 665837 74701 665893 74757
rect 665979 74701 666035 74757
rect 666121 74701 666177 74757
rect 666263 74701 666319 74757
rect 666405 74701 666461 74757
rect 666547 74701 666603 74757
rect 666689 74701 666745 74757
rect 666831 74701 666887 74757
rect 666973 74701 667029 74757
rect 667115 74701 667171 74757
rect 665269 74559 665325 74615
rect 665411 74559 665467 74615
rect 665553 74559 665609 74615
rect 665695 74559 665751 74615
rect 665837 74559 665893 74615
rect 665979 74559 666035 74615
rect 666121 74559 666177 74615
rect 666263 74559 666319 74615
rect 666405 74559 666461 74615
rect 666547 74559 666603 74615
rect 666689 74559 666745 74615
rect 666831 74559 666887 74615
rect 666973 74559 667029 74615
rect 667115 74559 667171 74615
rect 667899 75979 667955 76035
rect 668041 75979 668097 76035
rect 668893 75979 668949 76035
rect 669035 75979 669091 76035
rect 669177 75979 669233 76035
rect 669319 75979 669375 76035
rect 669461 75979 669517 76035
rect 669603 75979 669659 76035
rect 667899 75837 667955 75893
rect 668041 75837 668097 75893
rect 668893 75837 668949 75893
rect 669035 75837 669091 75893
rect 669177 75837 669233 75893
rect 669319 75837 669375 75893
rect 669461 75837 669517 75893
rect 669603 75837 669659 75893
rect 667899 75695 667955 75751
rect 668041 75695 668097 75751
rect 668893 75695 668949 75751
rect 669035 75695 669091 75751
rect 669177 75695 669233 75751
rect 669319 75695 669375 75751
rect 669461 75695 669517 75751
rect 669603 75695 669659 75751
rect 667899 75553 667955 75609
rect 668041 75553 668097 75609
rect 668893 75553 668949 75609
rect 669035 75553 669091 75609
rect 669177 75553 669233 75609
rect 669319 75553 669375 75609
rect 669461 75553 669517 75609
rect 669603 75553 669659 75609
rect 667899 75411 667955 75467
rect 668041 75411 668097 75467
rect 668893 75411 668949 75467
rect 669035 75411 669091 75467
rect 669177 75411 669233 75467
rect 669319 75411 669375 75467
rect 669461 75411 669517 75467
rect 669603 75411 669659 75467
rect 667899 75269 667955 75325
rect 668041 75269 668097 75325
rect 668893 75269 668949 75325
rect 669035 75269 669091 75325
rect 669177 75269 669233 75325
rect 669319 75269 669375 75325
rect 669461 75269 669517 75325
rect 669603 75269 669659 75325
rect 667899 75127 667955 75183
rect 668041 75127 668097 75183
rect 668893 75127 668949 75183
rect 669035 75127 669091 75183
rect 669177 75127 669233 75183
rect 669319 75127 669375 75183
rect 669461 75127 669517 75183
rect 669603 75127 669659 75183
rect 667899 74985 667955 75041
rect 668041 74985 668097 75041
rect 668893 74985 668949 75041
rect 669035 74985 669091 75041
rect 669177 74985 669233 75041
rect 669319 74985 669375 75041
rect 669461 74985 669517 75041
rect 669603 74985 669659 75041
rect 667899 74843 667955 74899
rect 668041 74843 668097 74899
rect 668893 74843 668949 74899
rect 669035 74843 669091 74899
rect 669177 74843 669233 74899
rect 669319 74843 669375 74899
rect 669461 74843 669517 74899
rect 669603 74843 669659 74899
rect 667899 74701 667955 74757
rect 668041 74701 668097 74757
rect 668893 74701 668949 74757
rect 669035 74701 669091 74757
rect 669177 74701 669233 74757
rect 669319 74701 669375 74757
rect 669461 74701 669517 74757
rect 669603 74701 669659 74757
rect 667899 74559 667955 74615
rect 668041 74559 668097 74615
rect 668893 74559 668949 74615
rect 669035 74559 669091 74615
rect 669177 74559 669233 74615
rect 669319 74559 669375 74615
rect 669461 74559 669517 74615
rect 669603 74559 669659 74615
rect 105343 73979 105399 74035
rect 105485 73979 105541 74035
rect 105627 73979 105683 74035
rect 105769 73979 105825 74035
rect 105911 73979 105967 74035
rect 106053 73979 106109 74035
rect 106195 73979 106251 74035
rect 106337 73979 106393 74035
rect 106479 73979 106535 74035
rect 106621 73979 106677 74035
rect 106763 73979 106819 74035
rect 106905 73979 106961 74035
rect 107047 73979 107103 74035
rect 105343 73837 105399 73893
rect 105485 73837 105541 73893
rect 105627 73837 105683 73893
rect 105769 73837 105825 73893
rect 105911 73837 105967 73893
rect 106053 73837 106109 73893
rect 106195 73837 106251 73893
rect 106337 73837 106393 73893
rect 106479 73837 106535 73893
rect 106621 73837 106677 73893
rect 106763 73837 106819 73893
rect 106905 73837 106961 73893
rect 107047 73837 107103 73893
rect 105343 73695 105399 73751
rect 105485 73695 105541 73751
rect 105627 73695 105683 73751
rect 105769 73695 105825 73751
rect 105911 73695 105967 73751
rect 106053 73695 106109 73751
rect 106195 73695 106251 73751
rect 106337 73695 106393 73751
rect 106479 73695 106535 73751
rect 106621 73695 106677 73751
rect 106763 73695 106819 73751
rect 106905 73695 106961 73751
rect 107047 73695 107103 73751
rect 105343 73553 105399 73609
rect 105485 73553 105541 73609
rect 105627 73553 105683 73609
rect 105769 73553 105825 73609
rect 105911 73553 105967 73609
rect 106053 73553 106109 73609
rect 106195 73553 106251 73609
rect 106337 73553 106393 73609
rect 106479 73553 106535 73609
rect 106621 73553 106677 73609
rect 106763 73553 106819 73609
rect 106905 73553 106961 73609
rect 107047 73553 107103 73609
rect 105343 73411 105399 73467
rect 105485 73411 105541 73467
rect 105627 73411 105683 73467
rect 105769 73411 105825 73467
rect 105911 73411 105967 73467
rect 106053 73411 106109 73467
rect 106195 73411 106251 73467
rect 106337 73411 106393 73467
rect 106479 73411 106535 73467
rect 106621 73411 106677 73467
rect 106763 73411 106819 73467
rect 106905 73411 106961 73467
rect 107047 73411 107103 73467
rect 105343 73269 105399 73325
rect 105485 73269 105541 73325
rect 105627 73269 105683 73325
rect 105769 73269 105825 73325
rect 105911 73269 105967 73325
rect 106053 73269 106109 73325
rect 106195 73269 106251 73325
rect 106337 73269 106393 73325
rect 106479 73269 106535 73325
rect 106621 73269 106677 73325
rect 106763 73269 106819 73325
rect 106905 73269 106961 73325
rect 107047 73269 107103 73325
rect 105343 73127 105399 73183
rect 105485 73127 105541 73183
rect 105627 73127 105683 73183
rect 105769 73127 105825 73183
rect 105911 73127 105967 73183
rect 106053 73127 106109 73183
rect 106195 73127 106251 73183
rect 106337 73127 106393 73183
rect 106479 73127 106535 73183
rect 106621 73127 106677 73183
rect 106763 73127 106819 73183
rect 106905 73127 106961 73183
rect 107047 73127 107103 73183
rect 105343 72985 105399 73041
rect 105485 72985 105541 73041
rect 105627 72985 105683 73041
rect 105769 72985 105825 73041
rect 105911 72985 105967 73041
rect 106053 72985 106109 73041
rect 106195 72985 106251 73041
rect 106337 72985 106393 73041
rect 106479 72985 106535 73041
rect 106621 72985 106677 73041
rect 106763 72985 106819 73041
rect 106905 72985 106961 73041
rect 107047 72985 107103 73041
rect 105343 72843 105399 72899
rect 105485 72843 105541 72899
rect 105627 72843 105683 72899
rect 105769 72843 105825 72899
rect 105911 72843 105967 72899
rect 106053 72843 106109 72899
rect 106195 72843 106251 72899
rect 106337 72843 106393 72899
rect 106479 72843 106535 72899
rect 106621 72843 106677 72899
rect 106763 72843 106819 72899
rect 106905 72843 106961 72899
rect 107047 72843 107103 72899
rect 105343 72701 105399 72757
rect 105485 72701 105541 72757
rect 105627 72701 105683 72757
rect 105769 72701 105825 72757
rect 105911 72701 105967 72757
rect 106053 72701 106109 72757
rect 106195 72701 106251 72757
rect 106337 72701 106393 72757
rect 106479 72701 106535 72757
rect 106621 72701 106677 72757
rect 106763 72701 106819 72757
rect 106905 72701 106961 72757
rect 107047 72701 107103 72757
rect 105343 72559 105399 72615
rect 105485 72559 105541 72615
rect 105627 72559 105683 72615
rect 105769 72559 105825 72615
rect 105911 72559 105967 72615
rect 106053 72559 106109 72615
rect 106195 72559 106251 72615
rect 106337 72559 106393 72615
rect 106479 72559 106535 72615
rect 106621 72559 106677 72615
rect 106763 72559 106819 72615
rect 106905 72559 106961 72615
rect 107047 72559 107103 72615
rect 105343 72417 105399 72473
rect 105485 72417 105541 72473
rect 105627 72417 105683 72473
rect 105769 72417 105825 72473
rect 105911 72417 105967 72473
rect 106053 72417 106109 72473
rect 106195 72417 106251 72473
rect 106337 72417 106393 72473
rect 106479 72417 106535 72473
rect 106621 72417 106677 72473
rect 106763 72417 106819 72473
rect 106905 72417 106961 72473
rect 107047 72417 107103 72473
rect 105343 72275 105399 72331
rect 105485 72275 105541 72331
rect 105627 72275 105683 72331
rect 105769 72275 105825 72331
rect 105911 72275 105967 72331
rect 106053 72275 106109 72331
rect 106195 72275 106251 72331
rect 106337 72275 106393 72331
rect 106479 72275 106535 72331
rect 106621 72275 106677 72331
rect 106763 72275 106819 72331
rect 106905 72275 106961 72331
rect 107047 72275 107103 72331
rect 105343 72133 105399 72189
rect 105485 72133 105541 72189
rect 105627 72133 105683 72189
rect 105769 72133 105825 72189
rect 105911 72133 105967 72189
rect 106053 72133 106109 72189
rect 106195 72133 106251 72189
rect 106337 72133 106393 72189
rect 106479 72133 106535 72189
rect 106621 72133 106677 72189
rect 106763 72133 106819 72189
rect 106905 72133 106961 72189
rect 107047 72133 107103 72189
rect 108995 73979 109051 74035
rect 109137 73979 109193 74035
rect 109279 73979 109335 74035
rect 109421 73979 109477 74035
rect 109563 73979 109619 74035
rect 109705 73979 109761 74035
rect 108995 73837 109051 73893
rect 109137 73837 109193 73893
rect 109279 73837 109335 73893
rect 109421 73837 109477 73893
rect 109563 73837 109619 73893
rect 109705 73837 109761 73893
rect 108995 73695 109051 73751
rect 109137 73695 109193 73751
rect 109279 73695 109335 73751
rect 109421 73695 109477 73751
rect 109563 73695 109619 73751
rect 109705 73695 109761 73751
rect 108995 73553 109051 73609
rect 109137 73553 109193 73609
rect 109279 73553 109335 73609
rect 109421 73553 109477 73609
rect 109563 73553 109619 73609
rect 109705 73553 109761 73609
rect 108995 73411 109051 73467
rect 109137 73411 109193 73467
rect 109279 73411 109335 73467
rect 109421 73411 109477 73467
rect 109563 73411 109619 73467
rect 109705 73411 109761 73467
rect 108995 73269 109051 73325
rect 109137 73269 109193 73325
rect 109279 73269 109335 73325
rect 109421 73269 109477 73325
rect 109563 73269 109619 73325
rect 109705 73269 109761 73325
rect 108995 73127 109051 73183
rect 109137 73127 109193 73183
rect 109279 73127 109335 73183
rect 109421 73127 109477 73183
rect 109563 73127 109619 73183
rect 109705 73127 109761 73183
rect 108995 72985 109051 73041
rect 109137 72985 109193 73041
rect 109279 72985 109335 73041
rect 109421 72985 109477 73041
rect 109563 72985 109619 73041
rect 109705 72985 109761 73041
rect 108995 72843 109051 72899
rect 109137 72843 109193 72899
rect 109279 72843 109335 72899
rect 109421 72843 109477 72899
rect 109563 72843 109619 72899
rect 109705 72843 109761 72899
rect 108995 72701 109051 72757
rect 109137 72701 109193 72757
rect 109279 72701 109335 72757
rect 109421 72701 109477 72757
rect 109563 72701 109619 72757
rect 109705 72701 109761 72757
rect 108995 72559 109051 72615
rect 109137 72559 109193 72615
rect 109279 72559 109335 72615
rect 109421 72559 109477 72615
rect 109563 72559 109619 72615
rect 109705 72559 109761 72615
rect 108995 72417 109051 72473
rect 109137 72417 109193 72473
rect 109279 72417 109335 72473
rect 109421 72417 109477 72473
rect 109563 72417 109619 72473
rect 109705 72417 109761 72473
rect 108995 72275 109051 72331
rect 109137 72275 109193 72331
rect 109279 72275 109335 72331
rect 109421 72275 109477 72331
rect 109563 72275 109619 72331
rect 109705 72275 109761 72331
rect 108995 72133 109051 72189
rect 109137 72133 109193 72189
rect 109279 72133 109335 72189
rect 109421 72133 109477 72189
rect 109563 72133 109619 72189
rect 109705 72133 109761 72189
rect 110193 73979 110249 74035
rect 110335 73979 110391 74035
rect 110477 73979 110533 74035
rect 110619 73979 110675 74035
rect 110761 73979 110817 74035
rect 110903 73979 110959 74035
rect 111045 73979 111101 74035
rect 111187 73979 111243 74035
rect 111329 73979 111385 74035
rect 111471 73979 111527 74035
rect 111613 73979 111669 74035
rect 111755 73979 111811 74035
rect 111897 73979 111953 74035
rect 112039 73979 112095 74035
rect 110193 73837 110249 73893
rect 110335 73837 110391 73893
rect 110477 73837 110533 73893
rect 110619 73837 110675 73893
rect 110761 73837 110817 73893
rect 110903 73837 110959 73893
rect 111045 73837 111101 73893
rect 111187 73837 111243 73893
rect 111329 73837 111385 73893
rect 111471 73837 111527 73893
rect 111613 73837 111669 73893
rect 111755 73837 111811 73893
rect 111897 73837 111953 73893
rect 112039 73837 112095 73893
rect 110193 73695 110249 73751
rect 110335 73695 110391 73751
rect 110477 73695 110533 73751
rect 110619 73695 110675 73751
rect 110761 73695 110817 73751
rect 110903 73695 110959 73751
rect 111045 73695 111101 73751
rect 111187 73695 111243 73751
rect 111329 73695 111385 73751
rect 111471 73695 111527 73751
rect 111613 73695 111669 73751
rect 111755 73695 111811 73751
rect 111897 73695 111953 73751
rect 112039 73695 112095 73751
rect 110193 73553 110249 73609
rect 110335 73553 110391 73609
rect 110477 73553 110533 73609
rect 110619 73553 110675 73609
rect 110761 73553 110817 73609
rect 110903 73553 110959 73609
rect 111045 73553 111101 73609
rect 111187 73553 111243 73609
rect 111329 73553 111385 73609
rect 111471 73553 111527 73609
rect 111613 73553 111669 73609
rect 111755 73553 111811 73609
rect 111897 73553 111953 73609
rect 112039 73553 112095 73609
rect 110193 73411 110249 73467
rect 110335 73411 110391 73467
rect 110477 73411 110533 73467
rect 110619 73411 110675 73467
rect 110761 73411 110817 73467
rect 110903 73411 110959 73467
rect 111045 73411 111101 73467
rect 111187 73411 111243 73467
rect 111329 73411 111385 73467
rect 111471 73411 111527 73467
rect 111613 73411 111669 73467
rect 111755 73411 111811 73467
rect 111897 73411 111953 73467
rect 112039 73411 112095 73467
rect 110193 73269 110249 73325
rect 110335 73269 110391 73325
rect 110477 73269 110533 73325
rect 110619 73269 110675 73325
rect 110761 73269 110817 73325
rect 110903 73269 110959 73325
rect 111045 73269 111101 73325
rect 111187 73269 111243 73325
rect 111329 73269 111385 73325
rect 111471 73269 111527 73325
rect 111613 73269 111669 73325
rect 111755 73269 111811 73325
rect 111897 73269 111953 73325
rect 112039 73269 112095 73325
rect 110193 73127 110249 73183
rect 110335 73127 110391 73183
rect 110477 73127 110533 73183
rect 110619 73127 110675 73183
rect 110761 73127 110817 73183
rect 110903 73127 110959 73183
rect 111045 73127 111101 73183
rect 111187 73127 111243 73183
rect 111329 73127 111385 73183
rect 111471 73127 111527 73183
rect 111613 73127 111669 73183
rect 111755 73127 111811 73183
rect 111897 73127 111953 73183
rect 112039 73127 112095 73183
rect 110193 72985 110249 73041
rect 110335 72985 110391 73041
rect 110477 72985 110533 73041
rect 110619 72985 110675 73041
rect 110761 72985 110817 73041
rect 110903 72985 110959 73041
rect 111045 72985 111101 73041
rect 111187 72985 111243 73041
rect 111329 72985 111385 73041
rect 111471 72985 111527 73041
rect 111613 72985 111669 73041
rect 111755 72985 111811 73041
rect 111897 72985 111953 73041
rect 112039 72985 112095 73041
rect 110193 72843 110249 72899
rect 110335 72843 110391 72899
rect 110477 72843 110533 72899
rect 110619 72843 110675 72899
rect 110761 72843 110817 72899
rect 110903 72843 110959 72899
rect 111045 72843 111101 72899
rect 111187 72843 111243 72899
rect 111329 72843 111385 72899
rect 111471 72843 111527 72899
rect 111613 72843 111669 72899
rect 111755 72843 111811 72899
rect 111897 72843 111953 72899
rect 112039 72843 112095 72899
rect 110193 72701 110249 72757
rect 110335 72701 110391 72757
rect 110477 72701 110533 72757
rect 110619 72701 110675 72757
rect 110761 72701 110817 72757
rect 110903 72701 110959 72757
rect 111045 72701 111101 72757
rect 111187 72701 111243 72757
rect 111329 72701 111385 72757
rect 111471 72701 111527 72757
rect 111613 72701 111669 72757
rect 111755 72701 111811 72757
rect 111897 72701 111953 72757
rect 112039 72701 112095 72757
rect 110193 72559 110249 72615
rect 110335 72559 110391 72615
rect 110477 72559 110533 72615
rect 110619 72559 110675 72615
rect 110761 72559 110817 72615
rect 110903 72559 110959 72615
rect 111045 72559 111101 72615
rect 111187 72559 111243 72615
rect 111329 72559 111385 72615
rect 111471 72559 111527 72615
rect 111613 72559 111669 72615
rect 111755 72559 111811 72615
rect 111897 72559 111953 72615
rect 112039 72559 112095 72615
rect 110193 72417 110249 72473
rect 110335 72417 110391 72473
rect 110477 72417 110533 72473
rect 110619 72417 110675 72473
rect 110761 72417 110817 72473
rect 110903 72417 110959 72473
rect 111045 72417 111101 72473
rect 111187 72417 111243 72473
rect 111329 72417 111385 72473
rect 111471 72417 111527 72473
rect 111613 72417 111669 72473
rect 111755 72417 111811 72473
rect 111897 72417 111953 72473
rect 112039 72417 112095 72473
rect 110193 72275 110249 72331
rect 110335 72275 110391 72331
rect 110477 72275 110533 72331
rect 110619 72275 110675 72331
rect 110761 72275 110817 72331
rect 110903 72275 110959 72331
rect 111045 72275 111101 72331
rect 111187 72275 111243 72331
rect 111329 72275 111385 72331
rect 111471 72275 111527 72331
rect 111613 72275 111669 72331
rect 111755 72275 111811 72331
rect 111897 72275 111953 72331
rect 112039 72275 112095 72331
rect 110193 72133 110249 72189
rect 110335 72133 110391 72189
rect 110477 72133 110533 72189
rect 110619 72133 110675 72189
rect 110761 72133 110817 72189
rect 110903 72133 110959 72189
rect 111045 72133 111101 72189
rect 111187 72133 111243 72189
rect 111329 72133 111385 72189
rect 111471 72133 111527 72189
rect 111613 72133 111669 72189
rect 111755 72133 111811 72189
rect 111897 72133 111953 72189
rect 112039 72133 112095 72189
rect 113325 73979 113381 74035
rect 113467 73979 113523 74035
rect 113609 73979 113665 74035
rect 113751 73979 113807 74035
rect 113893 73979 113949 74035
rect 114035 73979 114091 74035
rect 114177 73979 114233 74035
rect 114319 73979 114375 74035
rect 114461 73979 114517 74035
rect 114603 73979 114659 74035
rect 114745 73979 114801 74035
rect 113325 73837 113381 73893
rect 113467 73837 113523 73893
rect 113609 73837 113665 73893
rect 113751 73837 113807 73893
rect 113893 73837 113949 73893
rect 114035 73837 114091 73893
rect 114177 73837 114233 73893
rect 114319 73837 114375 73893
rect 114461 73837 114517 73893
rect 114603 73837 114659 73893
rect 114745 73837 114801 73893
rect 113325 73695 113381 73751
rect 113467 73695 113523 73751
rect 113609 73695 113665 73751
rect 113751 73695 113807 73751
rect 113893 73695 113949 73751
rect 114035 73695 114091 73751
rect 114177 73695 114233 73751
rect 114319 73695 114375 73751
rect 114461 73695 114517 73751
rect 114603 73695 114659 73751
rect 114745 73695 114801 73751
rect 113325 73553 113381 73609
rect 113467 73553 113523 73609
rect 113609 73553 113665 73609
rect 113751 73553 113807 73609
rect 113893 73553 113949 73609
rect 114035 73553 114091 73609
rect 114177 73553 114233 73609
rect 114319 73553 114375 73609
rect 114461 73553 114517 73609
rect 114603 73553 114659 73609
rect 114745 73553 114801 73609
rect 113325 73411 113381 73467
rect 113467 73411 113523 73467
rect 113609 73411 113665 73467
rect 113751 73411 113807 73467
rect 113893 73411 113949 73467
rect 114035 73411 114091 73467
rect 114177 73411 114233 73467
rect 114319 73411 114375 73467
rect 114461 73411 114517 73467
rect 114603 73411 114659 73467
rect 114745 73411 114801 73467
rect 113325 73269 113381 73325
rect 113467 73269 113523 73325
rect 113609 73269 113665 73325
rect 113751 73269 113807 73325
rect 113893 73269 113949 73325
rect 114035 73269 114091 73325
rect 114177 73269 114233 73325
rect 114319 73269 114375 73325
rect 114461 73269 114517 73325
rect 114603 73269 114659 73325
rect 114745 73269 114801 73325
rect 113325 73127 113381 73183
rect 113467 73127 113523 73183
rect 113609 73127 113665 73183
rect 113751 73127 113807 73183
rect 113893 73127 113949 73183
rect 114035 73127 114091 73183
rect 114177 73127 114233 73183
rect 114319 73127 114375 73183
rect 114461 73127 114517 73183
rect 114603 73127 114659 73183
rect 114745 73127 114801 73183
rect 113325 72985 113381 73041
rect 113467 72985 113523 73041
rect 113609 72985 113665 73041
rect 113751 72985 113807 73041
rect 113893 72985 113949 73041
rect 114035 72985 114091 73041
rect 114177 72985 114233 73041
rect 114319 72985 114375 73041
rect 114461 72985 114517 73041
rect 114603 72985 114659 73041
rect 114745 72985 114801 73041
rect 113325 72843 113381 72899
rect 113467 72843 113523 72899
rect 113609 72843 113665 72899
rect 113751 72843 113807 72899
rect 113893 72843 113949 72899
rect 114035 72843 114091 72899
rect 114177 72843 114233 72899
rect 114319 72843 114375 72899
rect 114461 72843 114517 72899
rect 114603 72843 114659 72899
rect 114745 72843 114801 72899
rect 113325 72701 113381 72757
rect 113467 72701 113523 72757
rect 113609 72701 113665 72757
rect 113751 72701 113807 72757
rect 113893 72701 113949 72757
rect 114035 72701 114091 72757
rect 114177 72701 114233 72757
rect 114319 72701 114375 72757
rect 114461 72701 114517 72757
rect 114603 72701 114659 72757
rect 114745 72701 114801 72757
rect 113325 72559 113381 72615
rect 113467 72559 113523 72615
rect 113609 72559 113665 72615
rect 113751 72559 113807 72615
rect 113893 72559 113949 72615
rect 114035 72559 114091 72615
rect 114177 72559 114233 72615
rect 114319 72559 114375 72615
rect 114461 72559 114517 72615
rect 114603 72559 114659 72615
rect 114745 72559 114801 72615
rect 113325 72417 113381 72473
rect 113467 72417 113523 72473
rect 113609 72417 113665 72473
rect 113751 72417 113807 72473
rect 113893 72417 113949 72473
rect 114035 72417 114091 72473
rect 114177 72417 114233 72473
rect 114319 72417 114375 72473
rect 114461 72417 114517 72473
rect 114603 72417 114659 72473
rect 114745 72417 114801 72473
rect 113325 72275 113381 72331
rect 113467 72275 113523 72331
rect 113609 72275 113665 72331
rect 113751 72275 113807 72331
rect 113893 72275 113949 72331
rect 114035 72275 114091 72331
rect 114177 72275 114233 72331
rect 114319 72275 114375 72331
rect 114461 72275 114517 72331
rect 114603 72275 114659 72331
rect 114745 72275 114801 72331
rect 113325 72133 113381 72189
rect 113467 72133 113523 72189
rect 113609 72133 113665 72189
rect 113751 72133 113807 72189
rect 113893 72133 113949 72189
rect 114035 72133 114091 72189
rect 114177 72133 114233 72189
rect 114319 72133 114375 72189
rect 114461 72133 114517 72189
rect 114603 72133 114659 72189
rect 114745 72133 114801 72189
rect 115269 73979 115325 74035
rect 115411 73979 115467 74035
rect 115553 73979 115609 74035
rect 115695 73979 115751 74035
rect 115837 73979 115893 74035
rect 115979 73979 116035 74035
rect 116121 73979 116177 74035
rect 116263 73979 116319 74035
rect 116405 73979 116461 74035
rect 116547 73979 116603 74035
rect 116689 73979 116745 74035
rect 116831 73979 116887 74035
rect 116973 73979 117029 74035
rect 117115 73979 117171 74035
rect 115269 73837 115325 73893
rect 115411 73837 115467 73893
rect 115553 73837 115609 73893
rect 115695 73837 115751 73893
rect 115837 73837 115893 73893
rect 115979 73837 116035 73893
rect 116121 73837 116177 73893
rect 116263 73837 116319 73893
rect 116405 73837 116461 73893
rect 116547 73837 116603 73893
rect 116689 73837 116745 73893
rect 116831 73837 116887 73893
rect 116973 73837 117029 73893
rect 117115 73837 117171 73893
rect 115269 73695 115325 73751
rect 115411 73695 115467 73751
rect 115553 73695 115609 73751
rect 115695 73695 115751 73751
rect 115837 73695 115893 73751
rect 115979 73695 116035 73751
rect 116121 73695 116177 73751
rect 116263 73695 116319 73751
rect 116405 73695 116461 73751
rect 116547 73695 116603 73751
rect 116689 73695 116745 73751
rect 116831 73695 116887 73751
rect 116973 73695 117029 73751
rect 117115 73695 117171 73751
rect 115269 73553 115325 73609
rect 115411 73553 115467 73609
rect 115553 73553 115609 73609
rect 115695 73553 115751 73609
rect 115837 73553 115893 73609
rect 115979 73553 116035 73609
rect 116121 73553 116177 73609
rect 116263 73553 116319 73609
rect 116405 73553 116461 73609
rect 116547 73553 116603 73609
rect 116689 73553 116745 73609
rect 116831 73553 116887 73609
rect 116973 73553 117029 73609
rect 117115 73553 117171 73609
rect 115269 73411 115325 73467
rect 115411 73411 115467 73467
rect 115553 73411 115609 73467
rect 115695 73411 115751 73467
rect 115837 73411 115893 73467
rect 115979 73411 116035 73467
rect 116121 73411 116177 73467
rect 116263 73411 116319 73467
rect 116405 73411 116461 73467
rect 116547 73411 116603 73467
rect 116689 73411 116745 73467
rect 116831 73411 116887 73467
rect 116973 73411 117029 73467
rect 117115 73411 117171 73467
rect 115269 73269 115325 73325
rect 115411 73269 115467 73325
rect 115553 73269 115609 73325
rect 115695 73269 115751 73325
rect 115837 73269 115893 73325
rect 115979 73269 116035 73325
rect 116121 73269 116177 73325
rect 116263 73269 116319 73325
rect 116405 73269 116461 73325
rect 116547 73269 116603 73325
rect 116689 73269 116745 73325
rect 116831 73269 116887 73325
rect 116973 73269 117029 73325
rect 117115 73269 117171 73325
rect 115269 73127 115325 73183
rect 115411 73127 115467 73183
rect 115553 73127 115609 73183
rect 115695 73127 115751 73183
rect 115837 73127 115893 73183
rect 115979 73127 116035 73183
rect 116121 73127 116177 73183
rect 116263 73127 116319 73183
rect 116405 73127 116461 73183
rect 116547 73127 116603 73183
rect 116689 73127 116745 73183
rect 116831 73127 116887 73183
rect 116973 73127 117029 73183
rect 117115 73127 117171 73183
rect 115269 72985 115325 73041
rect 115411 72985 115467 73041
rect 115553 72985 115609 73041
rect 115695 72985 115751 73041
rect 115837 72985 115893 73041
rect 115979 72985 116035 73041
rect 116121 72985 116177 73041
rect 116263 72985 116319 73041
rect 116405 72985 116461 73041
rect 116547 72985 116603 73041
rect 116689 72985 116745 73041
rect 116831 72985 116887 73041
rect 116973 72985 117029 73041
rect 117115 72985 117171 73041
rect 115269 72843 115325 72899
rect 115411 72843 115467 72899
rect 115553 72843 115609 72899
rect 115695 72843 115751 72899
rect 115837 72843 115893 72899
rect 115979 72843 116035 72899
rect 116121 72843 116177 72899
rect 116263 72843 116319 72899
rect 116405 72843 116461 72899
rect 116547 72843 116603 72899
rect 116689 72843 116745 72899
rect 116831 72843 116887 72899
rect 116973 72843 117029 72899
rect 117115 72843 117171 72899
rect 115269 72701 115325 72757
rect 115411 72701 115467 72757
rect 115553 72701 115609 72757
rect 115695 72701 115751 72757
rect 115837 72701 115893 72757
rect 115979 72701 116035 72757
rect 116121 72701 116177 72757
rect 116263 72701 116319 72757
rect 116405 72701 116461 72757
rect 116547 72701 116603 72757
rect 116689 72701 116745 72757
rect 116831 72701 116887 72757
rect 116973 72701 117029 72757
rect 117115 72701 117171 72757
rect 115269 72559 115325 72615
rect 115411 72559 115467 72615
rect 115553 72559 115609 72615
rect 115695 72559 115751 72615
rect 115837 72559 115893 72615
rect 115979 72559 116035 72615
rect 116121 72559 116177 72615
rect 116263 72559 116319 72615
rect 116405 72559 116461 72615
rect 116547 72559 116603 72615
rect 116689 72559 116745 72615
rect 116831 72559 116887 72615
rect 116973 72559 117029 72615
rect 117115 72559 117171 72615
rect 115269 72417 115325 72473
rect 115411 72417 115467 72473
rect 115553 72417 115609 72473
rect 115695 72417 115751 72473
rect 115837 72417 115893 72473
rect 115979 72417 116035 72473
rect 116121 72417 116177 72473
rect 116263 72417 116319 72473
rect 116405 72417 116461 72473
rect 116547 72417 116603 72473
rect 116689 72417 116745 72473
rect 116831 72417 116887 72473
rect 116973 72417 117029 72473
rect 117115 72417 117171 72473
rect 115269 72275 115325 72331
rect 115411 72275 115467 72331
rect 115553 72275 115609 72331
rect 115695 72275 115751 72331
rect 115837 72275 115893 72331
rect 115979 72275 116035 72331
rect 116121 72275 116177 72331
rect 116263 72275 116319 72331
rect 116405 72275 116461 72331
rect 116547 72275 116603 72331
rect 116689 72275 116745 72331
rect 116831 72275 116887 72331
rect 116973 72275 117029 72331
rect 117115 72275 117171 72331
rect 115269 72133 115325 72189
rect 115411 72133 115467 72189
rect 115553 72133 115609 72189
rect 115695 72133 115751 72189
rect 115837 72133 115893 72189
rect 115979 72133 116035 72189
rect 116121 72133 116177 72189
rect 116263 72133 116319 72189
rect 116405 72133 116461 72189
rect 116547 72133 116603 72189
rect 116689 72133 116745 72189
rect 116831 72133 116887 72189
rect 116973 72133 117029 72189
rect 117115 72133 117171 72189
rect 117899 73979 117955 74035
rect 118041 73979 118097 74035
rect 118183 73979 118239 74035
rect 118325 73979 118381 74035
rect 118467 73979 118523 74035
rect 118609 73979 118665 74035
rect 118751 73979 118807 74035
rect 118893 73979 118949 74035
rect 119035 73979 119091 74035
rect 119177 73979 119233 74035
rect 119319 73979 119375 74035
rect 119461 73979 119517 74035
rect 119603 73979 119659 74035
rect 117899 73837 117955 73893
rect 118041 73837 118097 73893
rect 118183 73837 118239 73893
rect 118325 73837 118381 73893
rect 118467 73837 118523 73893
rect 118609 73837 118665 73893
rect 118751 73837 118807 73893
rect 118893 73837 118949 73893
rect 119035 73837 119091 73893
rect 119177 73837 119233 73893
rect 119319 73837 119375 73893
rect 119461 73837 119517 73893
rect 119603 73837 119659 73893
rect 117899 73695 117955 73751
rect 118041 73695 118097 73751
rect 118183 73695 118239 73751
rect 118325 73695 118381 73751
rect 118467 73695 118523 73751
rect 118609 73695 118665 73751
rect 118751 73695 118807 73751
rect 118893 73695 118949 73751
rect 119035 73695 119091 73751
rect 119177 73695 119233 73751
rect 119319 73695 119375 73751
rect 119461 73695 119517 73751
rect 119603 73695 119659 73751
rect 117899 73553 117955 73609
rect 118041 73553 118097 73609
rect 118183 73553 118239 73609
rect 118325 73553 118381 73609
rect 118467 73553 118523 73609
rect 118609 73553 118665 73609
rect 118751 73553 118807 73609
rect 118893 73553 118949 73609
rect 119035 73553 119091 73609
rect 119177 73553 119233 73609
rect 119319 73553 119375 73609
rect 119461 73553 119517 73609
rect 119603 73553 119659 73609
rect 117899 73411 117955 73467
rect 118041 73411 118097 73467
rect 118183 73411 118239 73467
rect 118325 73411 118381 73467
rect 118467 73411 118523 73467
rect 118609 73411 118665 73467
rect 118751 73411 118807 73467
rect 118893 73411 118949 73467
rect 119035 73411 119091 73467
rect 119177 73411 119233 73467
rect 119319 73411 119375 73467
rect 119461 73411 119517 73467
rect 119603 73411 119659 73467
rect 117899 73269 117955 73325
rect 118041 73269 118097 73325
rect 118183 73269 118239 73325
rect 118325 73269 118381 73325
rect 118467 73269 118523 73325
rect 118609 73269 118665 73325
rect 118751 73269 118807 73325
rect 118893 73269 118949 73325
rect 119035 73269 119091 73325
rect 119177 73269 119233 73325
rect 119319 73269 119375 73325
rect 119461 73269 119517 73325
rect 119603 73269 119659 73325
rect 117899 73127 117955 73183
rect 118041 73127 118097 73183
rect 118183 73127 118239 73183
rect 118325 73127 118381 73183
rect 118467 73127 118523 73183
rect 118609 73127 118665 73183
rect 118751 73127 118807 73183
rect 118893 73127 118949 73183
rect 119035 73127 119091 73183
rect 119177 73127 119233 73183
rect 119319 73127 119375 73183
rect 119461 73127 119517 73183
rect 119603 73127 119659 73183
rect 117899 72985 117955 73041
rect 118041 72985 118097 73041
rect 118183 72985 118239 73041
rect 118325 72985 118381 73041
rect 118467 72985 118523 73041
rect 118609 72985 118665 73041
rect 118751 72985 118807 73041
rect 118893 72985 118949 73041
rect 119035 72985 119091 73041
rect 119177 72985 119233 73041
rect 119319 72985 119375 73041
rect 119461 72985 119517 73041
rect 119603 72985 119659 73041
rect 117899 72843 117955 72899
rect 118041 72843 118097 72899
rect 118183 72843 118239 72899
rect 118325 72843 118381 72899
rect 118467 72843 118523 72899
rect 118609 72843 118665 72899
rect 118751 72843 118807 72899
rect 118893 72843 118949 72899
rect 119035 72843 119091 72899
rect 119177 72843 119233 72899
rect 119319 72843 119375 72899
rect 119461 72843 119517 72899
rect 119603 72843 119659 72899
rect 117899 72701 117955 72757
rect 118041 72701 118097 72757
rect 118183 72701 118239 72757
rect 118325 72701 118381 72757
rect 118467 72701 118523 72757
rect 118609 72701 118665 72757
rect 118751 72701 118807 72757
rect 118893 72701 118949 72757
rect 119035 72701 119091 72757
rect 119177 72701 119233 72757
rect 119319 72701 119375 72757
rect 119461 72701 119517 72757
rect 119603 72701 119659 72757
rect 117899 72559 117955 72615
rect 118041 72559 118097 72615
rect 118183 72559 118239 72615
rect 118325 72559 118381 72615
rect 118467 72559 118523 72615
rect 118609 72559 118665 72615
rect 118751 72559 118807 72615
rect 118893 72559 118949 72615
rect 119035 72559 119091 72615
rect 119177 72559 119233 72615
rect 119319 72559 119375 72615
rect 119461 72559 119517 72615
rect 119603 72559 119659 72615
rect 117899 72417 117955 72473
rect 118041 72417 118097 72473
rect 118183 72417 118239 72473
rect 118325 72417 118381 72473
rect 118467 72417 118523 72473
rect 118609 72417 118665 72473
rect 118751 72417 118807 72473
rect 118893 72417 118949 72473
rect 119035 72417 119091 72473
rect 119177 72417 119233 72473
rect 119319 72417 119375 72473
rect 119461 72417 119517 72473
rect 119603 72417 119659 72473
rect 117899 72275 117955 72331
rect 118041 72275 118097 72331
rect 118183 72275 118239 72331
rect 118325 72275 118381 72331
rect 118467 72275 118523 72331
rect 118609 72275 118665 72331
rect 118751 72275 118807 72331
rect 118893 72275 118949 72331
rect 119035 72275 119091 72331
rect 119177 72275 119233 72331
rect 119319 72275 119375 72331
rect 119461 72275 119517 72331
rect 119603 72275 119659 72331
rect 117899 72133 117955 72189
rect 118041 72133 118097 72189
rect 118183 72133 118239 72189
rect 118325 72133 118381 72189
rect 118467 72133 118523 72189
rect 118609 72133 118665 72189
rect 118751 72133 118807 72189
rect 118893 72133 118949 72189
rect 119035 72133 119091 72189
rect 119177 72133 119233 72189
rect 119319 72133 119375 72189
rect 119461 72133 119517 72189
rect 119603 72133 119659 72189
rect 270343 73979 270399 74035
rect 270485 73979 270541 74035
rect 270627 73979 270683 74035
rect 270769 73979 270825 74035
rect 270911 73979 270967 74035
rect 271053 73979 271109 74035
rect 271195 73979 271251 74035
rect 271337 73979 271393 74035
rect 271479 73979 271535 74035
rect 271621 73979 271677 74035
rect 271763 73979 271819 74035
rect 271905 73979 271961 74035
rect 272047 73979 272103 74035
rect 270343 73837 270399 73893
rect 270485 73837 270541 73893
rect 270627 73837 270683 73893
rect 270769 73837 270825 73893
rect 270911 73837 270967 73893
rect 271053 73837 271109 73893
rect 271195 73837 271251 73893
rect 271337 73837 271393 73893
rect 271479 73837 271535 73893
rect 271621 73837 271677 73893
rect 271763 73837 271819 73893
rect 271905 73837 271961 73893
rect 272047 73837 272103 73893
rect 270343 73695 270399 73751
rect 270485 73695 270541 73751
rect 270627 73695 270683 73751
rect 270769 73695 270825 73751
rect 270911 73695 270967 73751
rect 271053 73695 271109 73751
rect 271195 73695 271251 73751
rect 271337 73695 271393 73751
rect 271479 73695 271535 73751
rect 271621 73695 271677 73751
rect 271763 73695 271819 73751
rect 271905 73695 271961 73751
rect 272047 73695 272103 73751
rect 270343 73553 270399 73609
rect 270485 73553 270541 73609
rect 270627 73553 270683 73609
rect 270769 73553 270825 73609
rect 270911 73553 270967 73609
rect 271053 73553 271109 73609
rect 271195 73553 271251 73609
rect 271337 73553 271393 73609
rect 271479 73553 271535 73609
rect 271621 73553 271677 73609
rect 271763 73553 271819 73609
rect 271905 73553 271961 73609
rect 272047 73553 272103 73609
rect 270343 73411 270399 73467
rect 270485 73411 270541 73467
rect 270627 73411 270683 73467
rect 270769 73411 270825 73467
rect 270911 73411 270967 73467
rect 271053 73411 271109 73467
rect 271195 73411 271251 73467
rect 271337 73411 271393 73467
rect 271479 73411 271535 73467
rect 271621 73411 271677 73467
rect 271763 73411 271819 73467
rect 271905 73411 271961 73467
rect 272047 73411 272103 73467
rect 270343 73269 270399 73325
rect 270485 73269 270541 73325
rect 270627 73269 270683 73325
rect 270769 73269 270825 73325
rect 270911 73269 270967 73325
rect 271053 73269 271109 73325
rect 271195 73269 271251 73325
rect 271337 73269 271393 73325
rect 271479 73269 271535 73325
rect 271621 73269 271677 73325
rect 271763 73269 271819 73325
rect 271905 73269 271961 73325
rect 272047 73269 272103 73325
rect 270343 73127 270399 73183
rect 270485 73127 270541 73183
rect 270627 73127 270683 73183
rect 270769 73127 270825 73183
rect 270911 73127 270967 73183
rect 271053 73127 271109 73183
rect 271195 73127 271251 73183
rect 271337 73127 271393 73183
rect 271479 73127 271535 73183
rect 271621 73127 271677 73183
rect 271763 73127 271819 73183
rect 271905 73127 271961 73183
rect 272047 73127 272103 73183
rect 270343 72985 270399 73041
rect 270485 72985 270541 73041
rect 270627 72985 270683 73041
rect 270769 72985 270825 73041
rect 270911 72985 270967 73041
rect 271053 72985 271109 73041
rect 271195 72985 271251 73041
rect 271337 72985 271393 73041
rect 271479 72985 271535 73041
rect 271621 72985 271677 73041
rect 271763 72985 271819 73041
rect 271905 72985 271961 73041
rect 272047 72985 272103 73041
rect 270343 72843 270399 72899
rect 270485 72843 270541 72899
rect 270627 72843 270683 72899
rect 270769 72843 270825 72899
rect 270911 72843 270967 72899
rect 271053 72843 271109 72899
rect 271195 72843 271251 72899
rect 271337 72843 271393 72899
rect 271479 72843 271535 72899
rect 271621 72843 271677 72899
rect 271763 72843 271819 72899
rect 271905 72843 271961 72899
rect 272047 72843 272103 72899
rect 270343 72701 270399 72757
rect 270485 72701 270541 72757
rect 270627 72701 270683 72757
rect 270769 72701 270825 72757
rect 270911 72701 270967 72757
rect 271053 72701 271109 72757
rect 271195 72701 271251 72757
rect 271337 72701 271393 72757
rect 271479 72701 271535 72757
rect 271621 72701 271677 72757
rect 271763 72701 271819 72757
rect 271905 72701 271961 72757
rect 272047 72701 272103 72757
rect 270343 72559 270399 72615
rect 270485 72559 270541 72615
rect 270627 72559 270683 72615
rect 270769 72559 270825 72615
rect 270911 72559 270967 72615
rect 271053 72559 271109 72615
rect 271195 72559 271251 72615
rect 271337 72559 271393 72615
rect 271479 72559 271535 72615
rect 271621 72559 271677 72615
rect 271763 72559 271819 72615
rect 271905 72559 271961 72615
rect 272047 72559 272103 72615
rect 270343 72417 270399 72473
rect 270485 72417 270541 72473
rect 270627 72417 270683 72473
rect 270769 72417 270825 72473
rect 270911 72417 270967 72473
rect 271053 72417 271109 72473
rect 271195 72417 271251 72473
rect 271337 72417 271393 72473
rect 271479 72417 271535 72473
rect 271621 72417 271677 72473
rect 271763 72417 271819 72473
rect 271905 72417 271961 72473
rect 272047 72417 272103 72473
rect 270343 72275 270399 72331
rect 270485 72275 270541 72331
rect 270627 72275 270683 72331
rect 270769 72275 270825 72331
rect 270911 72275 270967 72331
rect 271053 72275 271109 72331
rect 271195 72275 271251 72331
rect 271337 72275 271393 72331
rect 271479 72275 271535 72331
rect 271621 72275 271677 72331
rect 271763 72275 271819 72331
rect 271905 72275 271961 72331
rect 272047 72275 272103 72331
rect 270343 72133 270399 72189
rect 270485 72133 270541 72189
rect 270627 72133 270683 72189
rect 270769 72133 270825 72189
rect 270911 72133 270967 72189
rect 271053 72133 271109 72189
rect 271195 72133 271251 72189
rect 271337 72133 271393 72189
rect 271479 72133 271535 72189
rect 271621 72133 271677 72189
rect 271763 72133 271819 72189
rect 271905 72133 271961 72189
rect 272047 72133 272103 72189
rect 273249 73979 273305 74035
rect 273391 73979 273447 74035
rect 273533 73979 273589 74035
rect 273675 73979 273731 74035
rect 273817 73979 273873 74035
rect 273959 73979 274015 74035
rect 274101 73979 274157 74035
rect 274243 73979 274299 74035
rect 274385 73979 274441 74035
rect 274527 73979 274583 74035
rect 274669 73979 274725 74035
rect 273249 73837 273305 73893
rect 273391 73837 273447 73893
rect 273533 73837 273589 73893
rect 273675 73837 273731 73893
rect 273817 73837 273873 73893
rect 273959 73837 274015 73893
rect 274101 73837 274157 73893
rect 274243 73837 274299 73893
rect 274385 73837 274441 73893
rect 274527 73837 274583 73893
rect 274669 73837 274725 73893
rect 273249 73695 273305 73751
rect 273391 73695 273447 73751
rect 273533 73695 273589 73751
rect 273675 73695 273731 73751
rect 273817 73695 273873 73751
rect 273959 73695 274015 73751
rect 274101 73695 274157 73751
rect 274243 73695 274299 73751
rect 274385 73695 274441 73751
rect 274527 73695 274583 73751
rect 274669 73695 274725 73751
rect 273249 73553 273305 73609
rect 273391 73553 273447 73609
rect 273533 73553 273589 73609
rect 273675 73553 273731 73609
rect 273817 73553 273873 73609
rect 273959 73553 274015 73609
rect 274101 73553 274157 73609
rect 274243 73553 274299 73609
rect 274385 73553 274441 73609
rect 274527 73553 274583 73609
rect 274669 73553 274725 73609
rect 273249 73411 273305 73467
rect 273391 73411 273447 73467
rect 273533 73411 273589 73467
rect 273675 73411 273731 73467
rect 273817 73411 273873 73467
rect 273959 73411 274015 73467
rect 274101 73411 274157 73467
rect 274243 73411 274299 73467
rect 274385 73411 274441 73467
rect 274527 73411 274583 73467
rect 274669 73411 274725 73467
rect 273249 73269 273305 73325
rect 273391 73269 273447 73325
rect 273533 73269 273589 73325
rect 273675 73269 273731 73325
rect 273817 73269 273873 73325
rect 273959 73269 274015 73325
rect 274101 73269 274157 73325
rect 274243 73269 274299 73325
rect 274385 73269 274441 73325
rect 274527 73269 274583 73325
rect 274669 73269 274725 73325
rect 273249 73127 273305 73183
rect 273391 73127 273447 73183
rect 273533 73127 273589 73183
rect 273675 73127 273731 73183
rect 273817 73127 273873 73183
rect 273959 73127 274015 73183
rect 274101 73127 274157 73183
rect 274243 73127 274299 73183
rect 274385 73127 274441 73183
rect 274527 73127 274583 73183
rect 274669 73127 274725 73183
rect 273249 72985 273305 73041
rect 273391 72985 273447 73041
rect 273533 72985 273589 73041
rect 273675 72985 273731 73041
rect 273817 72985 273873 73041
rect 273959 72985 274015 73041
rect 274101 72985 274157 73041
rect 274243 72985 274299 73041
rect 274385 72985 274441 73041
rect 274527 72985 274583 73041
rect 274669 72985 274725 73041
rect 273249 72843 273305 72899
rect 273391 72843 273447 72899
rect 273533 72843 273589 72899
rect 273675 72843 273731 72899
rect 273817 72843 273873 72899
rect 273959 72843 274015 72899
rect 274101 72843 274157 72899
rect 274243 72843 274299 72899
rect 274385 72843 274441 72899
rect 274527 72843 274583 72899
rect 274669 72843 274725 72899
rect 273249 72701 273305 72757
rect 273391 72701 273447 72757
rect 273533 72701 273589 72757
rect 273675 72701 273731 72757
rect 273817 72701 273873 72757
rect 273959 72701 274015 72757
rect 274101 72701 274157 72757
rect 274243 72701 274299 72757
rect 274385 72701 274441 72757
rect 274527 72701 274583 72757
rect 274669 72701 274725 72757
rect 273249 72559 273305 72615
rect 273391 72559 273447 72615
rect 273533 72559 273589 72615
rect 273675 72559 273731 72615
rect 273817 72559 273873 72615
rect 273959 72559 274015 72615
rect 274101 72559 274157 72615
rect 274243 72559 274299 72615
rect 274385 72559 274441 72615
rect 274527 72559 274583 72615
rect 274669 72559 274725 72615
rect 273249 72417 273305 72473
rect 273391 72417 273447 72473
rect 273533 72417 273589 72473
rect 273675 72417 273731 72473
rect 273817 72417 273873 72473
rect 273959 72417 274015 72473
rect 274101 72417 274157 72473
rect 274243 72417 274299 72473
rect 274385 72417 274441 72473
rect 274527 72417 274583 72473
rect 274669 72417 274725 72473
rect 273249 72275 273305 72331
rect 273391 72275 273447 72331
rect 273533 72275 273589 72331
rect 273675 72275 273731 72331
rect 273817 72275 273873 72331
rect 273959 72275 274015 72331
rect 274101 72275 274157 72331
rect 274243 72275 274299 72331
rect 274385 72275 274441 72331
rect 274527 72275 274583 72331
rect 274669 72275 274725 72331
rect 273249 72133 273305 72189
rect 273391 72133 273447 72189
rect 273533 72133 273589 72189
rect 273675 72133 273731 72189
rect 273817 72133 273873 72189
rect 273959 72133 274015 72189
rect 274101 72133 274157 72189
rect 274243 72133 274299 72189
rect 274385 72133 274441 72189
rect 274527 72133 274583 72189
rect 274669 72133 274725 72189
rect 275193 73979 275249 74035
rect 275335 73979 275391 74035
rect 275477 73979 275533 74035
rect 275619 73979 275675 74035
rect 275761 73979 275817 74035
rect 275903 73979 275959 74035
rect 276045 73979 276101 74035
rect 276187 73979 276243 74035
rect 276329 73979 276385 74035
rect 276471 73979 276527 74035
rect 276613 73979 276669 74035
rect 276755 73979 276811 74035
rect 276897 73979 276953 74035
rect 277039 73979 277095 74035
rect 275193 73837 275249 73893
rect 275335 73837 275391 73893
rect 275477 73837 275533 73893
rect 275619 73837 275675 73893
rect 275761 73837 275817 73893
rect 275903 73837 275959 73893
rect 276045 73837 276101 73893
rect 276187 73837 276243 73893
rect 276329 73837 276385 73893
rect 276471 73837 276527 73893
rect 276613 73837 276669 73893
rect 276755 73837 276811 73893
rect 276897 73837 276953 73893
rect 277039 73837 277095 73893
rect 275193 73695 275249 73751
rect 275335 73695 275391 73751
rect 275477 73695 275533 73751
rect 275619 73695 275675 73751
rect 275761 73695 275817 73751
rect 275903 73695 275959 73751
rect 276045 73695 276101 73751
rect 276187 73695 276243 73751
rect 276329 73695 276385 73751
rect 276471 73695 276527 73751
rect 276613 73695 276669 73751
rect 276755 73695 276811 73751
rect 276897 73695 276953 73751
rect 277039 73695 277095 73751
rect 275193 73553 275249 73609
rect 275335 73553 275391 73609
rect 275477 73553 275533 73609
rect 275619 73553 275675 73609
rect 275761 73553 275817 73609
rect 275903 73553 275959 73609
rect 276045 73553 276101 73609
rect 276187 73553 276243 73609
rect 276329 73553 276385 73609
rect 276471 73553 276527 73609
rect 276613 73553 276669 73609
rect 276755 73553 276811 73609
rect 276897 73553 276953 73609
rect 277039 73553 277095 73609
rect 275193 73411 275249 73467
rect 275335 73411 275391 73467
rect 275477 73411 275533 73467
rect 275619 73411 275675 73467
rect 275761 73411 275817 73467
rect 275903 73411 275959 73467
rect 276045 73411 276101 73467
rect 276187 73411 276243 73467
rect 276329 73411 276385 73467
rect 276471 73411 276527 73467
rect 276613 73411 276669 73467
rect 276755 73411 276811 73467
rect 276897 73411 276953 73467
rect 277039 73411 277095 73467
rect 275193 73269 275249 73325
rect 275335 73269 275391 73325
rect 275477 73269 275533 73325
rect 275619 73269 275675 73325
rect 275761 73269 275817 73325
rect 275903 73269 275959 73325
rect 276045 73269 276101 73325
rect 276187 73269 276243 73325
rect 276329 73269 276385 73325
rect 276471 73269 276527 73325
rect 276613 73269 276669 73325
rect 276755 73269 276811 73325
rect 276897 73269 276953 73325
rect 277039 73269 277095 73325
rect 275193 73127 275249 73183
rect 275335 73127 275391 73183
rect 275477 73127 275533 73183
rect 275619 73127 275675 73183
rect 275761 73127 275817 73183
rect 275903 73127 275959 73183
rect 276045 73127 276101 73183
rect 276187 73127 276243 73183
rect 276329 73127 276385 73183
rect 276471 73127 276527 73183
rect 276613 73127 276669 73183
rect 276755 73127 276811 73183
rect 276897 73127 276953 73183
rect 277039 73127 277095 73183
rect 275193 72985 275249 73041
rect 275335 72985 275391 73041
rect 275477 72985 275533 73041
rect 275619 72985 275675 73041
rect 275761 72985 275817 73041
rect 275903 72985 275959 73041
rect 276045 72985 276101 73041
rect 276187 72985 276243 73041
rect 276329 72985 276385 73041
rect 276471 72985 276527 73041
rect 276613 72985 276669 73041
rect 276755 72985 276811 73041
rect 276897 72985 276953 73041
rect 277039 72985 277095 73041
rect 275193 72843 275249 72899
rect 275335 72843 275391 72899
rect 275477 72843 275533 72899
rect 275619 72843 275675 72899
rect 275761 72843 275817 72899
rect 275903 72843 275959 72899
rect 276045 72843 276101 72899
rect 276187 72843 276243 72899
rect 276329 72843 276385 72899
rect 276471 72843 276527 72899
rect 276613 72843 276669 72899
rect 276755 72843 276811 72899
rect 276897 72843 276953 72899
rect 277039 72843 277095 72899
rect 275193 72701 275249 72757
rect 275335 72701 275391 72757
rect 275477 72701 275533 72757
rect 275619 72701 275675 72757
rect 275761 72701 275817 72757
rect 275903 72701 275959 72757
rect 276045 72701 276101 72757
rect 276187 72701 276243 72757
rect 276329 72701 276385 72757
rect 276471 72701 276527 72757
rect 276613 72701 276669 72757
rect 276755 72701 276811 72757
rect 276897 72701 276953 72757
rect 277039 72701 277095 72757
rect 275193 72559 275249 72615
rect 275335 72559 275391 72615
rect 275477 72559 275533 72615
rect 275619 72559 275675 72615
rect 275761 72559 275817 72615
rect 275903 72559 275959 72615
rect 276045 72559 276101 72615
rect 276187 72559 276243 72615
rect 276329 72559 276385 72615
rect 276471 72559 276527 72615
rect 276613 72559 276669 72615
rect 276755 72559 276811 72615
rect 276897 72559 276953 72615
rect 277039 72559 277095 72615
rect 275193 72417 275249 72473
rect 275335 72417 275391 72473
rect 275477 72417 275533 72473
rect 275619 72417 275675 72473
rect 275761 72417 275817 72473
rect 275903 72417 275959 72473
rect 276045 72417 276101 72473
rect 276187 72417 276243 72473
rect 276329 72417 276385 72473
rect 276471 72417 276527 72473
rect 276613 72417 276669 72473
rect 276755 72417 276811 72473
rect 276897 72417 276953 72473
rect 277039 72417 277095 72473
rect 275193 72275 275249 72331
rect 275335 72275 275391 72331
rect 275477 72275 275533 72331
rect 275619 72275 275675 72331
rect 275761 72275 275817 72331
rect 275903 72275 275959 72331
rect 276045 72275 276101 72331
rect 276187 72275 276243 72331
rect 276329 72275 276385 72331
rect 276471 72275 276527 72331
rect 276613 72275 276669 72331
rect 276755 72275 276811 72331
rect 276897 72275 276953 72331
rect 277039 72275 277095 72331
rect 275193 72133 275249 72189
rect 275335 72133 275391 72189
rect 275477 72133 275533 72189
rect 275619 72133 275675 72189
rect 275761 72133 275817 72189
rect 275903 72133 275959 72189
rect 276045 72133 276101 72189
rect 276187 72133 276243 72189
rect 276329 72133 276385 72189
rect 276471 72133 276527 72189
rect 276613 72133 276669 72189
rect 276755 72133 276811 72189
rect 276897 72133 276953 72189
rect 277039 72133 277095 72189
rect 277899 73979 277955 74035
rect 278041 73979 278097 74035
rect 278183 73979 278239 74035
rect 278325 73979 278381 74035
rect 278467 73979 278523 74035
rect 278609 73979 278665 74035
rect 278751 73979 278807 74035
rect 278893 73979 278949 74035
rect 279035 73979 279091 74035
rect 279177 73979 279233 74035
rect 279319 73979 279375 74035
rect 279461 73979 279517 74035
rect 279603 73979 279659 74035
rect 279745 73979 279801 74035
rect 277899 73837 277955 73893
rect 278041 73837 278097 73893
rect 278183 73837 278239 73893
rect 278325 73837 278381 73893
rect 278467 73837 278523 73893
rect 278609 73837 278665 73893
rect 278751 73837 278807 73893
rect 278893 73837 278949 73893
rect 279035 73837 279091 73893
rect 279177 73837 279233 73893
rect 279319 73837 279375 73893
rect 279461 73837 279517 73893
rect 279603 73837 279659 73893
rect 279745 73837 279801 73893
rect 277899 73695 277955 73751
rect 278041 73695 278097 73751
rect 278183 73695 278239 73751
rect 278325 73695 278381 73751
rect 278467 73695 278523 73751
rect 278609 73695 278665 73751
rect 278751 73695 278807 73751
rect 278893 73695 278949 73751
rect 279035 73695 279091 73751
rect 279177 73695 279233 73751
rect 279319 73695 279375 73751
rect 279461 73695 279517 73751
rect 279603 73695 279659 73751
rect 279745 73695 279801 73751
rect 277899 73553 277955 73609
rect 278041 73553 278097 73609
rect 278183 73553 278239 73609
rect 278325 73553 278381 73609
rect 278467 73553 278523 73609
rect 278609 73553 278665 73609
rect 278751 73553 278807 73609
rect 278893 73553 278949 73609
rect 279035 73553 279091 73609
rect 279177 73553 279233 73609
rect 279319 73553 279375 73609
rect 279461 73553 279517 73609
rect 279603 73553 279659 73609
rect 279745 73553 279801 73609
rect 277899 73411 277955 73467
rect 278041 73411 278097 73467
rect 278183 73411 278239 73467
rect 278325 73411 278381 73467
rect 278467 73411 278523 73467
rect 278609 73411 278665 73467
rect 278751 73411 278807 73467
rect 278893 73411 278949 73467
rect 279035 73411 279091 73467
rect 279177 73411 279233 73467
rect 279319 73411 279375 73467
rect 279461 73411 279517 73467
rect 279603 73411 279659 73467
rect 279745 73411 279801 73467
rect 277899 73269 277955 73325
rect 278041 73269 278097 73325
rect 278183 73269 278239 73325
rect 278325 73269 278381 73325
rect 278467 73269 278523 73325
rect 278609 73269 278665 73325
rect 278751 73269 278807 73325
rect 278893 73269 278949 73325
rect 279035 73269 279091 73325
rect 279177 73269 279233 73325
rect 279319 73269 279375 73325
rect 279461 73269 279517 73325
rect 279603 73269 279659 73325
rect 279745 73269 279801 73325
rect 277899 73127 277955 73183
rect 278041 73127 278097 73183
rect 278183 73127 278239 73183
rect 278325 73127 278381 73183
rect 278467 73127 278523 73183
rect 278609 73127 278665 73183
rect 278751 73127 278807 73183
rect 278893 73127 278949 73183
rect 279035 73127 279091 73183
rect 279177 73127 279233 73183
rect 279319 73127 279375 73183
rect 279461 73127 279517 73183
rect 279603 73127 279659 73183
rect 279745 73127 279801 73183
rect 277899 72985 277955 73041
rect 278041 72985 278097 73041
rect 278183 72985 278239 73041
rect 278325 72985 278381 73041
rect 278467 72985 278523 73041
rect 278609 72985 278665 73041
rect 278751 72985 278807 73041
rect 278893 72985 278949 73041
rect 279035 72985 279091 73041
rect 279177 72985 279233 73041
rect 279319 72985 279375 73041
rect 279461 72985 279517 73041
rect 279603 72985 279659 73041
rect 279745 72985 279801 73041
rect 277899 72843 277955 72899
rect 278041 72843 278097 72899
rect 278183 72843 278239 72899
rect 278325 72843 278381 72899
rect 278467 72843 278523 72899
rect 278609 72843 278665 72899
rect 278751 72843 278807 72899
rect 278893 72843 278949 72899
rect 279035 72843 279091 72899
rect 279177 72843 279233 72899
rect 279319 72843 279375 72899
rect 279461 72843 279517 72899
rect 279603 72843 279659 72899
rect 279745 72843 279801 72899
rect 277899 72701 277955 72757
rect 278041 72701 278097 72757
rect 278183 72701 278239 72757
rect 278325 72701 278381 72757
rect 278467 72701 278523 72757
rect 278609 72701 278665 72757
rect 278751 72701 278807 72757
rect 278893 72701 278949 72757
rect 279035 72701 279091 72757
rect 279177 72701 279233 72757
rect 279319 72701 279375 72757
rect 279461 72701 279517 72757
rect 279603 72701 279659 72757
rect 279745 72701 279801 72757
rect 277899 72559 277955 72615
rect 278041 72559 278097 72615
rect 278183 72559 278239 72615
rect 278325 72559 278381 72615
rect 278467 72559 278523 72615
rect 278609 72559 278665 72615
rect 278751 72559 278807 72615
rect 278893 72559 278949 72615
rect 279035 72559 279091 72615
rect 279177 72559 279233 72615
rect 279319 72559 279375 72615
rect 279461 72559 279517 72615
rect 279603 72559 279659 72615
rect 279745 72559 279801 72615
rect 277899 72417 277955 72473
rect 278041 72417 278097 72473
rect 278183 72417 278239 72473
rect 278325 72417 278381 72473
rect 278467 72417 278523 72473
rect 278609 72417 278665 72473
rect 278751 72417 278807 72473
rect 278893 72417 278949 72473
rect 279035 72417 279091 72473
rect 279177 72417 279233 72473
rect 279319 72417 279375 72473
rect 279461 72417 279517 72473
rect 279603 72417 279659 72473
rect 279745 72417 279801 72473
rect 277899 72275 277955 72331
rect 278041 72275 278097 72331
rect 278183 72275 278239 72331
rect 278325 72275 278381 72331
rect 278467 72275 278523 72331
rect 278609 72275 278665 72331
rect 278751 72275 278807 72331
rect 278893 72275 278949 72331
rect 279035 72275 279091 72331
rect 279177 72275 279233 72331
rect 279319 72275 279375 72331
rect 279461 72275 279517 72331
rect 279603 72275 279659 72331
rect 279745 72275 279801 72331
rect 277899 72133 277955 72189
rect 278041 72133 278097 72189
rect 278183 72133 278239 72189
rect 278325 72133 278381 72189
rect 278467 72133 278523 72189
rect 278609 72133 278665 72189
rect 278751 72133 278807 72189
rect 278893 72133 278949 72189
rect 279035 72133 279091 72189
rect 279177 72133 279233 72189
rect 279319 72133 279375 72189
rect 279461 72133 279517 72189
rect 279603 72133 279659 72189
rect 279745 72133 279801 72189
rect 280269 73979 280325 74035
rect 280411 73979 280467 74035
rect 280553 73979 280609 74035
rect 280695 73979 280751 74035
rect 280837 73979 280893 74035
rect 280979 73979 281035 74035
rect 281121 73979 281177 74035
rect 281263 73979 281319 74035
rect 281405 73979 281461 74035
rect 281547 73979 281603 74035
rect 281689 73979 281745 74035
rect 281831 73979 281887 74035
rect 281973 73979 282029 74035
rect 282115 73979 282171 74035
rect 280269 73837 280325 73893
rect 280411 73837 280467 73893
rect 280553 73837 280609 73893
rect 280695 73837 280751 73893
rect 280837 73837 280893 73893
rect 280979 73837 281035 73893
rect 281121 73837 281177 73893
rect 281263 73837 281319 73893
rect 281405 73837 281461 73893
rect 281547 73837 281603 73893
rect 281689 73837 281745 73893
rect 281831 73837 281887 73893
rect 281973 73837 282029 73893
rect 282115 73837 282171 73893
rect 280269 73695 280325 73751
rect 280411 73695 280467 73751
rect 280553 73695 280609 73751
rect 280695 73695 280751 73751
rect 280837 73695 280893 73751
rect 280979 73695 281035 73751
rect 281121 73695 281177 73751
rect 281263 73695 281319 73751
rect 281405 73695 281461 73751
rect 281547 73695 281603 73751
rect 281689 73695 281745 73751
rect 281831 73695 281887 73751
rect 281973 73695 282029 73751
rect 282115 73695 282171 73751
rect 280269 73553 280325 73609
rect 280411 73553 280467 73609
rect 280553 73553 280609 73609
rect 280695 73553 280751 73609
rect 280837 73553 280893 73609
rect 280979 73553 281035 73609
rect 281121 73553 281177 73609
rect 281263 73553 281319 73609
rect 281405 73553 281461 73609
rect 281547 73553 281603 73609
rect 281689 73553 281745 73609
rect 281831 73553 281887 73609
rect 281973 73553 282029 73609
rect 282115 73553 282171 73609
rect 280269 73411 280325 73467
rect 280411 73411 280467 73467
rect 280553 73411 280609 73467
rect 280695 73411 280751 73467
rect 280837 73411 280893 73467
rect 280979 73411 281035 73467
rect 281121 73411 281177 73467
rect 281263 73411 281319 73467
rect 281405 73411 281461 73467
rect 281547 73411 281603 73467
rect 281689 73411 281745 73467
rect 281831 73411 281887 73467
rect 281973 73411 282029 73467
rect 282115 73411 282171 73467
rect 280269 73269 280325 73325
rect 280411 73269 280467 73325
rect 280553 73269 280609 73325
rect 280695 73269 280751 73325
rect 280837 73269 280893 73325
rect 280979 73269 281035 73325
rect 281121 73269 281177 73325
rect 281263 73269 281319 73325
rect 281405 73269 281461 73325
rect 281547 73269 281603 73325
rect 281689 73269 281745 73325
rect 281831 73269 281887 73325
rect 281973 73269 282029 73325
rect 282115 73269 282171 73325
rect 280269 73127 280325 73183
rect 280411 73127 280467 73183
rect 280553 73127 280609 73183
rect 280695 73127 280751 73183
rect 280837 73127 280893 73183
rect 280979 73127 281035 73183
rect 281121 73127 281177 73183
rect 281263 73127 281319 73183
rect 281405 73127 281461 73183
rect 281547 73127 281603 73183
rect 281689 73127 281745 73183
rect 281831 73127 281887 73183
rect 281973 73127 282029 73183
rect 282115 73127 282171 73183
rect 280269 72985 280325 73041
rect 280411 72985 280467 73041
rect 280553 72985 280609 73041
rect 280695 72985 280751 73041
rect 280837 72985 280893 73041
rect 280979 72985 281035 73041
rect 281121 72985 281177 73041
rect 281263 72985 281319 73041
rect 281405 72985 281461 73041
rect 281547 72985 281603 73041
rect 281689 72985 281745 73041
rect 281831 72985 281887 73041
rect 281973 72985 282029 73041
rect 282115 72985 282171 73041
rect 280269 72843 280325 72899
rect 280411 72843 280467 72899
rect 280553 72843 280609 72899
rect 280695 72843 280751 72899
rect 280837 72843 280893 72899
rect 280979 72843 281035 72899
rect 281121 72843 281177 72899
rect 281263 72843 281319 72899
rect 281405 72843 281461 72899
rect 281547 72843 281603 72899
rect 281689 72843 281745 72899
rect 281831 72843 281887 72899
rect 281973 72843 282029 72899
rect 282115 72843 282171 72899
rect 280269 72701 280325 72757
rect 280411 72701 280467 72757
rect 280553 72701 280609 72757
rect 280695 72701 280751 72757
rect 280837 72701 280893 72757
rect 280979 72701 281035 72757
rect 281121 72701 281177 72757
rect 281263 72701 281319 72757
rect 281405 72701 281461 72757
rect 281547 72701 281603 72757
rect 281689 72701 281745 72757
rect 281831 72701 281887 72757
rect 281973 72701 282029 72757
rect 282115 72701 282171 72757
rect 280269 72559 280325 72615
rect 280411 72559 280467 72615
rect 280553 72559 280609 72615
rect 280695 72559 280751 72615
rect 280837 72559 280893 72615
rect 280979 72559 281035 72615
rect 281121 72559 281177 72615
rect 281263 72559 281319 72615
rect 281405 72559 281461 72615
rect 281547 72559 281603 72615
rect 281689 72559 281745 72615
rect 281831 72559 281887 72615
rect 281973 72559 282029 72615
rect 282115 72559 282171 72615
rect 280269 72417 280325 72473
rect 280411 72417 280467 72473
rect 280553 72417 280609 72473
rect 280695 72417 280751 72473
rect 280837 72417 280893 72473
rect 280979 72417 281035 72473
rect 281121 72417 281177 72473
rect 281263 72417 281319 72473
rect 281405 72417 281461 72473
rect 281547 72417 281603 72473
rect 281689 72417 281745 72473
rect 281831 72417 281887 72473
rect 281973 72417 282029 72473
rect 282115 72417 282171 72473
rect 280269 72275 280325 72331
rect 280411 72275 280467 72331
rect 280553 72275 280609 72331
rect 280695 72275 280751 72331
rect 280837 72275 280893 72331
rect 280979 72275 281035 72331
rect 281121 72275 281177 72331
rect 281263 72275 281319 72331
rect 281405 72275 281461 72331
rect 281547 72275 281603 72331
rect 281689 72275 281745 72331
rect 281831 72275 281887 72331
rect 281973 72275 282029 72331
rect 282115 72275 282171 72331
rect 280269 72133 280325 72189
rect 280411 72133 280467 72189
rect 280553 72133 280609 72189
rect 280695 72133 280751 72189
rect 280837 72133 280893 72189
rect 280979 72133 281035 72189
rect 281121 72133 281177 72189
rect 281263 72133 281319 72189
rect 281405 72133 281461 72189
rect 281547 72133 281603 72189
rect 281689 72133 281745 72189
rect 281831 72133 281887 72189
rect 281973 72133 282029 72189
rect 282115 72133 282171 72189
rect 282899 73979 282955 74035
rect 283041 73979 283097 74035
rect 283183 73979 283239 74035
rect 283325 73979 283381 74035
rect 283467 73979 283523 74035
rect 283609 73979 283665 74035
rect 283751 73979 283807 74035
rect 283893 73979 283949 74035
rect 282899 73837 282955 73893
rect 283041 73837 283097 73893
rect 283183 73837 283239 73893
rect 283325 73837 283381 73893
rect 283467 73837 283523 73893
rect 283609 73837 283665 73893
rect 283751 73837 283807 73893
rect 283893 73837 283949 73893
rect 282899 73695 282955 73751
rect 283041 73695 283097 73751
rect 283183 73695 283239 73751
rect 283325 73695 283381 73751
rect 283467 73695 283523 73751
rect 283609 73695 283665 73751
rect 283751 73695 283807 73751
rect 283893 73695 283949 73751
rect 282899 73553 282955 73609
rect 283041 73553 283097 73609
rect 283183 73553 283239 73609
rect 283325 73553 283381 73609
rect 283467 73553 283523 73609
rect 283609 73553 283665 73609
rect 283751 73553 283807 73609
rect 283893 73553 283949 73609
rect 282899 73411 282955 73467
rect 283041 73411 283097 73467
rect 283183 73411 283239 73467
rect 283325 73411 283381 73467
rect 283467 73411 283523 73467
rect 283609 73411 283665 73467
rect 283751 73411 283807 73467
rect 283893 73411 283949 73467
rect 282899 73269 282955 73325
rect 283041 73269 283097 73325
rect 283183 73269 283239 73325
rect 283325 73269 283381 73325
rect 283467 73269 283523 73325
rect 283609 73269 283665 73325
rect 283751 73269 283807 73325
rect 283893 73269 283949 73325
rect 282899 73127 282955 73183
rect 283041 73127 283097 73183
rect 283183 73127 283239 73183
rect 283325 73127 283381 73183
rect 283467 73127 283523 73183
rect 283609 73127 283665 73183
rect 283751 73127 283807 73183
rect 283893 73127 283949 73183
rect 282899 72985 282955 73041
rect 283041 72985 283097 73041
rect 283183 72985 283239 73041
rect 283325 72985 283381 73041
rect 283467 72985 283523 73041
rect 283609 72985 283665 73041
rect 283751 72985 283807 73041
rect 283893 72985 283949 73041
rect 282899 72843 282955 72899
rect 283041 72843 283097 72899
rect 283183 72843 283239 72899
rect 283325 72843 283381 72899
rect 283467 72843 283523 72899
rect 283609 72843 283665 72899
rect 283751 72843 283807 72899
rect 283893 72843 283949 72899
rect 282899 72701 282955 72757
rect 283041 72701 283097 72757
rect 283183 72701 283239 72757
rect 283325 72701 283381 72757
rect 283467 72701 283523 72757
rect 283609 72701 283665 72757
rect 283751 72701 283807 72757
rect 283893 72701 283949 72757
rect 282899 72559 282955 72615
rect 283041 72559 283097 72615
rect 283183 72559 283239 72615
rect 283325 72559 283381 72615
rect 283467 72559 283523 72615
rect 283609 72559 283665 72615
rect 283751 72559 283807 72615
rect 283893 72559 283949 72615
rect 282899 72417 282955 72473
rect 283041 72417 283097 72473
rect 283183 72417 283239 72473
rect 283325 72417 283381 72473
rect 283467 72417 283523 72473
rect 283609 72417 283665 72473
rect 283751 72417 283807 72473
rect 283893 72417 283949 72473
rect 282899 72275 282955 72331
rect 283041 72275 283097 72331
rect 283183 72275 283239 72331
rect 283325 72275 283381 72331
rect 283467 72275 283523 72331
rect 283609 72275 283665 72331
rect 283751 72275 283807 72331
rect 283893 72275 283949 72331
rect 282899 72133 282955 72189
rect 283041 72133 283097 72189
rect 283183 72133 283239 72189
rect 283325 72133 283381 72189
rect 283467 72133 283523 72189
rect 283609 72133 283665 72189
rect 283751 72133 283807 72189
rect 283893 72133 283949 72189
rect 600343 73979 600399 74035
rect 600485 73979 600541 74035
rect 600627 73979 600683 74035
rect 600769 73979 600825 74035
rect 600911 73979 600967 74035
rect 601053 73979 601109 74035
rect 601195 73979 601251 74035
rect 601337 73979 601393 74035
rect 601479 73979 601535 74035
rect 601621 73979 601677 74035
rect 601763 73979 601819 74035
rect 601905 73979 601961 74035
rect 602047 73979 602103 74035
rect 600343 73837 600399 73893
rect 600485 73837 600541 73893
rect 600627 73837 600683 73893
rect 600769 73837 600825 73893
rect 600911 73837 600967 73893
rect 601053 73837 601109 73893
rect 601195 73837 601251 73893
rect 601337 73837 601393 73893
rect 601479 73837 601535 73893
rect 601621 73837 601677 73893
rect 601763 73837 601819 73893
rect 601905 73837 601961 73893
rect 602047 73837 602103 73893
rect 600343 73695 600399 73751
rect 600485 73695 600541 73751
rect 600627 73695 600683 73751
rect 600769 73695 600825 73751
rect 600911 73695 600967 73751
rect 601053 73695 601109 73751
rect 601195 73695 601251 73751
rect 601337 73695 601393 73751
rect 601479 73695 601535 73751
rect 601621 73695 601677 73751
rect 601763 73695 601819 73751
rect 601905 73695 601961 73751
rect 602047 73695 602103 73751
rect 600343 73553 600399 73609
rect 600485 73553 600541 73609
rect 600627 73553 600683 73609
rect 600769 73553 600825 73609
rect 600911 73553 600967 73609
rect 601053 73553 601109 73609
rect 601195 73553 601251 73609
rect 601337 73553 601393 73609
rect 601479 73553 601535 73609
rect 601621 73553 601677 73609
rect 601763 73553 601819 73609
rect 601905 73553 601961 73609
rect 602047 73553 602103 73609
rect 600343 73411 600399 73467
rect 600485 73411 600541 73467
rect 600627 73411 600683 73467
rect 600769 73411 600825 73467
rect 600911 73411 600967 73467
rect 601053 73411 601109 73467
rect 601195 73411 601251 73467
rect 601337 73411 601393 73467
rect 601479 73411 601535 73467
rect 601621 73411 601677 73467
rect 601763 73411 601819 73467
rect 601905 73411 601961 73467
rect 602047 73411 602103 73467
rect 600343 73269 600399 73325
rect 600485 73269 600541 73325
rect 600627 73269 600683 73325
rect 600769 73269 600825 73325
rect 600911 73269 600967 73325
rect 601053 73269 601109 73325
rect 601195 73269 601251 73325
rect 601337 73269 601393 73325
rect 601479 73269 601535 73325
rect 601621 73269 601677 73325
rect 601763 73269 601819 73325
rect 601905 73269 601961 73325
rect 602047 73269 602103 73325
rect 600343 73127 600399 73183
rect 600485 73127 600541 73183
rect 600627 73127 600683 73183
rect 600769 73127 600825 73183
rect 600911 73127 600967 73183
rect 601053 73127 601109 73183
rect 601195 73127 601251 73183
rect 601337 73127 601393 73183
rect 601479 73127 601535 73183
rect 601621 73127 601677 73183
rect 601763 73127 601819 73183
rect 601905 73127 601961 73183
rect 602047 73127 602103 73183
rect 600343 72985 600399 73041
rect 600485 72985 600541 73041
rect 600627 72985 600683 73041
rect 600769 72985 600825 73041
rect 600911 72985 600967 73041
rect 601053 72985 601109 73041
rect 601195 72985 601251 73041
rect 601337 72985 601393 73041
rect 601479 72985 601535 73041
rect 601621 72985 601677 73041
rect 601763 72985 601819 73041
rect 601905 72985 601961 73041
rect 602047 72985 602103 73041
rect 600343 72843 600399 72899
rect 600485 72843 600541 72899
rect 600627 72843 600683 72899
rect 600769 72843 600825 72899
rect 600911 72843 600967 72899
rect 601053 72843 601109 72899
rect 601195 72843 601251 72899
rect 601337 72843 601393 72899
rect 601479 72843 601535 72899
rect 601621 72843 601677 72899
rect 601763 72843 601819 72899
rect 601905 72843 601961 72899
rect 602047 72843 602103 72899
rect 600343 72701 600399 72757
rect 600485 72701 600541 72757
rect 600627 72701 600683 72757
rect 600769 72701 600825 72757
rect 600911 72701 600967 72757
rect 601053 72701 601109 72757
rect 601195 72701 601251 72757
rect 601337 72701 601393 72757
rect 601479 72701 601535 72757
rect 601621 72701 601677 72757
rect 601763 72701 601819 72757
rect 601905 72701 601961 72757
rect 602047 72701 602103 72757
rect 600343 72559 600399 72615
rect 600485 72559 600541 72615
rect 600627 72559 600683 72615
rect 600769 72559 600825 72615
rect 600911 72559 600967 72615
rect 601053 72559 601109 72615
rect 601195 72559 601251 72615
rect 601337 72559 601393 72615
rect 601479 72559 601535 72615
rect 601621 72559 601677 72615
rect 601763 72559 601819 72615
rect 601905 72559 601961 72615
rect 602047 72559 602103 72615
rect 600343 72417 600399 72473
rect 600485 72417 600541 72473
rect 600627 72417 600683 72473
rect 600769 72417 600825 72473
rect 600911 72417 600967 72473
rect 601053 72417 601109 72473
rect 601195 72417 601251 72473
rect 601337 72417 601393 72473
rect 601479 72417 601535 72473
rect 601621 72417 601677 72473
rect 601763 72417 601819 72473
rect 601905 72417 601961 72473
rect 602047 72417 602103 72473
rect 600343 72275 600399 72331
rect 600485 72275 600541 72331
rect 600627 72275 600683 72331
rect 600769 72275 600825 72331
rect 600911 72275 600967 72331
rect 601053 72275 601109 72331
rect 601195 72275 601251 72331
rect 601337 72275 601393 72331
rect 601479 72275 601535 72331
rect 601621 72275 601677 72331
rect 601763 72275 601819 72331
rect 601905 72275 601961 72331
rect 602047 72275 602103 72331
rect 600343 72133 600399 72189
rect 600485 72133 600541 72189
rect 600627 72133 600683 72189
rect 600769 72133 600825 72189
rect 600911 72133 600967 72189
rect 601053 72133 601109 72189
rect 601195 72133 601251 72189
rect 601337 72133 601393 72189
rect 601479 72133 601535 72189
rect 601621 72133 601677 72189
rect 601763 72133 601819 72189
rect 601905 72133 601961 72189
rect 602047 72133 602103 72189
rect 602823 73979 602879 74035
rect 602965 73979 603021 74035
rect 603107 73979 603163 74035
rect 603249 73979 603305 74035
rect 603391 73979 603447 74035
rect 603533 73979 603589 74035
rect 603675 73979 603731 74035
rect 603817 73979 603873 74035
rect 603959 73979 604015 74035
rect 602823 73837 602879 73893
rect 602965 73837 603021 73893
rect 603107 73837 603163 73893
rect 603249 73837 603305 73893
rect 603391 73837 603447 73893
rect 603533 73837 603589 73893
rect 603675 73837 603731 73893
rect 603817 73837 603873 73893
rect 603959 73837 604015 73893
rect 602823 73695 602879 73751
rect 602965 73695 603021 73751
rect 603107 73695 603163 73751
rect 603249 73695 603305 73751
rect 603391 73695 603447 73751
rect 603533 73695 603589 73751
rect 603675 73695 603731 73751
rect 603817 73695 603873 73751
rect 603959 73695 604015 73751
rect 602823 73553 602879 73609
rect 602965 73553 603021 73609
rect 603107 73553 603163 73609
rect 603249 73553 603305 73609
rect 603391 73553 603447 73609
rect 603533 73553 603589 73609
rect 603675 73553 603731 73609
rect 603817 73553 603873 73609
rect 603959 73553 604015 73609
rect 602823 73411 602879 73467
rect 602965 73411 603021 73467
rect 603107 73411 603163 73467
rect 603249 73411 603305 73467
rect 603391 73411 603447 73467
rect 603533 73411 603589 73467
rect 603675 73411 603731 73467
rect 603817 73411 603873 73467
rect 603959 73411 604015 73467
rect 602823 73269 602879 73325
rect 602965 73269 603021 73325
rect 603107 73269 603163 73325
rect 603249 73269 603305 73325
rect 603391 73269 603447 73325
rect 603533 73269 603589 73325
rect 603675 73269 603731 73325
rect 603817 73269 603873 73325
rect 603959 73269 604015 73325
rect 602823 73127 602879 73183
rect 602965 73127 603021 73183
rect 603107 73127 603163 73183
rect 603249 73127 603305 73183
rect 603391 73127 603447 73183
rect 603533 73127 603589 73183
rect 603675 73127 603731 73183
rect 603817 73127 603873 73183
rect 603959 73127 604015 73183
rect 602823 72985 602879 73041
rect 602965 72985 603021 73041
rect 603107 72985 603163 73041
rect 603249 72985 603305 73041
rect 603391 72985 603447 73041
rect 603533 72985 603589 73041
rect 603675 72985 603731 73041
rect 603817 72985 603873 73041
rect 603959 72985 604015 73041
rect 602823 72843 602879 72899
rect 602965 72843 603021 72899
rect 603107 72843 603163 72899
rect 603249 72843 603305 72899
rect 603391 72843 603447 72899
rect 603533 72843 603589 72899
rect 603675 72843 603731 72899
rect 603817 72843 603873 72899
rect 603959 72843 604015 72899
rect 602823 72701 602879 72757
rect 602965 72701 603021 72757
rect 603107 72701 603163 72757
rect 603249 72701 603305 72757
rect 603391 72701 603447 72757
rect 603533 72701 603589 72757
rect 603675 72701 603731 72757
rect 603817 72701 603873 72757
rect 603959 72701 604015 72757
rect 602823 72559 602879 72615
rect 602965 72559 603021 72615
rect 603107 72559 603163 72615
rect 603249 72559 603305 72615
rect 603391 72559 603447 72615
rect 603533 72559 603589 72615
rect 603675 72559 603731 72615
rect 603817 72559 603873 72615
rect 603959 72559 604015 72615
rect 602823 72417 602879 72473
rect 602965 72417 603021 72473
rect 603107 72417 603163 72473
rect 603249 72417 603305 72473
rect 603391 72417 603447 72473
rect 603533 72417 603589 72473
rect 603675 72417 603731 72473
rect 603817 72417 603873 72473
rect 603959 72417 604015 72473
rect 602823 72275 602879 72331
rect 602965 72275 603021 72331
rect 603107 72275 603163 72331
rect 603249 72275 603305 72331
rect 603391 72275 603447 72331
rect 603533 72275 603589 72331
rect 603675 72275 603731 72331
rect 603817 72275 603873 72331
rect 603959 72275 604015 72331
rect 602823 72133 602879 72189
rect 602965 72133 603021 72189
rect 603107 72133 603163 72189
rect 603249 72133 603305 72189
rect 603391 72133 603447 72189
rect 603533 72133 603589 72189
rect 603675 72133 603731 72189
rect 603817 72133 603873 72189
rect 603959 72133 604015 72189
rect 605193 73979 605249 74035
rect 605335 73979 605391 74035
rect 605477 73979 605533 74035
rect 605619 73979 605675 74035
rect 605761 73979 605817 74035
rect 605903 73979 605959 74035
rect 606045 73979 606101 74035
rect 606187 73979 606243 74035
rect 606329 73979 606385 74035
rect 606471 73979 606527 74035
rect 606613 73979 606669 74035
rect 606755 73979 606811 74035
rect 606897 73979 606953 74035
rect 607039 73979 607095 74035
rect 605193 73837 605249 73893
rect 605335 73837 605391 73893
rect 605477 73837 605533 73893
rect 605619 73837 605675 73893
rect 605761 73837 605817 73893
rect 605903 73837 605959 73893
rect 606045 73837 606101 73893
rect 606187 73837 606243 73893
rect 606329 73837 606385 73893
rect 606471 73837 606527 73893
rect 606613 73837 606669 73893
rect 606755 73837 606811 73893
rect 606897 73837 606953 73893
rect 607039 73837 607095 73893
rect 605193 73695 605249 73751
rect 605335 73695 605391 73751
rect 605477 73695 605533 73751
rect 605619 73695 605675 73751
rect 605761 73695 605817 73751
rect 605903 73695 605959 73751
rect 606045 73695 606101 73751
rect 606187 73695 606243 73751
rect 606329 73695 606385 73751
rect 606471 73695 606527 73751
rect 606613 73695 606669 73751
rect 606755 73695 606811 73751
rect 606897 73695 606953 73751
rect 607039 73695 607095 73751
rect 605193 73553 605249 73609
rect 605335 73553 605391 73609
rect 605477 73553 605533 73609
rect 605619 73553 605675 73609
rect 605761 73553 605817 73609
rect 605903 73553 605959 73609
rect 606045 73553 606101 73609
rect 606187 73553 606243 73609
rect 606329 73553 606385 73609
rect 606471 73553 606527 73609
rect 606613 73553 606669 73609
rect 606755 73553 606811 73609
rect 606897 73553 606953 73609
rect 607039 73553 607095 73609
rect 605193 73411 605249 73467
rect 605335 73411 605391 73467
rect 605477 73411 605533 73467
rect 605619 73411 605675 73467
rect 605761 73411 605817 73467
rect 605903 73411 605959 73467
rect 606045 73411 606101 73467
rect 606187 73411 606243 73467
rect 606329 73411 606385 73467
rect 606471 73411 606527 73467
rect 606613 73411 606669 73467
rect 606755 73411 606811 73467
rect 606897 73411 606953 73467
rect 607039 73411 607095 73467
rect 605193 73269 605249 73325
rect 605335 73269 605391 73325
rect 605477 73269 605533 73325
rect 605619 73269 605675 73325
rect 605761 73269 605817 73325
rect 605903 73269 605959 73325
rect 606045 73269 606101 73325
rect 606187 73269 606243 73325
rect 606329 73269 606385 73325
rect 606471 73269 606527 73325
rect 606613 73269 606669 73325
rect 606755 73269 606811 73325
rect 606897 73269 606953 73325
rect 607039 73269 607095 73325
rect 605193 73127 605249 73183
rect 605335 73127 605391 73183
rect 605477 73127 605533 73183
rect 605619 73127 605675 73183
rect 605761 73127 605817 73183
rect 605903 73127 605959 73183
rect 606045 73127 606101 73183
rect 606187 73127 606243 73183
rect 606329 73127 606385 73183
rect 606471 73127 606527 73183
rect 606613 73127 606669 73183
rect 606755 73127 606811 73183
rect 606897 73127 606953 73183
rect 607039 73127 607095 73183
rect 605193 72985 605249 73041
rect 605335 72985 605391 73041
rect 605477 72985 605533 73041
rect 605619 72985 605675 73041
rect 605761 72985 605817 73041
rect 605903 72985 605959 73041
rect 606045 72985 606101 73041
rect 606187 72985 606243 73041
rect 606329 72985 606385 73041
rect 606471 72985 606527 73041
rect 606613 72985 606669 73041
rect 606755 72985 606811 73041
rect 606897 72985 606953 73041
rect 607039 72985 607095 73041
rect 605193 72843 605249 72899
rect 605335 72843 605391 72899
rect 605477 72843 605533 72899
rect 605619 72843 605675 72899
rect 605761 72843 605817 72899
rect 605903 72843 605959 72899
rect 606045 72843 606101 72899
rect 606187 72843 606243 72899
rect 606329 72843 606385 72899
rect 606471 72843 606527 72899
rect 606613 72843 606669 72899
rect 606755 72843 606811 72899
rect 606897 72843 606953 72899
rect 607039 72843 607095 72899
rect 605193 72701 605249 72757
rect 605335 72701 605391 72757
rect 605477 72701 605533 72757
rect 605619 72701 605675 72757
rect 605761 72701 605817 72757
rect 605903 72701 605959 72757
rect 606045 72701 606101 72757
rect 606187 72701 606243 72757
rect 606329 72701 606385 72757
rect 606471 72701 606527 72757
rect 606613 72701 606669 72757
rect 606755 72701 606811 72757
rect 606897 72701 606953 72757
rect 607039 72701 607095 72757
rect 605193 72559 605249 72615
rect 605335 72559 605391 72615
rect 605477 72559 605533 72615
rect 605619 72559 605675 72615
rect 605761 72559 605817 72615
rect 605903 72559 605959 72615
rect 606045 72559 606101 72615
rect 606187 72559 606243 72615
rect 606329 72559 606385 72615
rect 606471 72559 606527 72615
rect 606613 72559 606669 72615
rect 606755 72559 606811 72615
rect 606897 72559 606953 72615
rect 607039 72559 607095 72615
rect 605193 72417 605249 72473
rect 605335 72417 605391 72473
rect 605477 72417 605533 72473
rect 605619 72417 605675 72473
rect 605761 72417 605817 72473
rect 605903 72417 605959 72473
rect 606045 72417 606101 72473
rect 606187 72417 606243 72473
rect 606329 72417 606385 72473
rect 606471 72417 606527 72473
rect 606613 72417 606669 72473
rect 606755 72417 606811 72473
rect 606897 72417 606953 72473
rect 607039 72417 607095 72473
rect 605193 72275 605249 72331
rect 605335 72275 605391 72331
rect 605477 72275 605533 72331
rect 605619 72275 605675 72331
rect 605761 72275 605817 72331
rect 605903 72275 605959 72331
rect 606045 72275 606101 72331
rect 606187 72275 606243 72331
rect 606329 72275 606385 72331
rect 606471 72275 606527 72331
rect 606613 72275 606669 72331
rect 606755 72275 606811 72331
rect 606897 72275 606953 72331
rect 607039 72275 607095 72331
rect 605193 72133 605249 72189
rect 605335 72133 605391 72189
rect 605477 72133 605533 72189
rect 605619 72133 605675 72189
rect 605761 72133 605817 72189
rect 605903 72133 605959 72189
rect 606045 72133 606101 72189
rect 606187 72133 606243 72189
rect 606329 72133 606385 72189
rect 606471 72133 606527 72189
rect 606613 72133 606669 72189
rect 606755 72133 606811 72189
rect 606897 72133 606953 72189
rect 607039 72133 607095 72189
rect 607899 73979 607955 74035
rect 608041 73979 608097 74035
rect 608183 73979 608239 74035
rect 608325 73979 608381 74035
rect 608467 73979 608523 74035
rect 609319 73979 609375 74035
rect 609461 73979 609517 74035
rect 609603 73979 609659 74035
rect 609745 73979 609801 74035
rect 607899 73837 607955 73893
rect 608041 73837 608097 73893
rect 608183 73837 608239 73893
rect 608325 73837 608381 73893
rect 608467 73837 608523 73893
rect 609319 73837 609375 73893
rect 609461 73837 609517 73893
rect 609603 73837 609659 73893
rect 609745 73837 609801 73893
rect 607899 73695 607955 73751
rect 608041 73695 608097 73751
rect 608183 73695 608239 73751
rect 608325 73695 608381 73751
rect 608467 73695 608523 73751
rect 609319 73695 609375 73751
rect 609461 73695 609517 73751
rect 609603 73695 609659 73751
rect 609745 73695 609801 73751
rect 607899 73553 607955 73609
rect 608041 73553 608097 73609
rect 608183 73553 608239 73609
rect 608325 73553 608381 73609
rect 608467 73553 608523 73609
rect 609319 73553 609375 73609
rect 609461 73553 609517 73609
rect 609603 73553 609659 73609
rect 609745 73553 609801 73609
rect 607899 73411 607955 73467
rect 608041 73411 608097 73467
rect 608183 73411 608239 73467
rect 608325 73411 608381 73467
rect 608467 73411 608523 73467
rect 609319 73411 609375 73467
rect 609461 73411 609517 73467
rect 609603 73411 609659 73467
rect 609745 73411 609801 73467
rect 607899 73269 607955 73325
rect 608041 73269 608097 73325
rect 608183 73269 608239 73325
rect 608325 73269 608381 73325
rect 608467 73269 608523 73325
rect 609319 73269 609375 73325
rect 609461 73269 609517 73325
rect 609603 73269 609659 73325
rect 609745 73269 609801 73325
rect 607899 73127 607955 73183
rect 608041 73127 608097 73183
rect 608183 73127 608239 73183
rect 608325 73127 608381 73183
rect 608467 73127 608523 73183
rect 609319 73127 609375 73183
rect 609461 73127 609517 73183
rect 609603 73127 609659 73183
rect 609745 73127 609801 73183
rect 607899 72985 607955 73041
rect 608041 72985 608097 73041
rect 608183 72985 608239 73041
rect 608325 72985 608381 73041
rect 608467 72985 608523 73041
rect 609319 72985 609375 73041
rect 609461 72985 609517 73041
rect 609603 72985 609659 73041
rect 609745 72985 609801 73041
rect 607899 72843 607955 72899
rect 608041 72843 608097 72899
rect 608183 72843 608239 72899
rect 608325 72843 608381 72899
rect 608467 72843 608523 72899
rect 609319 72843 609375 72899
rect 609461 72843 609517 72899
rect 609603 72843 609659 72899
rect 609745 72843 609801 72899
rect 607899 72701 607955 72757
rect 608041 72701 608097 72757
rect 608183 72701 608239 72757
rect 608325 72701 608381 72757
rect 608467 72701 608523 72757
rect 609319 72701 609375 72757
rect 609461 72701 609517 72757
rect 609603 72701 609659 72757
rect 609745 72701 609801 72757
rect 607899 72559 607955 72615
rect 608041 72559 608097 72615
rect 608183 72559 608239 72615
rect 608325 72559 608381 72615
rect 608467 72559 608523 72615
rect 609319 72559 609375 72615
rect 609461 72559 609517 72615
rect 609603 72559 609659 72615
rect 609745 72559 609801 72615
rect 607899 72417 607955 72473
rect 608041 72417 608097 72473
rect 608183 72417 608239 72473
rect 608325 72417 608381 72473
rect 608467 72417 608523 72473
rect 609319 72417 609375 72473
rect 609461 72417 609517 72473
rect 609603 72417 609659 72473
rect 609745 72417 609801 72473
rect 607899 72275 607955 72331
rect 608041 72275 608097 72331
rect 608183 72275 608239 72331
rect 608325 72275 608381 72331
rect 608467 72275 608523 72331
rect 609319 72275 609375 72331
rect 609461 72275 609517 72331
rect 609603 72275 609659 72331
rect 609745 72275 609801 72331
rect 607899 72133 607955 72189
rect 608041 72133 608097 72189
rect 608183 72133 608239 72189
rect 608325 72133 608381 72189
rect 608467 72133 608523 72189
rect 609319 72133 609375 72189
rect 609461 72133 609517 72189
rect 609603 72133 609659 72189
rect 609745 72133 609801 72189
rect 610269 73979 610325 74035
rect 610411 73979 610467 74035
rect 610553 73979 610609 74035
rect 610695 73979 610751 74035
rect 610837 73979 610893 74035
rect 610979 73979 611035 74035
rect 611121 73979 611177 74035
rect 611263 73979 611319 74035
rect 611405 73979 611461 74035
rect 611547 73979 611603 74035
rect 611689 73979 611745 74035
rect 611831 73979 611887 74035
rect 611973 73979 612029 74035
rect 612115 73979 612171 74035
rect 610269 73837 610325 73893
rect 610411 73837 610467 73893
rect 610553 73837 610609 73893
rect 610695 73837 610751 73893
rect 610837 73837 610893 73893
rect 610979 73837 611035 73893
rect 611121 73837 611177 73893
rect 611263 73837 611319 73893
rect 611405 73837 611461 73893
rect 611547 73837 611603 73893
rect 611689 73837 611745 73893
rect 611831 73837 611887 73893
rect 611973 73837 612029 73893
rect 612115 73837 612171 73893
rect 610269 73695 610325 73751
rect 610411 73695 610467 73751
rect 610553 73695 610609 73751
rect 610695 73695 610751 73751
rect 610837 73695 610893 73751
rect 610979 73695 611035 73751
rect 611121 73695 611177 73751
rect 611263 73695 611319 73751
rect 611405 73695 611461 73751
rect 611547 73695 611603 73751
rect 611689 73695 611745 73751
rect 611831 73695 611887 73751
rect 611973 73695 612029 73751
rect 612115 73695 612171 73751
rect 610269 73553 610325 73609
rect 610411 73553 610467 73609
rect 610553 73553 610609 73609
rect 610695 73553 610751 73609
rect 610837 73553 610893 73609
rect 610979 73553 611035 73609
rect 611121 73553 611177 73609
rect 611263 73553 611319 73609
rect 611405 73553 611461 73609
rect 611547 73553 611603 73609
rect 611689 73553 611745 73609
rect 611831 73553 611887 73609
rect 611973 73553 612029 73609
rect 612115 73553 612171 73609
rect 610269 73411 610325 73467
rect 610411 73411 610467 73467
rect 610553 73411 610609 73467
rect 610695 73411 610751 73467
rect 610837 73411 610893 73467
rect 610979 73411 611035 73467
rect 611121 73411 611177 73467
rect 611263 73411 611319 73467
rect 611405 73411 611461 73467
rect 611547 73411 611603 73467
rect 611689 73411 611745 73467
rect 611831 73411 611887 73467
rect 611973 73411 612029 73467
rect 612115 73411 612171 73467
rect 610269 73269 610325 73325
rect 610411 73269 610467 73325
rect 610553 73269 610609 73325
rect 610695 73269 610751 73325
rect 610837 73269 610893 73325
rect 610979 73269 611035 73325
rect 611121 73269 611177 73325
rect 611263 73269 611319 73325
rect 611405 73269 611461 73325
rect 611547 73269 611603 73325
rect 611689 73269 611745 73325
rect 611831 73269 611887 73325
rect 611973 73269 612029 73325
rect 612115 73269 612171 73325
rect 610269 73127 610325 73183
rect 610411 73127 610467 73183
rect 610553 73127 610609 73183
rect 610695 73127 610751 73183
rect 610837 73127 610893 73183
rect 610979 73127 611035 73183
rect 611121 73127 611177 73183
rect 611263 73127 611319 73183
rect 611405 73127 611461 73183
rect 611547 73127 611603 73183
rect 611689 73127 611745 73183
rect 611831 73127 611887 73183
rect 611973 73127 612029 73183
rect 612115 73127 612171 73183
rect 610269 72985 610325 73041
rect 610411 72985 610467 73041
rect 610553 72985 610609 73041
rect 610695 72985 610751 73041
rect 610837 72985 610893 73041
rect 610979 72985 611035 73041
rect 611121 72985 611177 73041
rect 611263 72985 611319 73041
rect 611405 72985 611461 73041
rect 611547 72985 611603 73041
rect 611689 72985 611745 73041
rect 611831 72985 611887 73041
rect 611973 72985 612029 73041
rect 612115 72985 612171 73041
rect 610269 72843 610325 72899
rect 610411 72843 610467 72899
rect 610553 72843 610609 72899
rect 610695 72843 610751 72899
rect 610837 72843 610893 72899
rect 610979 72843 611035 72899
rect 611121 72843 611177 72899
rect 611263 72843 611319 72899
rect 611405 72843 611461 72899
rect 611547 72843 611603 72899
rect 611689 72843 611745 72899
rect 611831 72843 611887 72899
rect 611973 72843 612029 72899
rect 612115 72843 612171 72899
rect 610269 72701 610325 72757
rect 610411 72701 610467 72757
rect 610553 72701 610609 72757
rect 610695 72701 610751 72757
rect 610837 72701 610893 72757
rect 610979 72701 611035 72757
rect 611121 72701 611177 72757
rect 611263 72701 611319 72757
rect 611405 72701 611461 72757
rect 611547 72701 611603 72757
rect 611689 72701 611745 72757
rect 611831 72701 611887 72757
rect 611973 72701 612029 72757
rect 612115 72701 612171 72757
rect 610269 72559 610325 72615
rect 610411 72559 610467 72615
rect 610553 72559 610609 72615
rect 610695 72559 610751 72615
rect 610837 72559 610893 72615
rect 610979 72559 611035 72615
rect 611121 72559 611177 72615
rect 611263 72559 611319 72615
rect 611405 72559 611461 72615
rect 611547 72559 611603 72615
rect 611689 72559 611745 72615
rect 611831 72559 611887 72615
rect 611973 72559 612029 72615
rect 612115 72559 612171 72615
rect 610269 72417 610325 72473
rect 610411 72417 610467 72473
rect 610553 72417 610609 72473
rect 610695 72417 610751 72473
rect 610837 72417 610893 72473
rect 610979 72417 611035 72473
rect 611121 72417 611177 72473
rect 611263 72417 611319 72473
rect 611405 72417 611461 72473
rect 611547 72417 611603 72473
rect 611689 72417 611745 72473
rect 611831 72417 611887 72473
rect 611973 72417 612029 72473
rect 612115 72417 612171 72473
rect 610269 72275 610325 72331
rect 610411 72275 610467 72331
rect 610553 72275 610609 72331
rect 610695 72275 610751 72331
rect 610837 72275 610893 72331
rect 610979 72275 611035 72331
rect 611121 72275 611177 72331
rect 611263 72275 611319 72331
rect 611405 72275 611461 72331
rect 611547 72275 611603 72331
rect 611689 72275 611745 72331
rect 611831 72275 611887 72331
rect 611973 72275 612029 72331
rect 612115 72275 612171 72331
rect 610269 72133 610325 72189
rect 610411 72133 610467 72189
rect 610553 72133 610609 72189
rect 610695 72133 610751 72189
rect 610837 72133 610893 72189
rect 610979 72133 611035 72189
rect 611121 72133 611177 72189
rect 611263 72133 611319 72189
rect 611405 72133 611461 72189
rect 611547 72133 611603 72189
rect 611689 72133 611745 72189
rect 611831 72133 611887 72189
rect 611973 72133 612029 72189
rect 612115 72133 612171 72189
rect 612899 73979 612955 74035
rect 613041 73979 613097 74035
rect 613183 73979 613239 74035
rect 613325 73979 613381 74035
rect 613467 73979 613523 74035
rect 613609 73979 613665 74035
rect 613751 73979 613807 74035
rect 613893 73979 613949 74035
rect 614035 73979 614091 74035
rect 614177 73979 614233 74035
rect 614319 73979 614375 74035
rect 614461 73979 614517 74035
rect 614603 73979 614659 74035
rect 612899 73837 612955 73893
rect 613041 73837 613097 73893
rect 613183 73837 613239 73893
rect 613325 73837 613381 73893
rect 613467 73837 613523 73893
rect 613609 73837 613665 73893
rect 613751 73837 613807 73893
rect 613893 73837 613949 73893
rect 614035 73837 614091 73893
rect 614177 73837 614233 73893
rect 614319 73837 614375 73893
rect 614461 73837 614517 73893
rect 614603 73837 614659 73893
rect 612899 73695 612955 73751
rect 613041 73695 613097 73751
rect 613183 73695 613239 73751
rect 613325 73695 613381 73751
rect 613467 73695 613523 73751
rect 613609 73695 613665 73751
rect 613751 73695 613807 73751
rect 613893 73695 613949 73751
rect 614035 73695 614091 73751
rect 614177 73695 614233 73751
rect 614319 73695 614375 73751
rect 614461 73695 614517 73751
rect 614603 73695 614659 73751
rect 612899 73553 612955 73609
rect 613041 73553 613097 73609
rect 613183 73553 613239 73609
rect 613325 73553 613381 73609
rect 613467 73553 613523 73609
rect 613609 73553 613665 73609
rect 613751 73553 613807 73609
rect 613893 73553 613949 73609
rect 614035 73553 614091 73609
rect 614177 73553 614233 73609
rect 614319 73553 614375 73609
rect 614461 73553 614517 73609
rect 614603 73553 614659 73609
rect 612899 73411 612955 73467
rect 613041 73411 613097 73467
rect 613183 73411 613239 73467
rect 613325 73411 613381 73467
rect 613467 73411 613523 73467
rect 613609 73411 613665 73467
rect 613751 73411 613807 73467
rect 613893 73411 613949 73467
rect 614035 73411 614091 73467
rect 614177 73411 614233 73467
rect 614319 73411 614375 73467
rect 614461 73411 614517 73467
rect 614603 73411 614659 73467
rect 612899 73269 612955 73325
rect 613041 73269 613097 73325
rect 613183 73269 613239 73325
rect 613325 73269 613381 73325
rect 613467 73269 613523 73325
rect 613609 73269 613665 73325
rect 613751 73269 613807 73325
rect 613893 73269 613949 73325
rect 614035 73269 614091 73325
rect 614177 73269 614233 73325
rect 614319 73269 614375 73325
rect 614461 73269 614517 73325
rect 614603 73269 614659 73325
rect 612899 73127 612955 73183
rect 613041 73127 613097 73183
rect 613183 73127 613239 73183
rect 613325 73127 613381 73183
rect 613467 73127 613523 73183
rect 613609 73127 613665 73183
rect 613751 73127 613807 73183
rect 613893 73127 613949 73183
rect 614035 73127 614091 73183
rect 614177 73127 614233 73183
rect 614319 73127 614375 73183
rect 614461 73127 614517 73183
rect 614603 73127 614659 73183
rect 612899 72985 612955 73041
rect 613041 72985 613097 73041
rect 613183 72985 613239 73041
rect 613325 72985 613381 73041
rect 613467 72985 613523 73041
rect 613609 72985 613665 73041
rect 613751 72985 613807 73041
rect 613893 72985 613949 73041
rect 614035 72985 614091 73041
rect 614177 72985 614233 73041
rect 614319 72985 614375 73041
rect 614461 72985 614517 73041
rect 614603 72985 614659 73041
rect 612899 72843 612955 72899
rect 613041 72843 613097 72899
rect 613183 72843 613239 72899
rect 613325 72843 613381 72899
rect 613467 72843 613523 72899
rect 613609 72843 613665 72899
rect 613751 72843 613807 72899
rect 613893 72843 613949 72899
rect 614035 72843 614091 72899
rect 614177 72843 614233 72899
rect 614319 72843 614375 72899
rect 614461 72843 614517 72899
rect 614603 72843 614659 72899
rect 612899 72701 612955 72757
rect 613041 72701 613097 72757
rect 613183 72701 613239 72757
rect 613325 72701 613381 72757
rect 613467 72701 613523 72757
rect 613609 72701 613665 72757
rect 613751 72701 613807 72757
rect 613893 72701 613949 72757
rect 614035 72701 614091 72757
rect 614177 72701 614233 72757
rect 614319 72701 614375 72757
rect 614461 72701 614517 72757
rect 614603 72701 614659 72757
rect 612899 72559 612955 72615
rect 613041 72559 613097 72615
rect 613183 72559 613239 72615
rect 613325 72559 613381 72615
rect 613467 72559 613523 72615
rect 613609 72559 613665 72615
rect 613751 72559 613807 72615
rect 613893 72559 613949 72615
rect 614035 72559 614091 72615
rect 614177 72559 614233 72615
rect 614319 72559 614375 72615
rect 614461 72559 614517 72615
rect 614603 72559 614659 72615
rect 612899 72417 612955 72473
rect 613041 72417 613097 72473
rect 613183 72417 613239 72473
rect 613325 72417 613381 72473
rect 613467 72417 613523 72473
rect 613609 72417 613665 72473
rect 613751 72417 613807 72473
rect 613893 72417 613949 72473
rect 614035 72417 614091 72473
rect 614177 72417 614233 72473
rect 614319 72417 614375 72473
rect 614461 72417 614517 72473
rect 614603 72417 614659 72473
rect 612899 72275 612955 72331
rect 613041 72275 613097 72331
rect 613183 72275 613239 72331
rect 613325 72275 613381 72331
rect 613467 72275 613523 72331
rect 613609 72275 613665 72331
rect 613751 72275 613807 72331
rect 613893 72275 613949 72331
rect 614035 72275 614091 72331
rect 614177 72275 614233 72331
rect 614319 72275 614375 72331
rect 614461 72275 614517 72331
rect 614603 72275 614659 72331
rect 612899 72133 612955 72189
rect 613041 72133 613097 72189
rect 613183 72133 613239 72189
rect 613325 72133 613381 72189
rect 613467 72133 613523 72189
rect 613609 72133 613665 72189
rect 613751 72133 613807 72189
rect 613893 72133 613949 72189
rect 614035 72133 614091 72189
rect 614177 72133 614233 72189
rect 614319 72133 614375 72189
rect 614461 72133 614517 72189
rect 614603 72133 614659 72189
<< properties >>
string FIXED_BBOX 0 0 3880 5070
<< end >>
