magic
tech gf180mcuC
magscale 1 10
timestamp 1654780538
<< metal1 >>
rect 3882 12854 3894 12906
rect 3946 12903 3958 12906
rect 7242 12903 7254 12906
rect 3946 12857 7254 12903
rect 3946 12854 3958 12857
rect 7242 12854 7254 12857
rect 7306 12854 7318 12906
rect 1120 11786 13776 11820
rect 1120 11734 2585 11786
rect 2637 11734 2689 11786
rect 2741 11734 2793 11786
rect 2845 11734 5775 11786
rect 5827 11734 5879 11786
rect 5931 11734 5983 11786
rect 6035 11734 8965 11786
rect 9017 11734 9069 11786
rect 9121 11734 9173 11786
rect 9225 11734 12155 11786
rect 12207 11734 12259 11786
rect 12311 11734 12363 11786
rect 12415 11734 13776 11786
rect 1120 11700 13776 11734
rect 13850 11622 13862 11674
rect 13914 11671 13926 11674
rect 14746 11671 14758 11674
rect 13914 11625 14758 11671
rect 13914 11622 13926 11625
rect 14746 11622 14758 11625
rect 14810 11622 14822 11674
rect 7982 11282 8034 11294
rect 7982 11218 8034 11230
rect 12350 11170 12402 11182
rect 12350 11106 12402 11118
rect 1120 11002 13776 11036
rect 1120 10950 4180 11002
rect 4232 10950 4284 11002
rect 4336 10950 4388 11002
rect 4440 10950 7370 11002
rect 7422 10950 7474 11002
rect 7526 10950 7578 11002
rect 7630 10950 10560 11002
rect 10612 10950 10664 11002
rect 10716 10950 10768 11002
rect 10820 10950 13776 11002
rect 1120 10916 13776 10950
rect 3166 10834 3218 10846
rect 3166 10770 3218 10782
rect 11230 10722 11282 10734
rect 1766 10666 1818 10678
rect 2426 10670 2438 10722
rect 2490 10670 2502 10722
rect 1766 10602 1818 10614
rect 7982 10666 8034 10678
rect 11230 10658 11282 10670
rect 11946 10660 11958 10712
rect 12010 10660 12022 10712
rect 12294 10666 12346 10678
rect 2314 10558 2326 10610
rect 2378 10558 2390 10610
rect 7410 10558 7422 10610
rect 7474 10558 7486 10610
rect 7982 10602 8034 10614
rect 8138 10552 8150 10604
rect 8202 10552 8214 10604
rect 12294 10602 12346 10614
rect 12686 10610 12738 10622
rect 12686 10546 12738 10558
rect 7130 10440 7142 10492
rect 7194 10440 7206 10492
rect 13022 10442 13074 10454
rect 13850 10390 13862 10442
rect 13914 10439 13926 10442
rect 14746 10439 14758 10442
rect 13914 10393 14758 10439
rect 13914 10390 13926 10393
rect 14746 10390 14758 10393
rect 14810 10390 14822 10442
rect 13022 10378 13074 10390
rect 1120 10218 13776 10252
rect 1120 10166 2585 10218
rect 2637 10166 2689 10218
rect 2741 10166 2793 10218
rect 2845 10166 5775 10218
rect 5827 10166 5879 10218
rect 5931 10166 5983 10218
rect 6035 10166 8965 10218
rect 9017 10166 9069 10218
rect 9121 10166 9173 10218
rect 9225 10166 12155 10218
rect 12207 10166 12259 10218
rect 12311 10166 12363 10218
rect 12415 10166 13776 10218
rect 1120 10132 13776 10166
rect 2158 10050 2210 10062
rect 2158 9986 2210 9998
rect 7982 9714 8034 9726
rect 7982 9650 8034 9662
rect 12126 9714 12178 9726
rect 12126 9650 12178 9662
rect 1120 9434 13776 9468
rect 1120 9382 4180 9434
rect 4232 9382 4284 9434
rect 4336 9382 4388 9434
rect 4440 9382 7370 9434
rect 7422 9382 7474 9434
rect 7526 9382 7578 9434
rect 7630 9382 10560 9434
rect 10612 9382 10664 9434
rect 10716 9382 10768 9434
rect 10820 9382 13776 9434
rect 1120 9348 13776 9382
rect 2830 9266 2882 9278
rect 2830 9202 2882 9214
rect 7086 9266 7138 9278
rect 7086 9202 7138 9214
rect 2158 8874 2210 8886
rect 2158 8810 2210 8822
rect 1120 8650 13776 8684
rect 1120 8598 2585 8650
rect 2637 8598 2689 8650
rect 2741 8598 2793 8650
rect 2845 8598 5775 8650
rect 5827 8598 5879 8650
rect 5931 8598 5983 8650
rect 6035 8598 8965 8650
rect 9017 8598 9069 8650
rect 9121 8598 9173 8650
rect 9225 8598 12155 8650
rect 12207 8598 12259 8650
rect 12311 8598 12363 8650
rect 12415 8598 13776 8650
rect 1120 8564 13776 8598
rect 8094 8426 8146 8438
rect 8094 8362 8146 8374
rect 7758 8258 7810 8270
rect 7366 8202 7418 8214
rect 7758 8194 7810 8206
rect 7130 8090 7142 8142
rect 7194 8090 7206 8142
rect 7366 8138 7418 8150
rect 8878 8090 8930 8102
rect 8878 8026 8930 8038
rect 11342 8034 11394 8046
rect 11342 7970 11394 7982
rect 1120 7866 13776 7900
rect 1120 7814 4180 7866
rect 4232 7814 4284 7866
rect 4336 7814 4388 7866
rect 4440 7814 7370 7866
rect 7422 7814 7474 7866
rect 7526 7814 7578 7866
rect 7630 7814 10560 7866
rect 10612 7814 10664 7866
rect 10716 7814 10768 7866
rect 10820 7814 13776 7866
rect 1120 7780 13776 7814
rect 6526 7642 6578 7654
rect 5854 7586 5906 7598
rect 6526 7578 6578 7590
rect 7758 7586 7810 7598
rect 5854 7522 5906 7534
rect 7758 7522 7810 7534
rect 9550 7586 9602 7598
rect 9550 7522 9602 7534
rect 10378 7422 10390 7474
rect 10442 7422 10454 7474
rect 10826 7422 10838 7474
rect 10890 7422 10902 7474
rect 10938 7254 10950 7306
rect 11002 7254 11014 7306
rect 1120 7082 13776 7116
rect 1120 7030 2585 7082
rect 2637 7030 2689 7082
rect 2741 7030 2793 7082
rect 2845 7030 5775 7082
rect 5827 7030 5879 7082
rect 5931 7030 5983 7082
rect 6035 7030 8965 7082
rect 9017 7030 9069 7082
rect 9121 7030 9173 7082
rect 9225 7030 12155 7082
rect 12207 7030 12259 7082
rect 12311 7030 12363 7082
rect 12415 7030 13776 7082
rect 1120 6996 13776 7030
rect 6570 6638 6582 6690
rect 6634 6638 6646 6690
rect 8822 6522 8874 6534
rect 8822 6458 8874 6470
rect 1120 6298 13776 6332
rect 1120 6246 4180 6298
rect 4232 6246 4284 6298
rect 4336 6246 4388 6298
rect 4440 6246 7370 6298
rect 7422 6246 7474 6298
rect 7526 6246 7578 6298
rect 7630 6246 10560 6298
rect 10612 6246 10664 6298
rect 10716 6246 10768 6298
rect 10820 6246 13776 6298
rect 1120 6212 13776 6246
rect 6862 5850 6914 5862
rect 7186 5854 7198 5906
rect 7250 5854 7262 5906
rect 6862 5786 6914 5798
rect 1120 5514 13776 5548
rect 1120 5462 2585 5514
rect 2637 5462 2689 5514
rect 2741 5462 2793 5514
rect 2845 5462 5775 5514
rect 5827 5462 5879 5514
rect 5931 5462 5983 5514
rect 6035 5462 8965 5514
rect 9017 5462 9069 5514
rect 9121 5462 9173 5514
rect 9225 5462 12155 5514
rect 12207 5462 12259 5514
rect 12311 5462 12363 5514
rect 12415 5462 13776 5514
rect 1120 5428 13776 5462
rect 3278 5010 3330 5022
rect 3278 4946 3330 4958
rect 1120 4730 13776 4764
rect 1120 4678 4180 4730
rect 4232 4678 4284 4730
rect 4336 4678 4388 4730
rect 4440 4678 7370 4730
rect 7422 4678 7474 4730
rect 7526 4678 7578 4730
rect 7630 4678 10560 4730
rect 10612 4678 10664 4730
rect 10716 4678 10768 4730
rect 10820 4678 13776 4730
rect 1120 4644 13776 4678
rect 2158 4562 2210 4574
rect 2158 4498 2210 4510
rect 10670 4506 10722 4518
rect 10670 4442 10722 4454
rect 12686 4226 12738 4238
rect 12686 4162 12738 4174
rect 1120 3946 13776 3980
rect 1120 3894 2585 3946
rect 2637 3894 2689 3946
rect 2741 3894 2793 3946
rect 2845 3894 5775 3946
rect 5827 3894 5879 3946
rect 5931 3894 5983 3946
rect 6035 3894 8965 3946
rect 9017 3894 9069 3946
rect 9121 3894 9173 3946
rect 9225 3894 12155 3946
rect 12207 3894 12259 3946
rect 12311 3894 12363 3946
rect 12415 3894 13776 3946
rect 1120 3860 13776 3894
rect 11958 3722 12010 3734
rect 2538 3614 2550 3666
rect 2602 3614 2614 3666
rect 11958 3658 12010 3670
rect 2874 3502 2886 3554
rect 2938 3502 2950 3554
rect 7802 3490 7814 3542
rect 7866 3490 7878 3542
rect 8418 3502 8430 3554
rect 8482 3502 8494 3554
rect 10714 3514 10726 3566
rect 10778 3514 10790 3566
rect 11162 3493 11174 3545
rect 11226 3493 11238 3545
rect 2438 3386 2490 3398
rect 2438 3322 2490 3334
rect 6078 3386 6130 3398
rect 6078 3322 6130 3334
rect 7310 3386 7362 3398
rect 7310 3322 7362 3334
rect 1120 3162 13776 3196
rect 1120 3110 4180 3162
rect 4232 3110 4284 3162
rect 4336 3110 4388 3162
rect 4440 3110 7370 3162
rect 7422 3110 7474 3162
rect 7526 3110 7578 3162
rect 7630 3110 10560 3162
rect 10612 3110 10664 3162
rect 10716 3110 10768 3162
rect 10820 3110 13776 3162
rect 1120 3076 13776 3110
rect 9438 2994 9490 3006
rect 9438 2930 9490 2942
rect 6974 2882 7026 2894
rect 10222 2882 10274 2894
rect 8250 2830 8262 2882
rect 8314 2830 8326 2882
rect 6974 2818 7026 2830
rect 10222 2818 10274 2830
rect 1922 2718 1934 2770
rect 1986 2718 1998 2770
rect 2258 2718 2270 2770
rect 2322 2718 2334 2770
rect 4778 2706 4790 2758
rect 4842 2706 4854 2758
rect 5226 2727 5238 2779
rect 5290 2727 5302 2779
rect 7914 2718 7926 2770
rect 7978 2718 7990 2770
rect 5910 2602 5962 2614
rect 7802 2550 7814 2602
rect 7866 2550 7878 2602
rect 5910 2538 5962 2550
rect 1120 2378 13776 2412
rect 1120 2326 2585 2378
rect 2637 2326 2689 2378
rect 2741 2326 2793 2378
rect 2845 2326 5775 2378
rect 5827 2326 5879 2378
rect 5931 2326 5983 2378
rect 6035 2326 8965 2378
rect 9017 2326 9069 2378
rect 9121 2326 9173 2378
rect 9225 2326 12155 2378
rect 12207 2326 12259 2378
rect 12311 2326 12363 2378
rect 12415 2326 13776 2378
rect 1120 2292 13776 2326
rect 3950 2098 4002 2110
rect 3950 2034 4002 2046
rect 7690 1909 7702 1961
rect 7754 1909 7766 1961
rect 2718 1874 2770 1886
rect 2718 1810 2770 1822
rect 5518 1874 5570 1886
rect 9326 1874 9378 1886
rect 5518 1810 5570 1822
rect 7914 1811 7926 1863
rect 7978 1811 7990 1863
rect 9326 1810 9378 1822
rect 2046 1762 2098 1774
rect 2046 1698 2098 1710
rect 6190 1762 6242 1774
rect 6190 1698 6242 1710
rect 1120 1594 13776 1628
rect 1120 1542 4180 1594
rect 4232 1542 4284 1594
rect 4336 1542 4388 1594
rect 4440 1542 7370 1594
rect 7422 1542 7474 1594
rect 7526 1542 7578 1594
rect 7630 1542 10560 1594
rect 10612 1542 10664 1594
rect 10716 1542 10768 1594
rect 10820 1542 13776 1594
rect 1120 1508 13776 1542
rect 4666 1318 4678 1370
rect 4730 1367 4742 1370
rect 6178 1367 6190 1370
rect 4730 1321 6190 1367
rect 4730 1318 4742 1321
rect 6178 1318 6190 1321
rect 6242 1318 6254 1370
<< via1 >>
rect 3894 12854 3946 12906
rect 7254 12854 7306 12906
rect 2585 11734 2637 11786
rect 2689 11734 2741 11786
rect 2793 11734 2845 11786
rect 5775 11734 5827 11786
rect 5879 11734 5931 11786
rect 5983 11734 6035 11786
rect 8965 11734 9017 11786
rect 9069 11734 9121 11786
rect 9173 11734 9225 11786
rect 12155 11734 12207 11786
rect 12259 11734 12311 11786
rect 12363 11734 12415 11786
rect 13862 11622 13914 11674
rect 14758 11622 14810 11674
rect 7982 11230 8034 11282
rect 12350 11118 12402 11170
rect 4180 10950 4232 11002
rect 4284 10950 4336 11002
rect 4388 10950 4440 11002
rect 7370 10950 7422 11002
rect 7474 10950 7526 11002
rect 7578 10950 7630 11002
rect 10560 10950 10612 11002
rect 10664 10950 10716 11002
rect 10768 10950 10820 11002
rect 3166 10782 3218 10834
rect 2438 10670 2490 10722
rect 1766 10614 1818 10666
rect 7982 10614 8034 10666
rect 11230 10670 11282 10722
rect 11958 10660 12010 10712
rect 2326 10558 2378 10610
rect 7422 10558 7474 10610
rect 12294 10614 12346 10666
rect 8150 10552 8202 10604
rect 12686 10558 12738 10610
rect 7142 10440 7194 10492
rect 13022 10390 13074 10442
rect 13862 10390 13914 10442
rect 14758 10390 14810 10442
rect 2585 10166 2637 10218
rect 2689 10166 2741 10218
rect 2793 10166 2845 10218
rect 5775 10166 5827 10218
rect 5879 10166 5931 10218
rect 5983 10166 6035 10218
rect 8965 10166 9017 10218
rect 9069 10166 9121 10218
rect 9173 10166 9225 10218
rect 12155 10166 12207 10218
rect 12259 10166 12311 10218
rect 12363 10166 12415 10218
rect 2158 9998 2210 10050
rect 7982 9662 8034 9714
rect 12126 9662 12178 9714
rect 4180 9382 4232 9434
rect 4284 9382 4336 9434
rect 4388 9382 4440 9434
rect 7370 9382 7422 9434
rect 7474 9382 7526 9434
rect 7578 9382 7630 9434
rect 10560 9382 10612 9434
rect 10664 9382 10716 9434
rect 10768 9382 10820 9434
rect 2830 9214 2882 9266
rect 7086 9214 7138 9266
rect 2158 8822 2210 8874
rect 2585 8598 2637 8650
rect 2689 8598 2741 8650
rect 2793 8598 2845 8650
rect 5775 8598 5827 8650
rect 5879 8598 5931 8650
rect 5983 8598 6035 8650
rect 8965 8598 9017 8650
rect 9069 8598 9121 8650
rect 9173 8598 9225 8650
rect 12155 8598 12207 8650
rect 12259 8598 12311 8650
rect 12363 8598 12415 8650
rect 8094 8374 8146 8426
rect 7366 8150 7418 8202
rect 7758 8206 7810 8258
rect 7142 8090 7194 8142
rect 8878 8038 8930 8090
rect 11342 7982 11394 8034
rect 4180 7814 4232 7866
rect 4284 7814 4336 7866
rect 4388 7814 4440 7866
rect 7370 7814 7422 7866
rect 7474 7814 7526 7866
rect 7578 7814 7630 7866
rect 10560 7814 10612 7866
rect 10664 7814 10716 7866
rect 10768 7814 10820 7866
rect 5854 7534 5906 7586
rect 6526 7590 6578 7642
rect 7758 7534 7810 7586
rect 9550 7534 9602 7586
rect 10390 7422 10442 7474
rect 10838 7422 10890 7474
rect 10950 7254 11002 7306
rect 2585 7030 2637 7082
rect 2689 7030 2741 7082
rect 2793 7030 2845 7082
rect 5775 7030 5827 7082
rect 5879 7030 5931 7082
rect 5983 7030 6035 7082
rect 8965 7030 9017 7082
rect 9069 7030 9121 7082
rect 9173 7030 9225 7082
rect 12155 7030 12207 7082
rect 12259 7030 12311 7082
rect 12363 7030 12415 7082
rect 6582 6638 6634 6690
rect 8822 6470 8874 6522
rect 4180 6246 4232 6298
rect 4284 6246 4336 6298
rect 4388 6246 4440 6298
rect 7370 6246 7422 6298
rect 7474 6246 7526 6298
rect 7578 6246 7630 6298
rect 10560 6246 10612 6298
rect 10664 6246 10716 6298
rect 10768 6246 10820 6298
rect 7198 5854 7250 5906
rect 6862 5798 6914 5850
rect 2585 5462 2637 5514
rect 2689 5462 2741 5514
rect 2793 5462 2845 5514
rect 5775 5462 5827 5514
rect 5879 5462 5931 5514
rect 5983 5462 6035 5514
rect 8965 5462 9017 5514
rect 9069 5462 9121 5514
rect 9173 5462 9225 5514
rect 12155 5462 12207 5514
rect 12259 5462 12311 5514
rect 12363 5462 12415 5514
rect 3278 4958 3330 5010
rect 4180 4678 4232 4730
rect 4284 4678 4336 4730
rect 4388 4678 4440 4730
rect 7370 4678 7422 4730
rect 7474 4678 7526 4730
rect 7578 4678 7630 4730
rect 10560 4678 10612 4730
rect 10664 4678 10716 4730
rect 10768 4678 10820 4730
rect 2158 4510 2210 4562
rect 10670 4454 10722 4506
rect 12686 4174 12738 4226
rect 2585 3894 2637 3946
rect 2689 3894 2741 3946
rect 2793 3894 2845 3946
rect 5775 3894 5827 3946
rect 5879 3894 5931 3946
rect 5983 3894 6035 3946
rect 8965 3894 9017 3946
rect 9069 3894 9121 3946
rect 9173 3894 9225 3946
rect 12155 3894 12207 3946
rect 12259 3894 12311 3946
rect 12363 3894 12415 3946
rect 11958 3670 12010 3722
rect 2550 3614 2602 3666
rect 2886 3502 2938 3554
rect 7814 3490 7866 3542
rect 8430 3502 8482 3554
rect 10726 3514 10778 3566
rect 11174 3493 11226 3545
rect 2438 3334 2490 3386
rect 6078 3334 6130 3386
rect 7310 3334 7362 3386
rect 4180 3110 4232 3162
rect 4284 3110 4336 3162
rect 4388 3110 4440 3162
rect 7370 3110 7422 3162
rect 7474 3110 7526 3162
rect 7578 3110 7630 3162
rect 10560 3110 10612 3162
rect 10664 3110 10716 3162
rect 10768 3110 10820 3162
rect 9438 2942 9490 2994
rect 6974 2830 7026 2882
rect 8262 2830 8314 2882
rect 10222 2830 10274 2882
rect 1934 2718 1986 2770
rect 2270 2718 2322 2770
rect 4790 2706 4842 2758
rect 5238 2727 5290 2779
rect 7926 2718 7978 2770
rect 5910 2550 5962 2602
rect 7814 2550 7866 2602
rect 2585 2326 2637 2378
rect 2689 2326 2741 2378
rect 2793 2326 2845 2378
rect 5775 2326 5827 2378
rect 5879 2326 5931 2378
rect 5983 2326 6035 2378
rect 8965 2326 9017 2378
rect 9069 2326 9121 2378
rect 9173 2326 9225 2378
rect 12155 2326 12207 2378
rect 12259 2326 12311 2378
rect 12363 2326 12415 2378
rect 3950 2046 4002 2098
rect 7702 1909 7754 1961
rect 2718 1822 2770 1874
rect 5518 1822 5570 1874
rect 7926 1811 7978 1863
rect 9326 1822 9378 1874
rect 2046 1710 2098 1762
rect 6190 1710 6242 1762
rect 4180 1542 4232 1594
rect 4284 1542 4336 1594
rect 4388 1542 4440 1594
rect 7370 1542 7422 1594
rect 7474 1542 7526 1594
rect 7578 1542 7630 1594
rect 10560 1542 10612 1594
rect 10664 1542 10716 1594
rect 10768 1542 10820 1594
rect 4678 1318 4730 1370
rect 6190 1318 6242 1370
<< metal2 >>
rect -56 13200 56 14000
rect 1288 13200 1400 14000
rect 2632 13200 2744 14000
rect 2884 13300 3388 13356
rect -28 12796 28 13200
rect -28 12740 140 12796
rect 84 10892 140 12740
rect 84 10826 140 10836
rect 1316 8428 1372 13200
rect 2660 13132 2716 13200
rect 2884 13132 2940 13300
rect 2660 13076 2940 13132
rect 2583 11788 2847 11798
rect 2639 11732 2687 11788
rect 2743 11732 2791 11788
rect 2583 11722 2847 11732
rect 2100 11564 2156 11574
rect 1764 10892 1820 10902
rect 1764 10666 1820 10836
rect 1764 10614 1766 10666
rect 1818 10614 1820 10666
rect 1764 10602 1820 10614
rect 2100 10556 2156 11508
rect 2436 10892 2492 10902
rect 2436 10722 2492 10836
rect 3164 10892 3220 10902
rect 3164 10834 3220 10836
rect 3164 10782 3166 10834
rect 3218 10782 3220 10834
rect 3164 10770 3220 10782
rect 2436 10670 2438 10722
rect 2490 10670 2492 10722
rect 2436 10658 2492 10670
rect 2324 10610 2380 10622
rect 2324 10558 2326 10610
rect 2378 10558 2380 10610
rect 2100 10500 2212 10556
rect 2156 10050 2212 10500
rect 2156 9998 2158 10050
rect 2210 9998 2212 10050
rect 2156 9986 2212 9998
rect 2324 9436 2380 10558
rect 2583 10220 2847 10230
rect 2639 10164 2687 10220
rect 2743 10164 2791 10220
rect 2583 10154 2847 10164
rect 2324 9380 2884 9436
rect 2828 9266 2884 9380
rect 2828 9214 2830 9266
rect 2882 9214 2884 9266
rect 3332 9324 3388 13300
rect 3976 13200 4088 14000
rect 5320 13200 5432 14000
rect 6664 13200 6776 14000
rect 8008 13200 8120 14000
rect 8484 13300 9212 13356
rect 3892 12908 3948 12918
rect 3892 12814 3948 12852
rect 3332 9258 3388 9268
rect 2828 9212 2884 9214
rect 2828 9156 3052 9212
rect 2156 8876 2212 8886
rect 2156 8782 2212 8820
rect 2583 8652 2847 8662
rect 2639 8596 2687 8652
rect 2743 8596 2791 8652
rect 2583 8586 2847 8596
rect 1316 8372 2156 8428
rect 2100 5068 2156 8372
rect 2583 7084 2847 7094
rect 2639 7028 2687 7084
rect 2743 7028 2791 7084
rect 2583 7018 2847 7028
rect 2996 6188 3052 9156
rect 4004 8540 4060 13200
rect 4178 11004 4442 11014
rect 4234 10948 4282 11004
rect 4338 10948 4386 11004
rect 4178 10938 4442 10948
rect 5348 10892 5404 13200
rect 5773 11788 6037 11798
rect 5829 11732 5877 11788
rect 5933 11732 5981 11788
rect 5773 11722 6037 11732
rect 5348 10826 5404 10836
rect 6692 10668 6748 13200
rect 6692 10602 6748 10612
rect 7252 12906 7308 12918
rect 7252 12854 7254 12906
rect 7306 12854 7308 12906
rect 7140 10492 7196 10504
rect 7140 10440 7142 10492
rect 7194 10440 7196 10492
rect 7140 10332 7196 10440
rect 7140 10266 7196 10276
rect 5773 10220 6037 10230
rect 5829 10164 5877 10220
rect 5933 10164 5981 10220
rect 5773 10154 6037 10164
rect 7252 9548 7308 12854
rect 8036 11788 8092 13200
rect 8036 11732 8204 11788
rect 7980 11564 8036 11574
rect 7980 11282 8036 11508
rect 7980 11230 7982 11282
rect 8034 11230 8036 11282
rect 7980 11228 8036 11230
rect 7700 11172 8036 11228
rect 7368 11004 7632 11014
rect 7424 10948 7472 11004
rect 7528 10948 7576 11004
rect 7368 10938 7632 10948
rect 7700 10780 7756 11172
rect 8148 10892 8204 11732
rect 7476 10724 7756 10780
rect 7812 10836 8204 10892
rect 7476 10668 7532 10724
rect 7420 10612 7532 10668
rect 7420 10610 7476 10612
rect 7420 10558 7422 10610
rect 7474 10558 7476 10610
rect 7420 10546 7476 10558
rect 7252 9482 7308 9492
rect 4178 9436 4442 9446
rect 4234 9380 4282 9436
rect 4338 9380 4386 9436
rect 4178 9370 4442 9380
rect 7368 9436 7632 9446
rect 7424 9380 7472 9436
rect 7528 9380 7576 9436
rect 7368 9370 7632 9380
rect 7084 9324 7140 9334
rect 7084 9266 7140 9268
rect 7084 9214 7086 9266
rect 7138 9214 7140 9266
rect 7084 9212 7140 9214
rect 7812 9212 7868 10836
rect 7924 10668 8036 10678
rect 7980 10666 8036 10668
rect 7980 10614 7982 10666
rect 8034 10614 8036 10666
rect 7980 10612 8036 10614
rect 7924 10602 8036 10612
rect 8148 10604 8204 10616
rect 8148 10552 8150 10604
rect 8202 10552 8204 10604
rect 8148 10108 8204 10552
rect 8372 10332 8428 10342
rect 7980 10052 8148 10108
rect 7980 9714 8036 10052
rect 8148 9976 8204 10052
rect 8260 10276 8372 10332
rect 7980 9662 7982 9714
rect 8034 9662 8036 9714
rect 7980 9650 8036 9662
rect 7084 9156 7420 9212
rect 5773 8652 6037 8662
rect 5829 8596 5877 8652
rect 5933 8596 5981 8652
rect 5773 8586 6037 8596
rect 4004 8474 4060 8484
rect 5796 8316 5852 8326
rect 5796 8204 5852 8260
rect 6580 8316 6636 8326
rect 5796 8148 5908 8204
rect 4178 7868 4442 7878
rect 4234 7812 4282 7868
rect 4338 7812 4386 7868
rect 4178 7802 4442 7812
rect 5012 7644 5068 7654
rect 4178 6300 4442 6310
rect 4234 6244 4282 6300
rect 4338 6244 4386 6300
rect 4178 6234 4442 6244
rect 2996 6122 3052 6132
rect 2583 5516 2847 5526
rect 2639 5460 2687 5516
rect 2743 5460 2791 5516
rect 2583 5450 2847 5460
rect 3276 5068 3332 5078
rect 2100 5012 2212 5068
rect 2156 4562 2212 5012
rect 3276 5010 3332 5012
rect 3276 4958 3278 5010
rect 3330 4958 3332 5010
rect 3276 4956 3332 4958
rect 2156 4510 2158 4562
rect 2210 4510 2212 4562
rect 2156 3836 2212 4510
rect 2996 4900 3332 4956
rect 2583 3948 2847 3958
rect 2639 3892 2687 3948
rect 2743 3892 2791 3948
rect 2583 3882 2847 3892
rect 1988 3780 2212 3836
rect 1988 2828 2044 3780
rect 2548 3666 2604 3678
rect 2548 3614 2550 3666
rect 2602 3614 2604 3666
rect 2436 3388 2492 3398
rect 2436 3294 2492 3332
rect 1932 2772 2044 2828
rect 1932 2770 1988 2772
rect 1932 2718 1934 2770
rect 1986 2718 1988 2770
rect 1932 2706 1988 2718
rect 2268 2770 2324 2782
rect 2268 2718 2270 2770
rect 2322 2718 2324 2770
rect 2268 2716 2324 2718
rect 2212 2660 2324 2716
rect 2212 2380 2268 2660
rect 2548 2604 2604 3614
rect 2884 3556 2940 3566
rect 2996 3556 3052 4900
rect 4178 4732 4442 4742
rect 4234 4676 4282 4732
rect 4338 4676 4386 4732
rect 4178 4666 4442 4676
rect 2884 3554 3052 3556
rect 2884 3502 2886 3554
rect 2938 3502 3052 3554
rect 2884 3500 3052 3502
rect 2884 3490 2940 3500
rect 4178 3164 4442 3174
rect 4234 3108 4282 3164
rect 4338 3108 4386 3164
rect 4178 3098 4442 3108
rect 2044 2324 2268 2380
rect 2436 2548 2604 2604
rect 4788 2758 4844 2770
rect 4788 2706 4790 2758
rect 4842 2706 4844 2758
rect 2044 1762 2100 2324
rect 2436 1932 2492 2548
rect 2583 2380 2847 2390
rect 2639 2324 2687 2380
rect 2743 2324 2791 2380
rect 2583 2314 2847 2324
rect 4788 2156 4844 2706
rect 5012 2268 5068 7588
rect 5852 7586 5908 8148
rect 6580 7654 6636 8260
rect 7364 8202 7420 9156
rect 7140 8142 7196 8154
rect 7140 8092 7142 8142
rect 7194 8092 7196 8142
rect 7364 8150 7366 8202
rect 7418 8150 7420 8202
rect 7364 8138 7420 8150
rect 7588 9156 7868 9212
rect 7924 9548 7980 9558
rect 7588 8092 7644 9156
rect 7700 8316 7756 8326
rect 7756 8260 7812 8316
rect 7700 8258 7812 8260
rect 7700 8250 7758 8258
rect 7756 8206 7758 8250
rect 7810 8206 7812 8258
rect 7756 8194 7812 8206
rect 7588 8036 7812 8092
rect 7140 8026 7196 8036
rect 7368 7868 7632 7878
rect 7424 7812 7472 7868
rect 7528 7812 7576 7868
rect 7368 7802 7632 7812
rect 5852 7534 5854 7586
rect 5906 7534 5908 7586
rect 6524 7644 6636 7654
rect 6580 7588 6636 7644
rect 6524 7550 6580 7588
rect 7756 7586 7812 8036
rect 5852 7420 5908 7534
rect 7756 7534 7758 7586
rect 7810 7534 7812 7586
rect 5852 7364 6636 7420
rect 5773 7084 6037 7094
rect 5829 7028 5877 7084
rect 5933 7028 5981 7084
rect 5773 7018 6037 7028
rect 6580 6690 6636 7364
rect 7756 7308 7812 7534
rect 6580 6638 6582 6690
rect 6634 6638 6636 6690
rect 6580 6626 6636 6638
rect 7700 7252 7812 7308
rect 7368 6300 7632 6310
rect 7424 6244 7472 6300
rect 7528 6244 7576 6300
rect 7368 6234 7632 6244
rect 7700 5964 7756 7252
rect 7196 5908 7756 5964
rect 7196 5906 7252 5908
rect 6860 5852 6916 5862
rect 6692 5850 6916 5852
rect 6692 5798 6862 5850
rect 6914 5798 6916 5850
rect 7196 5854 7198 5906
rect 7250 5854 7252 5906
rect 7196 5842 7252 5854
rect 6692 5796 6916 5798
rect 5773 5516 6037 5526
rect 5829 5460 5877 5516
rect 5933 5460 5981 5516
rect 5773 5450 6037 5460
rect 5572 4844 5628 4854
rect 5236 3388 5292 3398
rect 5236 2779 5292 3332
rect 5236 2727 5238 2779
rect 5290 2727 5292 2779
rect 5236 2715 5292 2727
rect 5572 2604 5628 4788
rect 5773 3948 6037 3958
rect 5829 3892 5877 3948
rect 5933 3892 5981 3948
rect 5773 3882 6037 3892
rect 6244 3500 6300 3510
rect 6076 3388 6132 3398
rect 6076 3294 6132 3332
rect 5908 2604 5964 2614
rect 5572 2602 5964 2604
rect 5572 2550 5910 2602
rect 5962 2550 5964 2602
rect 5572 2548 5964 2550
rect 5908 2538 5964 2548
rect 5773 2380 6037 2390
rect 6244 2380 6300 3444
rect 5829 2324 5877 2380
rect 5933 2324 5981 2380
rect 5773 2314 6037 2324
rect 6188 2324 6300 2380
rect 5012 2202 5068 2212
rect 3948 2098 4004 2110
rect 3948 2046 3950 2098
rect 4002 2046 4004 2098
rect 4788 2090 4844 2100
rect 5516 2156 5572 2166
rect 2436 1876 2772 1932
rect 2044 1710 2046 1762
rect 2098 1710 2100 1762
rect 2044 1708 2100 1710
rect 1652 1652 2100 1708
rect 2660 1874 2772 1876
rect 2660 1822 2718 1874
rect 2770 1822 2772 1874
rect 2660 1810 2772 1822
rect 1652 1484 1708 1652
rect 1092 1428 1708 1484
rect 0 28 800 56
rect 1092 28 1148 1428
rect 1316 1260 1372 1270
rect 1316 800 1372 1204
rect 2660 800 2716 1810
rect 3948 1484 4004 2046
rect 5516 1874 5572 2100
rect 5516 1822 5518 1874
rect 5570 1822 5572 1874
rect 5516 1810 5572 1822
rect 6188 1762 6244 2324
rect 6692 2044 6748 5796
rect 6860 5786 6916 5796
rect 7368 4732 7632 4742
rect 7424 4676 7472 4732
rect 7528 4676 7576 4732
rect 7368 4666 7632 4676
rect 7924 4060 7980 9492
rect 8092 8428 8148 8438
rect 8260 8428 8316 10276
rect 8372 10266 8428 10276
rect 8092 8426 8316 8428
rect 8092 8374 8094 8426
rect 8146 8374 8316 8426
rect 8092 8372 8316 8374
rect 8092 8362 8148 8372
rect 8484 8204 8540 13300
rect 9156 13132 9212 13300
rect 9352 13200 9464 14000
rect 10696 13200 10808 14000
rect 12040 13200 12152 14000
rect 13384 13200 13496 14000
rect 14728 13200 14840 14000
rect 9380 13132 9436 13200
rect 9156 13076 9436 13132
rect 8963 11788 9227 11798
rect 9019 11732 9067 11788
rect 9123 11732 9171 11788
rect 8963 11722 9227 11732
rect 9716 11452 9772 11462
rect 8963 10220 9227 10230
rect 9019 10164 9067 10220
rect 9123 10164 9171 10220
rect 8963 10154 9227 10164
rect 9716 10108 9772 11396
rect 10724 11228 10780 13200
rect 12068 13020 12124 13200
rect 12404 13076 12684 13132
rect 12404 13020 12460 13076
rect 12068 12964 12460 13020
rect 12516 12908 12572 12918
rect 12153 11788 12417 11798
rect 12209 11732 12257 11788
rect 12313 11732 12361 11788
rect 12153 11722 12417 11732
rect 9716 10042 9772 10052
rect 10388 11172 10780 11228
rect 8963 8652 9227 8662
rect 9019 8596 9067 8652
rect 9123 8596 9171 8652
rect 8963 8586 9227 8596
rect 8484 8138 8540 8148
rect 9380 8540 9436 8550
rect 8876 8092 8932 8102
rect 8876 7998 8932 8036
rect 8963 7084 9227 7094
rect 9019 7028 9067 7084
rect 9123 7028 9171 7084
rect 8963 7018 9227 7028
rect 8820 6524 8876 6534
rect 8820 6430 8876 6468
rect 8963 5516 9227 5526
rect 9019 5460 9067 5516
rect 9123 5460 9171 5516
rect 8963 5450 9227 5460
rect 7308 4004 7980 4060
rect 7308 3386 7364 4004
rect 7812 3542 7868 3554
rect 7812 3500 7814 3542
rect 7866 3500 7868 3542
rect 7812 3434 7868 3444
rect 7308 3334 7310 3386
rect 7362 3334 7364 3386
rect 7308 3322 7364 3334
rect 7368 3164 7632 3174
rect 7424 3108 7472 3164
rect 7528 3108 7576 3164
rect 7368 3098 7632 3108
rect 6972 2882 7028 2894
rect 6972 2830 6974 2882
rect 7026 2830 7028 2882
rect 6972 2828 7028 2830
rect 6188 1710 6190 1762
rect 6242 1710 6244 1762
rect 4178 1596 4442 1606
rect 4234 1540 4282 1596
rect 4338 1540 4386 1596
rect 4178 1530 4442 1540
rect 3948 1428 4060 1484
rect 4004 800 4060 1428
rect 4676 1370 4732 1382
rect 4676 1318 4678 1370
rect 4730 1318 4732 1370
rect 4676 812 4732 1318
rect 6188 1370 6244 1710
rect 6188 1318 6190 1370
rect 6242 1318 6244 1370
rect 6188 1306 6244 1318
rect 6356 1988 6748 2044
rect 6804 2772 7028 2828
rect 0 -28 1148 28
rect 1288 0 1400 800
rect 2632 0 2744 800
rect 3976 0 4088 800
rect 5348 868 5628 924
rect 5348 800 5404 868
rect 4676 746 4732 756
rect 5320 0 5432 800
rect 5572 700 5628 868
rect 6356 812 6412 1988
rect 6804 1932 6860 2772
rect 7924 2770 7980 4004
rect 8963 3948 9227 3958
rect 9019 3892 9067 3948
rect 9123 3892 9171 3948
rect 8963 3882 9227 3892
rect 9380 3612 9436 8484
rect 10388 7644 10444 11172
rect 12348 11170 12404 11182
rect 12348 11118 12350 11170
rect 12402 11118 12404 11170
rect 10558 11004 10822 11014
rect 10614 10948 10662 11004
rect 10718 10948 10766 11004
rect 10558 10938 10822 10948
rect 11844 10892 11900 10902
rect 12348 10892 12404 11118
rect 11228 10722 11284 10734
rect 11228 10670 11230 10722
rect 11282 10670 11284 10722
rect 11228 10668 11284 10670
rect 11228 10602 11284 10612
rect 10558 9436 10822 9446
rect 10614 9380 10662 9436
rect 10718 9380 10766 9436
rect 10558 9370 10822 9380
rect 11340 8034 11396 8046
rect 11340 7982 11342 8034
rect 11394 7982 11396 8034
rect 11340 7980 11396 7982
rect 11844 7980 11900 10836
rect 11956 10836 12404 10892
rect 11956 10712 12012 10836
rect 12516 10780 12572 12852
rect 12628 11116 12684 13076
rect 12628 11060 12740 11116
rect 11956 10660 11958 10712
rect 12010 10660 12012 10712
rect 11956 8204 12012 10660
rect 12292 10724 12572 10780
rect 12292 10668 12348 10724
rect 12292 10536 12348 10612
rect 12684 10610 12740 11060
rect 13412 10892 13468 13200
rect 13860 11674 13916 11686
rect 13860 11622 13862 11674
rect 13914 11622 13916 11674
rect 13860 11564 13916 11622
rect 14756 11674 14812 13200
rect 14756 11622 14758 11674
rect 14810 11622 14812 11674
rect 14756 11610 14812 11622
rect 13860 11498 13916 11508
rect 13412 10826 13468 10836
rect 12684 10558 12686 10610
rect 12738 10558 12740 10610
rect 12153 10220 12417 10230
rect 12209 10164 12257 10220
rect 12313 10164 12361 10220
rect 12153 10154 12417 10164
rect 12684 9996 12740 10558
rect 13020 10444 13076 10454
rect 13860 10444 13916 10454
rect 13020 10442 13916 10444
rect 13020 10390 13022 10442
rect 13074 10390 13862 10442
rect 13914 10390 13916 10442
rect 13020 10388 13916 10390
rect 13020 10378 13076 10388
rect 13860 10378 13916 10388
rect 14756 10442 14812 10454
rect 14756 10390 14758 10442
rect 14810 10390 14812 10442
rect 12124 9940 12740 9996
rect 12124 9714 12180 9940
rect 12124 9662 12126 9714
rect 12178 9662 12180 9714
rect 12124 9650 12180 9662
rect 12153 8652 12417 8662
rect 12209 8596 12257 8652
rect 12313 8596 12361 8652
rect 12153 8586 12417 8596
rect 11956 8138 12012 8148
rect 11340 7924 11900 7980
rect 10558 7868 10822 7878
rect 10614 7812 10662 7868
rect 10718 7812 10766 7868
rect 10558 7802 10822 7812
rect 9548 7586 9604 7598
rect 10388 7588 10556 7644
rect 9548 7534 9550 7586
rect 9602 7534 9604 7586
rect 9548 7532 9604 7534
rect 9548 7466 9604 7476
rect 10276 7532 10332 7542
rect 10332 7476 10444 7532
rect 10276 7466 10332 7476
rect 10388 7474 10444 7476
rect 10388 7422 10390 7474
rect 10442 7422 10444 7474
rect 10388 7410 10444 7422
rect 9604 6524 9660 6534
rect 10500 6524 10556 7588
rect 11340 7532 11396 7924
rect 10836 7476 11396 7532
rect 10836 7474 10892 7476
rect 10836 7422 10838 7474
rect 10890 7422 10892 7474
rect 10836 7410 10892 7422
rect 8428 3556 9492 3612
rect 8428 3554 8484 3556
rect 8428 3502 8430 3554
rect 8482 3502 8484 3554
rect 8428 3490 8484 3502
rect 9436 2994 9492 3556
rect 9436 2942 9438 2994
rect 9490 2942 9492 2994
rect 9436 2930 9492 2942
rect 8260 2882 8316 2894
rect 8260 2830 8262 2882
rect 8314 2830 8316 2882
rect 8260 2828 8316 2830
rect 8260 2772 8876 2828
rect 7924 2718 7926 2770
rect 7978 2718 7980 2770
rect 7924 2706 7980 2718
rect 7812 2604 7868 2614
rect 7812 2602 8092 2604
rect 7812 2550 7814 2602
rect 7866 2550 8092 2602
rect 7812 2548 8092 2550
rect 7812 2538 7868 2548
rect 7700 1961 7756 1973
rect 7700 1932 7702 1961
rect 6132 756 6412 812
rect 6692 1909 7702 1932
rect 7754 1909 7756 1961
rect 6692 1876 7756 1909
rect 6692 800 6748 1876
rect 7924 1863 7980 1875
rect 7924 1811 7926 1863
rect 7978 1811 7980 1863
rect 7924 1708 7980 1811
rect 7924 1642 7980 1652
rect 7368 1596 7632 1606
rect 7424 1540 7472 1596
rect 7528 1540 7576 1596
rect 7368 1530 7632 1540
rect 8036 800 8092 2548
rect 8820 1932 8876 2772
rect 8963 2380 9227 2390
rect 9019 2324 9067 2380
rect 9123 2324 9171 2380
rect 8963 2314 9227 2324
rect 8820 1876 9380 1932
rect 9324 1874 9380 1876
rect 9324 1822 9326 1874
rect 9378 1822 9380 1874
rect 9324 1596 9380 1822
rect 9324 1540 9436 1596
rect 9380 800 9436 1540
rect 9604 812 9660 6468
rect 10388 6468 10556 6524
rect 10948 7306 11004 7318
rect 10948 7254 10950 7306
rect 11002 7254 11004 7306
rect 10052 6188 10108 6198
rect 10052 5068 10108 6132
rect 10052 5002 10108 5012
rect 10388 4508 10444 6468
rect 10558 6300 10822 6310
rect 10614 6244 10662 6300
rect 10718 6244 10766 6300
rect 10558 6234 10822 6244
rect 10558 4732 10822 4742
rect 10614 4676 10662 4732
rect 10718 4676 10766 4732
rect 10558 4666 10822 4676
rect 10668 4508 10724 4518
rect 10388 4506 10780 4508
rect 10388 4454 10670 4506
rect 10722 4454 10780 4506
rect 10388 4452 10780 4454
rect 10668 4442 10780 4452
rect 10724 3566 10780 4442
rect 10724 3514 10726 3566
rect 10778 3514 10780 3566
rect 10724 3502 10780 3514
rect 10220 3388 10276 3398
rect 10220 2884 10276 3332
rect 10558 3164 10822 3174
rect 10614 3108 10662 3164
rect 10718 3108 10766 3164
rect 10558 3098 10822 3108
rect 10164 2882 10276 2884
rect 10164 2830 10222 2882
rect 10274 2830 10276 2882
rect 10164 2818 10276 2830
rect 10164 1372 10220 2818
rect 10558 1596 10822 1606
rect 10614 1540 10662 1596
rect 10718 1540 10766 1596
rect 10558 1530 10822 1540
rect 10948 1372 11004 7254
rect 12153 7084 12417 7094
rect 12209 7028 12257 7084
rect 12313 7028 12361 7084
rect 12153 7018 12417 7028
rect 12153 5516 12417 5526
rect 12209 5460 12257 5516
rect 12313 5460 12361 5516
rect 12153 5450 12417 5460
rect 12740 4844 12796 4854
rect 12684 4788 12740 4844
rect 12684 4778 12796 4788
rect 12684 4226 12740 4778
rect 12684 4174 12686 4226
rect 12738 4174 12740 4226
rect 12684 4162 12740 4174
rect 12153 3948 12417 3958
rect 12209 3892 12257 3948
rect 12313 3892 12361 3948
rect 12153 3882 12417 3892
rect 11956 3724 12012 3734
rect 11956 3630 12012 3668
rect 13412 3724 13468 3734
rect 11172 3545 11228 3557
rect 11172 3493 11174 3545
rect 11226 3493 11228 3545
rect 11172 3388 11228 3493
rect 11172 3322 11228 3332
rect 12153 2380 12417 2390
rect 12209 2324 12257 2380
rect 12313 2324 12361 2380
rect 12153 2314 12417 2324
rect 10164 1306 10220 1316
rect 10724 1316 11004 1372
rect 12068 2156 12124 2166
rect 6132 700 6188 756
rect 5572 644 6188 700
rect 6664 0 6776 800
rect 8008 0 8120 800
rect 9352 0 9464 800
rect 10724 800 10780 1316
rect 12068 800 12124 2100
rect 13412 800 13468 3668
rect 14756 800 14812 10390
rect 9604 746 9660 756
rect 10696 0 10808 800
rect 12040 0 12152 800
rect 13384 0 13496 800
rect 14728 0 14840 800
rect 0 -56 800 -28
<< via2 >>
rect 84 10836 140 10892
rect 2583 11786 2639 11788
rect 2583 11734 2585 11786
rect 2585 11734 2637 11786
rect 2637 11734 2639 11786
rect 2583 11732 2639 11734
rect 2687 11786 2743 11788
rect 2687 11734 2689 11786
rect 2689 11734 2741 11786
rect 2741 11734 2743 11786
rect 2687 11732 2743 11734
rect 2791 11786 2847 11788
rect 2791 11734 2793 11786
rect 2793 11734 2845 11786
rect 2845 11734 2847 11786
rect 2791 11732 2847 11734
rect 2100 11508 2156 11564
rect 1764 10836 1820 10892
rect 2436 10836 2492 10892
rect 3164 10836 3220 10892
rect 2583 10218 2639 10220
rect 2583 10166 2585 10218
rect 2585 10166 2637 10218
rect 2637 10166 2639 10218
rect 2583 10164 2639 10166
rect 2687 10218 2743 10220
rect 2687 10166 2689 10218
rect 2689 10166 2741 10218
rect 2741 10166 2743 10218
rect 2687 10164 2743 10166
rect 2791 10218 2847 10220
rect 2791 10166 2793 10218
rect 2793 10166 2845 10218
rect 2845 10166 2847 10218
rect 2791 10164 2847 10166
rect 3892 12906 3948 12908
rect 3892 12854 3894 12906
rect 3894 12854 3946 12906
rect 3946 12854 3948 12906
rect 3892 12852 3948 12854
rect 3332 9268 3388 9324
rect 2156 8874 2212 8876
rect 2156 8822 2158 8874
rect 2158 8822 2210 8874
rect 2210 8822 2212 8874
rect 2156 8820 2212 8822
rect 2583 8650 2639 8652
rect 2583 8598 2585 8650
rect 2585 8598 2637 8650
rect 2637 8598 2639 8650
rect 2583 8596 2639 8598
rect 2687 8650 2743 8652
rect 2687 8598 2689 8650
rect 2689 8598 2741 8650
rect 2741 8598 2743 8650
rect 2687 8596 2743 8598
rect 2791 8650 2847 8652
rect 2791 8598 2793 8650
rect 2793 8598 2845 8650
rect 2845 8598 2847 8650
rect 2791 8596 2847 8598
rect 2583 7082 2639 7084
rect 2583 7030 2585 7082
rect 2585 7030 2637 7082
rect 2637 7030 2639 7082
rect 2583 7028 2639 7030
rect 2687 7082 2743 7084
rect 2687 7030 2689 7082
rect 2689 7030 2741 7082
rect 2741 7030 2743 7082
rect 2687 7028 2743 7030
rect 2791 7082 2847 7084
rect 2791 7030 2793 7082
rect 2793 7030 2845 7082
rect 2845 7030 2847 7082
rect 2791 7028 2847 7030
rect 4178 11002 4234 11004
rect 4178 10950 4180 11002
rect 4180 10950 4232 11002
rect 4232 10950 4234 11002
rect 4178 10948 4234 10950
rect 4282 11002 4338 11004
rect 4282 10950 4284 11002
rect 4284 10950 4336 11002
rect 4336 10950 4338 11002
rect 4282 10948 4338 10950
rect 4386 11002 4442 11004
rect 4386 10950 4388 11002
rect 4388 10950 4440 11002
rect 4440 10950 4442 11002
rect 4386 10948 4442 10950
rect 5773 11786 5829 11788
rect 5773 11734 5775 11786
rect 5775 11734 5827 11786
rect 5827 11734 5829 11786
rect 5773 11732 5829 11734
rect 5877 11786 5933 11788
rect 5877 11734 5879 11786
rect 5879 11734 5931 11786
rect 5931 11734 5933 11786
rect 5877 11732 5933 11734
rect 5981 11786 6037 11788
rect 5981 11734 5983 11786
rect 5983 11734 6035 11786
rect 6035 11734 6037 11786
rect 5981 11732 6037 11734
rect 5348 10836 5404 10892
rect 6692 10612 6748 10668
rect 7140 10276 7196 10332
rect 5773 10218 5829 10220
rect 5773 10166 5775 10218
rect 5775 10166 5827 10218
rect 5827 10166 5829 10218
rect 5773 10164 5829 10166
rect 5877 10218 5933 10220
rect 5877 10166 5879 10218
rect 5879 10166 5931 10218
rect 5931 10166 5933 10218
rect 5877 10164 5933 10166
rect 5981 10218 6037 10220
rect 5981 10166 5983 10218
rect 5983 10166 6035 10218
rect 6035 10166 6037 10218
rect 5981 10164 6037 10166
rect 7980 11508 8036 11564
rect 7368 11002 7424 11004
rect 7368 10950 7370 11002
rect 7370 10950 7422 11002
rect 7422 10950 7424 11002
rect 7368 10948 7424 10950
rect 7472 11002 7528 11004
rect 7472 10950 7474 11002
rect 7474 10950 7526 11002
rect 7526 10950 7528 11002
rect 7472 10948 7528 10950
rect 7576 11002 7632 11004
rect 7576 10950 7578 11002
rect 7578 10950 7630 11002
rect 7630 10950 7632 11002
rect 7576 10948 7632 10950
rect 7252 9492 7308 9548
rect 4178 9434 4234 9436
rect 4178 9382 4180 9434
rect 4180 9382 4232 9434
rect 4232 9382 4234 9434
rect 4178 9380 4234 9382
rect 4282 9434 4338 9436
rect 4282 9382 4284 9434
rect 4284 9382 4336 9434
rect 4336 9382 4338 9434
rect 4282 9380 4338 9382
rect 4386 9434 4442 9436
rect 4386 9382 4388 9434
rect 4388 9382 4440 9434
rect 4440 9382 4442 9434
rect 4386 9380 4442 9382
rect 7368 9434 7424 9436
rect 7368 9382 7370 9434
rect 7370 9382 7422 9434
rect 7422 9382 7424 9434
rect 7368 9380 7424 9382
rect 7472 9434 7528 9436
rect 7472 9382 7474 9434
rect 7474 9382 7526 9434
rect 7526 9382 7528 9434
rect 7472 9380 7528 9382
rect 7576 9434 7632 9436
rect 7576 9382 7578 9434
rect 7578 9382 7630 9434
rect 7630 9382 7632 9434
rect 7576 9380 7632 9382
rect 7084 9268 7140 9324
rect 7924 10612 7980 10668
rect 8148 10052 8204 10108
rect 8372 10276 8428 10332
rect 5773 8650 5829 8652
rect 5773 8598 5775 8650
rect 5775 8598 5827 8650
rect 5827 8598 5829 8650
rect 5773 8596 5829 8598
rect 5877 8650 5933 8652
rect 5877 8598 5879 8650
rect 5879 8598 5931 8650
rect 5931 8598 5933 8650
rect 5877 8596 5933 8598
rect 5981 8650 6037 8652
rect 5981 8598 5983 8650
rect 5983 8598 6035 8650
rect 6035 8598 6037 8650
rect 5981 8596 6037 8598
rect 4004 8484 4060 8540
rect 5796 8260 5852 8316
rect 6580 8260 6636 8316
rect 4178 7866 4234 7868
rect 4178 7814 4180 7866
rect 4180 7814 4232 7866
rect 4232 7814 4234 7866
rect 4178 7812 4234 7814
rect 4282 7866 4338 7868
rect 4282 7814 4284 7866
rect 4284 7814 4336 7866
rect 4336 7814 4338 7866
rect 4282 7812 4338 7814
rect 4386 7866 4442 7868
rect 4386 7814 4388 7866
rect 4388 7814 4440 7866
rect 4440 7814 4442 7866
rect 4386 7812 4442 7814
rect 5012 7588 5068 7644
rect 4178 6298 4234 6300
rect 4178 6246 4180 6298
rect 4180 6246 4232 6298
rect 4232 6246 4234 6298
rect 4178 6244 4234 6246
rect 4282 6298 4338 6300
rect 4282 6246 4284 6298
rect 4284 6246 4336 6298
rect 4336 6246 4338 6298
rect 4282 6244 4338 6246
rect 4386 6298 4442 6300
rect 4386 6246 4388 6298
rect 4388 6246 4440 6298
rect 4440 6246 4442 6298
rect 4386 6244 4442 6246
rect 2996 6132 3052 6188
rect 2583 5514 2639 5516
rect 2583 5462 2585 5514
rect 2585 5462 2637 5514
rect 2637 5462 2639 5514
rect 2583 5460 2639 5462
rect 2687 5514 2743 5516
rect 2687 5462 2689 5514
rect 2689 5462 2741 5514
rect 2741 5462 2743 5514
rect 2687 5460 2743 5462
rect 2791 5514 2847 5516
rect 2791 5462 2793 5514
rect 2793 5462 2845 5514
rect 2845 5462 2847 5514
rect 2791 5460 2847 5462
rect 3276 5012 3332 5068
rect 2583 3946 2639 3948
rect 2583 3894 2585 3946
rect 2585 3894 2637 3946
rect 2637 3894 2639 3946
rect 2583 3892 2639 3894
rect 2687 3946 2743 3948
rect 2687 3894 2689 3946
rect 2689 3894 2741 3946
rect 2741 3894 2743 3946
rect 2687 3892 2743 3894
rect 2791 3946 2847 3948
rect 2791 3894 2793 3946
rect 2793 3894 2845 3946
rect 2845 3894 2847 3946
rect 2791 3892 2847 3894
rect 2436 3386 2492 3388
rect 2436 3334 2438 3386
rect 2438 3334 2490 3386
rect 2490 3334 2492 3386
rect 2436 3332 2492 3334
rect 4178 4730 4234 4732
rect 4178 4678 4180 4730
rect 4180 4678 4232 4730
rect 4232 4678 4234 4730
rect 4178 4676 4234 4678
rect 4282 4730 4338 4732
rect 4282 4678 4284 4730
rect 4284 4678 4336 4730
rect 4336 4678 4338 4730
rect 4282 4676 4338 4678
rect 4386 4730 4442 4732
rect 4386 4678 4388 4730
rect 4388 4678 4440 4730
rect 4440 4678 4442 4730
rect 4386 4676 4442 4678
rect 4178 3162 4234 3164
rect 4178 3110 4180 3162
rect 4180 3110 4232 3162
rect 4232 3110 4234 3162
rect 4178 3108 4234 3110
rect 4282 3162 4338 3164
rect 4282 3110 4284 3162
rect 4284 3110 4336 3162
rect 4336 3110 4338 3162
rect 4282 3108 4338 3110
rect 4386 3162 4442 3164
rect 4386 3110 4388 3162
rect 4388 3110 4440 3162
rect 4440 3110 4442 3162
rect 4386 3108 4442 3110
rect 2583 2378 2639 2380
rect 2583 2326 2585 2378
rect 2585 2326 2637 2378
rect 2637 2326 2639 2378
rect 2583 2324 2639 2326
rect 2687 2378 2743 2380
rect 2687 2326 2689 2378
rect 2689 2326 2741 2378
rect 2741 2326 2743 2378
rect 2687 2324 2743 2326
rect 2791 2378 2847 2380
rect 2791 2326 2793 2378
rect 2793 2326 2845 2378
rect 2845 2326 2847 2378
rect 2791 2324 2847 2326
rect 7924 9492 7980 9548
rect 7140 8090 7142 8092
rect 7142 8090 7194 8092
rect 7194 8090 7196 8092
rect 7140 8036 7196 8090
rect 7700 8260 7756 8316
rect 7368 7866 7424 7868
rect 7368 7814 7370 7866
rect 7370 7814 7422 7866
rect 7422 7814 7424 7866
rect 7368 7812 7424 7814
rect 7472 7866 7528 7868
rect 7472 7814 7474 7866
rect 7474 7814 7526 7866
rect 7526 7814 7528 7866
rect 7472 7812 7528 7814
rect 7576 7866 7632 7868
rect 7576 7814 7578 7866
rect 7578 7814 7630 7866
rect 7630 7814 7632 7866
rect 7576 7812 7632 7814
rect 6524 7642 6580 7644
rect 6524 7590 6526 7642
rect 6526 7590 6578 7642
rect 6578 7590 6580 7642
rect 6524 7588 6580 7590
rect 5773 7082 5829 7084
rect 5773 7030 5775 7082
rect 5775 7030 5827 7082
rect 5827 7030 5829 7082
rect 5773 7028 5829 7030
rect 5877 7082 5933 7084
rect 5877 7030 5879 7082
rect 5879 7030 5931 7082
rect 5931 7030 5933 7082
rect 5877 7028 5933 7030
rect 5981 7082 6037 7084
rect 5981 7030 5983 7082
rect 5983 7030 6035 7082
rect 6035 7030 6037 7082
rect 5981 7028 6037 7030
rect 7368 6298 7424 6300
rect 7368 6246 7370 6298
rect 7370 6246 7422 6298
rect 7422 6246 7424 6298
rect 7368 6244 7424 6246
rect 7472 6298 7528 6300
rect 7472 6246 7474 6298
rect 7474 6246 7526 6298
rect 7526 6246 7528 6298
rect 7472 6244 7528 6246
rect 7576 6298 7632 6300
rect 7576 6246 7578 6298
rect 7578 6246 7630 6298
rect 7630 6246 7632 6298
rect 7576 6244 7632 6246
rect 5773 5514 5829 5516
rect 5773 5462 5775 5514
rect 5775 5462 5827 5514
rect 5827 5462 5829 5514
rect 5773 5460 5829 5462
rect 5877 5514 5933 5516
rect 5877 5462 5879 5514
rect 5879 5462 5931 5514
rect 5931 5462 5933 5514
rect 5877 5460 5933 5462
rect 5981 5514 6037 5516
rect 5981 5462 5983 5514
rect 5983 5462 6035 5514
rect 6035 5462 6037 5514
rect 5981 5460 6037 5462
rect 5572 4788 5628 4844
rect 5236 3332 5292 3388
rect 5773 3946 5829 3948
rect 5773 3894 5775 3946
rect 5775 3894 5827 3946
rect 5827 3894 5829 3946
rect 5773 3892 5829 3894
rect 5877 3946 5933 3948
rect 5877 3894 5879 3946
rect 5879 3894 5931 3946
rect 5931 3894 5933 3946
rect 5877 3892 5933 3894
rect 5981 3946 6037 3948
rect 5981 3894 5983 3946
rect 5983 3894 6035 3946
rect 6035 3894 6037 3946
rect 5981 3892 6037 3894
rect 6244 3444 6300 3500
rect 6076 3386 6132 3388
rect 6076 3334 6078 3386
rect 6078 3334 6130 3386
rect 6130 3334 6132 3386
rect 6076 3332 6132 3334
rect 5773 2378 5829 2380
rect 5773 2326 5775 2378
rect 5775 2326 5827 2378
rect 5827 2326 5829 2378
rect 5773 2324 5829 2326
rect 5877 2378 5933 2380
rect 5877 2326 5879 2378
rect 5879 2326 5931 2378
rect 5931 2326 5933 2378
rect 5877 2324 5933 2326
rect 5981 2378 6037 2380
rect 5981 2326 5983 2378
rect 5983 2326 6035 2378
rect 6035 2326 6037 2378
rect 5981 2324 6037 2326
rect 5012 2212 5068 2268
rect 4788 2100 4844 2156
rect 5516 2100 5572 2156
rect 1316 1204 1372 1260
rect 7368 4730 7424 4732
rect 7368 4678 7370 4730
rect 7370 4678 7422 4730
rect 7422 4678 7424 4730
rect 7368 4676 7424 4678
rect 7472 4730 7528 4732
rect 7472 4678 7474 4730
rect 7474 4678 7526 4730
rect 7526 4678 7528 4730
rect 7472 4676 7528 4678
rect 7576 4730 7632 4732
rect 7576 4678 7578 4730
rect 7578 4678 7630 4730
rect 7630 4678 7632 4730
rect 7576 4676 7632 4678
rect 8963 11786 9019 11788
rect 8963 11734 8965 11786
rect 8965 11734 9017 11786
rect 9017 11734 9019 11786
rect 8963 11732 9019 11734
rect 9067 11786 9123 11788
rect 9067 11734 9069 11786
rect 9069 11734 9121 11786
rect 9121 11734 9123 11786
rect 9067 11732 9123 11734
rect 9171 11786 9227 11788
rect 9171 11734 9173 11786
rect 9173 11734 9225 11786
rect 9225 11734 9227 11786
rect 9171 11732 9227 11734
rect 9716 11396 9772 11452
rect 8963 10218 9019 10220
rect 8963 10166 8965 10218
rect 8965 10166 9017 10218
rect 9017 10166 9019 10218
rect 8963 10164 9019 10166
rect 9067 10218 9123 10220
rect 9067 10166 9069 10218
rect 9069 10166 9121 10218
rect 9121 10166 9123 10218
rect 9067 10164 9123 10166
rect 9171 10218 9227 10220
rect 9171 10166 9173 10218
rect 9173 10166 9225 10218
rect 9225 10166 9227 10218
rect 9171 10164 9227 10166
rect 12516 12852 12572 12908
rect 12153 11786 12209 11788
rect 12153 11734 12155 11786
rect 12155 11734 12207 11786
rect 12207 11734 12209 11786
rect 12153 11732 12209 11734
rect 12257 11786 12313 11788
rect 12257 11734 12259 11786
rect 12259 11734 12311 11786
rect 12311 11734 12313 11786
rect 12257 11732 12313 11734
rect 12361 11786 12417 11788
rect 12361 11734 12363 11786
rect 12363 11734 12415 11786
rect 12415 11734 12417 11786
rect 12361 11732 12417 11734
rect 9716 10052 9772 10108
rect 8963 8650 9019 8652
rect 8963 8598 8965 8650
rect 8965 8598 9017 8650
rect 9017 8598 9019 8650
rect 8963 8596 9019 8598
rect 9067 8650 9123 8652
rect 9067 8598 9069 8650
rect 9069 8598 9121 8650
rect 9121 8598 9123 8650
rect 9067 8596 9123 8598
rect 9171 8650 9227 8652
rect 9171 8598 9173 8650
rect 9173 8598 9225 8650
rect 9225 8598 9227 8650
rect 9171 8596 9227 8598
rect 8484 8148 8540 8204
rect 9380 8484 9436 8540
rect 8876 8090 8932 8092
rect 8876 8038 8878 8090
rect 8878 8038 8930 8090
rect 8930 8038 8932 8090
rect 8876 8036 8932 8038
rect 8963 7082 9019 7084
rect 8963 7030 8965 7082
rect 8965 7030 9017 7082
rect 9017 7030 9019 7082
rect 8963 7028 9019 7030
rect 9067 7082 9123 7084
rect 9067 7030 9069 7082
rect 9069 7030 9121 7082
rect 9121 7030 9123 7082
rect 9067 7028 9123 7030
rect 9171 7082 9227 7084
rect 9171 7030 9173 7082
rect 9173 7030 9225 7082
rect 9225 7030 9227 7082
rect 9171 7028 9227 7030
rect 8820 6522 8876 6524
rect 8820 6470 8822 6522
rect 8822 6470 8874 6522
rect 8874 6470 8876 6522
rect 8820 6468 8876 6470
rect 8963 5514 9019 5516
rect 8963 5462 8965 5514
rect 8965 5462 9017 5514
rect 9017 5462 9019 5514
rect 8963 5460 9019 5462
rect 9067 5514 9123 5516
rect 9067 5462 9069 5514
rect 9069 5462 9121 5514
rect 9121 5462 9123 5514
rect 9067 5460 9123 5462
rect 9171 5514 9227 5516
rect 9171 5462 9173 5514
rect 9173 5462 9225 5514
rect 9225 5462 9227 5514
rect 9171 5460 9227 5462
rect 7812 3490 7814 3500
rect 7814 3490 7866 3500
rect 7866 3490 7868 3500
rect 7812 3444 7868 3490
rect 7368 3162 7424 3164
rect 7368 3110 7370 3162
rect 7370 3110 7422 3162
rect 7422 3110 7424 3162
rect 7368 3108 7424 3110
rect 7472 3162 7528 3164
rect 7472 3110 7474 3162
rect 7474 3110 7526 3162
rect 7526 3110 7528 3162
rect 7472 3108 7528 3110
rect 7576 3162 7632 3164
rect 7576 3110 7578 3162
rect 7578 3110 7630 3162
rect 7630 3110 7632 3162
rect 7576 3108 7632 3110
rect 4178 1594 4234 1596
rect 4178 1542 4180 1594
rect 4180 1542 4232 1594
rect 4232 1542 4234 1594
rect 4178 1540 4234 1542
rect 4282 1594 4338 1596
rect 4282 1542 4284 1594
rect 4284 1542 4336 1594
rect 4336 1542 4338 1594
rect 4282 1540 4338 1542
rect 4386 1594 4442 1596
rect 4386 1542 4388 1594
rect 4388 1542 4440 1594
rect 4440 1542 4442 1594
rect 4386 1540 4442 1542
rect 4676 756 4732 812
rect 8963 3946 9019 3948
rect 8963 3894 8965 3946
rect 8965 3894 9017 3946
rect 9017 3894 9019 3946
rect 8963 3892 9019 3894
rect 9067 3946 9123 3948
rect 9067 3894 9069 3946
rect 9069 3894 9121 3946
rect 9121 3894 9123 3946
rect 9067 3892 9123 3894
rect 9171 3946 9227 3948
rect 9171 3894 9173 3946
rect 9173 3894 9225 3946
rect 9225 3894 9227 3946
rect 9171 3892 9227 3894
rect 10558 11002 10614 11004
rect 10558 10950 10560 11002
rect 10560 10950 10612 11002
rect 10612 10950 10614 11002
rect 10558 10948 10614 10950
rect 10662 11002 10718 11004
rect 10662 10950 10664 11002
rect 10664 10950 10716 11002
rect 10716 10950 10718 11002
rect 10662 10948 10718 10950
rect 10766 11002 10822 11004
rect 10766 10950 10768 11002
rect 10768 10950 10820 11002
rect 10820 10950 10822 11002
rect 10766 10948 10822 10950
rect 11844 10836 11900 10892
rect 11228 10612 11284 10668
rect 10558 9434 10614 9436
rect 10558 9382 10560 9434
rect 10560 9382 10612 9434
rect 10612 9382 10614 9434
rect 10558 9380 10614 9382
rect 10662 9434 10718 9436
rect 10662 9382 10664 9434
rect 10664 9382 10716 9434
rect 10716 9382 10718 9434
rect 10662 9380 10718 9382
rect 10766 9434 10822 9436
rect 10766 9382 10768 9434
rect 10768 9382 10820 9434
rect 10820 9382 10822 9434
rect 10766 9380 10822 9382
rect 12292 10666 12348 10668
rect 12292 10614 12294 10666
rect 12294 10614 12346 10666
rect 12346 10614 12348 10666
rect 12292 10612 12348 10614
rect 13860 11508 13916 11564
rect 13412 10836 13468 10892
rect 12153 10218 12209 10220
rect 12153 10166 12155 10218
rect 12155 10166 12207 10218
rect 12207 10166 12209 10218
rect 12153 10164 12209 10166
rect 12257 10218 12313 10220
rect 12257 10166 12259 10218
rect 12259 10166 12311 10218
rect 12311 10166 12313 10218
rect 12257 10164 12313 10166
rect 12361 10218 12417 10220
rect 12361 10166 12363 10218
rect 12363 10166 12415 10218
rect 12415 10166 12417 10218
rect 12361 10164 12417 10166
rect 12153 8650 12209 8652
rect 12153 8598 12155 8650
rect 12155 8598 12207 8650
rect 12207 8598 12209 8650
rect 12153 8596 12209 8598
rect 12257 8650 12313 8652
rect 12257 8598 12259 8650
rect 12259 8598 12311 8650
rect 12311 8598 12313 8650
rect 12257 8596 12313 8598
rect 12361 8650 12417 8652
rect 12361 8598 12363 8650
rect 12363 8598 12415 8650
rect 12415 8598 12417 8650
rect 12361 8596 12417 8598
rect 11956 8148 12012 8204
rect 10558 7866 10614 7868
rect 10558 7814 10560 7866
rect 10560 7814 10612 7866
rect 10612 7814 10614 7866
rect 10558 7812 10614 7814
rect 10662 7866 10718 7868
rect 10662 7814 10664 7866
rect 10664 7814 10716 7866
rect 10716 7814 10718 7866
rect 10662 7812 10718 7814
rect 10766 7866 10822 7868
rect 10766 7814 10768 7866
rect 10768 7814 10820 7866
rect 10820 7814 10822 7866
rect 10766 7812 10822 7814
rect 9548 7476 9604 7532
rect 10276 7476 10332 7532
rect 9604 6468 9660 6524
rect 7924 1652 7980 1708
rect 7368 1594 7424 1596
rect 7368 1542 7370 1594
rect 7370 1542 7422 1594
rect 7422 1542 7424 1594
rect 7368 1540 7424 1542
rect 7472 1594 7528 1596
rect 7472 1542 7474 1594
rect 7474 1542 7526 1594
rect 7526 1542 7528 1594
rect 7472 1540 7528 1542
rect 7576 1594 7632 1596
rect 7576 1542 7578 1594
rect 7578 1542 7630 1594
rect 7630 1542 7632 1594
rect 7576 1540 7632 1542
rect 8963 2378 9019 2380
rect 8963 2326 8965 2378
rect 8965 2326 9017 2378
rect 9017 2326 9019 2378
rect 8963 2324 9019 2326
rect 9067 2378 9123 2380
rect 9067 2326 9069 2378
rect 9069 2326 9121 2378
rect 9121 2326 9123 2378
rect 9067 2324 9123 2326
rect 9171 2378 9227 2380
rect 9171 2326 9173 2378
rect 9173 2326 9225 2378
rect 9225 2326 9227 2378
rect 9171 2324 9227 2326
rect 10052 6132 10108 6188
rect 10052 5012 10108 5068
rect 10558 6298 10614 6300
rect 10558 6246 10560 6298
rect 10560 6246 10612 6298
rect 10612 6246 10614 6298
rect 10558 6244 10614 6246
rect 10662 6298 10718 6300
rect 10662 6246 10664 6298
rect 10664 6246 10716 6298
rect 10716 6246 10718 6298
rect 10662 6244 10718 6246
rect 10766 6298 10822 6300
rect 10766 6246 10768 6298
rect 10768 6246 10820 6298
rect 10820 6246 10822 6298
rect 10766 6244 10822 6246
rect 10558 4730 10614 4732
rect 10558 4678 10560 4730
rect 10560 4678 10612 4730
rect 10612 4678 10614 4730
rect 10558 4676 10614 4678
rect 10662 4730 10718 4732
rect 10662 4678 10664 4730
rect 10664 4678 10716 4730
rect 10716 4678 10718 4730
rect 10662 4676 10718 4678
rect 10766 4730 10822 4732
rect 10766 4678 10768 4730
rect 10768 4678 10820 4730
rect 10820 4678 10822 4730
rect 10766 4676 10822 4678
rect 10220 3332 10276 3388
rect 10558 3162 10614 3164
rect 10558 3110 10560 3162
rect 10560 3110 10612 3162
rect 10612 3110 10614 3162
rect 10558 3108 10614 3110
rect 10662 3162 10718 3164
rect 10662 3110 10664 3162
rect 10664 3110 10716 3162
rect 10716 3110 10718 3162
rect 10662 3108 10718 3110
rect 10766 3162 10822 3164
rect 10766 3110 10768 3162
rect 10768 3110 10820 3162
rect 10820 3110 10822 3162
rect 10766 3108 10822 3110
rect 10558 1594 10614 1596
rect 10558 1542 10560 1594
rect 10560 1542 10612 1594
rect 10612 1542 10614 1594
rect 10558 1540 10614 1542
rect 10662 1594 10718 1596
rect 10662 1542 10664 1594
rect 10664 1542 10716 1594
rect 10716 1542 10718 1594
rect 10662 1540 10718 1542
rect 10766 1594 10822 1596
rect 10766 1542 10768 1594
rect 10768 1542 10820 1594
rect 10820 1542 10822 1594
rect 10766 1540 10822 1542
rect 12153 7082 12209 7084
rect 12153 7030 12155 7082
rect 12155 7030 12207 7082
rect 12207 7030 12209 7082
rect 12153 7028 12209 7030
rect 12257 7082 12313 7084
rect 12257 7030 12259 7082
rect 12259 7030 12311 7082
rect 12311 7030 12313 7082
rect 12257 7028 12313 7030
rect 12361 7082 12417 7084
rect 12361 7030 12363 7082
rect 12363 7030 12415 7082
rect 12415 7030 12417 7082
rect 12361 7028 12417 7030
rect 12153 5514 12209 5516
rect 12153 5462 12155 5514
rect 12155 5462 12207 5514
rect 12207 5462 12209 5514
rect 12153 5460 12209 5462
rect 12257 5514 12313 5516
rect 12257 5462 12259 5514
rect 12259 5462 12311 5514
rect 12311 5462 12313 5514
rect 12257 5460 12313 5462
rect 12361 5514 12417 5516
rect 12361 5462 12363 5514
rect 12363 5462 12415 5514
rect 12415 5462 12417 5514
rect 12361 5460 12417 5462
rect 12740 4788 12796 4844
rect 12153 3946 12209 3948
rect 12153 3894 12155 3946
rect 12155 3894 12207 3946
rect 12207 3894 12209 3946
rect 12153 3892 12209 3894
rect 12257 3946 12313 3948
rect 12257 3894 12259 3946
rect 12259 3894 12311 3946
rect 12311 3894 12313 3946
rect 12257 3892 12313 3894
rect 12361 3946 12417 3948
rect 12361 3894 12363 3946
rect 12363 3894 12415 3946
rect 12415 3894 12417 3946
rect 12361 3892 12417 3894
rect 11956 3722 12012 3724
rect 11956 3670 11958 3722
rect 11958 3670 12010 3722
rect 12010 3670 12012 3722
rect 11956 3668 12012 3670
rect 13412 3668 13468 3724
rect 11172 3332 11228 3388
rect 12153 2378 12209 2380
rect 12153 2326 12155 2378
rect 12155 2326 12207 2378
rect 12207 2326 12209 2378
rect 12153 2324 12209 2326
rect 12257 2378 12313 2380
rect 12257 2326 12259 2378
rect 12259 2326 12311 2378
rect 12311 2326 12313 2378
rect 12257 2324 12313 2326
rect 12361 2378 12417 2380
rect 12361 2326 12363 2378
rect 12363 2326 12415 2378
rect 12415 2326 12417 2378
rect 12361 2324 12417 2326
rect 10164 1316 10220 1372
rect 12068 2100 12124 2156
rect 9604 756 9660 812
<< metal3 >>
rect 0 12908 800 12936
rect 14200 12908 15000 12936
rect 0 12852 3892 12908
rect 3948 12852 3958 12908
rect 12506 12852 12516 12908
rect 12572 12852 15000 12908
rect 0 12824 800 12852
rect 14200 12824 15000 12852
rect 2573 11732 2583 11788
rect 2639 11732 2687 11788
rect 2743 11732 2791 11788
rect 2847 11732 2857 11788
rect 5763 11732 5773 11788
rect 5829 11732 5877 11788
rect 5933 11732 5981 11788
rect 6037 11732 6047 11788
rect 8953 11732 8963 11788
rect 9019 11732 9067 11788
rect 9123 11732 9171 11788
rect 9227 11732 9237 11788
rect 12143 11732 12153 11788
rect 12209 11732 12257 11788
rect 12313 11732 12361 11788
rect 12417 11732 12427 11788
rect 0 11564 800 11592
rect 14200 11564 15000 11592
rect 0 11508 2100 11564
rect 2156 11508 2166 11564
rect 7970 11508 7980 11564
rect 8036 11508 13860 11564
rect 13916 11508 13926 11564
rect 14084 11508 15000 11564
rect 0 11480 800 11508
rect 14084 11452 14140 11508
rect 14200 11480 15000 11508
rect 9706 11396 9716 11452
rect 9772 11396 14140 11452
rect 4168 10948 4178 11004
rect 4234 10948 4282 11004
rect 4338 10948 4386 11004
rect 4442 10948 4452 11004
rect 7358 10948 7368 11004
rect 7424 10948 7472 11004
rect 7528 10948 7576 11004
rect 7632 10948 7642 11004
rect 10548 10948 10558 11004
rect 10614 10948 10662 11004
rect 10718 10948 10766 11004
rect 10822 10948 10832 11004
rect 74 10836 84 10892
rect 140 10836 1764 10892
rect 1820 10836 1830 10892
rect 2426 10836 2436 10892
rect 2492 10836 3164 10892
rect 3220 10836 5348 10892
rect 5404 10836 5414 10892
rect 11834 10836 11844 10892
rect 11900 10836 13412 10892
rect 13468 10836 13478 10892
rect 6682 10612 6692 10668
rect 6748 10612 7924 10668
rect 7980 10612 7990 10668
rect 11218 10612 11228 10668
rect 11284 10612 12292 10668
rect 12348 10612 12358 10668
rect 2436 10276 7140 10332
rect 7196 10276 7206 10332
rect 8362 10276 8372 10332
rect 8428 10276 12572 10332
rect 0 10220 800 10248
rect 2436 10220 2492 10276
rect 12516 10220 12572 10276
rect 14200 10220 15000 10248
rect 0 10164 2492 10220
rect 2573 10164 2583 10220
rect 2639 10164 2687 10220
rect 2743 10164 2791 10220
rect 2847 10164 2857 10220
rect 5763 10164 5773 10220
rect 5829 10164 5877 10220
rect 5933 10164 5981 10220
rect 6037 10164 6047 10220
rect 8953 10164 8963 10220
rect 9019 10164 9067 10220
rect 9123 10164 9171 10220
rect 9227 10164 9237 10220
rect 12143 10164 12153 10220
rect 12209 10164 12257 10220
rect 12313 10164 12361 10220
rect 12417 10164 12427 10220
rect 12516 10164 15000 10220
rect 0 10136 800 10164
rect 14200 10136 15000 10164
rect 8138 10052 8148 10108
rect 8204 10052 9716 10108
rect 9772 10052 9782 10108
rect 7242 9492 7252 9548
rect 7308 9492 7924 9548
rect 7980 9492 7990 9548
rect 4168 9380 4178 9436
rect 4234 9380 4282 9436
rect 4338 9380 4386 9436
rect 4442 9380 4452 9436
rect 7358 9380 7368 9436
rect 7424 9380 7472 9436
rect 7528 9380 7576 9436
rect 7632 9380 7642 9436
rect 10548 9380 10558 9436
rect 10614 9380 10662 9436
rect 10718 9380 10766 9436
rect 10822 9380 10832 9436
rect 3322 9268 3332 9324
rect 3388 9268 7084 9324
rect 7140 9268 7150 9324
rect 0 8876 800 8904
rect 14200 8876 15000 8904
rect 0 8820 2156 8876
rect 2212 8820 2222 8876
rect 14084 8820 15000 8876
rect 0 8792 800 8820
rect 2573 8596 2583 8652
rect 2639 8596 2687 8652
rect 2743 8596 2791 8652
rect 2847 8596 2857 8652
rect 5763 8596 5773 8652
rect 5829 8596 5877 8652
rect 5933 8596 5981 8652
rect 6037 8596 6047 8652
rect 8953 8596 8963 8652
rect 9019 8596 9067 8652
rect 9123 8596 9171 8652
rect 9227 8596 9237 8652
rect 12143 8596 12153 8652
rect 12209 8596 12257 8652
rect 12313 8596 12361 8652
rect 12417 8596 12427 8652
rect 14084 8540 14140 8820
rect 14200 8792 15000 8820
rect 3444 8484 4004 8540
rect 4060 8484 4070 8540
rect 9370 8484 9380 8540
rect 9436 8484 11788 8540
rect 14084 8484 14364 8540
rect 3444 8316 3500 8484
rect 11732 8316 11788 8484
rect 14308 8316 14364 8484
rect 3444 8260 5796 8316
rect 5852 8260 5862 8316
rect 6570 8260 6580 8316
rect 6636 8260 7700 8316
rect 7756 8260 7766 8316
rect 11732 8260 14364 8316
rect 8474 8148 8484 8204
rect 8540 8148 11956 8204
rect 12012 8148 12022 8204
rect 7130 8036 7140 8092
rect 7196 8036 8876 8092
rect 8932 8036 14364 8092
rect 4168 7812 4178 7868
rect 4234 7812 4282 7868
rect 4338 7812 4386 7868
rect 4442 7812 4452 7868
rect 7358 7812 7368 7868
rect 7424 7812 7472 7868
rect 7528 7812 7576 7868
rect 7632 7812 7642 7868
rect 10548 7812 10558 7868
rect 10614 7812 10662 7868
rect 10718 7812 10766 7868
rect 10822 7812 10832 7868
rect 14308 7756 14364 8036
rect 14084 7700 14364 7756
rect 5002 7588 5012 7644
rect 5068 7588 6524 7644
rect 6580 7588 6590 7644
rect 0 7532 800 7560
rect 14084 7532 14140 7700
rect 14200 7532 15000 7560
rect 0 7476 9548 7532
rect 9604 7476 10276 7532
rect 10332 7476 10342 7532
rect 14084 7476 15000 7532
rect 0 7448 800 7476
rect 14200 7448 15000 7476
rect 2573 7028 2583 7084
rect 2639 7028 2687 7084
rect 2743 7028 2791 7084
rect 2847 7028 2857 7084
rect 5763 7028 5773 7084
rect 5829 7028 5877 7084
rect 5933 7028 5981 7084
rect 6037 7028 6047 7084
rect 8953 7028 8963 7084
rect 9019 7028 9067 7084
rect 9123 7028 9171 7084
rect 9227 7028 9237 7084
rect 12143 7028 12153 7084
rect 12209 7028 12257 7084
rect 12313 7028 12361 7084
rect 12417 7028 12427 7084
rect 8810 6468 8820 6524
rect 8876 6468 9604 6524
rect 9660 6468 9670 6524
rect 4168 6244 4178 6300
rect 4234 6244 4282 6300
rect 4338 6244 4386 6300
rect 4442 6244 4452 6300
rect 7358 6244 7368 6300
rect 7424 6244 7472 6300
rect 7528 6244 7576 6300
rect 7632 6244 7642 6300
rect 10548 6244 10558 6300
rect 10614 6244 10662 6300
rect 10718 6244 10766 6300
rect 10822 6244 10832 6300
rect 0 6188 800 6216
rect 14200 6188 15000 6216
rect 0 6132 2996 6188
rect 3052 6132 3062 6188
rect 10042 6132 10052 6188
rect 10108 6132 15000 6188
rect 0 6104 800 6132
rect 14200 6104 15000 6132
rect 2573 5460 2583 5516
rect 2639 5460 2687 5516
rect 2743 5460 2791 5516
rect 2847 5460 2857 5516
rect 5763 5460 5773 5516
rect 5829 5460 5877 5516
rect 5933 5460 5981 5516
rect 6037 5460 6047 5516
rect 8953 5460 8963 5516
rect 9019 5460 9067 5516
rect 9123 5460 9171 5516
rect 9227 5460 9237 5516
rect 12143 5460 12153 5516
rect 12209 5460 12257 5516
rect 12313 5460 12361 5516
rect 12417 5460 12427 5516
rect 3266 5012 3276 5068
rect 3332 5012 10052 5068
rect 10108 5012 10118 5068
rect 0 4844 800 4872
rect 14200 4844 15000 4872
rect 0 4788 5572 4844
rect 5628 4788 5638 4844
rect 12730 4788 12740 4844
rect 12796 4788 15000 4844
rect 0 4760 800 4788
rect 14200 4760 15000 4788
rect 4168 4676 4178 4732
rect 4234 4676 4282 4732
rect 4338 4676 4386 4732
rect 4442 4676 4452 4732
rect 7358 4676 7368 4732
rect 7424 4676 7472 4732
rect 7528 4676 7576 4732
rect 7632 4676 7642 4732
rect 10548 4676 10558 4732
rect 10614 4676 10662 4732
rect 10718 4676 10766 4732
rect 10822 4676 10832 4732
rect 2573 3892 2583 3948
rect 2639 3892 2687 3948
rect 2743 3892 2791 3948
rect 2847 3892 2857 3948
rect 5763 3892 5773 3948
rect 5829 3892 5877 3948
rect 5933 3892 5981 3948
rect 6037 3892 6047 3948
rect 8953 3892 8963 3948
rect 9019 3892 9067 3948
rect 9123 3892 9171 3948
rect 9227 3892 9237 3948
rect 12143 3892 12153 3948
rect 12209 3892 12257 3948
rect 12313 3892 12361 3948
rect 12417 3892 12427 3948
rect 11946 3668 11956 3724
rect 12012 3668 13412 3724
rect 13468 3668 13478 3724
rect 0 3500 800 3528
rect 14200 3500 15000 3528
rect 0 3444 2492 3500
rect 6234 3444 6244 3500
rect 6300 3444 7812 3500
rect 7868 3444 7878 3500
rect 8372 3444 15000 3500
rect 0 3416 800 3444
rect 2436 3388 2492 3444
rect 8372 3388 8428 3444
rect 14200 3416 15000 3444
rect 2426 3332 2436 3388
rect 2492 3332 2502 3388
rect 5226 3332 5236 3388
rect 5292 3332 6076 3388
rect 6132 3332 8428 3388
rect 10210 3332 10220 3388
rect 10276 3332 11172 3388
rect 11228 3332 11238 3388
rect 4168 3108 4178 3164
rect 4234 3108 4282 3164
rect 4338 3108 4386 3164
rect 4442 3108 4452 3164
rect 7358 3108 7368 3164
rect 7424 3108 7472 3164
rect 7528 3108 7576 3164
rect 7632 3108 7642 3164
rect 10548 3108 10558 3164
rect 10614 3108 10662 3164
rect 10718 3108 10766 3164
rect 10822 3108 10832 3164
rect 2573 2324 2583 2380
rect 2639 2324 2687 2380
rect 2743 2324 2791 2380
rect 2847 2324 2857 2380
rect 5763 2324 5773 2380
rect 5829 2324 5877 2380
rect 5933 2324 5981 2380
rect 6037 2324 6047 2380
rect 8953 2324 8963 2380
rect 9019 2324 9067 2380
rect 9123 2324 9171 2380
rect 9227 2324 9237 2380
rect 12143 2324 12153 2380
rect 12209 2324 12257 2380
rect 12313 2324 12361 2380
rect 12417 2324 12427 2380
rect 4564 2212 5012 2268
rect 5068 2212 5078 2268
rect 0 2156 800 2184
rect 4564 2156 4620 2212
rect 14200 2156 15000 2184
rect 0 2100 4620 2156
rect 4778 2100 4788 2156
rect 4844 2100 5516 2156
rect 5572 2100 12068 2156
rect 12124 2100 12134 2156
rect 12292 2100 15000 2156
rect 0 2072 800 2100
rect 12292 1708 12348 2100
rect 14200 2072 15000 2100
rect 7914 1652 7924 1708
rect 7980 1652 12348 1708
rect 4168 1540 4178 1596
rect 4234 1540 4282 1596
rect 4338 1540 4386 1596
rect 4442 1540 4452 1596
rect 7358 1540 7368 1596
rect 7424 1540 7472 1596
rect 7528 1540 7576 1596
rect 7632 1540 7642 1596
rect 10548 1540 10558 1596
rect 10614 1540 10662 1596
rect 10718 1540 10766 1596
rect 10822 1540 10832 1596
rect 1316 1316 10164 1372
rect 10220 1316 10230 1372
rect 1316 1260 1372 1316
rect 1306 1204 1316 1260
rect 1372 1204 1382 1260
rect 0 812 800 840
rect 14200 812 15000 840
rect 0 756 4676 812
rect 4732 756 4742 812
rect 9594 756 9604 812
rect 9660 756 15000 812
rect 0 728 800 756
rect 14200 728 15000 756
<< via3 >>
rect 2583 11732 2639 11788
rect 2687 11732 2743 11788
rect 2791 11732 2847 11788
rect 5773 11732 5829 11788
rect 5877 11732 5933 11788
rect 5981 11732 6037 11788
rect 8963 11732 9019 11788
rect 9067 11732 9123 11788
rect 9171 11732 9227 11788
rect 12153 11732 12209 11788
rect 12257 11732 12313 11788
rect 12361 11732 12417 11788
rect 4178 10948 4234 11004
rect 4282 10948 4338 11004
rect 4386 10948 4442 11004
rect 7368 10948 7424 11004
rect 7472 10948 7528 11004
rect 7576 10948 7632 11004
rect 10558 10948 10614 11004
rect 10662 10948 10718 11004
rect 10766 10948 10822 11004
rect 2583 10164 2639 10220
rect 2687 10164 2743 10220
rect 2791 10164 2847 10220
rect 5773 10164 5829 10220
rect 5877 10164 5933 10220
rect 5981 10164 6037 10220
rect 8963 10164 9019 10220
rect 9067 10164 9123 10220
rect 9171 10164 9227 10220
rect 12153 10164 12209 10220
rect 12257 10164 12313 10220
rect 12361 10164 12417 10220
rect 4178 9380 4234 9436
rect 4282 9380 4338 9436
rect 4386 9380 4442 9436
rect 7368 9380 7424 9436
rect 7472 9380 7528 9436
rect 7576 9380 7632 9436
rect 10558 9380 10614 9436
rect 10662 9380 10718 9436
rect 10766 9380 10822 9436
rect 2583 8596 2639 8652
rect 2687 8596 2743 8652
rect 2791 8596 2847 8652
rect 5773 8596 5829 8652
rect 5877 8596 5933 8652
rect 5981 8596 6037 8652
rect 8963 8596 9019 8652
rect 9067 8596 9123 8652
rect 9171 8596 9227 8652
rect 12153 8596 12209 8652
rect 12257 8596 12313 8652
rect 12361 8596 12417 8652
rect 4178 7812 4234 7868
rect 4282 7812 4338 7868
rect 4386 7812 4442 7868
rect 7368 7812 7424 7868
rect 7472 7812 7528 7868
rect 7576 7812 7632 7868
rect 10558 7812 10614 7868
rect 10662 7812 10718 7868
rect 10766 7812 10822 7868
rect 2583 7028 2639 7084
rect 2687 7028 2743 7084
rect 2791 7028 2847 7084
rect 5773 7028 5829 7084
rect 5877 7028 5933 7084
rect 5981 7028 6037 7084
rect 8963 7028 9019 7084
rect 9067 7028 9123 7084
rect 9171 7028 9227 7084
rect 12153 7028 12209 7084
rect 12257 7028 12313 7084
rect 12361 7028 12417 7084
rect 4178 6244 4234 6300
rect 4282 6244 4338 6300
rect 4386 6244 4442 6300
rect 7368 6244 7424 6300
rect 7472 6244 7528 6300
rect 7576 6244 7632 6300
rect 10558 6244 10614 6300
rect 10662 6244 10718 6300
rect 10766 6244 10822 6300
rect 2583 5460 2639 5516
rect 2687 5460 2743 5516
rect 2791 5460 2847 5516
rect 5773 5460 5829 5516
rect 5877 5460 5933 5516
rect 5981 5460 6037 5516
rect 8963 5460 9019 5516
rect 9067 5460 9123 5516
rect 9171 5460 9227 5516
rect 12153 5460 12209 5516
rect 12257 5460 12313 5516
rect 12361 5460 12417 5516
rect 4178 4676 4234 4732
rect 4282 4676 4338 4732
rect 4386 4676 4442 4732
rect 7368 4676 7424 4732
rect 7472 4676 7528 4732
rect 7576 4676 7632 4732
rect 10558 4676 10614 4732
rect 10662 4676 10718 4732
rect 10766 4676 10822 4732
rect 2583 3892 2639 3948
rect 2687 3892 2743 3948
rect 2791 3892 2847 3948
rect 5773 3892 5829 3948
rect 5877 3892 5933 3948
rect 5981 3892 6037 3948
rect 8963 3892 9019 3948
rect 9067 3892 9123 3948
rect 9171 3892 9227 3948
rect 12153 3892 12209 3948
rect 12257 3892 12313 3948
rect 12361 3892 12417 3948
rect 4178 3108 4234 3164
rect 4282 3108 4338 3164
rect 4386 3108 4442 3164
rect 7368 3108 7424 3164
rect 7472 3108 7528 3164
rect 7576 3108 7632 3164
rect 10558 3108 10614 3164
rect 10662 3108 10718 3164
rect 10766 3108 10822 3164
rect 2583 2324 2639 2380
rect 2687 2324 2743 2380
rect 2791 2324 2847 2380
rect 5773 2324 5829 2380
rect 5877 2324 5933 2380
rect 5981 2324 6037 2380
rect 8963 2324 9019 2380
rect 9067 2324 9123 2380
rect 9171 2324 9227 2380
rect 12153 2324 12209 2380
rect 12257 2324 12313 2380
rect 12361 2324 12417 2380
rect 4178 1540 4234 1596
rect 4282 1540 4338 1596
rect 4386 1540 4442 1596
rect 7368 1540 7424 1596
rect 7472 1540 7528 1596
rect 7576 1540 7632 1596
rect 10558 1540 10614 1596
rect 10662 1540 10718 1596
rect 10766 1540 10822 1596
<< metal4 >>
rect 2555 11788 2875 11820
rect 2555 11732 2583 11788
rect 2639 11732 2687 11788
rect 2743 11732 2791 11788
rect 2847 11732 2875 11788
rect 2555 11206 2875 11732
rect 2555 11150 2583 11206
rect 2639 11150 2687 11206
rect 2743 11150 2791 11206
rect 2847 11150 2875 11206
rect 2555 11102 2875 11150
rect 2555 11046 2583 11102
rect 2639 11046 2687 11102
rect 2743 11046 2791 11102
rect 2847 11046 2875 11102
rect 2555 10998 2875 11046
rect 2555 10942 2583 10998
rect 2639 10942 2687 10998
rect 2743 10942 2791 10998
rect 2847 10942 2875 10998
rect 2555 10220 2875 10942
rect 2555 10164 2583 10220
rect 2639 10164 2687 10220
rect 2743 10164 2791 10220
rect 2847 10164 2875 10220
rect 2555 8652 2875 10164
rect 2555 8596 2583 8652
rect 2639 8596 2687 8652
rect 2743 8596 2791 8652
rect 2847 8596 2875 8652
rect 2555 8490 2875 8596
rect 2555 8434 2583 8490
rect 2639 8434 2687 8490
rect 2743 8434 2791 8490
rect 2847 8434 2875 8490
rect 2555 8386 2875 8434
rect 2555 8330 2583 8386
rect 2639 8330 2687 8386
rect 2743 8330 2791 8386
rect 2847 8330 2875 8386
rect 2555 8282 2875 8330
rect 2555 8226 2583 8282
rect 2639 8226 2687 8282
rect 2743 8226 2791 8282
rect 2847 8226 2875 8282
rect 2555 7084 2875 8226
rect 2555 7028 2583 7084
rect 2639 7028 2687 7084
rect 2743 7028 2791 7084
rect 2847 7028 2875 7084
rect 2555 5774 2875 7028
rect 2555 5718 2583 5774
rect 2639 5718 2687 5774
rect 2743 5718 2791 5774
rect 2847 5718 2875 5774
rect 2555 5670 2875 5718
rect 2555 5614 2583 5670
rect 2639 5614 2687 5670
rect 2743 5614 2791 5670
rect 2847 5614 2875 5670
rect 2555 5566 2875 5614
rect 2555 5460 2583 5566
rect 2639 5460 2687 5566
rect 2743 5460 2791 5566
rect 2847 5460 2875 5566
rect 2555 3948 2875 5460
rect 2555 3892 2583 3948
rect 2639 3892 2687 3948
rect 2743 3892 2791 3948
rect 2847 3892 2875 3948
rect 2555 3058 2875 3892
rect 2555 3002 2583 3058
rect 2639 3002 2687 3058
rect 2743 3002 2791 3058
rect 2847 3002 2875 3058
rect 2555 2954 2875 3002
rect 2555 2898 2583 2954
rect 2639 2898 2687 2954
rect 2743 2898 2791 2954
rect 2847 2898 2875 2954
rect 2555 2850 2875 2898
rect 2555 2794 2583 2850
rect 2639 2794 2687 2850
rect 2743 2794 2791 2850
rect 2847 2794 2875 2850
rect 2555 2380 2875 2794
rect 2555 2324 2583 2380
rect 2639 2324 2687 2380
rect 2743 2324 2791 2380
rect 2847 2324 2875 2380
rect 2555 1508 2875 2324
rect 4150 11004 4470 11820
rect 4150 10948 4178 11004
rect 4234 10948 4282 11004
rect 4338 10948 4386 11004
rect 4442 10948 4470 11004
rect 4150 9848 4470 10948
rect 4150 9792 4178 9848
rect 4234 9792 4282 9848
rect 4338 9792 4386 9848
rect 4442 9792 4470 9848
rect 4150 9744 4470 9792
rect 4150 9688 4178 9744
rect 4234 9688 4282 9744
rect 4338 9688 4386 9744
rect 4442 9688 4470 9744
rect 4150 9640 4470 9688
rect 4150 9584 4178 9640
rect 4234 9584 4282 9640
rect 4338 9584 4386 9640
rect 4442 9584 4470 9640
rect 4150 9436 4470 9584
rect 4150 9380 4178 9436
rect 4234 9380 4282 9436
rect 4338 9380 4386 9436
rect 4442 9380 4470 9436
rect 4150 7868 4470 9380
rect 4150 7812 4178 7868
rect 4234 7812 4282 7868
rect 4338 7812 4386 7868
rect 4442 7812 4470 7868
rect 4150 7132 4470 7812
rect 4150 7076 4178 7132
rect 4234 7076 4282 7132
rect 4338 7076 4386 7132
rect 4442 7076 4470 7132
rect 4150 7028 4470 7076
rect 4150 6972 4178 7028
rect 4234 6972 4282 7028
rect 4338 6972 4386 7028
rect 4442 6972 4470 7028
rect 4150 6924 4470 6972
rect 4150 6868 4178 6924
rect 4234 6868 4282 6924
rect 4338 6868 4386 6924
rect 4442 6868 4470 6924
rect 4150 6300 4470 6868
rect 4150 6244 4178 6300
rect 4234 6244 4282 6300
rect 4338 6244 4386 6300
rect 4442 6244 4470 6300
rect 4150 4732 4470 6244
rect 4150 4676 4178 4732
rect 4234 4676 4282 4732
rect 4338 4676 4386 4732
rect 4442 4676 4470 4732
rect 4150 4416 4470 4676
rect 4150 4360 4178 4416
rect 4234 4360 4282 4416
rect 4338 4360 4386 4416
rect 4442 4360 4470 4416
rect 4150 4312 4470 4360
rect 4150 4256 4178 4312
rect 4234 4256 4282 4312
rect 4338 4256 4386 4312
rect 4442 4256 4470 4312
rect 4150 4208 4470 4256
rect 4150 4152 4178 4208
rect 4234 4152 4282 4208
rect 4338 4152 4386 4208
rect 4442 4152 4470 4208
rect 4150 3164 4470 4152
rect 4150 3108 4178 3164
rect 4234 3108 4282 3164
rect 4338 3108 4386 3164
rect 4442 3108 4470 3164
rect 4150 1596 4470 3108
rect 4150 1540 4178 1596
rect 4234 1540 4282 1596
rect 4338 1540 4386 1596
rect 4442 1540 4470 1596
rect 4150 1508 4470 1540
rect 5745 11788 6065 11820
rect 5745 11732 5773 11788
rect 5829 11732 5877 11788
rect 5933 11732 5981 11788
rect 6037 11732 6065 11788
rect 5745 11206 6065 11732
rect 5745 11150 5773 11206
rect 5829 11150 5877 11206
rect 5933 11150 5981 11206
rect 6037 11150 6065 11206
rect 5745 11102 6065 11150
rect 5745 11046 5773 11102
rect 5829 11046 5877 11102
rect 5933 11046 5981 11102
rect 6037 11046 6065 11102
rect 5745 10998 6065 11046
rect 5745 10942 5773 10998
rect 5829 10942 5877 10998
rect 5933 10942 5981 10998
rect 6037 10942 6065 10998
rect 5745 10220 6065 10942
rect 5745 10164 5773 10220
rect 5829 10164 5877 10220
rect 5933 10164 5981 10220
rect 6037 10164 6065 10220
rect 5745 8652 6065 10164
rect 5745 8596 5773 8652
rect 5829 8596 5877 8652
rect 5933 8596 5981 8652
rect 6037 8596 6065 8652
rect 5745 8490 6065 8596
rect 5745 8434 5773 8490
rect 5829 8434 5877 8490
rect 5933 8434 5981 8490
rect 6037 8434 6065 8490
rect 5745 8386 6065 8434
rect 5745 8330 5773 8386
rect 5829 8330 5877 8386
rect 5933 8330 5981 8386
rect 6037 8330 6065 8386
rect 5745 8282 6065 8330
rect 5745 8226 5773 8282
rect 5829 8226 5877 8282
rect 5933 8226 5981 8282
rect 6037 8226 6065 8282
rect 5745 7084 6065 8226
rect 5745 7028 5773 7084
rect 5829 7028 5877 7084
rect 5933 7028 5981 7084
rect 6037 7028 6065 7084
rect 5745 5774 6065 7028
rect 5745 5718 5773 5774
rect 5829 5718 5877 5774
rect 5933 5718 5981 5774
rect 6037 5718 6065 5774
rect 5745 5670 6065 5718
rect 5745 5614 5773 5670
rect 5829 5614 5877 5670
rect 5933 5614 5981 5670
rect 6037 5614 6065 5670
rect 5745 5566 6065 5614
rect 5745 5460 5773 5566
rect 5829 5460 5877 5566
rect 5933 5460 5981 5566
rect 6037 5460 6065 5566
rect 5745 3948 6065 5460
rect 5745 3892 5773 3948
rect 5829 3892 5877 3948
rect 5933 3892 5981 3948
rect 6037 3892 6065 3948
rect 5745 3058 6065 3892
rect 5745 3002 5773 3058
rect 5829 3002 5877 3058
rect 5933 3002 5981 3058
rect 6037 3002 6065 3058
rect 5745 2954 6065 3002
rect 5745 2898 5773 2954
rect 5829 2898 5877 2954
rect 5933 2898 5981 2954
rect 6037 2898 6065 2954
rect 5745 2850 6065 2898
rect 5745 2794 5773 2850
rect 5829 2794 5877 2850
rect 5933 2794 5981 2850
rect 6037 2794 6065 2850
rect 5745 2380 6065 2794
rect 5745 2324 5773 2380
rect 5829 2324 5877 2380
rect 5933 2324 5981 2380
rect 6037 2324 6065 2380
rect 5745 1508 6065 2324
rect 7340 11004 7660 11820
rect 7340 10948 7368 11004
rect 7424 10948 7472 11004
rect 7528 10948 7576 11004
rect 7632 10948 7660 11004
rect 7340 9848 7660 10948
rect 7340 9792 7368 9848
rect 7424 9792 7472 9848
rect 7528 9792 7576 9848
rect 7632 9792 7660 9848
rect 7340 9744 7660 9792
rect 7340 9688 7368 9744
rect 7424 9688 7472 9744
rect 7528 9688 7576 9744
rect 7632 9688 7660 9744
rect 7340 9640 7660 9688
rect 7340 9584 7368 9640
rect 7424 9584 7472 9640
rect 7528 9584 7576 9640
rect 7632 9584 7660 9640
rect 7340 9436 7660 9584
rect 7340 9380 7368 9436
rect 7424 9380 7472 9436
rect 7528 9380 7576 9436
rect 7632 9380 7660 9436
rect 7340 7868 7660 9380
rect 7340 7812 7368 7868
rect 7424 7812 7472 7868
rect 7528 7812 7576 7868
rect 7632 7812 7660 7868
rect 7340 7132 7660 7812
rect 7340 7076 7368 7132
rect 7424 7076 7472 7132
rect 7528 7076 7576 7132
rect 7632 7076 7660 7132
rect 7340 7028 7660 7076
rect 7340 6972 7368 7028
rect 7424 6972 7472 7028
rect 7528 6972 7576 7028
rect 7632 6972 7660 7028
rect 7340 6924 7660 6972
rect 7340 6868 7368 6924
rect 7424 6868 7472 6924
rect 7528 6868 7576 6924
rect 7632 6868 7660 6924
rect 7340 6300 7660 6868
rect 7340 6244 7368 6300
rect 7424 6244 7472 6300
rect 7528 6244 7576 6300
rect 7632 6244 7660 6300
rect 7340 4732 7660 6244
rect 7340 4676 7368 4732
rect 7424 4676 7472 4732
rect 7528 4676 7576 4732
rect 7632 4676 7660 4732
rect 7340 4416 7660 4676
rect 7340 4360 7368 4416
rect 7424 4360 7472 4416
rect 7528 4360 7576 4416
rect 7632 4360 7660 4416
rect 7340 4312 7660 4360
rect 7340 4256 7368 4312
rect 7424 4256 7472 4312
rect 7528 4256 7576 4312
rect 7632 4256 7660 4312
rect 7340 4208 7660 4256
rect 7340 4152 7368 4208
rect 7424 4152 7472 4208
rect 7528 4152 7576 4208
rect 7632 4152 7660 4208
rect 7340 3164 7660 4152
rect 7340 3108 7368 3164
rect 7424 3108 7472 3164
rect 7528 3108 7576 3164
rect 7632 3108 7660 3164
rect 7340 1596 7660 3108
rect 7340 1540 7368 1596
rect 7424 1540 7472 1596
rect 7528 1540 7576 1596
rect 7632 1540 7660 1596
rect 7340 1508 7660 1540
rect 8935 11788 9255 11820
rect 8935 11732 8963 11788
rect 9019 11732 9067 11788
rect 9123 11732 9171 11788
rect 9227 11732 9255 11788
rect 8935 11206 9255 11732
rect 8935 11150 8963 11206
rect 9019 11150 9067 11206
rect 9123 11150 9171 11206
rect 9227 11150 9255 11206
rect 8935 11102 9255 11150
rect 8935 11046 8963 11102
rect 9019 11046 9067 11102
rect 9123 11046 9171 11102
rect 9227 11046 9255 11102
rect 8935 10998 9255 11046
rect 8935 10942 8963 10998
rect 9019 10942 9067 10998
rect 9123 10942 9171 10998
rect 9227 10942 9255 10998
rect 8935 10220 9255 10942
rect 8935 10164 8963 10220
rect 9019 10164 9067 10220
rect 9123 10164 9171 10220
rect 9227 10164 9255 10220
rect 8935 8652 9255 10164
rect 8935 8596 8963 8652
rect 9019 8596 9067 8652
rect 9123 8596 9171 8652
rect 9227 8596 9255 8652
rect 8935 8490 9255 8596
rect 8935 8434 8963 8490
rect 9019 8434 9067 8490
rect 9123 8434 9171 8490
rect 9227 8434 9255 8490
rect 8935 8386 9255 8434
rect 8935 8330 8963 8386
rect 9019 8330 9067 8386
rect 9123 8330 9171 8386
rect 9227 8330 9255 8386
rect 8935 8282 9255 8330
rect 8935 8226 8963 8282
rect 9019 8226 9067 8282
rect 9123 8226 9171 8282
rect 9227 8226 9255 8282
rect 8935 7084 9255 8226
rect 8935 7028 8963 7084
rect 9019 7028 9067 7084
rect 9123 7028 9171 7084
rect 9227 7028 9255 7084
rect 8935 5774 9255 7028
rect 8935 5718 8963 5774
rect 9019 5718 9067 5774
rect 9123 5718 9171 5774
rect 9227 5718 9255 5774
rect 8935 5670 9255 5718
rect 8935 5614 8963 5670
rect 9019 5614 9067 5670
rect 9123 5614 9171 5670
rect 9227 5614 9255 5670
rect 8935 5566 9255 5614
rect 8935 5460 8963 5566
rect 9019 5460 9067 5566
rect 9123 5460 9171 5566
rect 9227 5460 9255 5566
rect 8935 3948 9255 5460
rect 8935 3892 8963 3948
rect 9019 3892 9067 3948
rect 9123 3892 9171 3948
rect 9227 3892 9255 3948
rect 8935 3058 9255 3892
rect 8935 3002 8963 3058
rect 9019 3002 9067 3058
rect 9123 3002 9171 3058
rect 9227 3002 9255 3058
rect 8935 2954 9255 3002
rect 8935 2898 8963 2954
rect 9019 2898 9067 2954
rect 9123 2898 9171 2954
rect 9227 2898 9255 2954
rect 8935 2850 9255 2898
rect 8935 2794 8963 2850
rect 9019 2794 9067 2850
rect 9123 2794 9171 2850
rect 9227 2794 9255 2850
rect 8935 2380 9255 2794
rect 8935 2324 8963 2380
rect 9019 2324 9067 2380
rect 9123 2324 9171 2380
rect 9227 2324 9255 2380
rect 8935 1508 9255 2324
rect 10530 11004 10850 11820
rect 10530 10948 10558 11004
rect 10614 10948 10662 11004
rect 10718 10948 10766 11004
rect 10822 10948 10850 11004
rect 10530 9848 10850 10948
rect 10530 9792 10558 9848
rect 10614 9792 10662 9848
rect 10718 9792 10766 9848
rect 10822 9792 10850 9848
rect 10530 9744 10850 9792
rect 10530 9688 10558 9744
rect 10614 9688 10662 9744
rect 10718 9688 10766 9744
rect 10822 9688 10850 9744
rect 10530 9640 10850 9688
rect 10530 9584 10558 9640
rect 10614 9584 10662 9640
rect 10718 9584 10766 9640
rect 10822 9584 10850 9640
rect 10530 9436 10850 9584
rect 10530 9380 10558 9436
rect 10614 9380 10662 9436
rect 10718 9380 10766 9436
rect 10822 9380 10850 9436
rect 10530 7868 10850 9380
rect 10530 7812 10558 7868
rect 10614 7812 10662 7868
rect 10718 7812 10766 7868
rect 10822 7812 10850 7868
rect 10530 7132 10850 7812
rect 10530 7076 10558 7132
rect 10614 7076 10662 7132
rect 10718 7076 10766 7132
rect 10822 7076 10850 7132
rect 10530 7028 10850 7076
rect 10530 6972 10558 7028
rect 10614 6972 10662 7028
rect 10718 6972 10766 7028
rect 10822 6972 10850 7028
rect 10530 6924 10850 6972
rect 10530 6868 10558 6924
rect 10614 6868 10662 6924
rect 10718 6868 10766 6924
rect 10822 6868 10850 6924
rect 10530 6300 10850 6868
rect 10530 6244 10558 6300
rect 10614 6244 10662 6300
rect 10718 6244 10766 6300
rect 10822 6244 10850 6300
rect 10530 4732 10850 6244
rect 10530 4676 10558 4732
rect 10614 4676 10662 4732
rect 10718 4676 10766 4732
rect 10822 4676 10850 4732
rect 10530 4416 10850 4676
rect 10530 4360 10558 4416
rect 10614 4360 10662 4416
rect 10718 4360 10766 4416
rect 10822 4360 10850 4416
rect 10530 4312 10850 4360
rect 10530 4256 10558 4312
rect 10614 4256 10662 4312
rect 10718 4256 10766 4312
rect 10822 4256 10850 4312
rect 10530 4208 10850 4256
rect 10530 4152 10558 4208
rect 10614 4152 10662 4208
rect 10718 4152 10766 4208
rect 10822 4152 10850 4208
rect 10530 3164 10850 4152
rect 10530 3108 10558 3164
rect 10614 3108 10662 3164
rect 10718 3108 10766 3164
rect 10822 3108 10850 3164
rect 10530 1596 10850 3108
rect 10530 1540 10558 1596
rect 10614 1540 10662 1596
rect 10718 1540 10766 1596
rect 10822 1540 10850 1596
rect 10530 1508 10850 1540
rect 12125 11788 12445 11820
rect 12125 11732 12153 11788
rect 12209 11732 12257 11788
rect 12313 11732 12361 11788
rect 12417 11732 12445 11788
rect 12125 11206 12445 11732
rect 12125 11150 12153 11206
rect 12209 11150 12257 11206
rect 12313 11150 12361 11206
rect 12417 11150 12445 11206
rect 12125 11102 12445 11150
rect 12125 11046 12153 11102
rect 12209 11046 12257 11102
rect 12313 11046 12361 11102
rect 12417 11046 12445 11102
rect 12125 10998 12445 11046
rect 12125 10942 12153 10998
rect 12209 10942 12257 10998
rect 12313 10942 12361 10998
rect 12417 10942 12445 10998
rect 12125 10220 12445 10942
rect 12125 10164 12153 10220
rect 12209 10164 12257 10220
rect 12313 10164 12361 10220
rect 12417 10164 12445 10220
rect 12125 8652 12445 10164
rect 12125 8596 12153 8652
rect 12209 8596 12257 8652
rect 12313 8596 12361 8652
rect 12417 8596 12445 8652
rect 12125 8490 12445 8596
rect 12125 8434 12153 8490
rect 12209 8434 12257 8490
rect 12313 8434 12361 8490
rect 12417 8434 12445 8490
rect 12125 8386 12445 8434
rect 12125 8330 12153 8386
rect 12209 8330 12257 8386
rect 12313 8330 12361 8386
rect 12417 8330 12445 8386
rect 12125 8282 12445 8330
rect 12125 8226 12153 8282
rect 12209 8226 12257 8282
rect 12313 8226 12361 8282
rect 12417 8226 12445 8282
rect 12125 7084 12445 8226
rect 12125 7028 12153 7084
rect 12209 7028 12257 7084
rect 12313 7028 12361 7084
rect 12417 7028 12445 7084
rect 12125 5774 12445 7028
rect 12125 5718 12153 5774
rect 12209 5718 12257 5774
rect 12313 5718 12361 5774
rect 12417 5718 12445 5774
rect 12125 5670 12445 5718
rect 12125 5614 12153 5670
rect 12209 5614 12257 5670
rect 12313 5614 12361 5670
rect 12417 5614 12445 5670
rect 12125 5566 12445 5614
rect 12125 5460 12153 5566
rect 12209 5460 12257 5566
rect 12313 5460 12361 5566
rect 12417 5460 12445 5566
rect 12125 3948 12445 5460
rect 12125 3892 12153 3948
rect 12209 3892 12257 3948
rect 12313 3892 12361 3948
rect 12417 3892 12445 3948
rect 12125 3058 12445 3892
rect 12125 3002 12153 3058
rect 12209 3002 12257 3058
rect 12313 3002 12361 3058
rect 12417 3002 12445 3058
rect 12125 2954 12445 3002
rect 12125 2898 12153 2954
rect 12209 2898 12257 2954
rect 12313 2898 12361 2954
rect 12417 2898 12445 2954
rect 12125 2850 12445 2898
rect 12125 2794 12153 2850
rect 12209 2794 12257 2850
rect 12313 2794 12361 2850
rect 12417 2794 12445 2850
rect 12125 2380 12445 2794
rect 12125 2324 12153 2380
rect 12209 2324 12257 2380
rect 12313 2324 12361 2380
rect 12417 2324 12445 2380
rect 12125 1508 12445 2324
<< via4 >>
rect 2583 11150 2639 11206
rect 2687 11150 2743 11206
rect 2791 11150 2847 11206
rect 2583 11046 2639 11102
rect 2687 11046 2743 11102
rect 2791 11046 2847 11102
rect 2583 10942 2639 10998
rect 2687 10942 2743 10998
rect 2791 10942 2847 10998
rect 2583 8434 2639 8490
rect 2687 8434 2743 8490
rect 2791 8434 2847 8490
rect 2583 8330 2639 8386
rect 2687 8330 2743 8386
rect 2791 8330 2847 8386
rect 2583 8226 2639 8282
rect 2687 8226 2743 8282
rect 2791 8226 2847 8282
rect 2583 5718 2639 5774
rect 2687 5718 2743 5774
rect 2791 5718 2847 5774
rect 2583 5614 2639 5670
rect 2687 5614 2743 5670
rect 2791 5614 2847 5670
rect 2583 5516 2639 5566
rect 2583 5510 2639 5516
rect 2687 5516 2743 5566
rect 2687 5510 2743 5516
rect 2791 5516 2847 5566
rect 2791 5510 2847 5516
rect 2583 3002 2639 3058
rect 2687 3002 2743 3058
rect 2791 3002 2847 3058
rect 2583 2898 2639 2954
rect 2687 2898 2743 2954
rect 2791 2898 2847 2954
rect 2583 2794 2639 2850
rect 2687 2794 2743 2850
rect 2791 2794 2847 2850
rect 4178 9792 4234 9848
rect 4282 9792 4338 9848
rect 4386 9792 4442 9848
rect 4178 9688 4234 9744
rect 4282 9688 4338 9744
rect 4386 9688 4442 9744
rect 4178 9584 4234 9640
rect 4282 9584 4338 9640
rect 4386 9584 4442 9640
rect 4178 7076 4234 7132
rect 4282 7076 4338 7132
rect 4386 7076 4442 7132
rect 4178 6972 4234 7028
rect 4282 6972 4338 7028
rect 4386 6972 4442 7028
rect 4178 6868 4234 6924
rect 4282 6868 4338 6924
rect 4386 6868 4442 6924
rect 4178 4360 4234 4416
rect 4282 4360 4338 4416
rect 4386 4360 4442 4416
rect 4178 4256 4234 4312
rect 4282 4256 4338 4312
rect 4386 4256 4442 4312
rect 4178 4152 4234 4208
rect 4282 4152 4338 4208
rect 4386 4152 4442 4208
rect 5773 11150 5829 11206
rect 5877 11150 5933 11206
rect 5981 11150 6037 11206
rect 5773 11046 5829 11102
rect 5877 11046 5933 11102
rect 5981 11046 6037 11102
rect 5773 10942 5829 10998
rect 5877 10942 5933 10998
rect 5981 10942 6037 10998
rect 5773 8434 5829 8490
rect 5877 8434 5933 8490
rect 5981 8434 6037 8490
rect 5773 8330 5829 8386
rect 5877 8330 5933 8386
rect 5981 8330 6037 8386
rect 5773 8226 5829 8282
rect 5877 8226 5933 8282
rect 5981 8226 6037 8282
rect 5773 5718 5829 5774
rect 5877 5718 5933 5774
rect 5981 5718 6037 5774
rect 5773 5614 5829 5670
rect 5877 5614 5933 5670
rect 5981 5614 6037 5670
rect 5773 5516 5829 5566
rect 5773 5510 5829 5516
rect 5877 5516 5933 5566
rect 5877 5510 5933 5516
rect 5981 5516 6037 5566
rect 5981 5510 6037 5516
rect 5773 3002 5829 3058
rect 5877 3002 5933 3058
rect 5981 3002 6037 3058
rect 5773 2898 5829 2954
rect 5877 2898 5933 2954
rect 5981 2898 6037 2954
rect 5773 2794 5829 2850
rect 5877 2794 5933 2850
rect 5981 2794 6037 2850
rect 7368 9792 7424 9848
rect 7472 9792 7528 9848
rect 7576 9792 7632 9848
rect 7368 9688 7424 9744
rect 7472 9688 7528 9744
rect 7576 9688 7632 9744
rect 7368 9584 7424 9640
rect 7472 9584 7528 9640
rect 7576 9584 7632 9640
rect 7368 7076 7424 7132
rect 7472 7076 7528 7132
rect 7576 7076 7632 7132
rect 7368 6972 7424 7028
rect 7472 6972 7528 7028
rect 7576 6972 7632 7028
rect 7368 6868 7424 6924
rect 7472 6868 7528 6924
rect 7576 6868 7632 6924
rect 7368 4360 7424 4416
rect 7472 4360 7528 4416
rect 7576 4360 7632 4416
rect 7368 4256 7424 4312
rect 7472 4256 7528 4312
rect 7576 4256 7632 4312
rect 7368 4152 7424 4208
rect 7472 4152 7528 4208
rect 7576 4152 7632 4208
rect 8963 11150 9019 11206
rect 9067 11150 9123 11206
rect 9171 11150 9227 11206
rect 8963 11046 9019 11102
rect 9067 11046 9123 11102
rect 9171 11046 9227 11102
rect 8963 10942 9019 10998
rect 9067 10942 9123 10998
rect 9171 10942 9227 10998
rect 8963 8434 9019 8490
rect 9067 8434 9123 8490
rect 9171 8434 9227 8490
rect 8963 8330 9019 8386
rect 9067 8330 9123 8386
rect 9171 8330 9227 8386
rect 8963 8226 9019 8282
rect 9067 8226 9123 8282
rect 9171 8226 9227 8282
rect 8963 5718 9019 5774
rect 9067 5718 9123 5774
rect 9171 5718 9227 5774
rect 8963 5614 9019 5670
rect 9067 5614 9123 5670
rect 9171 5614 9227 5670
rect 8963 5516 9019 5566
rect 8963 5510 9019 5516
rect 9067 5516 9123 5566
rect 9067 5510 9123 5516
rect 9171 5516 9227 5566
rect 9171 5510 9227 5516
rect 8963 3002 9019 3058
rect 9067 3002 9123 3058
rect 9171 3002 9227 3058
rect 8963 2898 9019 2954
rect 9067 2898 9123 2954
rect 9171 2898 9227 2954
rect 8963 2794 9019 2850
rect 9067 2794 9123 2850
rect 9171 2794 9227 2850
rect 10558 9792 10614 9848
rect 10662 9792 10718 9848
rect 10766 9792 10822 9848
rect 10558 9688 10614 9744
rect 10662 9688 10718 9744
rect 10766 9688 10822 9744
rect 10558 9584 10614 9640
rect 10662 9584 10718 9640
rect 10766 9584 10822 9640
rect 10558 7076 10614 7132
rect 10662 7076 10718 7132
rect 10766 7076 10822 7132
rect 10558 6972 10614 7028
rect 10662 6972 10718 7028
rect 10766 6972 10822 7028
rect 10558 6868 10614 6924
rect 10662 6868 10718 6924
rect 10766 6868 10822 6924
rect 10558 4360 10614 4416
rect 10662 4360 10718 4416
rect 10766 4360 10822 4416
rect 10558 4256 10614 4312
rect 10662 4256 10718 4312
rect 10766 4256 10822 4312
rect 10558 4152 10614 4208
rect 10662 4152 10718 4208
rect 10766 4152 10822 4208
rect 12153 11150 12209 11206
rect 12257 11150 12313 11206
rect 12361 11150 12417 11206
rect 12153 11046 12209 11102
rect 12257 11046 12313 11102
rect 12361 11046 12417 11102
rect 12153 10942 12209 10998
rect 12257 10942 12313 10998
rect 12361 10942 12417 10998
rect 12153 8434 12209 8490
rect 12257 8434 12313 8490
rect 12361 8434 12417 8490
rect 12153 8330 12209 8386
rect 12257 8330 12313 8386
rect 12361 8330 12417 8386
rect 12153 8226 12209 8282
rect 12257 8226 12313 8282
rect 12361 8226 12417 8282
rect 12153 5718 12209 5774
rect 12257 5718 12313 5774
rect 12361 5718 12417 5774
rect 12153 5614 12209 5670
rect 12257 5614 12313 5670
rect 12361 5614 12417 5670
rect 12153 5516 12209 5566
rect 12153 5510 12209 5516
rect 12257 5516 12313 5566
rect 12257 5510 12313 5516
rect 12361 5516 12417 5566
rect 12361 5510 12417 5516
rect 12153 3002 12209 3058
rect 12257 3002 12313 3058
rect 12361 3002 12417 3058
rect 12153 2898 12209 2954
rect 12257 2898 12313 2954
rect 12361 2898 12417 2954
rect 12153 2794 12209 2850
rect 12257 2794 12313 2850
rect 12361 2794 12417 2850
<< metal5 >>
rect 1060 11206 13836 11234
rect 1060 11150 2583 11206
rect 2639 11150 2687 11206
rect 2743 11150 2791 11206
rect 2847 11150 5773 11206
rect 5829 11150 5877 11206
rect 5933 11150 5981 11206
rect 6037 11150 8963 11206
rect 9019 11150 9067 11206
rect 9123 11150 9171 11206
rect 9227 11150 12153 11206
rect 12209 11150 12257 11206
rect 12313 11150 12361 11206
rect 12417 11150 13836 11206
rect 1060 11102 13836 11150
rect 1060 11046 2583 11102
rect 2639 11046 2687 11102
rect 2743 11046 2791 11102
rect 2847 11046 5773 11102
rect 5829 11046 5877 11102
rect 5933 11046 5981 11102
rect 6037 11046 8963 11102
rect 9019 11046 9067 11102
rect 9123 11046 9171 11102
rect 9227 11046 12153 11102
rect 12209 11046 12257 11102
rect 12313 11046 12361 11102
rect 12417 11046 13836 11102
rect 1060 10998 13836 11046
rect 1060 10942 2583 10998
rect 2639 10942 2687 10998
rect 2743 10942 2791 10998
rect 2847 10942 5773 10998
rect 5829 10942 5877 10998
rect 5933 10942 5981 10998
rect 6037 10942 8963 10998
rect 9019 10942 9067 10998
rect 9123 10942 9171 10998
rect 9227 10942 12153 10998
rect 12209 10942 12257 10998
rect 12313 10942 12361 10998
rect 12417 10942 13836 10998
rect 1060 10914 13836 10942
rect 1060 9848 13836 9876
rect 1060 9792 4178 9848
rect 4234 9792 4282 9848
rect 4338 9792 4386 9848
rect 4442 9792 7368 9848
rect 7424 9792 7472 9848
rect 7528 9792 7576 9848
rect 7632 9792 10558 9848
rect 10614 9792 10662 9848
rect 10718 9792 10766 9848
rect 10822 9792 13836 9848
rect 1060 9744 13836 9792
rect 1060 9688 4178 9744
rect 4234 9688 4282 9744
rect 4338 9688 4386 9744
rect 4442 9688 7368 9744
rect 7424 9688 7472 9744
rect 7528 9688 7576 9744
rect 7632 9688 10558 9744
rect 10614 9688 10662 9744
rect 10718 9688 10766 9744
rect 10822 9688 13836 9744
rect 1060 9640 13836 9688
rect 1060 9584 4178 9640
rect 4234 9584 4282 9640
rect 4338 9584 4386 9640
rect 4442 9584 7368 9640
rect 7424 9584 7472 9640
rect 7528 9584 7576 9640
rect 7632 9584 10558 9640
rect 10614 9584 10662 9640
rect 10718 9584 10766 9640
rect 10822 9584 13836 9640
rect 1060 9556 13836 9584
rect 1060 8490 13836 8518
rect 1060 8434 2583 8490
rect 2639 8434 2687 8490
rect 2743 8434 2791 8490
rect 2847 8434 5773 8490
rect 5829 8434 5877 8490
rect 5933 8434 5981 8490
rect 6037 8434 8963 8490
rect 9019 8434 9067 8490
rect 9123 8434 9171 8490
rect 9227 8434 12153 8490
rect 12209 8434 12257 8490
rect 12313 8434 12361 8490
rect 12417 8434 13836 8490
rect 1060 8386 13836 8434
rect 1060 8330 2583 8386
rect 2639 8330 2687 8386
rect 2743 8330 2791 8386
rect 2847 8330 5773 8386
rect 5829 8330 5877 8386
rect 5933 8330 5981 8386
rect 6037 8330 8963 8386
rect 9019 8330 9067 8386
rect 9123 8330 9171 8386
rect 9227 8330 12153 8386
rect 12209 8330 12257 8386
rect 12313 8330 12361 8386
rect 12417 8330 13836 8386
rect 1060 8282 13836 8330
rect 1060 8226 2583 8282
rect 2639 8226 2687 8282
rect 2743 8226 2791 8282
rect 2847 8226 5773 8282
rect 5829 8226 5877 8282
rect 5933 8226 5981 8282
rect 6037 8226 8963 8282
rect 9019 8226 9067 8282
rect 9123 8226 9171 8282
rect 9227 8226 12153 8282
rect 12209 8226 12257 8282
rect 12313 8226 12361 8282
rect 12417 8226 13836 8282
rect 1060 8198 13836 8226
rect 1060 7132 13836 7160
rect 1060 7076 4178 7132
rect 4234 7076 4282 7132
rect 4338 7076 4386 7132
rect 4442 7076 7368 7132
rect 7424 7076 7472 7132
rect 7528 7076 7576 7132
rect 7632 7076 10558 7132
rect 10614 7076 10662 7132
rect 10718 7076 10766 7132
rect 10822 7076 13836 7132
rect 1060 7028 13836 7076
rect 1060 6972 4178 7028
rect 4234 6972 4282 7028
rect 4338 6972 4386 7028
rect 4442 6972 7368 7028
rect 7424 6972 7472 7028
rect 7528 6972 7576 7028
rect 7632 6972 10558 7028
rect 10614 6972 10662 7028
rect 10718 6972 10766 7028
rect 10822 6972 13836 7028
rect 1060 6924 13836 6972
rect 1060 6868 4178 6924
rect 4234 6868 4282 6924
rect 4338 6868 4386 6924
rect 4442 6868 7368 6924
rect 7424 6868 7472 6924
rect 7528 6868 7576 6924
rect 7632 6868 10558 6924
rect 10614 6868 10662 6924
rect 10718 6868 10766 6924
rect 10822 6868 13836 6924
rect 1060 6840 13836 6868
rect 1060 5774 13836 5802
rect 1060 5718 2583 5774
rect 2639 5718 2687 5774
rect 2743 5718 2791 5774
rect 2847 5718 5773 5774
rect 5829 5718 5877 5774
rect 5933 5718 5981 5774
rect 6037 5718 8963 5774
rect 9019 5718 9067 5774
rect 9123 5718 9171 5774
rect 9227 5718 12153 5774
rect 12209 5718 12257 5774
rect 12313 5718 12361 5774
rect 12417 5718 13836 5774
rect 1060 5670 13836 5718
rect 1060 5614 2583 5670
rect 2639 5614 2687 5670
rect 2743 5614 2791 5670
rect 2847 5614 5773 5670
rect 5829 5614 5877 5670
rect 5933 5614 5981 5670
rect 6037 5614 8963 5670
rect 9019 5614 9067 5670
rect 9123 5614 9171 5670
rect 9227 5614 12153 5670
rect 12209 5614 12257 5670
rect 12313 5614 12361 5670
rect 12417 5614 13836 5670
rect 1060 5566 13836 5614
rect 1060 5510 2583 5566
rect 2639 5510 2687 5566
rect 2743 5510 2791 5566
rect 2847 5510 5773 5566
rect 5829 5510 5877 5566
rect 5933 5510 5981 5566
rect 6037 5510 8963 5566
rect 9019 5510 9067 5566
rect 9123 5510 9171 5566
rect 9227 5510 12153 5566
rect 12209 5510 12257 5566
rect 12313 5510 12361 5566
rect 12417 5510 13836 5566
rect 1060 5482 13836 5510
rect 1060 4416 13836 4444
rect 1060 4360 4178 4416
rect 4234 4360 4282 4416
rect 4338 4360 4386 4416
rect 4442 4360 7368 4416
rect 7424 4360 7472 4416
rect 7528 4360 7576 4416
rect 7632 4360 10558 4416
rect 10614 4360 10662 4416
rect 10718 4360 10766 4416
rect 10822 4360 13836 4416
rect 1060 4312 13836 4360
rect 1060 4256 4178 4312
rect 4234 4256 4282 4312
rect 4338 4256 4386 4312
rect 4442 4256 7368 4312
rect 7424 4256 7472 4312
rect 7528 4256 7576 4312
rect 7632 4256 10558 4312
rect 10614 4256 10662 4312
rect 10718 4256 10766 4312
rect 10822 4256 13836 4312
rect 1060 4208 13836 4256
rect 1060 4152 4178 4208
rect 4234 4152 4282 4208
rect 4338 4152 4386 4208
rect 4442 4152 7368 4208
rect 7424 4152 7472 4208
rect 7528 4152 7576 4208
rect 7632 4152 10558 4208
rect 10614 4152 10662 4208
rect 10718 4152 10766 4208
rect 10822 4152 13836 4208
rect 1060 4124 13836 4152
rect 1060 3058 13836 3086
rect 1060 3002 2583 3058
rect 2639 3002 2687 3058
rect 2743 3002 2791 3058
rect 2847 3002 5773 3058
rect 5829 3002 5877 3058
rect 5933 3002 5981 3058
rect 6037 3002 8963 3058
rect 9019 3002 9067 3058
rect 9123 3002 9171 3058
rect 9227 3002 12153 3058
rect 12209 3002 12257 3058
rect 12313 3002 12361 3058
rect 12417 3002 13836 3058
rect 1060 2954 13836 3002
rect 1060 2898 2583 2954
rect 2639 2898 2687 2954
rect 2743 2898 2791 2954
rect 2847 2898 5773 2954
rect 5829 2898 5877 2954
rect 5933 2898 5981 2954
rect 6037 2898 8963 2954
rect 9019 2898 9067 2954
rect 9123 2898 9171 2954
rect 9227 2898 12153 2954
rect 12209 2898 12257 2954
rect 12313 2898 12361 2954
rect 12417 2898 13836 2954
rect 1060 2850 13836 2898
rect 1060 2794 2583 2850
rect 2639 2794 2687 2850
rect 2743 2794 2791 2850
rect 2847 2794 5773 2850
rect 5829 2794 5877 2850
rect 5933 2794 5981 2850
rect 6037 2794 8963 2850
rect 9019 2794 9067 2850
rect 9123 2794 9171 2850
rect 9227 2794 12153 2850
rect 12209 2794 12257 2850
rect 12313 2794 12361 2850
rect 12417 2794 13836 2850
rect 1060 2766 13836 2794
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 1344 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_10 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 2240 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 2912 0 1 1568
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28
timestamp 1654395037
transform 1 0 4256 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_32
timestamp 1654395037
transform 1 0 4704 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 4928 0 1 1568
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_41
timestamp 1654395037
transform 1 0 5712 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47
timestamp 1654395037
transform 1 0 6384 0 1 1568
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_55
timestamp 1654395037
transform 1 0 7280 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63
timestamp 1654395037
transform 1 0 8176 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_0_67
timestamp 1654395037
transform 1 0 8624 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1654395037
transform 1 0 8848 0 1 1568
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 9632 0 1 1568
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92
timestamp 1654395037
transform 1 0 11424 0 1 1568
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100
timestamp 1654395037
transform 1 0 12320 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1654395037
transform 1 0 12768 0 1 1568
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107
timestamp 1654395037
transform 1 0 13104 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_2
timestamp 1654395037
transform 1 0 1344 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_4
timestamp 1654395037
transform 1 0 1568 0 -1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_46
timestamp 1654395037
transform 1 0 6272 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_50
timestamp 1654395037
transform 1 0 6720 0 -1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_55
timestamp 1654395037
transform 1 0 7280 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1654395037
transform 1 0 8512 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1654395037
transform 1 0 8960 0 -1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_1_77
timestamp 1654395037
transform 1 0 9744 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_83
timestamp 1654395037
transform 1 0 10416 0 -1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_99
timestamp 1654395037
transform 1 0 12208 0 -1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_107
timestamp 1654395037
transform 1 0 13104 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_2
timestamp 1654395037
transform 1 0 1344 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_6
timestamp 1654395037
transform 1 0 1792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_8
timestamp 1654395037
transform 1 0 2016 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_19
timestamp 1654395037
transform 1 0 3248 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_37
timestamp 1654395037
transform 1 0 5264 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_41
timestamp 1654395037
transform 1 0 5712 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_46
timestamp 1654395037
transform 1 0 6272 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_50
timestamp 1654395037
transform 1 0 6720 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_52
timestamp 1654395037
transform 1 0 6944 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_57
timestamp 1654395037
transform 1 0 7504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_100
timestamp 1654395037
transform 1 0 12320 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_104
timestamp 1654395037
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_2_108
timestamp 1654395037
transform 1 0 13216 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_110
timestamp 1654395037
transform 1 0 13440 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_2
timestamp 1654395037
transform 1 0 1344 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_6
timestamp 1654395037
transform 1 0 1792 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_12 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 2464 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_44
timestamp 1654395037
transform 1 0 6048 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_60
timestamp 1654395037
transform 1 0 7840 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_68
timestamp 1654395037
transform 1 0 8736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1654395037
transform 1 0 8960 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_73
timestamp 1654395037
transform 1 0 9296 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_81
timestamp 1654395037
transform 1 0 10192 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_87
timestamp 1654395037
transform 1 0 10864 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_95
timestamp 1654395037
transform 1 0 11760 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_99
timestamp 1654395037
transform 1 0 12208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_105
timestamp 1654395037
transform 1 0 12880 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_3_109
timestamp 1654395037
transform 1 0 13328 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_2
timestamp 1654395037
transform 1 0 1344 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_10
timestamp 1654395037
transform 1 0 2240 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_14
timestamp 1654395037
transform 1 0 2688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_16
timestamp 1654395037
transform 1 0 2912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_21
timestamp 1654395037
transform 1 0 3472 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_29
timestamp 1654395037
transform 1 0 4368 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_33
timestamp 1654395037
transform 1 0 4816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 5264 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1654395037
transform 1 0 12432 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1654395037
transform 1 0 12880 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_4_108
timestamp 1654395037
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_110
timestamp 1654395037
transform 1 0 13440 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_2
timestamp 1654395037
transform 1 0 1344 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_34
timestamp 1654395037
transform 1 0 4928 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_56
timestamp 1654395037
transform 1 0 7392 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_64
timestamp 1654395037
transform 1 0 8288 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_68
timestamp 1654395037
transform 1 0 8736 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1654395037
transform 1 0 8960 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_73
timestamp 1654395037
transform 1 0 9296 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_105
timestamp 1654395037
transform 1 0 12880 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_5_109
timestamp 1654395037
transform 1 0 13328 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1654395037
transform 1 0 1344 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1654395037
transform 1 0 4928 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_37
timestamp 1654395037
transform 1 0 5264 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_45
timestamp 1654395037
transform 1 0 6160 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_72
timestamp 1654395037
transform 1 0 9184 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_104
timestamp 1654395037
transform 1 0 12768 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_6_108
timestamp 1654395037
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_110
timestamp 1654395037
transform 1 0 13440 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_2
timestamp 1654395037
transform 1 0 1344 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_34
timestamp 1654395037
transform 1 0 4928 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_7_38
timestamp 1654395037
transform 1 0 5376 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_7_44
timestamp 1654395037
transform 1 0 6048 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_50
timestamp 1654395037
transform 1 0 6720 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_7_54
timestamp 1654395037
transform 1 0 7168 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_56
timestamp 1654395037
transform 1 0 7392 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_61
timestamp 1654395037
transform 1 0 7952 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_7_69
timestamp 1654395037
transform 1 0 8848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_73
timestamp 1654395037
transform 1 0 9296 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_7_78
timestamp 1654395037
transform 1 0 9856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_90
timestamp 1654395037
transform 1 0 11200 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_106
timestamp 1654395037
transform 1 0 12992 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_110
timestamp 1654395037
transform 1 0 13440 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1654395037
transform 1 0 1344 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1654395037
transform 1 0 4928 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_37
timestamp 1654395037
transform 1 0 5264 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_45
timestamp 1654395037
transform 1 0 6160 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_49
timestamp 1654395037
transform 1 0 6608 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_8_65
timestamp 1654395037
transform 1 0 8400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_71
timestamp 1654395037
transform 1 0 9072 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_8_87
timestamp 1654395037
transform 1 0 10864 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_93
timestamp 1654395037
transform 1 0 11536 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1654395037
transform 1 0 12432 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1654395037
transform 1 0 12880 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_8_108
timestamp 1654395037
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_110
timestamp 1654395037
transform 1 0 13440 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_2
timestamp 1654395037
transform 1 0 1344 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_9_6
timestamp 1654395037
transform 1 0 1792 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_9_12
timestamp 1654395037
transform 1 0 2464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_18
timestamp 1654395037
transform 1 0 3136 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_50
timestamp 1654395037
transform 1 0 6720 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_55
timestamp 1654395037
transform 1 0 7280 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_73
timestamp 1654395037
transform 1 0 9296 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_105
timestamp 1654395037
transform 1 0 12880 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_9_109
timestamp 1654395037
transform 1 0 13328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_2
timestamp 1654395037
transform 1 0 1344 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_10_6
timestamp 1654395037
transform 1 0 1792 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_12
timestamp 1654395037
transform 1 0 2464 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_28
timestamp 1654395037
transform 1 0 4256 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_10_32
timestamp 1654395037
transform 1 0 4704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1654395037
transform 1 0 4928 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_37
timestamp 1654395037
transform 1 0 5264 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_53
timestamp 1654395037
transform 1 0 7056 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_10_57
timestamp 1654395037
transform 1 0 7504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_63
timestamp 1654395037
transform 1 0 8176 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_10_95
timestamp 1654395037
transform 1 0 11760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1654395037
transform 1 0 12432 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1654395037
transform 1 0 12880 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_10_108
timestamp 1654395037
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_110
timestamp 1654395037
transform 1 0 13440 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_11_2
timestamp 1654395037
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_4
timestamp 1654395037
transform 1 0 1568 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_11_14
timestamp 1654395037
transform 1 0 2688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_20
timestamp 1654395037
transform 1 0 3360 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_11_58
timestamp 1654395037
transform 1 0 7616 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1654395037
transform 1 0 8512 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1654395037
transform 1 0 8960 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_73
timestamp 1654395037
transform 1 0 9296 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_81
timestamp 1654395037
transform 1 0 10192 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_11_85
timestamp 1654395037
transform 1 0 10640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_87
timestamp 1654395037
transform 1 0 10864 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_11_92
timestamp 1654395037
transform 1 0 11424 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_11_109
timestamp 1654395037
transform 1 0 13328 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1654395037
transform 1 0 1344 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1654395037
transform 1 0 4928 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_37
timestamp 1654395037
transform 1 0 5264 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_53
timestamp 1654395037
transform 1 0 7056 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_12_57
timestamp 1654395037
transform 1 0 7504 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_63
timestamp 1654395037
transform 1 0 8176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_12_67
timestamp 1654395037
transform 1 0 8624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_69
timestamp 1654395037
transform 1 0 8848 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_72
timestamp 1654395037
transform 1 0 9184 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_88
timestamp 1654395037
transform 1 0 10976 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_12_96
timestamp 1654395037
transform 1 0 11872 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  FILLER_12_102
timestamp 1654395037
transform 1 0 12544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_104
timestamp 1654395037
transform 1 0 12768 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_107
timestamp 1654395037
transform 1 0 13104 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 1120 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1654395037
transform -1 0 13776 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1654395037
transform 1 0 1120 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1654395037
transform -1 0 13776 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1654395037
transform 1 0 1120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1654395037
transform -1 0 13776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1654395037
transform 1 0 1120 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1654395037
transform -1 0 13776 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1654395037
transform 1 0 1120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1654395037
transform -1 0 13776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1654395037
transform 1 0 1120 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1654395037
transform -1 0 13776 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1654395037
transform 1 0 1120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1654395037
transform -1 0 13776 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1654395037
transform 1 0 1120 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1654395037
transform -1 0 13776 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1654395037
transform 1 0 1120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1654395037
transform -1 0 13776 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1654395037
transform 1 0 1120 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1654395037
transform -1 0 13776 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1654395037
transform 1 0 1120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1654395037
transform -1 0 13776 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1654395037
transform 1 0 1120 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1654395037
transform -1 0 13776 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1654395037
transform 1 0 1120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1654395037
transform -1 0 13776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_26
timestamp 1654395037
transform 1 0 5040 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_27
timestamp 1654395037
transform 1 0 8960 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_28
timestamp 1654395037
transform 1 0 12880 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_29
timestamp 1654395037
transform 1 0 9072 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_30
timestamp 1654395037
transform 1 0 5040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_31
timestamp 1654395037
transform 1 0 12992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_32
timestamp 1654395037
transform 1 0 9072 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_33
timestamp 1654395037
transform 1 0 5040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_34
timestamp 1654395037
transform 1 0 12992 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_35
timestamp 1654395037
transform 1 0 9072 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_36
timestamp 1654395037
transform 1 0 5040 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_37
timestamp 1654395037
transform 1 0 12992 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_38
timestamp 1654395037
transform 1 0 9072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_39
timestamp 1654395037
transform 1 0 5040 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_40
timestamp 1654395037
transform 1 0 12992 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_41
timestamp 1654395037
transform 1 0 9072 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_42
timestamp 1654395037
transform 1 0 5040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_43
timestamp 1654395037
transform 1 0 12992 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_44
timestamp 1654395037
transform 1 0 9072 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_45
timestamp 1654395037
transform 1 0 5040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_46
timestamp 1654395037
transform 1 0 8960 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_47
timestamp 1654395037
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__inv_12  spare_logic_biginv pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 9184 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  spare_logic_const_one\[0\] pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 4256 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  spare_logic_const_one\[1\]
timestamp 1654395037
transform -1 0 2464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  spare_logic_const_one\[2\]
timestamp 1654395037
transform 1 0 12432 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  spare_logic_const_one\[3\]
timestamp 1654395037
transform -1 0 2464 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[0\] pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 7728 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[1\]
timestamp 1654395037
transform 1 0 7504 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[2\]
timestamp 1654395037
transform -1 0 7280 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[3\]
timestamp 1654395037
transform 1 0 7728 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[4\]
timestamp 1654395037
transform 1 0 5600 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[5\]
timestamp 1654395037
transform 1 0 2912 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[6\]
timestamp 1654395037
transform -1 0 9632 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[7\]
timestamp 1654395037
transform -1 0 3136 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[8\]
timestamp 1654395037
transform 1 0 7056 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[9\]
timestamp 1654395037
transform 1 0 3024 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[10\]
timestamp 1654395037
transform -1 0 9856 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[11\]
timestamp 1654395037
transform 1 0 2464 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[12\]
timestamp 1654395037
transform 1 0 11088 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[13\]
timestamp 1654395037
transform 1 0 12096 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[14\]
timestamp 1654395037
transform 1 0 8624 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[15\]
timestamp 1654395037
transform -1 0 12432 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[16\]
timestamp 1654395037
transform 1 0 6272 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[17\]
timestamp 1654395037
transform 1 0 10976 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[18\]
timestamp 1654395037
transform 1 0 6832 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[19\]
timestamp 1654395037
transform 1 0 1792 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[20\]
timestamp 1654395037
transform -1 0 9744 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[21\]
timestamp 1654395037
transform -1 0 2464 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[22\]
timestamp 1654395037
transform 1 0 5936 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[23\]
timestamp 1654395037
transform 1 0 5264 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[24\]
timestamp 1654395037
transform 1 0 10416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[25\]
timestamp 1654395037
transform 1 0 5824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spare_logic_const_zero\[26\]
timestamp 1654395037
transform 1 0 9968 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2  spare_logic_flop\[0\] pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform 1 0 1680 0 -1 3136
box -86 -86 4678 870
use gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2  spare_logic_flop\[1\]
timestamp 1654395037
transform 1 0 7728 0 1 3136
box -86 -86 4678 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  spare_logic_inv\[0\] pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 8512 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  spare_logic_inv\[1\]
timestamp 1654395037
transform -1 0 7392 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  spare_logic_inv\[2\]
timestamp 1654395037
transform 1 0 7504 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  spare_logic_inv\[3\]
timestamp 1654395037
transform -1 0 7616 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  spare_logic_mux\[0\] pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 13328 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  spare_logic_mux\[1\]
timestamp 1654395037
transform -1 0 8400 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  spare_logic_nand\[0\] pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 2688 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  spare_logic_nand\[1\]
timestamp 1654395037
transform -1 0 8512 0 -1 3136
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  spare_logic_nor\[0\] pdk/gf180mcuC/libs.ref/gf180mcu_sc7_hv/mag
timestamp 1654395037
transform -1 0 3248 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  spare_logic_nor\[1\]
timestamp 1654395037
transform 1 0 10080 0 -1 7840
box -86 -86 1206 870
<< labels >>
flabel metal4 s 2555 1508 2875 11820 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 5745 1508 6065 11820 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 8935 1508 9255 11820 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 12125 1508 12445 11820 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 1060 2766 13836 3086 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 1060 5482 13836 5802 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 1060 8198 13836 8518 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal5 s 1060 10914 13836 11234 0 FreeSans 2304 0 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 4150 1508 4470 11820 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 7340 1508 7660 11820 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 10530 1508 10850 11820 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 1060 4124 13836 4444 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 1060 6840 13836 7160 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal5 s 1060 9556 13836 9876 0 FreeSans 2304 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal3 s 0 4760 800 4872 0 FreeSans 448 0 0 0 spare_xfq[0]
port 2 nsew signal tristate
flabel metal2 s 13384 0 13496 800 0 FreeSans 448 90 0 0 spare_xfq[1]
port 3 nsew signal tristate
flabel metal2 s 6664 13200 6776 14000 0 FreeSans 448 90 0 0 spare_xi[0]
port 4 nsew signal tristate
flabel metal2 s 5320 0 5432 800 0 FreeSans 448 90 0 0 spare_xi[1]
port 5 nsew signal tristate
flabel metal3 s 14200 2072 15000 2184 0 FreeSans 448 0 0 0 spare_xi[2]
port 6 nsew signal tristate
flabel metal3 s 0 10136 800 10248 0 FreeSans 448 0 0 0 spare_xi[3]
port 7 nsew signal tristate
flabel metal3 s 14200 728 15000 840 0 FreeSans 448 0 0 0 spare_xib
port 8 nsew signal tristate
flabel metal2 s 14728 0 14840 800 0 FreeSans 448 90 0 0 spare_xmx[0]
port 9 nsew signal tristate
flabel metal3 s 14200 10136 15000 10248 0 FreeSans 448 0 0 0 spare_xmx[1]
port 10 nsew signal tristate
flabel metal2 s -56 13200 56 14000 0 FreeSans 448 90 0 0 spare_xna[0]
port 11 nsew signal tristate
flabel metal2 s 8008 0 8120 800 0 FreeSans 448 90 0 0 spare_xna[1]
port 12 nsew signal tristate
flabel metal3 s 0 3416 800 3528 0 FreeSans 448 0 0 0 spare_xno[0]
port 13 nsew signal tristate
flabel metal2 s 10696 0 10808 800 0 FreeSans 448 90 0 0 spare_xno[1]
port 14 nsew signal tristate
flabel metal3 s 14200 11480 15000 11592 0 FreeSans 448 0 0 0 spare_xz[0]
port 15 nsew signal tristate
flabel metal3 s 0 7448 800 7560 0 FreeSans 448 0 0 0 spare_xz[10]
port 16 nsew signal tristate
flabel metal2 s 2632 0 2744 800 0 FreeSans 448 90 0 0 spare_xz[11]
port 17 nsew signal tristate
flabel metal2 s 13384 13200 13496 14000 0 FreeSans 448 90 0 0 spare_xz[12]
port 18 nsew signal tristate
flabel metal2 s 9352 13200 9464 14000 0 FreeSans 448 90 0 0 spare_xz[13]
port 19 nsew signal tristate
flabel metal3 s 14200 7448 15000 7560 0 FreeSans 448 0 0 0 spare_xz[14]
port 20 nsew signal tristate
flabel metal2 s 12040 13200 12152 14000 0 FreeSans 448 90 0 0 spare_xz[15]
port 21 nsew signal tristate
flabel metal3 s 0 2072 800 2184 0 FreeSans 448 0 0 0 spare_xz[16]
port 22 nsew signal tristate
flabel metal3 s 14200 12824 15000 12936 0 FreeSans 448 0 0 0 spare_xz[17]
port 23 nsew signal tristate
flabel metal2 s 2632 13200 2744 14000 0 FreeSans 448 90 0 0 spare_xz[18]
port 24 nsew signal tristate
flabel metal2 s 0 -56 800 56 0 FreeSans 448 0 0 0 spare_xz[19]
port 25 nsew signal tristate
flabel metal2 s 8008 13200 8120 14000 0 FreeSans 448 90 0 0 spare_xz[1]
port 26 nsew signal tristate
flabel metal3 s 14200 8792 15000 8904 0 FreeSans 448 0 0 0 spare_xz[20]
port 27 nsew signal tristate
flabel metal2 s 1288 13200 1400 14000 0 FreeSans 448 90 0 0 spare_xz[21]
port 28 nsew signal tristate
flabel metal3 s 0 728 800 840 0 FreeSans 448 0 0 0 spare_xz[22]
port 29 nsew signal tristate
flabel metal2 s 12040 0 12152 800 0 FreeSans 448 90 0 0 spare_xz[23]
port 30 nsew signal tristate
flabel metal2 s 10696 13200 10808 14000 0 FreeSans 448 90 0 0 spare_xz[24]
port 31 nsew signal tristate
flabel metal3 s 14200 3416 15000 3528 0 FreeSans 448 0 0 0 spare_xz[25]
port 32 nsew signal tristate
flabel metal2 s 1288 0 1400 800 0 FreeSans 448 90 0 0 spare_xz[26]
port 33 nsew signal tristate
flabel metal2 s 3976 0 4088 800 0 FreeSans 448 90 0 0 spare_xz[27]
port 34 nsew signal tristate
flabel metal3 s 0 11480 800 11592 0 FreeSans 448 0 0 0 spare_xz[28]
port 35 nsew signal tristate
flabel metal3 s 14200 4760 15000 4872 0 FreeSans 448 0 0 0 spare_xz[29]
port 36 nsew signal tristate
flabel metal2 s 6664 0 6776 800 0 FreeSans 448 90 0 0 spare_xz[2]
port 37 nsew signal tristate
flabel metal3 s 0 8792 800 8904 0 FreeSans 448 0 0 0 spare_xz[30]
port 38 nsew signal tristate
flabel metal2 s 14728 13200 14840 14000 0 FreeSans 448 90 0 0 spare_xz[3]
port 39 nsew signal tristate
flabel metal2 s 3976 13200 4088 14000 0 FreeSans 448 90 0 0 spare_xz[4]
port 40 nsew signal tristate
flabel metal2 s 5320 13200 5432 14000 0 FreeSans 448 90 0 0 spare_xz[5]
port 41 nsew signal tristate
flabel metal2 s 9352 0 9464 800 0 FreeSans 448 90 0 0 spare_xz[6]
port 42 nsew signal tristate
flabel metal3 s 0 6104 800 6216 0 FreeSans 448 0 0 0 spare_xz[7]
port 43 nsew signal tristate
flabel metal3 s 0 12824 800 12936 0 FreeSans 448 0 0 0 spare_xz[8]
port 44 nsew signal tristate
flabel metal3 s 14200 6104 15000 6216 0 FreeSans 448 0 0 0 spare_xz[9]
port 45 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 15000 14000
<< end >>
