magic
tech gf180mcuC
magscale 1 10
timestamp 1655309791
<< metal1 >>
rect 3923 8654 6463 8714
rect 3923 7964 3963 8654
rect 6403 7964 6463 8654
rect 20890 8230 21090 8247
rect 20890 8066 20908 8230
rect 21071 8066 21090 8230
rect 20890 8047 21090 8066
rect 22253 8210 22453 8227
rect 3923 7914 6463 7964
rect 20642 7959 20643 7974
rect 20907 7959 21045 8047
rect 22253 8046 22271 8210
rect 22434 8046 22453 8210
rect 22253 8027 22453 8046
rect 20642 7831 21045 7959
rect 20907 6821 21045 7831
rect 22342 7592 22451 8027
rect 3953 6634 6493 6684
rect 3953 5944 4003 6634
rect 6443 5944 6493 6634
rect 22096 6567 22204 7023
rect 22342 6808 22452 7592
rect 24708 7000 24908 7017
rect 24708 6995 24727 7000
rect 24085 6832 24727 6995
rect 24889 6832 24908 7000
rect 24085 6826 24908 6832
rect 24708 6817 24908 6826
rect 22096 6550 22310 6567
rect 22096 6386 22128 6550
rect 22291 6386 22310 6550
rect 22096 6367 22310 6386
rect 23960 6529 24160 6544
rect 24709 6529 24909 6542
rect 23960 6527 24909 6529
rect 23960 6363 23978 6527
rect 24141 6363 24728 6527
rect 23960 6360 24728 6363
rect 23960 6344 24160 6360
rect 24709 6359 24728 6360
rect 24890 6359 24909 6527
rect 24709 6342 24909 6359
rect 3953 5884 6493 5944
<< via1 >>
rect 3963 7964 6403 8654
rect 20908 8066 21071 8230
rect 22271 8046 22434 8210
rect 4003 5944 6443 6634
rect 24727 6832 24889 7000
rect 22128 6386 22291 6550
rect 23978 6363 24141 6527
rect 24728 6359 24890 6527
<< metal2 >>
rect 3923 8654 6463 8714
rect 3923 7964 3963 8654
rect 6403 7964 6463 8654
rect 20948 8465 22404 8602
rect 20948 8247 21085 8465
rect 20890 8230 21090 8247
rect 20890 8066 20908 8230
rect 21071 8066 21090 8230
rect 22267 8227 22404 8465
rect 20890 8047 21090 8066
rect 22253 8210 22453 8227
rect 22253 8046 22271 8210
rect 22434 8046 22453 8210
rect 22253 8027 22453 8046
rect 3923 7914 6463 7964
rect 7152 7611 7520 7647
rect 3953 6634 6493 6684
rect 3953 5944 4003 6634
rect 6443 5944 6493 6634
rect 7152 6601 7192 7611
rect 7470 6601 7520 7611
rect 7152 6561 7520 6601
rect 17284 7474 17907 7555
rect 17284 6395 17352 7474
rect 17830 6857 17907 7474
rect 24708 7000 25108 7017
rect 17830 6659 18224 6857
rect 24708 6832 24727 7000
rect 24889 6832 25108 7000
rect 24708 6817 25108 6832
rect 17830 6395 17907 6659
rect 17284 6306 17907 6395
rect 22110 6550 22310 6567
rect 22110 6386 22128 6550
rect 22291 6386 22310 6550
rect 22110 6367 22310 6386
rect 23960 6527 24160 6544
rect 3953 5884 6493 5944
rect 22185 5910 22306 6367
rect 23960 6363 23978 6527
rect 24141 6363 24160 6527
rect 23960 6344 24160 6363
rect 24709 6527 25109 6542
rect 24709 6359 24728 6527
rect 24890 6359 25109 6527
rect 23989 5910 24125 6344
rect 24709 6342 25109 6359
rect 22185 5774 24125 5910
<< via2 >>
rect 3963 7964 6403 8654
rect 4003 5944 6443 6634
rect 7192 6601 7470 7611
rect 17352 6395 17830 7474
<< metal3 >>
rect 3923 8654 6463 8714
rect 3923 7964 3963 8654
rect 6403 7964 6463 8654
rect 3923 7914 6463 7964
rect 7045 7611 7520 7647
rect 3953 6634 6493 6684
rect 3953 5944 4003 6634
rect 6443 5944 6493 6634
rect 7045 6601 7086 7611
rect 7470 6601 7520 7611
rect 7045 6561 7520 6601
rect 17284 7474 17907 7555
rect 17284 6395 17352 7474
rect 17830 6395 17907 7474
rect 17284 6306 17907 6395
rect 3953 5884 6493 5944
<< via3 >>
rect 3963 7964 6403 8654
rect 4003 5944 6443 6634
rect 7086 6601 7192 7611
rect 7192 6601 7364 7611
rect 17352 6395 17830 7474
<< metal4 >>
rect 3923 8654 6463 8714
rect 3923 7964 3963 8654
rect 6403 7964 6463 8654
rect 3923 7914 6463 7964
rect 7046 7611 7414 7647
rect 3953 6634 6493 6684
rect 3953 5944 4003 6634
rect 6443 5944 6493 6634
rect 7046 6601 7086 7611
rect 7364 6601 7414 7611
rect 17284 7474 17907 7555
rect 7046 6561 7414 6601
rect 15694 7196 17016 7256
rect 3953 5884 6493 5944
rect 15694 5877 15771 7196
rect 16930 5877 17016 7196
rect 17284 6395 17352 7474
rect 17830 6395 17907 7474
rect 17284 6306 17907 6395
rect 15694 5808 17016 5877
<< via4 >>
rect 3963 7964 6403 8654
rect 4003 5944 6443 6634
rect 7086 6601 7364 7611
rect 15771 5877 16930 7196
rect 17352 6395 17830 7474
<< metal5 >>
rect 24 8654 6463 8714
rect 24 7964 3963 8654
rect 6403 7964 6463 8654
rect 24 7914 6463 7964
rect 7157 7735 17700 7983
rect 7157 7647 7414 7735
rect 7046 7611 7414 7647
rect 24 6634 6493 6684
rect 24 5944 4003 6634
rect 6443 5944 6493 6634
rect 7046 6601 7086 7611
rect 7364 6601 7414 7611
rect 17284 7619 17700 7735
rect 17284 7474 17907 7619
rect 7046 6561 7414 6601
rect 15454 7196 17016 7256
rect 24 5884 6493 5944
rect 15454 5877 15771 7196
rect 16930 5877 17016 7196
rect 17284 6395 17352 7474
rect 17830 6395 17907 7474
rect 17284 6306 17907 6395
rect 15454 5808 17016 5877
use reduction_mirror  X0
timestamp 1655309791
transform 1 0 -261 0 1 6308
box 261 -6308 25417 2408
use large_mimcap  X1
timestamp 1655309791
transform 1 0 11168 0 1 368
box -3514 -294 4286 7615
use schmitt_inverter  X2
timestamp 1655307388
transform 1 0 17635 0 1 8025
box 526 -2315 3059 685
use std_inverter  X3
timestamp 1655304105
transform 1 0 20638 0 -1 7361
box 265 -1350 1460 1650
use std_buffer  std_buffer_0
timestamp 1655304105
transform 1 0 21358 0 -1 8992
box 1094 292 2782 3292
<< labels >>
flabel metal2 s 24908 6817 25108 7017 0 FreeSans 1280 0 0 0 por
port 3 nsew
flabel metal2 s 24909 6342 25109 6542 0 FreeSans 1280 0 0 0 porb
port 2 nsew
flabel metal5 s 803 8147 1003 8347 0 FreeSans 1280 0 0 0 VDD
port 0 nsew
flabel metal5 s 803 6188 1003 6388 0 FreeSans 1280 0 0 0 VSS
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 25110 8710
string GDS_FILE ../gds/simple_por.gds.gz
string GDS_START 0
string LEFclass BLOCK
<< end >>
