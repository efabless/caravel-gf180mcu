VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_id_textblock
  CLASS BLOCK ;
  FOREIGN user_id_textblock ;
  ORIGIN 0.000 0.000 ;
  SIZE 207.200 BY 54.050 ;
  OBS
      LAYER Metal5 ;
        RECT 4.800 4.450 203.915 49.810 ;
  END
END user_id_textblock
END LIBRARY

