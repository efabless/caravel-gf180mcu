magic
tech gf180mcuC
magscale 1 10
timestamp 1655307388
<< error_p >>
rect -58 -155 -47 -109
<< nwell >>
rect -378 -386 368 386
<< mvpmos >>
rect -60 -76 50 124
<< mvpdiff >>
rect -148 111 -60 124
rect -148 -63 -135 111
rect -89 -63 -60 111
rect -148 -76 -60 -63
rect 50 111 138 124
rect 50 -63 79 111
rect 125 -63 138 111
rect 50 -76 138 -63
<< mvpdiffc >>
rect -135 -63 -89 111
rect 79 -63 125 111
<< mvnsubdiff >>
rect -292 228 282 300
rect -292 184 -220 228
rect -292 -184 -279 184
rect -233 -184 -220 184
rect 210 184 282 228
rect -292 -228 -220 -184
rect 210 -184 223 184
rect 269 -184 282 184
rect 210 -228 282 -184
rect -292 -300 282 -228
<< mvnsubdiffcont >>
rect -279 -184 -233 184
rect 223 -184 269 184
<< polysilicon >>
rect -60 124 50 168
rect -60 -109 50 -76
rect -60 -155 -47 -109
rect 37 -155 50 -109
rect -60 -168 50 -155
<< polycontact >>
rect -47 -155 37 -109
<< metal1 >>
rect -279 241 269 287
rect -279 184 -233 241
rect 223 184 269 241
rect -135 111 -89 122
rect -135 -74 -89 -63
rect 79 111 125 122
rect 79 -74 125 -63
rect -58 -155 -47 -109
rect 37 -155 48 -109
rect -279 -241 -233 -184
rect 223 -241 269 -184
rect -279 -287 269 -241
<< properties >>
string FIXED_BBOX -246 -264 246 264
string gencell pmos_6p0
string library gf180mcu
string parameters w 1 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.5 wmin 0.3 full_metal 1 compatible {pmos_3p3 pmos_6p0}
<< end >>
