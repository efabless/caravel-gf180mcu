magic
tech gf180mcuC
magscale 1 10
timestamp 1670147978
<< metal1 >>
rect 9090 11118 9102 11170
rect 9154 11167 9166 11170
rect 10546 11167 10558 11170
rect 9154 11121 10558 11167
rect 9154 11118 9166 11121
rect 10546 11118 10558 11121
rect 10610 11167 10622 11170
rect 11554 11167 11566 11170
rect 10610 11121 11566 11167
rect 10610 11118 10622 11121
rect 11554 11118 11566 11121
rect 11618 11118 11630 11170
rect 14466 11118 14478 11170
rect 14530 11167 14542 11170
rect 15138 11167 15150 11170
rect 14530 11121 15150 11167
rect 14530 11118 14542 11121
rect 15138 11118 15150 11121
rect 15202 11118 15214 11170
rect 224 11002 16848 11036
rect 224 10950 4210 11002
rect 4262 10950 4314 11002
rect 4366 10950 4418 11002
rect 4470 10950 8326 11002
rect 8378 10950 8430 11002
rect 8482 10950 8534 11002
rect 8586 10950 12442 11002
rect 12494 10950 12546 11002
rect 12598 10950 12650 11002
rect 12702 10950 16558 11002
rect 16610 10950 16662 11002
rect 16714 10950 16766 11002
rect 16818 10950 16848 11002
rect 224 10916 16848 10950
rect 11566 10834 11618 10846
rect 11566 10770 11618 10782
rect 12350 10722 12402 10734
rect 1474 10670 1486 10722
rect 1538 10670 1550 10722
rect 12350 10658 12402 10670
rect 4734 10610 4786 10622
rect 2706 10558 2718 10610
rect 2770 10558 2782 10610
rect 5730 10558 5742 10610
rect 5794 10558 5806 10610
rect 10546 10558 10558 10610
rect 10610 10558 10622 10610
rect 15138 10558 15150 10610
rect 15202 10558 15214 10610
rect 4734 10546 4786 10558
rect 3726 10498 3778 10510
rect 6850 10446 6862 10498
rect 6914 10446 6926 10498
rect 9090 10446 9102 10498
rect 9154 10446 9166 10498
rect 14242 10446 14254 10498
rect 14306 10446 14318 10498
rect 3726 10434 3778 10446
rect 224 10218 16688 10252
rect 224 10166 2152 10218
rect 2204 10166 2256 10218
rect 2308 10166 2360 10218
rect 2412 10166 6268 10218
rect 6320 10166 6372 10218
rect 6424 10166 6476 10218
rect 6528 10166 10384 10218
rect 10436 10166 10488 10218
rect 10540 10166 10592 10218
rect 10644 10166 14500 10218
rect 14552 10166 14604 10218
rect 14656 10166 14708 10218
rect 14760 10166 16688 10218
rect 224 10132 16688 10166
rect 15362 9998 15374 10050
rect 15426 10047 15438 10050
rect 16034 10047 16046 10050
rect 15426 10001 16046 10047
rect 15426 9998 15438 10001
rect 16034 9998 16046 10001
rect 16098 9998 16110 10050
rect 11790 9938 11842 9950
rect 15598 9938 15650 9950
rect 2482 9886 2494 9938
rect 2546 9886 2558 9938
rect 7074 9886 7086 9938
rect 7138 9886 7150 9938
rect 14354 9886 14366 9938
rect 14418 9886 14430 9938
rect 11790 9874 11842 9886
rect 15598 9874 15650 9886
rect 16046 9938 16098 9950
rect 16046 9874 16098 9886
rect 3378 9774 3390 9826
rect 3442 9774 3454 9826
rect 7746 9774 7758 9826
rect 7810 9774 7822 9826
rect 10770 9774 10782 9826
rect 10834 9774 10846 9826
rect 12562 9774 12574 9826
rect 12626 9774 12638 9826
rect 4510 9714 4562 9726
rect 9538 9662 9550 9714
rect 9602 9662 9614 9714
rect 4510 9650 4562 9662
rect 224 9434 16848 9468
rect 224 9382 4210 9434
rect 4262 9382 4314 9434
rect 4366 9382 4418 9434
rect 4470 9382 8326 9434
rect 8378 9382 8430 9434
rect 8482 9382 8534 9434
rect 8586 9382 12442 9434
rect 12494 9382 12546 9434
rect 12598 9382 12650 9434
rect 12702 9382 16558 9434
rect 16610 9382 16662 9434
rect 16714 9382 16766 9434
rect 16818 9382 16848 9434
rect 224 9348 16848 9382
rect 12014 9042 12066 9054
rect 2930 8990 2942 9042
rect 2994 8990 3006 9042
rect 7298 8990 7310 9042
rect 7362 8990 7374 9042
rect 10994 8990 11006 9042
rect 11058 8990 11070 9042
rect 15474 8990 15486 9042
rect 15538 8990 15550 9042
rect 12014 8978 12066 8990
rect 3950 8930 4002 8942
rect 1922 8878 1934 8930
rect 1986 8878 1998 8930
rect 6514 8878 6526 8930
rect 6578 8878 6590 8930
rect 9874 8878 9886 8930
rect 9938 8878 9950 8930
rect 14690 8878 14702 8930
rect 14754 8878 14766 8930
rect 3950 8866 4002 8878
rect 224 8650 16688 8684
rect 224 8598 2152 8650
rect 2204 8598 2256 8650
rect 2308 8598 2360 8650
rect 2412 8598 6268 8650
rect 6320 8598 6372 8650
rect 6424 8598 6476 8650
rect 6528 8598 10384 8650
rect 10436 8598 10488 8650
rect 10540 8598 10592 8650
rect 10644 8598 14500 8650
rect 14552 8598 14604 8650
rect 14656 8598 14708 8650
rect 14760 8598 16688 8650
rect 224 8564 16688 8598
rect 914 8318 926 8370
rect 978 8318 990 8370
rect 8754 8318 8766 8370
rect 8818 8318 8830 8370
rect 14914 8318 14926 8370
rect 14978 8318 14990 8370
rect 3726 8258 3778 8270
rect 10670 8258 10722 8270
rect 2706 8206 2718 8258
rect 2770 8206 2782 8258
rect 9650 8206 9662 8258
rect 9714 8206 9726 8258
rect 16146 8206 16158 8258
rect 16210 8206 16222 8258
rect 3726 8194 3778 8206
rect 10670 8194 10722 8206
rect 7086 8034 7138 8046
rect 7086 7970 7138 7982
rect 224 7866 16848 7900
rect 224 7814 4210 7866
rect 4262 7814 4314 7866
rect 4366 7814 4418 7866
rect 4470 7814 8326 7866
rect 8378 7814 8430 7866
rect 8482 7814 8534 7866
rect 8586 7814 12442 7866
rect 12494 7814 12546 7866
rect 12598 7814 12650 7866
rect 12702 7814 16558 7866
rect 16610 7814 16662 7866
rect 16714 7814 16766 7866
rect 16818 7814 16848 7866
rect 224 7780 16848 7814
rect 15486 7698 15538 7710
rect 15486 7634 15538 7646
rect 2706 7422 2718 7474
rect 2770 7422 2782 7474
rect 14466 7422 14478 7474
rect 14530 7422 14542 7474
rect 3726 7362 3778 7374
rect 1026 7310 1038 7362
rect 1090 7310 1102 7362
rect 3726 7298 3778 7310
rect 8542 7362 8594 7374
rect 13570 7310 13582 7362
rect 13634 7310 13646 7362
rect 8542 7298 8594 7310
rect 224 7082 16688 7116
rect 224 7030 2152 7082
rect 2204 7030 2256 7082
rect 2308 7030 2360 7082
rect 2412 7030 6268 7082
rect 6320 7030 6372 7082
rect 6424 7030 6476 7082
rect 6528 7030 10384 7082
rect 10436 7030 10488 7082
rect 10540 7030 10592 7082
rect 10644 7030 14500 7082
rect 14552 7030 14604 7082
rect 14656 7030 14708 7082
rect 14760 7030 16688 7082
rect 224 6996 16688 7030
rect 16270 6802 16322 6814
rect 8194 6750 8206 6802
rect 8258 6750 8270 6802
rect 14018 6750 14030 6802
rect 14082 6750 14094 6802
rect 16270 6738 16322 6750
rect 9202 6638 9214 6690
rect 9266 6638 9278 6690
rect 15474 6638 15486 6690
rect 15538 6638 15550 6690
rect 10222 6466 10274 6478
rect 10222 6402 10274 6414
rect 224 6298 16848 6332
rect 224 6246 4210 6298
rect 4262 6246 4314 6298
rect 4366 6246 4418 6298
rect 4470 6246 8326 6298
rect 8378 6246 8430 6298
rect 8482 6246 8534 6298
rect 8586 6246 12442 6298
rect 12494 6246 12546 6298
rect 12598 6246 12650 6298
rect 12702 6246 16558 6298
rect 16610 6246 16662 6298
rect 16714 6246 16766 6298
rect 16818 6246 16848 6298
rect 224 6212 16848 6246
rect 15026 5966 15038 6018
rect 15090 5966 15102 6018
rect 5742 5906 5794 5918
rect 4722 5854 4734 5906
rect 4786 5854 4798 5906
rect 12674 5854 12686 5906
rect 12738 5854 12750 5906
rect 13234 5854 13246 5906
rect 13298 5854 13310 5906
rect 5742 5842 5794 5854
rect 3602 5742 3614 5794
rect 3666 5742 3678 5794
rect 11554 5742 11566 5794
rect 11618 5742 11630 5794
rect 224 5514 16688 5548
rect 224 5462 2152 5514
rect 2204 5462 2256 5514
rect 2308 5462 2360 5514
rect 2412 5462 6268 5514
rect 6320 5462 6372 5514
rect 6424 5462 6476 5514
rect 6528 5462 10384 5514
rect 10436 5462 10488 5514
rect 10540 5462 10592 5514
rect 10644 5462 14500 5514
rect 14552 5462 14604 5514
rect 14656 5462 14708 5514
rect 14760 5462 16688 5514
rect 224 5428 16688 5462
rect 11342 5234 11394 5246
rect 11342 5170 11394 5182
rect 11790 5234 11842 5246
rect 11790 5170 11842 5182
rect 12574 5234 12626 5246
rect 12574 5170 12626 5182
rect 13022 5234 13074 5246
rect 14914 5182 14926 5234
rect 14978 5182 14990 5234
rect 13022 5170 13074 5182
rect 15586 5070 15598 5122
rect 15650 5070 15662 5122
rect 3838 4898 3890 4910
rect 3838 4834 3890 4846
rect 4510 4898 4562 4910
rect 4510 4834 4562 4846
rect 4958 4898 5010 4910
rect 4958 4834 5010 4846
rect 224 4730 16848 4764
rect 224 4678 4210 4730
rect 4262 4678 4314 4730
rect 4366 4678 4418 4730
rect 4470 4678 8326 4730
rect 8378 4678 8430 4730
rect 8482 4678 8534 4730
rect 8586 4678 12442 4730
rect 12494 4678 12546 4730
rect 12598 4678 12650 4730
rect 12702 4678 16558 4730
rect 16610 4678 16662 4730
rect 16714 4678 16766 4730
rect 16818 4678 16848 4730
rect 224 4644 16848 4678
rect 15710 4562 15762 4574
rect 15710 4498 15762 4510
rect 3938 4286 3950 4338
rect 4002 4286 4014 4338
rect 6962 4286 6974 4338
rect 7026 4286 7038 4338
rect 11666 4286 11678 4338
rect 11730 4286 11742 4338
rect 14578 4286 14590 4338
rect 14642 4286 14654 4338
rect 8542 4226 8594 4238
rect 2818 4174 2830 4226
rect 2882 4174 2894 4226
rect 5954 4174 5966 4226
rect 6018 4174 6030 4226
rect 10210 4174 10222 4226
rect 10274 4174 10286 4226
rect 12786 4174 12798 4226
rect 12850 4174 12862 4226
rect 8542 4162 8594 4174
rect 224 3946 16688 3980
rect 224 3894 2152 3946
rect 2204 3894 2256 3946
rect 2308 3894 2360 3946
rect 2412 3894 6268 3946
rect 6320 3894 6372 3946
rect 6424 3894 6476 3946
rect 6528 3894 10384 3946
rect 10436 3894 10488 3946
rect 10540 3894 10592 3946
rect 10644 3894 14500 3946
rect 14552 3894 14604 3946
rect 14656 3894 14708 3946
rect 14760 3894 16688 3946
rect 224 3860 16688 3894
rect 16046 3666 16098 3678
rect 2706 3614 2718 3666
rect 2770 3614 2782 3666
rect 5506 3614 5518 3666
rect 5570 3614 5582 3666
rect 10658 3614 10670 3666
rect 10722 3614 10734 3666
rect 12898 3614 12910 3666
rect 12962 3614 12974 3666
rect 16046 3602 16098 3614
rect 15598 3554 15650 3566
rect 3378 3502 3390 3554
rect 3442 3502 3454 3554
rect 6738 3502 6750 3554
rect 6802 3502 6814 3554
rect 11218 3502 11230 3554
rect 11282 3502 11294 3554
rect 14578 3502 14590 3554
rect 14642 3502 14654 3554
rect 15598 3490 15650 3502
rect 7646 3442 7698 3454
rect 7646 3378 7698 3390
rect 8430 3330 8482 3342
rect 8430 3266 8482 3278
rect 224 3162 16848 3196
rect 224 3110 4210 3162
rect 4262 3110 4314 3162
rect 4366 3110 4418 3162
rect 4470 3110 8326 3162
rect 8378 3110 8430 3162
rect 8482 3110 8534 3162
rect 8586 3110 12442 3162
rect 12494 3110 12546 3162
rect 12598 3110 12650 3162
rect 12702 3110 16558 3162
rect 16610 3110 16662 3162
rect 16714 3110 16766 3162
rect 16818 3110 16848 3162
rect 224 3076 16848 3110
rect 14814 2994 14866 3006
rect 14814 2930 14866 2942
rect 15262 2994 15314 3006
rect 15262 2930 15314 2942
rect 15822 2994 15874 3006
rect 15822 2930 15874 2942
rect 4722 2718 4734 2770
rect 4786 2718 4798 2770
rect 7410 2718 7422 2770
rect 7474 2718 7486 2770
rect 8642 2718 8654 2770
rect 8706 2718 8718 2770
rect 13794 2718 13806 2770
rect 13858 2718 13870 2770
rect 2594 2606 2606 2658
rect 2658 2606 2670 2658
rect 6514 2606 6526 2658
rect 6578 2606 6590 2658
rect 10994 2606 11006 2658
rect 11058 2606 11070 2658
rect 12002 2606 12014 2658
rect 12066 2606 12078 2658
rect 224 2378 16688 2412
rect 224 2326 2152 2378
rect 2204 2326 2256 2378
rect 2308 2326 2360 2378
rect 2412 2326 6268 2378
rect 6320 2326 6372 2378
rect 6424 2326 6476 2378
rect 6528 2326 10384 2378
rect 10436 2326 10488 2378
rect 10540 2326 10592 2378
rect 10644 2326 14500 2378
rect 14552 2326 14604 2378
rect 14656 2326 14708 2378
rect 14760 2326 16688 2378
rect 224 2292 16688 2326
rect 8430 2098 8482 2110
rect 15486 2098 15538 2110
rect 3154 2046 3166 2098
rect 3218 2046 3230 2098
rect 5058 2046 5070 2098
rect 5122 2046 5134 2098
rect 10546 2046 10558 2098
rect 10610 2046 10622 2098
rect 12674 2046 12686 2098
rect 12738 2046 12750 2098
rect 8430 2034 8482 2046
rect 15486 2034 15538 2046
rect 814 1986 866 1998
rect 1586 1934 1598 1986
rect 1650 1934 1662 1986
rect 6738 1934 6750 1986
rect 6802 1934 6814 1986
rect 11666 1934 11678 1986
rect 11730 1934 11742 1986
rect 15026 1934 15038 1986
rect 15090 1934 15102 1986
rect 814 1922 866 1934
rect 7646 1874 7698 1886
rect 7646 1810 7698 1822
rect 224 1594 16848 1628
rect 224 1542 4210 1594
rect 4262 1542 4314 1594
rect 4366 1542 4418 1594
rect 4470 1542 8326 1594
rect 8378 1542 8430 1594
rect 8482 1542 8534 1594
rect 8586 1542 12442 1594
rect 12494 1542 12546 1594
rect 12598 1542 12650 1594
rect 12702 1542 16558 1594
rect 16610 1542 16662 1594
rect 16714 1542 16766 1594
rect 16818 1542 16848 1594
rect 224 1508 16848 1542
<< via1 >>
rect 9102 11118 9154 11170
rect 10558 11118 10610 11170
rect 11566 11118 11618 11170
rect 14478 11118 14530 11170
rect 15150 11118 15202 11170
rect 4210 10950 4262 11002
rect 4314 10950 4366 11002
rect 4418 10950 4470 11002
rect 8326 10950 8378 11002
rect 8430 10950 8482 11002
rect 8534 10950 8586 11002
rect 12442 10950 12494 11002
rect 12546 10950 12598 11002
rect 12650 10950 12702 11002
rect 16558 10950 16610 11002
rect 16662 10950 16714 11002
rect 16766 10950 16818 11002
rect 11566 10782 11618 10834
rect 1486 10670 1538 10722
rect 12350 10670 12402 10722
rect 2718 10558 2770 10610
rect 4734 10558 4786 10610
rect 5742 10558 5794 10610
rect 10558 10558 10610 10610
rect 15150 10558 15202 10610
rect 3726 10446 3778 10498
rect 6862 10446 6914 10498
rect 9102 10446 9154 10498
rect 14254 10446 14306 10498
rect 2152 10166 2204 10218
rect 2256 10166 2308 10218
rect 2360 10166 2412 10218
rect 6268 10166 6320 10218
rect 6372 10166 6424 10218
rect 6476 10166 6528 10218
rect 10384 10166 10436 10218
rect 10488 10166 10540 10218
rect 10592 10166 10644 10218
rect 14500 10166 14552 10218
rect 14604 10166 14656 10218
rect 14708 10166 14760 10218
rect 15374 9998 15426 10050
rect 16046 9998 16098 10050
rect 2494 9886 2546 9938
rect 7086 9886 7138 9938
rect 11790 9886 11842 9938
rect 14366 9886 14418 9938
rect 15598 9886 15650 9938
rect 16046 9886 16098 9938
rect 3390 9774 3442 9826
rect 7758 9774 7810 9826
rect 10782 9774 10834 9826
rect 12574 9774 12626 9826
rect 4510 9662 4562 9714
rect 9550 9662 9602 9714
rect 4210 9382 4262 9434
rect 4314 9382 4366 9434
rect 4418 9382 4470 9434
rect 8326 9382 8378 9434
rect 8430 9382 8482 9434
rect 8534 9382 8586 9434
rect 12442 9382 12494 9434
rect 12546 9382 12598 9434
rect 12650 9382 12702 9434
rect 16558 9382 16610 9434
rect 16662 9382 16714 9434
rect 16766 9382 16818 9434
rect 2942 8990 2994 9042
rect 7310 8990 7362 9042
rect 11006 8990 11058 9042
rect 12014 8990 12066 9042
rect 15486 8990 15538 9042
rect 1934 8878 1986 8930
rect 3950 8878 4002 8930
rect 6526 8878 6578 8930
rect 9886 8878 9938 8930
rect 14702 8878 14754 8930
rect 2152 8598 2204 8650
rect 2256 8598 2308 8650
rect 2360 8598 2412 8650
rect 6268 8598 6320 8650
rect 6372 8598 6424 8650
rect 6476 8598 6528 8650
rect 10384 8598 10436 8650
rect 10488 8598 10540 8650
rect 10592 8598 10644 8650
rect 14500 8598 14552 8650
rect 14604 8598 14656 8650
rect 14708 8598 14760 8650
rect 926 8318 978 8370
rect 8766 8318 8818 8370
rect 14926 8318 14978 8370
rect 2718 8206 2770 8258
rect 3726 8206 3778 8258
rect 9662 8206 9714 8258
rect 10670 8206 10722 8258
rect 16158 8206 16210 8258
rect 7086 7982 7138 8034
rect 4210 7814 4262 7866
rect 4314 7814 4366 7866
rect 4418 7814 4470 7866
rect 8326 7814 8378 7866
rect 8430 7814 8482 7866
rect 8534 7814 8586 7866
rect 12442 7814 12494 7866
rect 12546 7814 12598 7866
rect 12650 7814 12702 7866
rect 16558 7814 16610 7866
rect 16662 7814 16714 7866
rect 16766 7814 16818 7866
rect 15486 7646 15538 7698
rect 2718 7422 2770 7474
rect 14478 7422 14530 7474
rect 1038 7310 1090 7362
rect 3726 7310 3778 7362
rect 8542 7310 8594 7362
rect 13582 7310 13634 7362
rect 2152 7030 2204 7082
rect 2256 7030 2308 7082
rect 2360 7030 2412 7082
rect 6268 7030 6320 7082
rect 6372 7030 6424 7082
rect 6476 7030 6528 7082
rect 10384 7030 10436 7082
rect 10488 7030 10540 7082
rect 10592 7030 10644 7082
rect 14500 7030 14552 7082
rect 14604 7030 14656 7082
rect 14708 7030 14760 7082
rect 8206 6750 8258 6802
rect 14030 6750 14082 6802
rect 16270 6750 16322 6802
rect 9214 6638 9266 6690
rect 15486 6638 15538 6690
rect 10222 6414 10274 6466
rect 4210 6246 4262 6298
rect 4314 6246 4366 6298
rect 4418 6246 4470 6298
rect 8326 6246 8378 6298
rect 8430 6246 8482 6298
rect 8534 6246 8586 6298
rect 12442 6246 12494 6298
rect 12546 6246 12598 6298
rect 12650 6246 12702 6298
rect 16558 6246 16610 6298
rect 16662 6246 16714 6298
rect 16766 6246 16818 6298
rect 15038 5966 15090 6018
rect 4734 5854 4786 5906
rect 5742 5854 5794 5906
rect 12686 5854 12738 5906
rect 13246 5854 13298 5906
rect 3614 5742 3666 5794
rect 11566 5742 11618 5794
rect 2152 5462 2204 5514
rect 2256 5462 2308 5514
rect 2360 5462 2412 5514
rect 6268 5462 6320 5514
rect 6372 5462 6424 5514
rect 6476 5462 6528 5514
rect 10384 5462 10436 5514
rect 10488 5462 10540 5514
rect 10592 5462 10644 5514
rect 14500 5462 14552 5514
rect 14604 5462 14656 5514
rect 14708 5462 14760 5514
rect 11342 5182 11394 5234
rect 11790 5182 11842 5234
rect 12574 5182 12626 5234
rect 13022 5182 13074 5234
rect 14926 5182 14978 5234
rect 15598 5070 15650 5122
rect 3838 4846 3890 4898
rect 4510 4846 4562 4898
rect 4958 4846 5010 4898
rect 4210 4678 4262 4730
rect 4314 4678 4366 4730
rect 4418 4678 4470 4730
rect 8326 4678 8378 4730
rect 8430 4678 8482 4730
rect 8534 4678 8586 4730
rect 12442 4678 12494 4730
rect 12546 4678 12598 4730
rect 12650 4678 12702 4730
rect 16558 4678 16610 4730
rect 16662 4678 16714 4730
rect 16766 4678 16818 4730
rect 15710 4510 15762 4562
rect 3950 4286 4002 4338
rect 6974 4286 7026 4338
rect 11678 4286 11730 4338
rect 14590 4286 14642 4338
rect 2830 4174 2882 4226
rect 5966 4174 6018 4226
rect 8542 4174 8594 4226
rect 10222 4174 10274 4226
rect 12798 4174 12850 4226
rect 2152 3894 2204 3946
rect 2256 3894 2308 3946
rect 2360 3894 2412 3946
rect 6268 3894 6320 3946
rect 6372 3894 6424 3946
rect 6476 3894 6528 3946
rect 10384 3894 10436 3946
rect 10488 3894 10540 3946
rect 10592 3894 10644 3946
rect 14500 3894 14552 3946
rect 14604 3894 14656 3946
rect 14708 3894 14760 3946
rect 2718 3614 2770 3666
rect 5518 3614 5570 3666
rect 10670 3614 10722 3666
rect 12910 3614 12962 3666
rect 16046 3614 16098 3666
rect 3390 3502 3442 3554
rect 6750 3502 6802 3554
rect 11230 3502 11282 3554
rect 14590 3502 14642 3554
rect 15598 3502 15650 3554
rect 7646 3390 7698 3442
rect 8430 3278 8482 3330
rect 4210 3110 4262 3162
rect 4314 3110 4366 3162
rect 4418 3110 4470 3162
rect 8326 3110 8378 3162
rect 8430 3110 8482 3162
rect 8534 3110 8586 3162
rect 12442 3110 12494 3162
rect 12546 3110 12598 3162
rect 12650 3110 12702 3162
rect 16558 3110 16610 3162
rect 16662 3110 16714 3162
rect 16766 3110 16818 3162
rect 14814 2942 14866 2994
rect 15262 2942 15314 2994
rect 15822 2942 15874 2994
rect 4734 2718 4786 2770
rect 7422 2718 7474 2770
rect 8654 2718 8706 2770
rect 13806 2718 13858 2770
rect 2606 2606 2658 2658
rect 6526 2606 6578 2658
rect 11006 2606 11058 2658
rect 12014 2606 12066 2658
rect 2152 2326 2204 2378
rect 2256 2326 2308 2378
rect 2360 2326 2412 2378
rect 6268 2326 6320 2378
rect 6372 2326 6424 2378
rect 6476 2326 6528 2378
rect 10384 2326 10436 2378
rect 10488 2326 10540 2378
rect 10592 2326 10644 2378
rect 14500 2326 14552 2378
rect 14604 2326 14656 2378
rect 14708 2326 14760 2378
rect 3166 2046 3218 2098
rect 5070 2046 5122 2098
rect 8430 2046 8482 2098
rect 10558 2046 10610 2098
rect 12686 2046 12738 2098
rect 15486 2046 15538 2098
rect 814 1934 866 1986
rect 1598 1934 1650 1986
rect 6750 1934 6802 1986
rect 11678 1934 11730 1986
rect 15038 1934 15090 1986
rect 7646 1822 7698 1874
rect 4210 1542 4262 1594
rect 4314 1542 4366 1594
rect 4418 1542 4470 1594
rect 8326 1542 8378 1594
rect 8430 1542 8482 1594
rect 8534 1542 8586 1594
rect 12442 1542 12494 1594
rect 12546 1542 12598 1594
rect 12650 1542 12702 1594
rect 16558 1542 16610 1594
rect 16662 1542 16714 1594
rect 16766 1542 16818 1594
<< metal2 >>
rect 560 12200 672 13000
rect 1008 12200 1120 13000
rect 1456 12200 1568 13000
rect 1904 12200 2016 13000
rect 2352 12200 2464 13000
rect 2800 12200 2912 13000
rect 3248 12200 3360 13000
rect 3696 12200 3808 13000
rect 4144 12200 4256 13000
rect 4592 12200 4704 13000
rect 5040 12200 5152 13000
rect 5488 12200 5600 13000
rect 5936 12200 6048 13000
rect 6384 12200 6496 13000
rect 6832 12200 6944 13000
rect 7280 12200 7392 13000
rect 7728 12200 7840 13000
rect 8176 12200 8288 13000
rect 8624 12200 8736 13000
rect 9072 12200 9184 13000
rect 9520 12200 9632 13000
rect 9968 12200 10080 13000
rect 10416 12200 10528 13000
rect 10864 12200 10976 13000
rect 11312 12200 11424 13000
rect 11760 12200 11872 13000
rect 12208 12200 12320 13000
rect 12656 12200 12768 13000
rect 13104 12200 13216 13000
rect 13552 12200 13664 13000
rect 14000 12200 14112 13000
rect 14448 12200 14560 13000
rect 14896 12200 15008 13000
rect 15344 12200 15456 13000
rect 15792 12200 15904 13000
rect 16240 12200 16352 13000
rect 588 8428 644 12200
rect 588 8372 980 8428
rect 924 8370 980 8372
rect 924 8318 926 8370
rect 978 8318 980 8370
rect 924 8306 980 8318
rect 588 8260 644 8270
rect 588 800 644 8204
rect 1036 7362 1092 12200
rect 1484 10722 1540 12200
rect 1484 10670 1486 10722
rect 1538 10670 1540 10722
rect 1484 10658 1540 10670
rect 1036 7310 1038 7362
rect 1090 7310 1092 7362
rect 1036 7298 1092 7310
rect 1372 10612 1428 10622
rect 1036 6916 1092 6926
rect 812 1988 868 1998
rect 812 1894 868 1932
rect 1036 800 1092 6860
rect 1372 4228 1428 10556
rect 1932 8930 1988 12200
rect 2380 10724 2436 12200
rect 2380 10668 2548 10724
rect 2150 10220 2414 10230
rect 2206 10164 2254 10220
rect 2310 10164 2358 10220
rect 2150 10154 2414 10164
rect 2492 9938 2548 10668
rect 2716 10612 2772 10622
rect 2716 10518 2772 10556
rect 2492 9886 2494 9938
rect 2546 9886 2548 9938
rect 2492 9874 2548 9886
rect 1932 8878 1934 8930
rect 1986 8878 1988 8930
rect 1932 8866 1988 8878
rect 2492 9716 2548 9726
rect 2150 8652 2414 8662
rect 2206 8596 2254 8652
rect 2310 8596 2358 8652
rect 2150 8586 2414 8596
rect 1932 8484 1988 8494
rect 1372 4172 1540 4228
rect 1484 800 1540 4172
rect 1596 1988 1652 1998
rect 1596 1894 1652 1932
rect 1932 800 1988 8428
rect 2150 7084 2414 7094
rect 2206 7028 2254 7084
rect 2310 7028 2358 7084
rect 2150 7018 2414 7028
rect 2150 5516 2414 5526
rect 2206 5460 2254 5516
rect 2310 5460 2358 5516
rect 2150 5450 2414 5460
rect 2150 3948 2414 3958
rect 2206 3892 2254 3948
rect 2310 3892 2358 3948
rect 2150 3882 2414 3892
rect 2150 2380 2414 2390
rect 2206 2324 2254 2380
rect 2310 2324 2358 2380
rect 2150 2314 2414 2324
rect 2492 2212 2548 9660
rect 2716 8260 2772 8270
rect 2716 8166 2772 8204
rect 2716 7474 2772 7486
rect 2716 7422 2718 7474
rect 2770 7422 2772 7474
rect 2716 7364 2772 7422
rect 2716 6916 2772 7308
rect 2716 6850 2772 6860
rect 2604 5572 2660 5582
rect 2604 2658 2660 5516
rect 2828 4226 2884 12200
rect 3276 10388 3332 12200
rect 3724 10724 3780 12200
rect 4172 11172 4228 12200
rect 3052 10332 3332 10388
rect 3612 10668 3780 10724
rect 4060 11116 4228 11172
rect 2940 9042 2996 9054
rect 2940 8990 2942 9042
rect 2994 8990 2996 9042
rect 2940 8932 2996 8990
rect 2940 8484 2996 8876
rect 2940 8418 2996 8428
rect 2828 4174 2830 4226
rect 2882 4174 2884 4226
rect 2828 4162 2884 4174
rect 2716 3668 2772 3678
rect 3052 3668 3108 10332
rect 3388 9826 3444 9838
rect 3388 9774 3390 9826
rect 3442 9774 3444 9826
rect 3388 9716 3444 9774
rect 3388 9650 3444 9660
rect 3612 5794 3668 10668
rect 3724 10500 3780 10510
rect 3724 10406 3780 10444
rect 3948 8932 4004 8942
rect 3948 8838 4004 8876
rect 3724 8260 3780 8270
rect 3724 8166 3780 8204
rect 3724 7364 3780 7374
rect 3724 7270 3780 7308
rect 3612 5742 3614 5794
rect 3666 5742 3668 5794
rect 3612 5730 3668 5742
rect 3724 5908 3780 5918
rect 2716 3666 3108 3668
rect 2716 3614 2718 3666
rect 2770 3614 3108 3666
rect 2716 3612 3108 3614
rect 3164 5124 3220 5134
rect 2716 3602 2772 3612
rect 2604 2606 2606 2658
rect 2658 2606 2660 2658
rect 2604 2594 2660 2606
rect 2828 3444 2884 3454
rect 2380 2156 2548 2212
rect 2380 800 2436 2156
rect 2828 800 2884 3388
rect 3164 2098 3220 5068
rect 3388 4788 3444 4798
rect 3388 3556 3444 4732
rect 3164 2046 3166 2098
rect 3218 2046 3220 2098
rect 3164 2034 3220 2046
rect 3276 3554 3444 3556
rect 3276 3502 3390 3554
rect 3442 3502 3444 3554
rect 3276 3500 3444 3502
rect 3276 800 3332 3500
rect 3388 3490 3444 3500
rect 3724 800 3780 5852
rect 4060 5124 4116 11116
rect 4208 11004 4472 11014
rect 4264 10948 4312 11004
rect 4368 10948 4416 11004
rect 4208 10938 4472 10948
rect 4508 9716 4564 9726
rect 4508 9622 4564 9660
rect 4208 9436 4472 9446
rect 4264 9380 4312 9436
rect 4368 9380 4416 9436
rect 4208 9370 4472 9380
rect 4208 7868 4472 7878
rect 4264 7812 4312 7868
rect 4368 7812 4416 7868
rect 4208 7802 4472 7812
rect 4208 6300 4472 6310
rect 4264 6244 4312 6300
rect 4368 6244 4416 6300
rect 4208 6234 4472 6244
rect 4620 5572 4676 12200
rect 4732 10612 4788 10622
rect 4732 10518 4788 10556
rect 4732 5908 4788 5918
rect 4732 5814 4788 5852
rect 4620 5506 4676 5516
rect 4060 5058 4116 5068
rect 3836 4898 3892 4910
rect 3836 4846 3838 4898
rect 3890 4846 3892 4898
rect 3836 4788 3892 4846
rect 3836 4722 3892 4732
rect 3948 4900 4004 4910
rect 3948 4338 4004 4844
rect 4508 4900 4564 4938
rect 4508 4834 4564 4844
rect 4956 4898 5012 4910
rect 4956 4846 4958 4898
rect 5010 4846 5012 4898
rect 4208 4732 4472 4742
rect 4264 4676 4312 4732
rect 4368 4676 4416 4732
rect 4208 4666 4472 4676
rect 3948 4286 3950 4338
rect 4002 4286 4004 4338
rect 3948 3444 4004 4286
rect 3948 3378 4004 3388
rect 4208 3164 4472 3174
rect 4264 3108 4312 3164
rect 4368 3108 4416 3164
rect 4208 3098 4472 3108
rect 4732 2772 4788 2782
rect 4956 2772 5012 4846
rect 4620 2770 5012 2772
rect 4620 2718 4734 2770
rect 4786 2718 5012 2770
rect 4620 2716 5012 2718
rect 4060 1988 4116 1998
rect 4060 1428 4116 1932
rect 4208 1596 4472 1606
rect 4264 1540 4312 1596
rect 4368 1540 4416 1596
rect 4208 1530 4472 1540
rect 4060 1372 4228 1428
rect 4172 800 4228 1372
rect 4620 800 4676 2716
rect 4732 2706 4788 2716
rect 5068 2098 5124 12200
rect 5516 3666 5572 12200
rect 5740 10612 5796 10622
rect 5740 10518 5796 10556
rect 5740 5908 5796 5918
rect 5740 5814 5796 5852
rect 5964 4226 6020 12200
rect 6412 10388 6468 12200
rect 6748 10612 6804 10622
rect 6412 10332 6692 10388
rect 6266 10220 6530 10230
rect 6322 10164 6370 10220
rect 6426 10164 6474 10220
rect 6266 10154 6530 10164
rect 6524 9268 6580 9278
rect 6524 8930 6580 9212
rect 6524 8878 6526 8930
rect 6578 8878 6580 8930
rect 6524 8866 6580 8878
rect 6266 8652 6530 8662
rect 6322 8596 6370 8652
rect 6426 8596 6474 8652
rect 6266 8586 6530 8596
rect 6266 7084 6530 7094
rect 6322 7028 6370 7084
rect 6426 7028 6474 7084
rect 6266 7018 6530 7028
rect 6266 5516 6530 5526
rect 6322 5460 6370 5516
rect 6426 5460 6474 5516
rect 6266 5450 6530 5460
rect 5964 4174 5966 4226
rect 6018 4174 6020 4226
rect 5964 4162 6020 4174
rect 6266 3948 6530 3958
rect 6322 3892 6370 3948
rect 6426 3892 6474 3948
rect 6266 3882 6530 3892
rect 5516 3614 5518 3666
rect 5570 3614 5572 3666
rect 5516 3602 5572 3614
rect 5964 3780 6020 3790
rect 6636 3780 6692 10332
rect 6748 8428 6804 10556
rect 6860 10498 6916 12200
rect 6860 10446 6862 10498
rect 6914 10446 6916 10498
rect 6860 10434 6916 10446
rect 7084 10052 7140 10062
rect 7084 9938 7140 9996
rect 7084 9886 7086 9938
rect 7138 9886 7140 9938
rect 7084 9874 7140 9886
rect 7308 9268 7364 12200
rect 7756 10052 7812 12200
rect 7756 9986 7812 9996
rect 7308 9202 7364 9212
rect 7756 9826 7812 9838
rect 7756 9774 7758 9826
rect 7810 9774 7812 9826
rect 7308 9042 7364 9054
rect 7308 8990 7310 9042
rect 7362 8990 7364 9042
rect 7308 8428 7364 8990
rect 6748 8372 6916 8428
rect 5068 2046 5070 2098
rect 5122 2046 5124 2098
rect 5068 2034 5124 2046
rect 5516 3444 5572 3454
rect 5068 1876 5124 1886
rect 5068 800 5124 1820
rect 5516 800 5572 3388
rect 5964 800 6020 3724
rect 6524 3724 6692 3780
rect 6524 2658 6580 3724
rect 6748 3554 6804 3566
rect 6748 3502 6750 3554
rect 6802 3502 6804 3554
rect 6748 3444 6804 3502
rect 6748 3378 6804 3388
rect 6524 2606 6526 2658
rect 6578 2606 6580 2658
rect 6524 2594 6580 2606
rect 6266 2380 6530 2390
rect 6322 2324 6370 2380
rect 6426 2324 6474 2380
rect 6266 2314 6530 2324
rect 6412 2100 6468 2110
rect 6412 800 6468 2044
rect 6748 1986 6804 1998
rect 6748 1934 6750 1986
rect 6802 1934 6804 1986
rect 6748 1876 6804 1934
rect 6748 1810 6804 1820
rect 6860 800 6916 8372
rect 7084 8372 7364 8428
rect 7084 8034 7140 8372
rect 7084 7982 7086 8034
rect 7138 7982 7140 8034
rect 6972 4338 7028 4350
rect 6972 4286 6974 4338
rect 7026 4286 7028 4338
rect 6972 4228 7028 4286
rect 6972 3780 7028 4172
rect 6972 3714 7028 3724
rect 7084 2548 7140 7982
rect 7756 7364 7812 9774
rect 7644 3444 7700 3454
rect 7644 3350 7700 3388
rect 7420 2770 7476 2782
rect 7420 2718 7422 2770
rect 7474 2718 7476 2770
rect 7084 2492 7364 2548
rect 7308 800 7364 2492
rect 7420 2100 7476 2718
rect 7420 2034 7476 2044
rect 7644 1876 7700 1886
rect 7644 1782 7700 1820
rect 7756 800 7812 7308
rect 8204 6802 8260 12200
rect 8324 11004 8588 11014
rect 8380 10948 8428 11004
rect 8484 10948 8532 11004
rect 8324 10938 8588 10948
rect 8324 9436 8588 9446
rect 8380 9380 8428 9436
rect 8484 9380 8532 9436
rect 8324 9370 8588 9380
rect 8652 8260 8708 12200
rect 9100 11170 9156 12200
rect 9100 11118 9102 11170
rect 9154 11118 9156 11170
rect 9100 11106 9156 11118
rect 9100 10498 9156 10510
rect 9100 10446 9102 10498
rect 9154 10446 9156 10498
rect 8652 8194 8708 8204
rect 8764 8370 8820 8382
rect 8764 8318 8766 8370
rect 8818 8318 8820 8370
rect 8324 7868 8588 7878
rect 8380 7812 8428 7868
rect 8484 7812 8532 7868
rect 8324 7802 8588 7812
rect 8540 7364 8596 7374
rect 8540 7270 8596 7308
rect 8204 6750 8206 6802
rect 8258 6750 8260 6802
rect 8204 6738 8260 6750
rect 8324 6300 8588 6310
rect 8380 6244 8428 6300
rect 8484 6244 8532 6300
rect 8324 6234 8588 6244
rect 8204 6020 8260 6030
rect 8204 800 8260 5964
rect 8324 4732 8588 4742
rect 8380 4676 8428 4732
rect 8484 4676 8532 4732
rect 8324 4666 8588 4676
rect 8540 4228 8596 4238
rect 8540 4134 8596 4172
rect 8428 3332 8484 3342
rect 8428 3330 8708 3332
rect 8428 3278 8430 3330
rect 8482 3278 8708 3330
rect 8428 3276 8708 3278
rect 8428 3266 8484 3276
rect 8324 3164 8588 3174
rect 8380 3108 8428 3164
rect 8484 3108 8532 3164
rect 8324 3098 8588 3108
rect 8652 2770 8708 3276
rect 8652 2718 8654 2770
rect 8706 2718 8708 2770
rect 8652 2212 8708 2718
rect 8652 2146 8708 2156
rect 8428 2100 8484 2110
rect 8428 2006 8484 2044
rect 8764 1988 8820 8318
rect 8652 1932 8820 1988
rect 8324 1596 8588 1606
rect 8380 1540 8428 1596
rect 8484 1540 8532 1596
rect 8324 1530 8588 1540
rect 8652 800 8708 1932
rect 9100 800 9156 10446
rect 9548 9940 9604 12200
rect 9548 9874 9604 9884
rect 9548 9714 9604 9726
rect 9548 9662 9550 9714
rect 9602 9662 9604 9714
rect 9212 6690 9268 6702
rect 9212 6638 9214 6690
rect 9266 6638 9268 6690
rect 9212 6468 9268 6638
rect 9212 6020 9268 6412
rect 9212 5954 9268 5964
rect 9548 800 9604 9662
rect 9996 9044 10052 12200
rect 10444 10388 10500 12200
rect 10556 11170 10612 11182
rect 10556 11118 10558 11170
rect 10610 11118 10612 11170
rect 10556 10610 10612 11118
rect 10556 10558 10558 10610
rect 10610 10558 10612 10610
rect 10556 10546 10612 10558
rect 9996 8978 10052 8988
rect 10108 10332 10500 10388
rect 9884 8930 9940 8942
rect 9884 8878 9886 8930
rect 9938 8878 9940 8930
rect 9660 8260 9716 8270
rect 9660 8166 9716 8204
rect 9884 3220 9940 8878
rect 10108 5236 10164 10332
rect 10382 10220 10646 10230
rect 10438 10164 10486 10220
rect 10542 10164 10590 10220
rect 10382 10154 10646 10164
rect 10780 9940 10836 9950
rect 10780 9826 10836 9884
rect 10780 9774 10782 9826
rect 10834 9774 10836 9826
rect 10780 9762 10836 9774
rect 10382 8652 10646 8662
rect 10438 8596 10486 8652
rect 10542 8596 10590 8652
rect 10382 8586 10646 8596
rect 10892 8428 10948 12200
rect 11004 9044 11060 9054
rect 11004 8950 11060 8988
rect 10892 8372 11284 8428
rect 10668 8260 10724 8270
rect 10668 8166 10724 8204
rect 10382 7084 10646 7094
rect 10438 7028 10486 7084
rect 10542 7028 10590 7084
rect 10382 7018 10646 7028
rect 10220 6468 10276 6478
rect 10220 6374 10276 6412
rect 10382 5516 10646 5526
rect 10438 5460 10486 5516
rect 10542 5460 10590 5516
rect 10382 5450 10646 5460
rect 10108 5170 10164 5180
rect 11228 5236 11284 8372
rect 11340 6804 11396 12200
rect 11564 11170 11620 11182
rect 11564 11118 11566 11170
rect 11618 11118 11620 11170
rect 11564 10834 11620 11118
rect 11564 10782 11566 10834
rect 11618 10782 11620 10834
rect 11564 10770 11620 10782
rect 11788 10388 11844 12200
rect 11788 10332 11956 10388
rect 11788 9940 11844 9950
rect 11788 9846 11844 9884
rect 11340 6738 11396 6748
rect 11564 5796 11620 5806
rect 11564 5702 11620 5740
rect 11340 5236 11396 5246
rect 11788 5236 11844 5246
rect 11228 5234 11396 5236
rect 11228 5182 11342 5234
rect 11394 5182 11396 5234
rect 11228 5180 11396 5182
rect 10220 4226 10276 4238
rect 10220 4174 10222 4226
rect 10274 4174 10276 4226
rect 9884 3164 10052 3220
rect 9996 800 10052 3164
rect 10220 2100 10276 4174
rect 10382 3948 10646 3958
rect 10438 3892 10486 3948
rect 10542 3892 10590 3948
rect 10382 3882 10646 3892
rect 10668 3668 10724 3678
rect 10668 3666 10948 3668
rect 10668 3614 10670 3666
rect 10722 3614 10948 3666
rect 10668 3612 10948 3614
rect 10668 3602 10724 3612
rect 10382 2380 10646 2390
rect 10438 2324 10486 2380
rect 10542 2324 10590 2380
rect 10382 2314 10646 2324
rect 10556 2100 10612 2110
rect 10220 2044 10500 2100
rect 10444 800 10500 2044
rect 10556 2006 10612 2044
rect 10892 800 10948 3612
rect 11228 3554 11284 5180
rect 11340 5170 11396 5180
rect 11676 5180 11788 5236
rect 11676 4338 11732 5180
rect 11788 5142 11844 5180
rect 11676 4286 11678 4338
rect 11730 4286 11732 4338
rect 11676 4274 11732 4286
rect 11228 3502 11230 3554
rect 11282 3502 11284 3554
rect 11228 3490 11284 3502
rect 11900 3332 11956 10332
rect 12012 9044 12068 9054
rect 12012 8950 12068 8988
rect 12236 3892 12292 12200
rect 12684 11172 12740 12200
rect 12684 11116 12852 11172
rect 12440 11004 12704 11014
rect 12496 10948 12544 11004
rect 12600 10948 12648 11004
rect 12440 10938 12704 10948
rect 12348 10724 12404 10734
rect 12348 9828 12404 10668
rect 12572 9828 12628 9838
rect 12348 9826 12628 9828
rect 12348 9774 12574 9826
rect 12626 9774 12628 9826
rect 12348 9772 12628 9774
rect 12572 9762 12628 9772
rect 12440 9436 12704 9446
rect 12496 9380 12544 9436
rect 12600 9380 12648 9436
rect 12440 9370 12704 9380
rect 12440 7868 12704 7878
rect 12496 7812 12544 7868
rect 12600 7812 12648 7868
rect 12440 7802 12704 7812
rect 12440 6300 12704 6310
rect 12496 6244 12544 6300
rect 12600 6244 12648 6300
rect 12440 6234 12704 6244
rect 12684 5908 12740 5918
rect 12684 5814 12740 5852
rect 12572 5684 12628 5694
rect 12572 5234 12628 5628
rect 12572 5182 12574 5234
rect 12626 5182 12628 5234
rect 12572 5170 12628 5182
rect 12796 4900 12852 11116
rect 13020 5908 13076 5918
rect 13020 5234 13076 5852
rect 13020 5182 13022 5234
rect 13074 5182 13076 5234
rect 13020 5170 13076 5182
rect 12796 4834 12852 4844
rect 12440 4732 12704 4742
rect 12496 4676 12544 4732
rect 12600 4676 12648 4732
rect 12440 4666 12704 4676
rect 12796 4226 12852 4238
rect 12796 4174 12798 4226
rect 12850 4174 12852 4226
rect 12236 3836 12404 3892
rect 11900 3266 11956 3276
rect 12236 3668 12292 3678
rect 11004 2658 11060 2670
rect 11004 2606 11006 2658
rect 11058 2606 11060 2658
rect 11004 2212 11060 2606
rect 11004 2146 11060 2156
rect 11340 2660 11396 2670
rect 11340 800 11396 2604
rect 12012 2660 12068 2670
rect 12012 2566 12068 2604
rect 11676 2324 11732 2334
rect 11676 1986 11732 2268
rect 11676 1934 11678 1986
rect 11730 1934 11732 1986
rect 11676 1922 11732 1934
rect 11788 1764 11844 1774
rect 11788 800 11844 1708
rect 12236 800 12292 3612
rect 12348 3556 12404 3836
rect 12348 3490 12404 3500
rect 12440 3164 12704 3174
rect 12496 3108 12544 3164
rect 12600 3108 12648 3164
rect 12440 3098 12704 3108
rect 12684 2098 12740 2110
rect 12684 2046 12686 2098
rect 12738 2046 12740 2098
rect 12684 1764 12740 2046
rect 12684 1698 12740 1708
rect 12440 1596 12704 1606
rect 12496 1540 12544 1596
rect 12600 1540 12648 1596
rect 12440 1530 12704 1540
rect 12796 1428 12852 4174
rect 12908 3668 12964 3678
rect 12908 3574 12964 3612
rect 13132 2548 13188 12200
rect 13580 7812 13636 12200
rect 14028 10388 14084 12200
rect 14476 11170 14532 12200
rect 14476 11118 14478 11170
rect 14530 11118 14532 11170
rect 14476 11106 14532 11118
rect 14364 10724 14420 10734
rect 14252 10498 14308 10510
rect 14252 10446 14254 10498
rect 14306 10446 14308 10498
rect 14028 10332 14196 10388
rect 13580 7746 13636 7756
rect 13580 7362 13636 7374
rect 13580 7310 13582 7362
rect 13634 7310 13636 7362
rect 13244 5906 13300 5918
rect 13244 5854 13246 5906
rect 13298 5854 13300 5906
rect 13244 5684 13300 5854
rect 13244 5618 13300 5628
rect 13132 2324 13188 2492
rect 13132 2258 13188 2268
rect 12684 1372 12852 1428
rect 13132 2100 13188 2110
rect 12684 800 12740 1372
rect 13132 800 13188 2044
rect 13580 800 13636 7310
rect 13804 6804 13860 6814
rect 13804 2996 13860 6748
rect 13804 2770 13860 2940
rect 13804 2718 13806 2770
rect 13858 2718 13860 2770
rect 13804 2706 13860 2718
rect 14028 6802 14084 6814
rect 14028 6750 14030 6802
rect 14082 6750 14084 6802
rect 14028 800 14084 6750
rect 14140 6580 14196 10332
rect 14140 6514 14196 6524
rect 14252 1764 14308 10446
rect 14364 9938 14420 10668
rect 14498 10220 14762 10230
rect 14554 10164 14602 10220
rect 14658 10164 14706 10220
rect 14498 10154 14762 10164
rect 14364 9886 14366 9938
rect 14418 9886 14420 9938
rect 14364 9874 14420 9886
rect 14924 9716 14980 12200
rect 15148 11170 15204 11182
rect 15148 11118 15150 11170
rect 15202 11118 15204 11170
rect 15148 10610 15204 11118
rect 15148 10558 15150 10610
rect 15202 10558 15204 10610
rect 15148 9940 15204 10558
rect 15372 10052 15428 12200
rect 15372 10050 15540 10052
rect 15372 9998 15374 10050
rect 15426 9998 15540 10050
rect 15372 9996 15540 9998
rect 15372 9986 15428 9996
rect 15148 9874 15204 9884
rect 14924 9660 15092 9716
rect 14700 8932 14756 8942
rect 14700 8838 14756 8876
rect 14498 8652 14762 8662
rect 14554 8596 14602 8652
rect 14658 8596 14706 8652
rect 14498 8586 14762 8596
rect 14924 8370 14980 8382
rect 14924 8318 14926 8370
rect 14978 8318 14980 8370
rect 14476 7812 14532 7822
rect 14476 7474 14532 7756
rect 14476 7422 14478 7474
rect 14530 7422 14532 7474
rect 14476 7410 14532 7422
rect 14498 7084 14762 7094
rect 14554 7028 14602 7084
rect 14658 7028 14706 7084
rect 14498 7018 14762 7028
rect 14498 5516 14762 5526
rect 14554 5460 14602 5516
rect 14658 5460 14706 5516
rect 14498 5450 14762 5460
rect 14924 5460 14980 8318
rect 15036 6692 15092 9660
rect 15484 9042 15540 9996
rect 15596 9940 15652 9950
rect 15596 9846 15652 9884
rect 15484 8990 15486 9042
rect 15538 8990 15540 9042
rect 15484 8978 15540 8990
rect 15036 6626 15092 6636
rect 15372 8932 15428 8942
rect 15036 6468 15092 6478
rect 15036 6018 15092 6412
rect 15036 5966 15038 6018
rect 15090 5966 15092 6018
rect 15036 5954 15092 5966
rect 14924 5394 14980 5404
rect 14924 5234 14980 5246
rect 14924 5182 14926 5234
rect 14978 5182 14980 5234
rect 14588 4900 14644 4910
rect 14588 4338 14644 4844
rect 14588 4286 14590 4338
rect 14642 4286 14644 4338
rect 14588 4116 14644 4286
rect 14588 4050 14644 4060
rect 14498 3948 14762 3958
rect 14554 3892 14602 3948
rect 14658 3892 14706 3948
rect 14498 3882 14762 3892
rect 14588 3556 14644 3566
rect 14588 3462 14644 3500
rect 14812 2996 14868 3006
rect 14812 2902 14868 2940
rect 14498 2380 14762 2390
rect 14554 2324 14602 2380
rect 14658 2324 14706 2380
rect 14498 2314 14762 2324
rect 14252 1708 14532 1764
rect 14476 800 14532 1708
rect 14924 800 14980 5182
rect 15260 3332 15316 3342
rect 15260 2994 15316 3276
rect 15260 2942 15262 2994
rect 15314 2942 15316 2994
rect 15036 1988 15092 1998
rect 15260 1988 15316 2942
rect 15036 1986 15316 1988
rect 15036 1934 15038 1986
rect 15090 1934 15316 1986
rect 15036 1932 15316 1934
rect 15036 1922 15092 1932
rect 15372 800 15428 8876
rect 15484 7812 15540 7822
rect 15484 7698 15540 7756
rect 15484 7646 15486 7698
rect 15538 7646 15540 7698
rect 15484 7634 15540 7646
rect 15484 6690 15540 6702
rect 15484 6638 15486 6690
rect 15538 6638 15540 6690
rect 15484 6580 15540 6638
rect 15484 4564 15540 6524
rect 15596 6692 15652 6702
rect 15596 5124 15652 6636
rect 15820 5908 15876 12200
rect 16044 10050 16100 10062
rect 16044 9998 16046 10050
rect 16098 9998 16100 10050
rect 16044 9938 16100 9998
rect 16044 9886 16046 9938
rect 16098 9886 16100 9938
rect 16044 9874 16100 9886
rect 16156 8260 16212 8270
rect 16268 8260 16324 12200
rect 16556 11004 16820 11014
rect 16612 10948 16660 11004
rect 16716 10948 16764 11004
rect 16556 10938 16820 10948
rect 16556 9436 16820 9446
rect 16612 9380 16660 9436
rect 16716 9380 16764 9436
rect 16556 9370 16820 9380
rect 16156 8258 16324 8260
rect 16156 8206 16158 8258
rect 16210 8206 16324 8258
rect 16156 8204 16324 8206
rect 16156 8194 16212 8204
rect 16268 6802 16324 8204
rect 16556 7868 16820 7878
rect 16612 7812 16660 7868
rect 16716 7812 16764 7868
rect 16556 7802 16820 7812
rect 16268 6750 16270 6802
rect 16322 6750 16324 6802
rect 16268 6738 16324 6750
rect 16556 6300 16820 6310
rect 16612 6244 16660 6300
rect 16716 6244 16764 6300
rect 16556 6234 16820 6244
rect 15820 5842 15876 5852
rect 15932 5796 15988 5806
rect 15596 5122 15876 5124
rect 15596 5070 15598 5122
rect 15650 5070 15876 5122
rect 15596 5068 15876 5070
rect 15596 5058 15652 5068
rect 15708 4564 15764 4574
rect 15484 4562 15764 4564
rect 15484 4510 15710 4562
rect 15762 4510 15764 4562
rect 15484 4508 15764 4510
rect 15708 4498 15764 4508
rect 15596 3556 15652 3566
rect 15596 3462 15652 3500
rect 15820 2994 15876 5068
rect 15820 2942 15822 2994
rect 15874 2942 15876 2994
rect 15820 2930 15876 2942
rect 15932 2772 15988 5740
rect 16268 5460 16324 5470
rect 16044 4116 16100 4126
rect 16044 3666 16100 4060
rect 16044 3614 16046 3666
rect 16098 3614 16100 3666
rect 16044 3602 16100 3614
rect 15820 2716 15988 2772
rect 15484 2548 15540 2558
rect 15484 2098 15540 2492
rect 15484 2046 15486 2098
rect 15538 2046 15540 2098
rect 15484 2034 15540 2046
rect 15820 800 15876 2716
rect 16268 800 16324 5404
rect 16556 4732 16820 4742
rect 16612 4676 16660 4732
rect 16716 4676 16764 4732
rect 16556 4666 16820 4676
rect 16556 3164 16820 3174
rect 16612 3108 16660 3164
rect 16716 3108 16764 3164
rect 16556 3098 16820 3108
rect 16556 1596 16820 1606
rect 16612 1540 16660 1596
rect 16716 1540 16764 1596
rect 16556 1530 16820 1540
rect 560 0 672 800
rect 1008 0 1120 800
rect 1456 0 1568 800
rect 1904 0 2016 800
rect 2352 0 2464 800
rect 2800 0 2912 800
rect 3248 0 3360 800
rect 3696 0 3808 800
rect 4144 0 4256 800
rect 4592 0 4704 800
rect 5040 0 5152 800
rect 5488 0 5600 800
rect 5936 0 6048 800
rect 6384 0 6496 800
rect 6832 0 6944 800
rect 7280 0 7392 800
rect 7728 0 7840 800
rect 8176 0 8288 800
rect 8624 0 8736 800
rect 9072 0 9184 800
rect 9520 0 9632 800
rect 9968 0 10080 800
rect 10416 0 10528 800
rect 10864 0 10976 800
rect 11312 0 11424 800
rect 11760 0 11872 800
rect 12208 0 12320 800
rect 12656 0 12768 800
rect 13104 0 13216 800
rect 13552 0 13664 800
rect 14000 0 14112 800
rect 14448 0 14560 800
rect 14896 0 15008 800
rect 15344 0 15456 800
rect 15792 0 15904 800
rect 16240 0 16352 800
<< via2 >>
rect 588 8204 644 8260
rect 1372 10556 1428 10612
rect 1036 6860 1092 6916
rect 812 1986 868 1988
rect 812 1934 814 1986
rect 814 1934 866 1986
rect 866 1934 868 1986
rect 812 1932 868 1934
rect 2150 10218 2206 10220
rect 2150 10166 2152 10218
rect 2152 10166 2204 10218
rect 2204 10166 2206 10218
rect 2150 10164 2206 10166
rect 2254 10218 2310 10220
rect 2254 10166 2256 10218
rect 2256 10166 2308 10218
rect 2308 10166 2310 10218
rect 2254 10164 2310 10166
rect 2358 10218 2414 10220
rect 2358 10166 2360 10218
rect 2360 10166 2412 10218
rect 2412 10166 2414 10218
rect 2358 10164 2414 10166
rect 2716 10610 2772 10612
rect 2716 10558 2718 10610
rect 2718 10558 2770 10610
rect 2770 10558 2772 10610
rect 2716 10556 2772 10558
rect 2492 9660 2548 9716
rect 2150 8650 2206 8652
rect 2150 8598 2152 8650
rect 2152 8598 2204 8650
rect 2204 8598 2206 8650
rect 2150 8596 2206 8598
rect 2254 8650 2310 8652
rect 2254 8598 2256 8650
rect 2256 8598 2308 8650
rect 2308 8598 2310 8650
rect 2254 8596 2310 8598
rect 2358 8650 2414 8652
rect 2358 8598 2360 8650
rect 2360 8598 2412 8650
rect 2412 8598 2414 8650
rect 2358 8596 2414 8598
rect 1932 8428 1988 8484
rect 1596 1986 1652 1988
rect 1596 1934 1598 1986
rect 1598 1934 1650 1986
rect 1650 1934 1652 1986
rect 1596 1932 1652 1934
rect 2150 7082 2206 7084
rect 2150 7030 2152 7082
rect 2152 7030 2204 7082
rect 2204 7030 2206 7082
rect 2150 7028 2206 7030
rect 2254 7082 2310 7084
rect 2254 7030 2256 7082
rect 2256 7030 2308 7082
rect 2308 7030 2310 7082
rect 2254 7028 2310 7030
rect 2358 7082 2414 7084
rect 2358 7030 2360 7082
rect 2360 7030 2412 7082
rect 2412 7030 2414 7082
rect 2358 7028 2414 7030
rect 2150 5514 2206 5516
rect 2150 5462 2152 5514
rect 2152 5462 2204 5514
rect 2204 5462 2206 5514
rect 2150 5460 2206 5462
rect 2254 5514 2310 5516
rect 2254 5462 2256 5514
rect 2256 5462 2308 5514
rect 2308 5462 2310 5514
rect 2254 5460 2310 5462
rect 2358 5514 2414 5516
rect 2358 5462 2360 5514
rect 2360 5462 2412 5514
rect 2412 5462 2414 5514
rect 2358 5460 2414 5462
rect 2150 3946 2206 3948
rect 2150 3894 2152 3946
rect 2152 3894 2204 3946
rect 2204 3894 2206 3946
rect 2150 3892 2206 3894
rect 2254 3946 2310 3948
rect 2254 3894 2256 3946
rect 2256 3894 2308 3946
rect 2308 3894 2310 3946
rect 2254 3892 2310 3894
rect 2358 3946 2414 3948
rect 2358 3894 2360 3946
rect 2360 3894 2412 3946
rect 2412 3894 2414 3946
rect 2358 3892 2414 3894
rect 2150 2378 2206 2380
rect 2150 2326 2152 2378
rect 2152 2326 2204 2378
rect 2204 2326 2206 2378
rect 2150 2324 2206 2326
rect 2254 2378 2310 2380
rect 2254 2326 2256 2378
rect 2256 2326 2308 2378
rect 2308 2326 2310 2378
rect 2254 2324 2310 2326
rect 2358 2378 2414 2380
rect 2358 2326 2360 2378
rect 2360 2326 2412 2378
rect 2412 2326 2414 2378
rect 2358 2324 2414 2326
rect 2716 8258 2772 8260
rect 2716 8206 2718 8258
rect 2718 8206 2770 8258
rect 2770 8206 2772 8258
rect 2716 8204 2772 8206
rect 2716 7308 2772 7364
rect 2716 6860 2772 6916
rect 2604 5516 2660 5572
rect 2940 8876 2996 8932
rect 2940 8428 2996 8484
rect 3388 9660 3444 9716
rect 3724 10498 3780 10500
rect 3724 10446 3726 10498
rect 3726 10446 3778 10498
rect 3778 10446 3780 10498
rect 3724 10444 3780 10446
rect 3948 8930 4004 8932
rect 3948 8878 3950 8930
rect 3950 8878 4002 8930
rect 4002 8878 4004 8930
rect 3948 8876 4004 8878
rect 3724 8258 3780 8260
rect 3724 8206 3726 8258
rect 3726 8206 3778 8258
rect 3778 8206 3780 8258
rect 3724 8204 3780 8206
rect 3724 7362 3780 7364
rect 3724 7310 3726 7362
rect 3726 7310 3778 7362
rect 3778 7310 3780 7362
rect 3724 7308 3780 7310
rect 3724 5852 3780 5908
rect 3164 5068 3220 5124
rect 2828 3388 2884 3444
rect 3388 4732 3444 4788
rect 4208 11002 4264 11004
rect 4208 10950 4210 11002
rect 4210 10950 4262 11002
rect 4262 10950 4264 11002
rect 4208 10948 4264 10950
rect 4312 11002 4368 11004
rect 4312 10950 4314 11002
rect 4314 10950 4366 11002
rect 4366 10950 4368 11002
rect 4312 10948 4368 10950
rect 4416 11002 4472 11004
rect 4416 10950 4418 11002
rect 4418 10950 4470 11002
rect 4470 10950 4472 11002
rect 4416 10948 4472 10950
rect 4508 9714 4564 9716
rect 4508 9662 4510 9714
rect 4510 9662 4562 9714
rect 4562 9662 4564 9714
rect 4508 9660 4564 9662
rect 4208 9434 4264 9436
rect 4208 9382 4210 9434
rect 4210 9382 4262 9434
rect 4262 9382 4264 9434
rect 4208 9380 4264 9382
rect 4312 9434 4368 9436
rect 4312 9382 4314 9434
rect 4314 9382 4366 9434
rect 4366 9382 4368 9434
rect 4312 9380 4368 9382
rect 4416 9434 4472 9436
rect 4416 9382 4418 9434
rect 4418 9382 4470 9434
rect 4470 9382 4472 9434
rect 4416 9380 4472 9382
rect 4208 7866 4264 7868
rect 4208 7814 4210 7866
rect 4210 7814 4262 7866
rect 4262 7814 4264 7866
rect 4208 7812 4264 7814
rect 4312 7866 4368 7868
rect 4312 7814 4314 7866
rect 4314 7814 4366 7866
rect 4366 7814 4368 7866
rect 4312 7812 4368 7814
rect 4416 7866 4472 7868
rect 4416 7814 4418 7866
rect 4418 7814 4470 7866
rect 4470 7814 4472 7866
rect 4416 7812 4472 7814
rect 4208 6298 4264 6300
rect 4208 6246 4210 6298
rect 4210 6246 4262 6298
rect 4262 6246 4264 6298
rect 4208 6244 4264 6246
rect 4312 6298 4368 6300
rect 4312 6246 4314 6298
rect 4314 6246 4366 6298
rect 4366 6246 4368 6298
rect 4312 6244 4368 6246
rect 4416 6298 4472 6300
rect 4416 6246 4418 6298
rect 4418 6246 4470 6298
rect 4470 6246 4472 6298
rect 4416 6244 4472 6246
rect 4732 10610 4788 10612
rect 4732 10558 4734 10610
rect 4734 10558 4786 10610
rect 4786 10558 4788 10610
rect 4732 10556 4788 10558
rect 4732 5906 4788 5908
rect 4732 5854 4734 5906
rect 4734 5854 4786 5906
rect 4786 5854 4788 5906
rect 4732 5852 4788 5854
rect 4620 5516 4676 5572
rect 4060 5068 4116 5124
rect 3836 4732 3892 4788
rect 3948 4844 4004 4900
rect 4508 4898 4564 4900
rect 4508 4846 4510 4898
rect 4510 4846 4562 4898
rect 4562 4846 4564 4898
rect 4508 4844 4564 4846
rect 4208 4730 4264 4732
rect 4208 4678 4210 4730
rect 4210 4678 4262 4730
rect 4262 4678 4264 4730
rect 4208 4676 4264 4678
rect 4312 4730 4368 4732
rect 4312 4678 4314 4730
rect 4314 4678 4366 4730
rect 4366 4678 4368 4730
rect 4312 4676 4368 4678
rect 4416 4730 4472 4732
rect 4416 4678 4418 4730
rect 4418 4678 4470 4730
rect 4470 4678 4472 4730
rect 4416 4676 4472 4678
rect 3948 3388 4004 3444
rect 4208 3162 4264 3164
rect 4208 3110 4210 3162
rect 4210 3110 4262 3162
rect 4262 3110 4264 3162
rect 4208 3108 4264 3110
rect 4312 3162 4368 3164
rect 4312 3110 4314 3162
rect 4314 3110 4366 3162
rect 4366 3110 4368 3162
rect 4312 3108 4368 3110
rect 4416 3162 4472 3164
rect 4416 3110 4418 3162
rect 4418 3110 4470 3162
rect 4470 3110 4472 3162
rect 4416 3108 4472 3110
rect 4060 1932 4116 1988
rect 4208 1594 4264 1596
rect 4208 1542 4210 1594
rect 4210 1542 4262 1594
rect 4262 1542 4264 1594
rect 4208 1540 4264 1542
rect 4312 1594 4368 1596
rect 4312 1542 4314 1594
rect 4314 1542 4366 1594
rect 4366 1542 4368 1594
rect 4312 1540 4368 1542
rect 4416 1594 4472 1596
rect 4416 1542 4418 1594
rect 4418 1542 4470 1594
rect 4470 1542 4472 1594
rect 4416 1540 4472 1542
rect 5740 10610 5796 10612
rect 5740 10558 5742 10610
rect 5742 10558 5794 10610
rect 5794 10558 5796 10610
rect 5740 10556 5796 10558
rect 5740 5906 5796 5908
rect 5740 5854 5742 5906
rect 5742 5854 5794 5906
rect 5794 5854 5796 5906
rect 5740 5852 5796 5854
rect 6748 10556 6804 10612
rect 6266 10218 6322 10220
rect 6266 10166 6268 10218
rect 6268 10166 6320 10218
rect 6320 10166 6322 10218
rect 6266 10164 6322 10166
rect 6370 10218 6426 10220
rect 6370 10166 6372 10218
rect 6372 10166 6424 10218
rect 6424 10166 6426 10218
rect 6370 10164 6426 10166
rect 6474 10218 6530 10220
rect 6474 10166 6476 10218
rect 6476 10166 6528 10218
rect 6528 10166 6530 10218
rect 6474 10164 6530 10166
rect 6524 9212 6580 9268
rect 6266 8650 6322 8652
rect 6266 8598 6268 8650
rect 6268 8598 6320 8650
rect 6320 8598 6322 8650
rect 6266 8596 6322 8598
rect 6370 8650 6426 8652
rect 6370 8598 6372 8650
rect 6372 8598 6424 8650
rect 6424 8598 6426 8650
rect 6370 8596 6426 8598
rect 6474 8650 6530 8652
rect 6474 8598 6476 8650
rect 6476 8598 6528 8650
rect 6528 8598 6530 8650
rect 6474 8596 6530 8598
rect 6266 7082 6322 7084
rect 6266 7030 6268 7082
rect 6268 7030 6320 7082
rect 6320 7030 6322 7082
rect 6266 7028 6322 7030
rect 6370 7082 6426 7084
rect 6370 7030 6372 7082
rect 6372 7030 6424 7082
rect 6424 7030 6426 7082
rect 6370 7028 6426 7030
rect 6474 7082 6530 7084
rect 6474 7030 6476 7082
rect 6476 7030 6528 7082
rect 6528 7030 6530 7082
rect 6474 7028 6530 7030
rect 6266 5514 6322 5516
rect 6266 5462 6268 5514
rect 6268 5462 6320 5514
rect 6320 5462 6322 5514
rect 6266 5460 6322 5462
rect 6370 5514 6426 5516
rect 6370 5462 6372 5514
rect 6372 5462 6424 5514
rect 6424 5462 6426 5514
rect 6370 5460 6426 5462
rect 6474 5514 6530 5516
rect 6474 5462 6476 5514
rect 6476 5462 6528 5514
rect 6528 5462 6530 5514
rect 6474 5460 6530 5462
rect 6266 3946 6322 3948
rect 6266 3894 6268 3946
rect 6268 3894 6320 3946
rect 6320 3894 6322 3946
rect 6266 3892 6322 3894
rect 6370 3946 6426 3948
rect 6370 3894 6372 3946
rect 6372 3894 6424 3946
rect 6424 3894 6426 3946
rect 6370 3892 6426 3894
rect 6474 3946 6530 3948
rect 6474 3894 6476 3946
rect 6476 3894 6528 3946
rect 6528 3894 6530 3946
rect 6474 3892 6530 3894
rect 7084 9996 7140 10052
rect 7756 9996 7812 10052
rect 7308 9212 7364 9268
rect 5964 3724 6020 3780
rect 5516 3388 5572 3444
rect 5068 1820 5124 1876
rect 6748 3388 6804 3444
rect 6266 2378 6322 2380
rect 6266 2326 6268 2378
rect 6268 2326 6320 2378
rect 6320 2326 6322 2378
rect 6266 2324 6322 2326
rect 6370 2378 6426 2380
rect 6370 2326 6372 2378
rect 6372 2326 6424 2378
rect 6424 2326 6426 2378
rect 6370 2324 6426 2326
rect 6474 2378 6530 2380
rect 6474 2326 6476 2378
rect 6476 2326 6528 2378
rect 6528 2326 6530 2378
rect 6474 2324 6530 2326
rect 6412 2044 6468 2100
rect 6748 1820 6804 1876
rect 6972 4172 7028 4228
rect 6972 3724 7028 3780
rect 7756 7308 7812 7364
rect 7644 3442 7700 3444
rect 7644 3390 7646 3442
rect 7646 3390 7698 3442
rect 7698 3390 7700 3442
rect 7644 3388 7700 3390
rect 7420 2044 7476 2100
rect 7644 1874 7700 1876
rect 7644 1822 7646 1874
rect 7646 1822 7698 1874
rect 7698 1822 7700 1874
rect 7644 1820 7700 1822
rect 8324 11002 8380 11004
rect 8324 10950 8326 11002
rect 8326 10950 8378 11002
rect 8378 10950 8380 11002
rect 8324 10948 8380 10950
rect 8428 11002 8484 11004
rect 8428 10950 8430 11002
rect 8430 10950 8482 11002
rect 8482 10950 8484 11002
rect 8428 10948 8484 10950
rect 8532 11002 8588 11004
rect 8532 10950 8534 11002
rect 8534 10950 8586 11002
rect 8586 10950 8588 11002
rect 8532 10948 8588 10950
rect 8324 9434 8380 9436
rect 8324 9382 8326 9434
rect 8326 9382 8378 9434
rect 8378 9382 8380 9434
rect 8324 9380 8380 9382
rect 8428 9434 8484 9436
rect 8428 9382 8430 9434
rect 8430 9382 8482 9434
rect 8482 9382 8484 9434
rect 8428 9380 8484 9382
rect 8532 9434 8588 9436
rect 8532 9382 8534 9434
rect 8534 9382 8586 9434
rect 8586 9382 8588 9434
rect 8532 9380 8588 9382
rect 8652 8204 8708 8260
rect 8324 7866 8380 7868
rect 8324 7814 8326 7866
rect 8326 7814 8378 7866
rect 8378 7814 8380 7866
rect 8324 7812 8380 7814
rect 8428 7866 8484 7868
rect 8428 7814 8430 7866
rect 8430 7814 8482 7866
rect 8482 7814 8484 7866
rect 8428 7812 8484 7814
rect 8532 7866 8588 7868
rect 8532 7814 8534 7866
rect 8534 7814 8586 7866
rect 8586 7814 8588 7866
rect 8532 7812 8588 7814
rect 8540 7362 8596 7364
rect 8540 7310 8542 7362
rect 8542 7310 8594 7362
rect 8594 7310 8596 7362
rect 8540 7308 8596 7310
rect 8324 6298 8380 6300
rect 8324 6246 8326 6298
rect 8326 6246 8378 6298
rect 8378 6246 8380 6298
rect 8324 6244 8380 6246
rect 8428 6298 8484 6300
rect 8428 6246 8430 6298
rect 8430 6246 8482 6298
rect 8482 6246 8484 6298
rect 8428 6244 8484 6246
rect 8532 6298 8588 6300
rect 8532 6246 8534 6298
rect 8534 6246 8586 6298
rect 8586 6246 8588 6298
rect 8532 6244 8588 6246
rect 8204 5964 8260 6020
rect 8324 4730 8380 4732
rect 8324 4678 8326 4730
rect 8326 4678 8378 4730
rect 8378 4678 8380 4730
rect 8324 4676 8380 4678
rect 8428 4730 8484 4732
rect 8428 4678 8430 4730
rect 8430 4678 8482 4730
rect 8482 4678 8484 4730
rect 8428 4676 8484 4678
rect 8532 4730 8588 4732
rect 8532 4678 8534 4730
rect 8534 4678 8586 4730
rect 8586 4678 8588 4730
rect 8532 4676 8588 4678
rect 8540 4226 8596 4228
rect 8540 4174 8542 4226
rect 8542 4174 8594 4226
rect 8594 4174 8596 4226
rect 8540 4172 8596 4174
rect 8324 3162 8380 3164
rect 8324 3110 8326 3162
rect 8326 3110 8378 3162
rect 8378 3110 8380 3162
rect 8324 3108 8380 3110
rect 8428 3162 8484 3164
rect 8428 3110 8430 3162
rect 8430 3110 8482 3162
rect 8482 3110 8484 3162
rect 8428 3108 8484 3110
rect 8532 3162 8588 3164
rect 8532 3110 8534 3162
rect 8534 3110 8586 3162
rect 8586 3110 8588 3162
rect 8532 3108 8588 3110
rect 8652 2156 8708 2212
rect 8428 2098 8484 2100
rect 8428 2046 8430 2098
rect 8430 2046 8482 2098
rect 8482 2046 8484 2098
rect 8428 2044 8484 2046
rect 8324 1594 8380 1596
rect 8324 1542 8326 1594
rect 8326 1542 8378 1594
rect 8378 1542 8380 1594
rect 8324 1540 8380 1542
rect 8428 1594 8484 1596
rect 8428 1542 8430 1594
rect 8430 1542 8482 1594
rect 8482 1542 8484 1594
rect 8428 1540 8484 1542
rect 8532 1594 8588 1596
rect 8532 1542 8534 1594
rect 8534 1542 8586 1594
rect 8586 1542 8588 1594
rect 8532 1540 8588 1542
rect 9548 9884 9604 9940
rect 9212 6412 9268 6468
rect 9212 5964 9268 6020
rect 9996 8988 10052 9044
rect 9660 8258 9716 8260
rect 9660 8206 9662 8258
rect 9662 8206 9714 8258
rect 9714 8206 9716 8258
rect 9660 8204 9716 8206
rect 10382 10218 10438 10220
rect 10382 10166 10384 10218
rect 10384 10166 10436 10218
rect 10436 10166 10438 10218
rect 10382 10164 10438 10166
rect 10486 10218 10542 10220
rect 10486 10166 10488 10218
rect 10488 10166 10540 10218
rect 10540 10166 10542 10218
rect 10486 10164 10542 10166
rect 10590 10218 10646 10220
rect 10590 10166 10592 10218
rect 10592 10166 10644 10218
rect 10644 10166 10646 10218
rect 10590 10164 10646 10166
rect 10780 9884 10836 9940
rect 10382 8650 10438 8652
rect 10382 8598 10384 8650
rect 10384 8598 10436 8650
rect 10436 8598 10438 8650
rect 10382 8596 10438 8598
rect 10486 8650 10542 8652
rect 10486 8598 10488 8650
rect 10488 8598 10540 8650
rect 10540 8598 10542 8650
rect 10486 8596 10542 8598
rect 10590 8650 10646 8652
rect 10590 8598 10592 8650
rect 10592 8598 10644 8650
rect 10644 8598 10646 8650
rect 10590 8596 10646 8598
rect 11004 9042 11060 9044
rect 11004 8990 11006 9042
rect 11006 8990 11058 9042
rect 11058 8990 11060 9042
rect 11004 8988 11060 8990
rect 10668 8258 10724 8260
rect 10668 8206 10670 8258
rect 10670 8206 10722 8258
rect 10722 8206 10724 8258
rect 10668 8204 10724 8206
rect 10382 7082 10438 7084
rect 10382 7030 10384 7082
rect 10384 7030 10436 7082
rect 10436 7030 10438 7082
rect 10382 7028 10438 7030
rect 10486 7082 10542 7084
rect 10486 7030 10488 7082
rect 10488 7030 10540 7082
rect 10540 7030 10542 7082
rect 10486 7028 10542 7030
rect 10590 7082 10646 7084
rect 10590 7030 10592 7082
rect 10592 7030 10644 7082
rect 10644 7030 10646 7082
rect 10590 7028 10646 7030
rect 10220 6466 10276 6468
rect 10220 6414 10222 6466
rect 10222 6414 10274 6466
rect 10274 6414 10276 6466
rect 10220 6412 10276 6414
rect 10382 5514 10438 5516
rect 10382 5462 10384 5514
rect 10384 5462 10436 5514
rect 10436 5462 10438 5514
rect 10382 5460 10438 5462
rect 10486 5514 10542 5516
rect 10486 5462 10488 5514
rect 10488 5462 10540 5514
rect 10540 5462 10542 5514
rect 10486 5460 10542 5462
rect 10590 5514 10646 5516
rect 10590 5462 10592 5514
rect 10592 5462 10644 5514
rect 10644 5462 10646 5514
rect 10590 5460 10646 5462
rect 10108 5180 10164 5236
rect 11788 9938 11844 9940
rect 11788 9886 11790 9938
rect 11790 9886 11842 9938
rect 11842 9886 11844 9938
rect 11788 9884 11844 9886
rect 11340 6748 11396 6804
rect 11564 5794 11620 5796
rect 11564 5742 11566 5794
rect 11566 5742 11618 5794
rect 11618 5742 11620 5794
rect 11564 5740 11620 5742
rect 10382 3946 10438 3948
rect 10382 3894 10384 3946
rect 10384 3894 10436 3946
rect 10436 3894 10438 3946
rect 10382 3892 10438 3894
rect 10486 3946 10542 3948
rect 10486 3894 10488 3946
rect 10488 3894 10540 3946
rect 10540 3894 10542 3946
rect 10486 3892 10542 3894
rect 10590 3946 10646 3948
rect 10590 3894 10592 3946
rect 10592 3894 10644 3946
rect 10644 3894 10646 3946
rect 10590 3892 10646 3894
rect 10382 2378 10438 2380
rect 10382 2326 10384 2378
rect 10384 2326 10436 2378
rect 10436 2326 10438 2378
rect 10382 2324 10438 2326
rect 10486 2378 10542 2380
rect 10486 2326 10488 2378
rect 10488 2326 10540 2378
rect 10540 2326 10542 2378
rect 10486 2324 10542 2326
rect 10590 2378 10646 2380
rect 10590 2326 10592 2378
rect 10592 2326 10644 2378
rect 10644 2326 10646 2378
rect 10590 2324 10646 2326
rect 10556 2098 10612 2100
rect 10556 2046 10558 2098
rect 10558 2046 10610 2098
rect 10610 2046 10612 2098
rect 10556 2044 10612 2046
rect 11788 5234 11844 5236
rect 11788 5182 11790 5234
rect 11790 5182 11842 5234
rect 11842 5182 11844 5234
rect 11788 5180 11844 5182
rect 12012 9042 12068 9044
rect 12012 8990 12014 9042
rect 12014 8990 12066 9042
rect 12066 8990 12068 9042
rect 12012 8988 12068 8990
rect 12440 11002 12496 11004
rect 12440 10950 12442 11002
rect 12442 10950 12494 11002
rect 12494 10950 12496 11002
rect 12440 10948 12496 10950
rect 12544 11002 12600 11004
rect 12544 10950 12546 11002
rect 12546 10950 12598 11002
rect 12598 10950 12600 11002
rect 12544 10948 12600 10950
rect 12648 11002 12704 11004
rect 12648 10950 12650 11002
rect 12650 10950 12702 11002
rect 12702 10950 12704 11002
rect 12648 10948 12704 10950
rect 12348 10722 12404 10724
rect 12348 10670 12350 10722
rect 12350 10670 12402 10722
rect 12402 10670 12404 10722
rect 12348 10668 12404 10670
rect 12440 9434 12496 9436
rect 12440 9382 12442 9434
rect 12442 9382 12494 9434
rect 12494 9382 12496 9434
rect 12440 9380 12496 9382
rect 12544 9434 12600 9436
rect 12544 9382 12546 9434
rect 12546 9382 12598 9434
rect 12598 9382 12600 9434
rect 12544 9380 12600 9382
rect 12648 9434 12704 9436
rect 12648 9382 12650 9434
rect 12650 9382 12702 9434
rect 12702 9382 12704 9434
rect 12648 9380 12704 9382
rect 12440 7866 12496 7868
rect 12440 7814 12442 7866
rect 12442 7814 12494 7866
rect 12494 7814 12496 7866
rect 12440 7812 12496 7814
rect 12544 7866 12600 7868
rect 12544 7814 12546 7866
rect 12546 7814 12598 7866
rect 12598 7814 12600 7866
rect 12544 7812 12600 7814
rect 12648 7866 12704 7868
rect 12648 7814 12650 7866
rect 12650 7814 12702 7866
rect 12702 7814 12704 7866
rect 12648 7812 12704 7814
rect 12440 6298 12496 6300
rect 12440 6246 12442 6298
rect 12442 6246 12494 6298
rect 12494 6246 12496 6298
rect 12440 6244 12496 6246
rect 12544 6298 12600 6300
rect 12544 6246 12546 6298
rect 12546 6246 12598 6298
rect 12598 6246 12600 6298
rect 12544 6244 12600 6246
rect 12648 6298 12704 6300
rect 12648 6246 12650 6298
rect 12650 6246 12702 6298
rect 12702 6246 12704 6298
rect 12648 6244 12704 6246
rect 12684 5906 12740 5908
rect 12684 5854 12686 5906
rect 12686 5854 12738 5906
rect 12738 5854 12740 5906
rect 12684 5852 12740 5854
rect 12572 5628 12628 5684
rect 13020 5852 13076 5908
rect 12796 4844 12852 4900
rect 12440 4730 12496 4732
rect 12440 4678 12442 4730
rect 12442 4678 12494 4730
rect 12494 4678 12496 4730
rect 12440 4676 12496 4678
rect 12544 4730 12600 4732
rect 12544 4678 12546 4730
rect 12546 4678 12598 4730
rect 12598 4678 12600 4730
rect 12544 4676 12600 4678
rect 12648 4730 12704 4732
rect 12648 4678 12650 4730
rect 12650 4678 12702 4730
rect 12702 4678 12704 4730
rect 12648 4676 12704 4678
rect 11900 3276 11956 3332
rect 12236 3612 12292 3668
rect 11004 2156 11060 2212
rect 11340 2604 11396 2660
rect 12012 2658 12068 2660
rect 12012 2606 12014 2658
rect 12014 2606 12066 2658
rect 12066 2606 12068 2658
rect 12012 2604 12068 2606
rect 11676 2268 11732 2324
rect 11788 1708 11844 1764
rect 12348 3500 12404 3556
rect 12440 3162 12496 3164
rect 12440 3110 12442 3162
rect 12442 3110 12494 3162
rect 12494 3110 12496 3162
rect 12440 3108 12496 3110
rect 12544 3162 12600 3164
rect 12544 3110 12546 3162
rect 12546 3110 12598 3162
rect 12598 3110 12600 3162
rect 12544 3108 12600 3110
rect 12648 3162 12704 3164
rect 12648 3110 12650 3162
rect 12650 3110 12702 3162
rect 12702 3110 12704 3162
rect 12648 3108 12704 3110
rect 12684 1708 12740 1764
rect 12440 1594 12496 1596
rect 12440 1542 12442 1594
rect 12442 1542 12494 1594
rect 12494 1542 12496 1594
rect 12440 1540 12496 1542
rect 12544 1594 12600 1596
rect 12544 1542 12546 1594
rect 12546 1542 12598 1594
rect 12598 1542 12600 1594
rect 12544 1540 12600 1542
rect 12648 1594 12704 1596
rect 12648 1542 12650 1594
rect 12650 1542 12702 1594
rect 12702 1542 12704 1594
rect 12648 1540 12704 1542
rect 12908 3666 12964 3668
rect 12908 3614 12910 3666
rect 12910 3614 12962 3666
rect 12962 3614 12964 3666
rect 12908 3612 12964 3614
rect 14364 10668 14420 10724
rect 13580 7756 13636 7812
rect 13244 5628 13300 5684
rect 13132 2492 13188 2548
rect 13132 2268 13188 2324
rect 13132 2044 13188 2100
rect 13804 6748 13860 6804
rect 13804 2940 13860 2996
rect 14140 6524 14196 6580
rect 14498 10218 14554 10220
rect 14498 10166 14500 10218
rect 14500 10166 14552 10218
rect 14552 10166 14554 10218
rect 14498 10164 14554 10166
rect 14602 10218 14658 10220
rect 14602 10166 14604 10218
rect 14604 10166 14656 10218
rect 14656 10166 14658 10218
rect 14602 10164 14658 10166
rect 14706 10218 14762 10220
rect 14706 10166 14708 10218
rect 14708 10166 14760 10218
rect 14760 10166 14762 10218
rect 14706 10164 14762 10166
rect 15148 9884 15204 9940
rect 14700 8930 14756 8932
rect 14700 8878 14702 8930
rect 14702 8878 14754 8930
rect 14754 8878 14756 8930
rect 14700 8876 14756 8878
rect 14498 8650 14554 8652
rect 14498 8598 14500 8650
rect 14500 8598 14552 8650
rect 14552 8598 14554 8650
rect 14498 8596 14554 8598
rect 14602 8650 14658 8652
rect 14602 8598 14604 8650
rect 14604 8598 14656 8650
rect 14656 8598 14658 8650
rect 14602 8596 14658 8598
rect 14706 8650 14762 8652
rect 14706 8598 14708 8650
rect 14708 8598 14760 8650
rect 14760 8598 14762 8650
rect 14706 8596 14762 8598
rect 14476 7756 14532 7812
rect 14498 7082 14554 7084
rect 14498 7030 14500 7082
rect 14500 7030 14552 7082
rect 14552 7030 14554 7082
rect 14498 7028 14554 7030
rect 14602 7082 14658 7084
rect 14602 7030 14604 7082
rect 14604 7030 14656 7082
rect 14656 7030 14658 7082
rect 14602 7028 14658 7030
rect 14706 7082 14762 7084
rect 14706 7030 14708 7082
rect 14708 7030 14760 7082
rect 14760 7030 14762 7082
rect 14706 7028 14762 7030
rect 14498 5514 14554 5516
rect 14498 5462 14500 5514
rect 14500 5462 14552 5514
rect 14552 5462 14554 5514
rect 14498 5460 14554 5462
rect 14602 5514 14658 5516
rect 14602 5462 14604 5514
rect 14604 5462 14656 5514
rect 14656 5462 14658 5514
rect 14602 5460 14658 5462
rect 14706 5514 14762 5516
rect 14706 5462 14708 5514
rect 14708 5462 14760 5514
rect 14760 5462 14762 5514
rect 14706 5460 14762 5462
rect 15596 9938 15652 9940
rect 15596 9886 15598 9938
rect 15598 9886 15650 9938
rect 15650 9886 15652 9938
rect 15596 9884 15652 9886
rect 15036 6636 15092 6692
rect 15372 8876 15428 8932
rect 15036 6412 15092 6468
rect 14924 5404 14980 5460
rect 14588 4844 14644 4900
rect 14588 4060 14644 4116
rect 14498 3946 14554 3948
rect 14498 3894 14500 3946
rect 14500 3894 14552 3946
rect 14552 3894 14554 3946
rect 14498 3892 14554 3894
rect 14602 3946 14658 3948
rect 14602 3894 14604 3946
rect 14604 3894 14656 3946
rect 14656 3894 14658 3946
rect 14602 3892 14658 3894
rect 14706 3946 14762 3948
rect 14706 3894 14708 3946
rect 14708 3894 14760 3946
rect 14760 3894 14762 3946
rect 14706 3892 14762 3894
rect 14588 3554 14644 3556
rect 14588 3502 14590 3554
rect 14590 3502 14642 3554
rect 14642 3502 14644 3554
rect 14588 3500 14644 3502
rect 14812 2994 14868 2996
rect 14812 2942 14814 2994
rect 14814 2942 14866 2994
rect 14866 2942 14868 2994
rect 14812 2940 14868 2942
rect 14498 2378 14554 2380
rect 14498 2326 14500 2378
rect 14500 2326 14552 2378
rect 14552 2326 14554 2378
rect 14498 2324 14554 2326
rect 14602 2378 14658 2380
rect 14602 2326 14604 2378
rect 14604 2326 14656 2378
rect 14656 2326 14658 2378
rect 14602 2324 14658 2326
rect 14706 2378 14762 2380
rect 14706 2326 14708 2378
rect 14708 2326 14760 2378
rect 14760 2326 14762 2378
rect 14706 2324 14762 2326
rect 15260 3276 15316 3332
rect 15484 7756 15540 7812
rect 15484 6524 15540 6580
rect 15596 6636 15652 6692
rect 16556 11002 16612 11004
rect 16556 10950 16558 11002
rect 16558 10950 16610 11002
rect 16610 10950 16612 11002
rect 16556 10948 16612 10950
rect 16660 11002 16716 11004
rect 16660 10950 16662 11002
rect 16662 10950 16714 11002
rect 16714 10950 16716 11002
rect 16660 10948 16716 10950
rect 16764 11002 16820 11004
rect 16764 10950 16766 11002
rect 16766 10950 16818 11002
rect 16818 10950 16820 11002
rect 16764 10948 16820 10950
rect 16556 9434 16612 9436
rect 16556 9382 16558 9434
rect 16558 9382 16610 9434
rect 16610 9382 16612 9434
rect 16556 9380 16612 9382
rect 16660 9434 16716 9436
rect 16660 9382 16662 9434
rect 16662 9382 16714 9434
rect 16714 9382 16716 9434
rect 16660 9380 16716 9382
rect 16764 9434 16820 9436
rect 16764 9382 16766 9434
rect 16766 9382 16818 9434
rect 16818 9382 16820 9434
rect 16764 9380 16820 9382
rect 16556 7866 16612 7868
rect 16556 7814 16558 7866
rect 16558 7814 16610 7866
rect 16610 7814 16612 7866
rect 16556 7812 16612 7814
rect 16660 7866 16716 7868
rect 16660 7814 16662 7866
rect 16662 7814 16714 7866
rect 16714 7814 16716 7866
rect 16660 7812 16716 7814
rect 16764 7866 16820 7868
rect 16764 7814 16766 7866
rect 16766 7814 16818 7866
rect 16818 7814 16820 7866
rect 16764 7812 16820 7814
rect 16556 6298 16612 6300
rect 16556 6246 16558 6298
rect 16558 6246 16610 6298
rect 16610 6246 16612 6298
rect 16556 6244 16612 6246
rect 16660 6298 16716 6300
rect 16660 6246 16662 6298
rect 16662 6246 16714 6298
rect 16714 6246 16716 6298
rect 16660 6244 16716 6246
rect 16764 6298 16820 6300
rect 16764 6246 16766 6298
rect 16766 6246 16818 6298
rect 16818 6246 16820 6298
rect 16764 6244 16820 6246
rect 15820 5852 15876 5908
rect 15932 5740 15988 5796
rect 15596 3554 15652 3556
rect 15596 3502 15598 3554
rect 15598 3502 15650 3554
rect 15650 3502 15652 3554
rect 15596 3500 15652 3502
rect 16268 5404 16324 5460
rect 16044 4060 16100 4116
rect 15484 2492 15540 2548
rect 16556 4730 16612 4732
rect 16556 4678 16558 4730
rect 16558 4678 16610 4730
rect 16610 4678 16612 4730
rect 16556 4676 16612 4678
rect 16660 4730 16716 4732
rect 16660 4678 16662 4730
rect 16662 4678 16714 4730
rect 16714 4678 16716 4730
rect 16660 4676 16716 4678
rect 16764 4730 16820 4732
rect 16764 4678 16766 4730
rect 16766 4678 16818 4730
rect 16818 4678 16820 4730
rect 16764 4676 16820 4678
rect 16556 3162 16612 3164
rect 16556 3110 16558 3162
rect 16558 3110 16610 3162
rect 16610 3110 16612 3162
rect 16556 3108 16612 3110
rect 16660 3162 16716 3164
rect 16660 3110 16662 3162
rect 16662 3110 16714 3162
rect 16714 3110 16716 3162
rect 16660 3108 16716 3110
rect 16764 3162 16820 3164
rect 16764 3110 16766 3162
rect 16766 3110 16818 3162
rect 16818 3110 16820 3162
rect 16764 3108 16820 3110
rect 16556 1594 16612 1596
rect 16556 1542 16558 1594
rect 16558 1542 16610 1594
rect 16610 1542 16612 1594
rect 16556 1540 16612 1542
rect 16660 1594 16716 1596
rect 16660 1542 16662 1594
rect 16662 1542 16714 1594
rect 16714 1542 16716 1594
rect 16660 1540 16716 1542
rect 16764 1594 16820 1596
rect 16764 1542 16766 1594
rect 16766 1542 16818 1594
rect 16818 1542 16820 1594
rect 16764 1540 16820 1542
<< metal3 >>
rect 4198 10948 4208 11004
rect 4264 10948 4312 11004
rect 4368 10948 4416 11004
rect 4472 10948 4482 11004
rect 8314 10948 8324 11004
rect 8380 10948 8428 11004
rect 8484 10948 8532 11004
rect 8588 10948 8598 11004
rect 12430 10948 12440 11004
rect 12496 10948 12544 11004
rect 12600 10948 12648 11004
rect 12704 10948 12714 11004
rect 16546 10948 16556 11004
rect 16612 10948 16660 11004
rect 16716 10948 16764 11004
rect 16820 10948 16830 11004
rect 0 10724 800 10752
rect 16200 10724 17000 10752
rect 0 10668 12348 10724
rect 12404 10668 12414 10724
rect 14354 10668 14364 10724
rect 14420 10668 17000 10724
rect 0 10640 800 10668
rect 16200 10640 17000 10668
rect 1362 10556 1372 10612
rect 1428 10556 2716 10612
rect 2772 10556 3780 10612
rect 4722 10556 4732 10612
rect 4788 10556 5740 10612
rect 5796 10556 6748 10612
rect 6804 10556 6814 10612
rect 3724 10500 3780 10556
rect 3714 10444 3724 10500
rect 3780 10444 3790 10500
rect 2140 10164 2150 10220
rect 2206 10164 2254 10220
rect 2310 10164 2358 10220
rect 2414 10164 2424 10220
rect 6256 10164 6266 10220
rect 6322 10164 6370 10220
rect 6426 10164 6474 10220
rect 6530 10164 6540 10220
rect 10372 10164 10382 10220
rect 10438 10164 10486 10220
rect 10542 10164 10590 10220
rect 10646 10164 10656 10220
rect 14488 10164 14498 10220
rect 14554 10164 14602 10220
rect 14658 10164 14706 10220
rect 14762 10164 14772 10220
rect 7074 9996 7084 10052
rect 7140 9996 7756 10052
rect 7812 9996 7822 10052
rect 9538 9884 9548 9940
rect 9604 9884 10780 9940
rect 10836 9884 11788 9940
rect 11844 9884 11854 9940
rect 15138 9884 15148 9940
rect 15204 9884 15596 9940
rect 15652 9884 15662 9940
rect 2482 9660 2492 9716
rect 2548 9660 3388 9716
rect 3444 9660 4508 9716
rect 4564 9660 4574 9716
rect 4198 9380 4208 9436
rect 4264 9380 4312 9436
rect 4368 9380 4416 9436
rect 4472 9380 4482 9436
rect 8314 9380 8324 9436
rect 8380 9380 8428 9436
rect 8484 9380 8532 9436
rect 8588 9380 8598 9436
rect 12430 9380 12440 9436
rect 12496 9380 12544 9436
rect 12600 9380 12648 9436
rect 12704 9380 12714 9436
rect 16546 9380 16556 9436
rect 16612 9380 16660 9436
rect 16716 9380 16764 9436
rect 16820 9380 16830 9436
rect 6514 9212 6524 9268
rect 6580 9212 7308 9268
rect 7364 9212 7374 9268
rect 9986 8988 9996 9044
rect 10052 8988 11004 9044
rect 11060 8988 12012 9044
rect 12068 8988 12078 9044
rect 2930 8876 2940 8932
rect 2996 8876 3948 8932
rect 4004 8876 4014 8932
rect 14690 8876 14700 8932
rect 14756 8876 15372 8932
rect 15428 8876 15438 8932
rect 2140 8596 2150 8652
rect 2206 8596 2254 8652
rect 2310 8596 2358 8652
rect 2414 8596 2424 8652
rect 6256 8596 6266 8652
rect 6322 8596 6370 8652
rect 6426 8596 6474 8652
rect 6530 8596 6540 8652
rect 10372 8596 10382 8652
rect 10438 8596 10486 8652
rect 10542 8596 10590 8652
rect 10646 8596 10656 8652
rect 14488 8596 14498 8652
rect 14554 8596 14602 8652
rect 14658 8596 14706 8652
rect 14762 8596 14772 8652
rect 1922 8428 1932 8484
rect 1988 8428 2940 8484
rect 2996 8428 3006 8484
rect 578 8204 588 8260
rect 644 8204 2716 8260
rect 2772 8204 3724 8260
rect 3780 8204 3790 8260
rect 8642 8204 8652 8260
rect 8708 8204 9660 8260
rect 9716 8204 10668 8260
rect 10724 8204 10734 8260
rect 4198 7812 4208 7868
rect 4264 7812 4312 7868
rect 4368 7812 4416 7868
rect 4472 7812 4482 7868
rect 8314 7812 8324 7868
rect 8380 7812 8428 7868
rect 8484 7812 8532 7868
rect 8588 7812 8598 7868
rect 12430 7812 12440 7868
rect 12496 7812 12544 7868
rect 12600 7812 12648 7868
rect 12704 7812 12714 7868
rect 16546 7812 16556 7868
rect 16612 7812 16660 7868
rect 16716 7812 16764 7868
rect 16820 7812 16830 7868
rect 13570 7756 13580 7812
rect 13636 7756 14476 7812
rect 14532 7756 15484 7812
rect 15540 7756 15550 7812
rect 2706 7308 2716 7364
rect 2772 7308 3724 7364
rect 3780 7308 3790 7364
rect 7746 7308 7756 7364
rect 7812 7308 8540 7364
rect 8596 7308 8606 7364
rect 2140 7028 2150 7084
rect 2206 7028 2254 7084
rect 2310 7028 2358 7084
rect 2414 7028 2424 7084
rect 6256 7028 6266 7084
rect 6322 7028 6370 7084
rect 6426 7028 6474 7084
rect 6530 7028 6540 7084
rect 10372 7028 10382 7084
rect 10438 7028 10486 7084
rect 10542 7028 10590 7084
rect 10646 7028 10656 7084
rect 14488 7028 14498 7084
rect 14554 7028 14602 7084
rect 14658 7028 14706 7084
rect 14762 7028 14772 7084
rect 1026 6860 1036 6916
rect 1092 6860 2716 6916
rect 2772 6860 2782 6916
rect 11330 6748 11340 6804
rect 11396 6748 13804 6804
rect 13860 6748 13870 6804
rect 15026 6636 15036 6692
rect 15092 6636 15596 6692
rect 15652 6636 15662 6692
rect 14130 6524 14140 6580
rect 14196 6524 15484 6580
rect 15540 6524 15550 6580
rect 0 6468 800 6496
rect 16200 6468 17000 6496
rect 0 6412 980 6468
rect 9202 6412 9212 6468
rect 9268 6412 10220 6468
rect 10276 6412 10286 6468
rect 15026 6412 15036 6468
rect 15092 6412 17000 6468
rect 0 6384 800 6412
rect 924 6132 980 6412
rect 16200 6384 17000 6412
rect 4198 6244 4208 6300
rect 4264 6244 4312 6300
rect 4368 6244 4416 6300
rect 4472 6244 4482 6300
rect 8314 6244 8324 6300
rect 8380 6244 8428 6300
rect 8484 6244 8532 6300
rect 8588 6244 8598 6300
rect 12430 6244 12440 6300
rect 12496 6244 12544 6300
rect 12600 6244 12648 6300
rect 12704 6244 12714 6300
rect 16546 6244 16556 6300
rect 16612 6244 16660 6300
rect 16716 6244 16764 6300
rect 16820 6244 16830 6300
rect 700 6076 980 6132
rect 700 5684 756 6076
rect 8194 5964 8204 6020
rect 8260 5964 9212 6020
rect 9268 5964 9278 6020
rect 3714 5852 3724 5908
rect 3780 5852 4732 5908
rect 4788 5852 5740 5908
rect 5796 5852 5806 5908
rect 12674 5852 12684 5908
rect 12740 5852 13020 5908
rect 13076 5852 15820 5908
rect 15876 5852 15886 5908
rect 11554 5740 11564 5796
rect 11620 5740 15932 5796
rect 15988 5740 15998 5796
rect 700 5628 12572 5684
rect 12628 5628 13244 5684
rect 13300 5628 13310 5684
rect 2594 5516 2604 5572
rect 2660 5516 4620 5572
rect 4676 5516 4686 5572
rect 2140 5460 2150 5516
rect 2206 5460 2254 5516
rect 2310 5460 2358 5516
rect 2414 5460 2424 5516
rect 6256 5460 6266 5516
rect 6322 5460 6370 5516
rect 6426 5460 6474 5516
rect 6530 5460 6540 5516
rect 10372 5460 10382 5516
rect 10438 5460 10486 5516
rect 10542 5460 10590 5516
rect 10646 5460 10656 5516
rect 14488 5460 14498 5516
rect 14554 5460 14602 5516
rect 14658 5460 14706 5516
rect 14762 5460 14772 5516
rect 14914 5404 14924 5460
rect 14980 5404 16268 5460
rect 16324 5404 16334 5460
rect 10098 5180 10108 5236
rect 10164 5180 11788 5236
rect 11844 5180 11854 5236
rect 3154 5068 3164 5124
rect 3220 5068 4060 5124
rect 4116 5068 4126 5124
rect 3938 4844 3948 4900
rect 4004 4844 4508 4900
rect 4564 4844 4574 4900
rect 12786 4844 12796 4900
rect 12852 4844 14588 4900
rect 14644 4844 14654 4900
rect 3378 4732 3388 4788
rect 3444 4732 3836 4788
rect 3892 4732 3902 4788
rect 4198 4676 4208 4732
rect 4264 4676 4312 4732
rect 4368 4676 4416 4732
rect 4472 4676 4482 4732
rect 8314 4676 8324 4732
rect 8380 4676 8428 4732
rect 8484 4676 8532 4732
rect 8588 4676 8598 4732
rect 12430 4676 12440 4732
rect 12496 4676 12544 4732
rect 12600 4676 12648 4732
rect 12704 4676 12714 4732
rect 16546 4676 16556 4732
rect 16612 4676 16660 4732
rect 16716 4676 16764 4732
rect 16820 4676 16830 4732
rect 6962 4172 6972 4228
rect 7028 4172 8540 4228
rect 8596 4172 8606 4228
rect 14578 4060 14588 4116
rect 14644 4060 16044 4116
rect 16100 4060 16110 4116
rect 2140 3892 2150 3948
rect 2206 3892 2254 3948
rect 2310 3892 2358 3948
rect 2414 3892 2424 3948
rect 6256 3892 6266 3948
rect 6322 3892 6370 3948
rect 6426 3892 6474 3948
rect 6530 3892 6540 3948
rect 10372 3892 10382 3948
rect 10438 3892 10486 3948
rect 10542 3892 10590 3948
rect 10646 3892 10656 3948
rect 14488 3892 14498 3948
rect 14554 3892 14602 3948
rect 14658 3892 14706 3948
rect 14762 3892 14772 3948
rect 5954 3724 5964 3780
rect 6020 3724 6972 3780
rect 7028 3724 7038 3780
rect 12226 3612 12236 3668
rect 12292 3612 12908 3668
rect 12964 3612 12974 3668
rect 12338 3500 12348 3556
rect 12404 3500 14588 3556
rect 14644 3500 15596 3556
rect 15652 3500 15662 3556
rect 2818 3388 2828 3444
rect 2884 3388 3948 3444
rect 4004 3388 4014 3444
rect 5506 3388 5516 3444
rect 5572 3388 6748 3444
rect 6804 3388 7644 3444
rect 7700 3388 7710 3444
rect 11890 3276 11900 3332
rect 11956 3276 15260 3332
rect 15316 3276 15326 3332
rect 4198 3108 4208 3164
rect 4264 3108 4312 3164
rect 4368 3108 4416 3164
rect 4472 3108 4482 3164
rect 8314 3108 8324 3164
rect 8380 3108 8428 3164
rect 8484 3108 8532 3164
rect 8588 3108 8598 3164
rect 12430 3108 12440 3164
rect 12496 3108 12544 3164
rect 12600 3108 12648 3164
rect 12704 3108 12714 3164
rect 16546 3108 16556 3164
rect 16612 3108 16660 3164
rect 16716 3108 16764 3164
rect 16820 3108 16830 3164
rect 13794 2940 13804 2996
rect 13860 2940 14812 2996
rect 14868 2940 14878 2996
rect 11330 2604 11340 2660
rect 11396 2604 12012 2660
rect 12068 2604 12078 2660
rect 13122 2492 13132 2548
rect 13188 2492 15484 2548
rect 15540 2492 15550 2548
rect 2140 2324 2150 2380
rect 2206 2324 2254 2380
rect 2310 2324 2358 2380
rect 2414 2324 2424 2380
rect 6256 2324 6266 2380
rect 6322 2324 6370 2380
rect 6426 2324 6474 2380
rect 6530 2324 6540 2380
rect 10372 2324 10382 2380
rect 10438 2324 10486 2380
rect 10542 2324 10590 2380
rect 10646 2324 10656 2380
rect 14488 2324 14498 2380
rect 14554 2324 14602 2380
rect 14658 2324 14706 2380
rect 14762 2324 14772 2380
rect 11666 2268 11676 2324
rect 11732 2268 13132 2324
rect 13188 2268 13198 2324
rect 0 2212 800 2240
rect 16200 2212 17000 2240
rect 0 2156 8652 2212
rect 8708 2156 8718 2212
rect 10994 2156 11004 2212
rect 11060 2156 17000 2212
rect 0 2128 800 2156
rect 16200 2128 17000 2156
rect 6402 2044 6412 2100
rect 6468 2044 7420 2100
rect 7476 2044 8428 2100
rect 8484 2044 8494 2100
rect 10546 2044 10556 2100
rect 10612 2044 13132 2100
rect 13188 2044 13198 2100
rect 802 1932 812 1988
rect 868 1932 1596 1988
rect 1652 1932 4060 1988
rect 4116 1932 4126 1988
rect 5058 1820 5068 1876
rect 5124 1820 6748 1876
rect 6804 1820 7644 1876
rect 7700 1820 7710 1876
rect 11778 1708 11788 1764
rect 11844 1708 12684 1764
rect 12740 1708 12750 1764
rect 4198 1540 4208 1596
rect 4264 1540 4312 1596
rect 4368 1540 4416 1596
rect 4472 1540 4482 1596
rect 8314 1540 8324 1596
rect 8380 1540 8428 1596
rect 8484 1540 8532 1596
rect 8588 1540 8598 1596
rect 12430 1540 12440 1596
rect 12496 1540 12544 1596
rect 12600 1540 12648 1596
rect 12704 1540 12714 1596
rect 16546 1540 16556 1596
rect 16612 1540 16660 1596
rect 16716 1540 16764 1596
rect 16820 1540 16830 1596
<< via3 >>
rect 4208 10948 4264 11004
rect 4312 10948 4368 11004
rect 4416 10948 4472 11004
rect 8324 10948 8380 11004
rect 8428 10948 8484 11004
rect 8532 10948 8588 11004
rect 12440 10948 12496 11004
rect 12544 10948 12600 11004
rect 12648 10948 12704 11004
rect 16556 10948 16612 11004
rect 16660 10948 16716 11004
rect 16764 10948 16820 11004
rect 2150 10164 2206 10220
rect 2254 10164 2310 10220
rect 2358 10164 2414 10220
rect 6266 10164 6322 10220
rect 6370 10164 6426 10220
rect 6474 10164 6530 10220
rect 10382 10164 10438 10220
rect 10486 10164 10542 10220
rect 10590 10164 10646 10220
rect 14498 10164 14554 10220
rect 14602 10164 14658 10220
rect 14706 10164 14762 10220
rect 4208 9380 4264 9436
rect 4312 9380 4368 9436
rect 4416 9380 4472 9436
rect 8324 9380 8380 9436
rect 8428 9380 8484 9436
rect 8532 9380 8588 9436
rect 12440 9380 12496 9436
rect 12544 9380 12600 9436
rect 12648 9380 12704 9436
rect 16556 9380 16612 9436
rect 16660 9380 16716 9436
rect 16764 9380 16820 9436
rect 2150 8596 2206 8652
rect 2254 8596 2310 8652
rect 2358 8596 2414 8652
rect 6266 8596 6322 8652
rect 6370 8596 6426 8652
rect 6474 8596 6530 8652
rect 10382 8596 10438 8652
rect 10486 8596 10542 8652
rect 10590 8596 10646 8652
rect 14498 8596 14554 8652
rect 14602 8596 14658 8652
rect 14706 8596 14762 8652
rect 4208 7812 4264 7868
rect 4312 7812 4368 7868
rect 4416 7812 4472 7868
rect 8324 7812 8380 7868
rect 8428 7812 8484 7868
rect 8532 7812 8588 7868
rect 12440 7812 12496 7868
rect 12544 7812 12600 7868
rect 12648 7812 12704 7868
rect 16556 7812 16612 7868
rect 16660 7812 16716 7868
rect 16764 7812 16820 7868
rect 2150 7028 2206 7084
rect 2254 7028 2310 7084
rect 2358 7028 2414 7084
rect 6266 7028 6322 7084
rect 6370 7028 6426 7084
rect 6474 7028 6530 7084
rect 10382 7028 10438 7084
rect 10486 7028 10542 7084
rect 10590 7028 10646 7084
rect 14498 7028 14554 7084
rect 14602 7028 14658 7084
rect 14706 7028 14762 7084
rect 4208 6244 4264 6300
rect 4312 6244 4368 6300
rect 4416 6244 4472 6300
rect 8324 6244 8380 6300
rect 8428 6244 8484 6300
rect 8532 6244 8588 6300
rect 12440 6244 12496 6300
rect 12544 6244 12600 6300
rect 12648 6244 12704 6300
rect 16556 6244 16612 6300
rect 16660 6244 16716 6300
rect 16764 6244 16820 6300
rect 2150 5460 2206 5516
rect 2254 5460 2310 5516
rect 2358 5460 2414 5516
rect 6266 5460 6322 5516
rect 6370 5460 6426 5516
rect 6474 5460 6530 5516
rect 10382 5460 10438 5516
rect 10486 5460 10542 5516
rect 10590 5460 10646 5516
rect 14498 5460 14554 5516
rect 14602 5460 14658 5516
rect 14706 5460 14762 5516
rect 4208 4676 4264 4732
rect 4312 4676 4368 4732
rect 4416 4676 4472 4732
rect 8324 4676 8380 4732
rect 8428 4676 8484 4732
rect 8532 4676 8588 4732
rect 12440 4676 12496 4732
rect 12544 4676 12600 4732
rect 12648 4676 12704 4732
rect 16556 4676 16612 4732
rect 16660 4676 16716 4732
rect 16764 4676 16820 4732
rect 2150 3892 2206 3948
rect 2254 3892 2310 3948
rect 2358 3892 2414 3948
rect 6266 3892 6322 3948
rect 6370 3892 6426 3948
rect 6474 3892 6530 3948
rect 10382 3892 10438 3948
rect 10486 3892 10542 3948
rect 10590 3892 10646 3948
rect 14498 3892 14554 3948
rect 14602 3892 14658 3948
rect 14706 3892 14762 3948
rect 4208 3108 4264 3164
rect 4312 3108 4368 3164
rect 4416 3108 4472 3164
rect 8324 3108 8380 3164
rect 8428 3108 8484 3164
rect 8532 3108 8588 3164
rect 12440 3108 12496 3164
rect 12544 3108 12600 3164
rect 12648 3108 12704 3164
rect 16556 3108 16612 3164
rect 16660 3108 16716 3164
rect 16764 3108 16820 3164
rect 2150 2324 2206 2380
rect 2254 2324 2310 2380
rect 2358 2324 2414 2380
rect 6266 2324 6322 2380
rect 6370 2324 6426 2380
rect 6474 2324 6530 2380
rect 10382 2324 10438 2380
rect 10486 2324 10542 2380
rect 10590 2324 10646 2380
rect 14498 2324 14554 2380
rect 14602 2324 14658 2380
rect 14706 2324 14762 2380
rect 4208 1540 4264 1596
rect 4312 1540 4368 1596
rect 4416 1540 4472 1596
rect 8324 1540 8380 1596
rect 8428 1540 8484 1596
rect 8532 1540 8588 1596
rect 12440 1540 12496 1596
rect 12544 1540 12600 1596
rect 12648 1540 12704 1596
rect 16556 1540 16612 1596
rect 16660 1540 16716 1596
rect 16764 1540 16820 1596
<< metal4 >>
rect 2122 10220 2442 11036
rect 2122 10164 2150 10220
rect 2206 10164 2254 10220
rect 2310 10164 2358 10220
rect 2414 10164 2442 10220
rect 2122 8652 2442 10164
rect 2122 8596 2150 8652
rect 2206 8596 2254 8652
rect 2310 8596 2358 8652
rect 2414 8596 2442 8652
rect 2122 7084 2442 8596
rect 2122 7028 2150 7084
rect 2206 7028 2254 7084
rect 2310 7028 2358 7084
rect 2414 7028 2442 7084
rect 2122 5516 2442 7028
rect 2122 5460 2150 5516
rect 2206 5460 2254 5516
rect 2310 5460 2358 5516
rect 2414 5460 2442 5516
rect 2122 3948 2442 5460
rect 2122 3892 2150 3948
rect 2206 3892 2254 3948
rect 2310 3892 2358 3948
rect 2414 3892 2442 3948
rect 2122 2380 2442 3892
rect 2122 2324 2150 2380
rect 2206 2324 2254 2380
rect 2310 2324 2358 2380
rect 2414 2324 2442 2380
rect 2122 1508 2442 2324
rect 4180 11004 4500 11036
rect 4180 10948 4208 11004
rect 4264 10948 4312 11004
rect 4368 10948 4416 11004
rect 4472 10948 4500 11004
rect 4180 9436 4500 10948
rect 4180 9380 4208 9436
rect 4264 9380 4312 9436
rect 4368 9380 4416 9436
rect 4472 9380 4500 9436
rect 4180 7868 4500 9380
rect 4180 7812 4208 7868
rect 4264 7812 4312 7868
rect 4368 7812 4416 7868
rect 4472 7812 4500 7868
rect 4180 6300 4500 7812
rect 4180 6244 4208 6300
rect 4264 6244 4312 6300
rect 4368 6244 4416 6300
rect 4472 6244 4500 6300
rect 4180 4732 4500 6244
rect 4180 4676 4208 4732
rect 4264 4676 4312 4732
rect 4368 4676 4416 4732
rect 4472 4676 4500 4732
rect 4180 3164 4500 4676
rect 4180 3108 4208 3164
rect 4264 3108 4312 3164
rect 4368 3108 4416 3164
rect 4472 3108 4500 3164
rect 4180 1596 4500 3108
rect 4180 1540 4208 1596
rect 4264 1540 4312 1596
rect 4368 1540 4416 1596
rect 4472 1540 4500 1596
rect 4180 1508 4500 1540
rect 6238 10220 6558 11036
rect 6238 10164 6266 10220
rect 6322 10164 6370 10220
rect 6426 10164 6474 10220
rect 6530 10164 6558 10220
rect 6238 8652 6558 10164
rect 6238 8596 6266 8652
rect 6322 8596 6370 8652
rect 6426 8596 6474 8652
rect 6530 8596 6558 8652
rect 6238 7084 6558 8596
rect 6238 7028 6266 7084
rect 6322 7028 6370 7084
rect 6426 7028 6474 7084
rect 6530 7028 6558 7084
rect 6238 5516 6558 7028
rect 6238 5460 6266 5516
rect 6322 5460 6370 5516
rect 6426 5460 6474 5516
rect 6530 5460 6558 5516
rect 6238 3948 6558 5460
rect 6238 3892 6266 3948
rect 6322 3892 6370 3948
rect 6426 3892 6474 3948
rect 6530 3892 6558 3948
rect 6238 2380 6558 3892
rect 6238 2324 6266 2380
rect 6322 2324 6370 2380
rect 6426 2324 6474 2380
rect 6530 2324 6558 2380
rect 6238 1508 6558 2324
rect 8296 11004 8616 11036
rect 8296 10948 8324 11004
rect 8380 10948 8428 11004
rect 8484 10948 8532 11004
rect 8588 10948 8616 11004
rect 8296 9436 8616 10948
rect 8296 9380 8324 9436
rect 8380 9380 8428 9436
rect 8484 9380 8532 9436
rect 8588 9380 8616 9436
rect 8296 7868 8616 9380
rect 8296 7812 8324 7868
rect 8380 7812 8428 7868
rect 8484 7812 8532 7868
rect 8588 7812 8616 7868
rect 8296 6300 8616 7812
rect 8296 6244 8324 6300
rect 8380 6244 8428 6300
rect 8484 6244 8532 6300
rect 8588 6244 8616 6300
rect 8296 4732 8616 6244
rect 8296 4676 8324 4732
rect 8380 4676 8428 4732
rect 8484 4676 8532 4732
rect 8588 4676 8616 4732
rect 8296 3164 8616 4676
rect 8296 3108 8324 3164
rect 8380 3108 8428 3164
rect 8484 3108 8532 3164
rect 8588 3108 8616 3164
rect 8296 1596 8616 3108
rect 8296 1540 8324 1596
rect 8380 1540 8428 1596
rect 8484 1540 8532 1596
rect 8588 1540 8616 1596
rect 8296 1508 8616 1540
rect 10354 10220 10674 11036
rect 10354 10164 10382 10220
rect 10438 10164 10486 10220
rect 10542 10164 10590 10220
rect 10646 10164 10674 10220
rect 10354 8652 10674 10164
rect 10354 8596 10382 8652
rect 10438 8596 10486 8652
rect 10542 8596 10590 8652
rect 10646 8596 10674 8652
rect 10354 7084 10674 8596
rect 10354 7028 10382 7084
rect 10438 7028 10486 7084
rect 10542 7028 10590 7084
rect 10646 7028 10674 7084
rect 10354 5516 10674 7028
rect 10354 5460 10382 5516
rect 10438 5460 10486 5516
rect 10542 5460 10590 5516
rect 10646 5460 10674 5516
rect 10354 3948 10674 5460
rect 10354 3892 10382 3948
rect 10438 3892 10486 3948
rect 10542 3892 10590 3948
rect 10646 3892 10674 3948
rect 10354 2380 10674 3892
rect 10354 2324 10382 2380
rect 10438 2324 10486 2380
rect 10542 2324 10590 2380
rect 10646 2324 10674 2380
rect 10354 1508 10674 2324
rect 12412 11004 12732 11036
rect 12412 10948 12440 11004
rect 12496 10948 12544 11004
rect 12600 10948 12648 11004
rect 12704 10948 12732 11004
rect 12412 9436 12732 10948
rect 12412 9380 12440 9436
rect 12496 9380 12544 9436
rect 12600 9380 12648 9436
rect 12704 9380 12732 9436
rect 12412 7868 12732 9380
rect 12412 7812 12440 7868
rect 12496 7812 12544 7868
rect 12600 7812 12648 7868
rect 12704 7812 12732 7868
rect 12412 6300 12732 7812
rect 12412 6244 12440 6300
rect 12496 6244 12544 6300
rect 12600 6244 12648 6300
rect 12704 6244 12732 6300
rect 12412 4732 12732 6244
rect 12412 4676 12440 4732
rect 12496 4676 12544 4732
rect 12600 4676 12648 4732
rect 12704 4676 12732 4732
rect 12412 3164 12732 4676
rect 12412 3108 12440 3164
rect 12496 3108 12544 3164
rect 12600 3108 12648 3164
rect 12704 3108 12732 3164
rect 12412 1596 12732 3108
rect 12412 1540 12440 1596
rect 12496 1540 12544 1596
rect 12600 1540 12648 1596
rect 12704 1540 12732 1596
rect 12412 1508 12732 1540
rect 14470 10220 14790 11036
rect 14470 10164 14498 10220
rect 14554 10164 14602 10220
rect 14658 10164 14706 10220
rect 14762 10164 14790 10220
rect 14470 8652 14790 10164
rect 14470 8596 14498 8652
rect 14554 8596 14602 8652
rect 14658 8596 14706 8652
rect 14762 8596 14790 8652
rect 14470 7084 14790 8596
rect 14470 7028 14498 7084
rect 14554 7028 14602 7084
rect 14658 7028 14706 7084
rect 14762 7028 14790 7084
rect 14470 5516 14790 7028
rect 14470 5460 14498 5516
rect 14554 5460 14602 5516
rect 14658 5460 14706 5516
rect 14762 5460 14790 5516
rect 14470 3948 14790 5460
rect 14470 3892 14498 3948
rect 14554 3892 14602 3948
rect 14658 3892 14706 3948
rect 14762 3892 14790 3948
rect 14470 2380 14790 3892
rect 14470 2324 14498 2380
rect 14554 2324 14602 2380
rect 14658 2324 14706 2380
rect 14762 2324 14790 2380
rect 14470 1508 14790 2324
rect 16528 11004 16848 11036
rect 16528 10948 16556 11004
rect 16612 10948 16660 11004
rect 16716 10948 16764 11004
rect 16820 10948 16848 11004
rect 16528 9436 16848 10948
rect 16528 9380 16556 9436
rect 16612 9380 16660 9436
rect 16716 9380 16764 9436
rect 16820 9380 16848 9436
rect 16528 7868 16848 9380
rect 16528 7812 16556 7868
rect 16612 7812 16660 7868
rect 16716 7812 16764 7868
rect 16820 7812 16848 7868
rect 16528 6300 16848 7812
rect 16528 6244 16556 6300
rect 16612 6244 16660 6300
rect 16716 6244 16764 6300
rect 16820 6244 16848 6300
rect 16528 4732 16848 6244
rect 16528 4676 16556 4732
rect 16612 4676 16660 4732
rect 16716 4676 16764 4732
rect 16820 4676 16848 4732
rect 16528 3164 16848 4676
rect 16528 3108 16556 3164
rect 16612 3108 16660 3164
rect 16716 3108 16764 3164
rect 16820 3108 16848 3164
rect 16528 1596 16848 3108
rect 16528 1540 16556 1596
rect 16612 1540 16660 1596
rect 16716 1540 16764 1596
rect 16820 1540 16848 1596
rect 16528 1508 16848 1540
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[0\]_I $PDK_ROOT/$PDK/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670092720
transform 1 0 10640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[1\]_I
timestamp 1670092720
transform 1 0 11536 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[2\]_I
timestamp 1670092720
transform 1 0 11760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[3\]_I
timestamp 1670092720
transform 1 0 11984 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[4\]_I
timestamp 1670092720
transform 1 0 11760 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[5\]_I
timestamp 1670092720
transform 1 0 11312 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[6\]_I
timestamp 1670092720
transform 1 0 14784 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[7\]_I
timestamp 1670092720
transform 1 0 15232 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[8\]_I
timestamp 1670092720
transform 1 0 15568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[9\]_I
timestamp 1670092720
transform 1 0 16016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[10\]_I
timestamp 1670092720
transform 1 0 15456 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[11\]_I
timestamp 1670092720
transform 1 0 15456 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[12\]_I
timestamp 1670092720
transform 1 0 15680 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[13\]_I
timestamp 1670092720
transform 1 0 15568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[14\]_I
timestamp 1670092720
transform 1 0 15792 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[15\]_I
timestamp 1670092720
transform 1 0 16016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[16\]_I
timestamp 1670092720
transform -1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[17\]_I
timestamp 1670092720
transform -1 0 16352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[18\]_I
timestamp 1670092720
transform -1 0 8512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[19\]_I
timestamp 1670092720
transform -1 0 12656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[20\]_I
timestamp 1670092720
transform 1 0 12320 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[21\]_I
timestamp 1670092720
transform 1 0 3696 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[22\]_I
timestamp 1670092720
transform 1 0 3696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[23\]_I
timestamp 1670092720
transform 1 0 3696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[24\]_I
timestamp 1670092720
transform 1 0 3920 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[25\]_I
timestamp 1670092720
transform 1 0 4480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[26\]_I
timestamp 1670092720
transform 1 0 4480 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[27\]_I
timestamp 1670092720
transform 1 0 3808 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[28\]_I
timestamp 1670092720
transform 1 0 5712 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[29\]_I
timestamp 1670092720
transform -1 0 896 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[30\]_I
timestamp 1670092720
transform 1 0 4928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[31\]_I
timestamp 1670092720
transform 1 0 7616 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[32\]_I
timestamp 1670092720
transform 1 0 7616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[33\]_I
timestamp 1670092720
transform 1 0 8512 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[34\]_I
timestamp 1670092720
transform 1 0 8400 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[35\]_I
timestamp 1670092720
transform -1 0 4816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[36\]_I
timestamp 1670092720
transform 1 0 7056 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[37\]_I
timestamp 1670092720
transform 1 0 8512 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_BUF\[38\]_I
timestamp 1670092720
transform 1 0 10192 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[0\] $PDK_ROOT/$PDK/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670092720
transform -1 0 10416 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[1\]
timestamp 1670092720
transform -1 0 11312 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[2\]
timestamp 1670092720
transform -1 0 11536 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[3\]
timestamp 1670092720
transform -1 0 11760 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[4\]
timestamp 1670092720
transform -1 0 12208 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[5\]
timestamp 1670092720
transform -1 0 11984 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[6\]
timestamp 1670092720
transform -1 0 14560 0 -1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[7\]
timestamp 1670092720
transform -1 0 15232 0 1 1568
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[8\]
timestamp 1670092720
transform -1 0 15344 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[9\]
timestamp 1670092720
transform -1 0 15344 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[10\]
timestamp 1670092720
transform -1 0 11872 0 1 1568
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[11\]
timestamp 1670092720
transform -1 0 15232 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[12\]
timestamp 1670092720
transform -1 0 15680 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[13\]
timestamp 1670092720
transform -1 0 15792 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[14\]
timestamp 1670092720
transform -1 0 16352 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[15\]
timestamp 1670092720
transform -1 0 16016 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[16\]
timestamp 1670092720
transform -1 0 12880 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[17\]
timestamp 1670092720
transform -1 0 16352 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[18\]
timestamp 1670092720
transform 1 0 8512 0 -1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[19\]
timestamp 1670092720
transform 1 0 13104 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[20\]
timestamp 1670092720
transform 1 0 12432 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[21\]
timestamp 1670092720
transform -1 0 3472 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[22\]
timestamp 1670092720
transform -1 0 3472 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[23\]
timestamp 1670092720
transform -1 0 3472 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[24\]
timestamp 1670092720
transform -1 0 3696 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[25\]
timestamp 1670092720
transform -1 0 4032 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[26\]
timestamp 1670092720
transform -1 0 4256 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[27\]
timestamp 1670092720
transform -1 0 4032 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[28\]
timestamp 1670092720
transform -1 0 5488 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[29\]
timestamp 1670092720
transform 1 0 1120 0 1 1568
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[30\]
timestamp 1670092720
transform -1 0 4928 0 -1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[31\]
timestamp 1670092720
transform -1 0 7392 0 1 1568
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[32\]
timestamp 1670092720
transform -1 0 7392 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[33\]
timestamp 1670092720
transform -1 0 7728 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[34\]
timestamp 1670092720
transform -1 0 8064 0 -1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[35\]
timestamp 1670092720
transform 1 0 5040 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[36\]
timestamp 1670092720
transform -1 0 8064 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[37\]
timestamp 1670092720
transform -1 0 8400 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  BUF\[38\]
timestamp 1670092720
transform -1 0 9968 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2 $PDK_ROOT/$PDK/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670092720
transform 1 0 448 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6
timestamp 1670092720
transform 1 0 896 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 $PDK_ROOT/$PDK/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670092720
transform 1 0 4032 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1670092720
transform 1 0 4368 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64
timestamp 1670092720
transform 1 0 7392 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68
timestamp 1670092720
transform 1 0 7840 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72
timestamp 1670092720
transform 1 0 8288 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75
timestamp 1670092720
transform 1 0 8624 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77
timestamp 1670092720
transform 1 0 8848 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1670092720
transform 1 0 11872 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107
timestamp 1670092720
transform 1 0 12208 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_134
timestamp 1670092720
transform 1 0 15232 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_138
timestamp 1670092720
transform 1 0 15680 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_142
timestamp 1670092720
transform 1 0 16128 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_144
timestamp 1670092720
transform 1 0 16352 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_2 $PDK_ROOT/$PDK/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670092720
transform 1 0 448 0 -1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_10 $PDK_ROOT/$PDK/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670092720
transform 1 0 1344 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_14
timestamp 1670092720
transform 1 0 1792 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_42
timestamp 1670092720
transform 1 0 4928 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1670092720
transform 1 0 8064 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_73
timestamp 1670092720
transform 1 0 8400 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_100
timestamp 1670092720
transform 1 0 11424 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_128
timestamp 1670092720
transform 1 0 14560 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_132
timestamp 1670092720
transform 1 0 15008 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_136
timestamp 1670092720
transform 1 0 15456 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_138
timestamp 1670092720
transform 1 0 15680 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1670092720
transform 1 0 16016 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_144
timestamp 1670092720
transform 1 0 16352 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_2
timestamp 1670092720
transform 1 0 448 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_6
timestamp 1670092720
transform 1 0 896 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1670092720
transform 1 0 4032 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_37
timestamp 1670092720
transform 1 0 4368 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_64
timestamp 1670092720
transform 1 0 7392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_68
timestamp 1670092720
transform 1 0 7840 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_74
timestamp 1670092720
transform 1 0 8512 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_78
timestamp 1670092720
transform 1 0 8960 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1670092720
transform 1 0 11984 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_108
timestamp 1670092720
transform 1 0 12320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_135
timestamp 1670092720
transform 1 0 15344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_139
timestamp 1670092720
transform 1 0 15792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_143
timestamp 1670092720
transform 1 0 16240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_2
timestamp 1670092720
transform 1 0 448 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_36
timestamp 1670092720
transform 1 0 4256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_40
timestamp 1670092720
transform 1 0 4704 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_67
timestamp 1670092720
transform 1 0 7728 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_73
timestamp 1670092720
transform 1 0 8400 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_76
timestamp 1670092720
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_80
timestamp 1670092720
transform 1 0 9184 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_107
timestamp 1670092720
transform 1 0 12208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_135
timestamp 1670092720
transform 1 0 15344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_137
timestamp 1670092720
transform 1 0 15568 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_140
timestamp 1670092720
transform 1 0 15904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_144
timestamp 1670092720
transform 1 0 16352 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_2 $PDK_ROOT/$PDK/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670092720
transform 1 0 448 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_18
timestamp 1670092720
transform 1 0 2240 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_26
timestamp 1670092720
transform 1 0 3136 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_30
timestamp 1670092720
transform 1 0 3584 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1670092720
transform 1 0 4032 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_37
timestamp 1670092720
transform 1 0 4368 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_40
timestamp 1670092720
transform 1 0 4704 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_44 $PDK_ROOT/$PDK/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670092720
transform 1 0 5152 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_76
timestamp 1670092720
transform 1 0 8736 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_92
timestamp 1670092720
transform 1 0 10528 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_96
timestamp 1670092720
transform 1 0 10976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_98
timestamp 1670092720
transform 1 0 11200 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_101
timestamp 1670092720
transform 1 0 11536 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1670092720
transform 1 0 11984 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_108
timestamp 1670092720
transform 1 0 12320 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_111
timestamp 1670092720
transform 1 0 12656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_115
timestamp 1670092720
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_117
timestamp 1670092720
transform 1 0 13328 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_144
timestamp 1670092720
transform 1 0 16352 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_2
timestamp 1670092720
transform 1 0 448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_18
timestamp 1670092720
transform 1 0 2240 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_20
timestamp 1670092720
transform 1 0 2464 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_47
timestamp 1670092720
transform 1 0 5488 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_51
timestamp 1670092720
transform 1 0 5936 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_67
timestamp 1670092720
transform 1 0 7728 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_73
timestamp 1670092720
transform 1 0 8400 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_81
timestamp 1670092720
transform 1 0 9296 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_85
timestamp 1670092720
transform 1 0 9744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_113
timestamp 1670092720
transform 1 0 12880 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1670092720
transform 1 0 16016 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_144
timestamp 1670092720
transform 1 0 16352 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1670092720
transform 1 0 448 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1670092720
transform 1 0 4032 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_37
timestamp 1670092720
transform 1 0 4368 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_53
timestamp 1670092720
transform 1 0 6160 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_87
timestamp 1670092720
transform 1 0 9968 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_91
timestamp 1670092720
transform 1 0 10416 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_99
timestamp 1670092720
transform 1 0 11312 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_103
timestamp 1670092720
transform 1 0 11760 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1670092720
transform 1 0 11984 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_108
timestamp 1670092720
transform 1 0 12320 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_138
timestamp 1670092720
transform 1 0 15680 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_144
timestamp 1670092720
transform 1 0 16352 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_2
timestamp 1670092720
transform 1 0 448 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_29
timestamp 1670092720
transform 1 0 3472 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_33
timestamp 1670092720
transform 1 0 3920 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_65
timestamp 1670092720
transform 1 0 7504 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_69
timestamp 1670092720
transform 1 0 7952 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_73
timestamp 1670092720
transform 1 0 8400 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_76
timestamp 1670092720
transform 1 0 8736 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_134
timestamp 1670092720
transform 1 0 15232 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_138
timestamp 1670092720
transform 1 0 15680 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_144
timestamp 1670092720
transform 1 0 16352 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_2
timestamp 1670092720
transform 1 0 448 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_29
timestamp 1670092720
transform 1 0 3472 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_33
timestamp 1670092720
transform 1 0 3920 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_37
timestamp 1670092720
transform 1 0 4368 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_53
timestamp 1670092720
transform 1 0 6160 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_63
timestamp 1670092720
transform 1 0 7280 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_91
timestamp 1670092720
transform 1 0 10416 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_95
timestamp 1670092720
transform 1 0 10864 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_103
timestamp 1670092720
transform 1 0 11760 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1670092720
transform 1 0 11984 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_108
timestamp 1670092720
transform 1 0 12320 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_116
timestamp 1670092720
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_144
timestamp 1670092720
transform 1 0 16352 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_2
timestamp 1670092720
transform 1 0 448 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_4
timestamp 1670092720
transform 1 0 672 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_31
timestamp 1670092720
transform 1 0 3696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_35
timestamp 1670092720
transform 1 0 4144 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_43
timestamp 1670092720
transform 1 0 5040 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1670092720
transform 1 0 8064 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_73
timestamp 1670092720
transform 1 0 8400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_103
timestamp 1670092720
transform 1 0 11760 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_107
timestamp 1670092720
transform 1 0 12208 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1670092720
transform 1 0 16016 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_144
timestamp 1670092720
transform 1 0 16352 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_2
timestamp 1670092720
transform 1 0 448 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_6
timestamp 1670092720
transform 1 0 896 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1670092720
transform 1 0 4032 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_37
timestamp 1670092720
transform 1 0 4368 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_40
timestamp 1670092720
transform 1 0 4704 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_44
timestamp 1670092720
transform 1 0 5152 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_46
timestamp 1670092720
transform 1 0 5376 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_73
timestamp 1670092720
transform 1 0 8400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_101
timestamp 1670092720
transform 1 0 11536 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1670092720
transform 1 0 11984 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_108
timestamp 1670092720
transform 1 0 12320 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_135
timestamp 1670092720
transform 1 0 15344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_139
timestamp 1670092720
transform 1 0 15792 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_143
timestamp 1670092720
transform 1 0 16240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_2
timestamp 1670092720
transform 1 0 448 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_29
timestamp 1670092720
transform 1 0 3472 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_33
timestamp 1670092720
transform 1 0 3920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_37
timestamp 1670092720
transform 1 0 4368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_41
timestamp 1670092720
transform 1 0 4816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_69
timestamp 1670092720
transform 1 0 7952 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_72
timestamp 1670092720
transform 1 0 8288 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_99
timestamp 1670092720
transform 1 0 11312 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_103
timestamp 1670092720
transform 1 0 11760 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_107
timestamp 1670092720
transform 1 0 12208 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_110
timestamp 1670092720
transform 1 0 12544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_112
timestamp 1670092720
transform 1 0 12768 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_139
timestamp 1670092720
transform 1 0 15792 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_142
timestamp 1670092720
transform 1 0 16128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_144
timestamp 1670092720
transform 1 0 16352 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 $PDK_ROOT/$PDK/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670092720
transform 1 0 224 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1670092720
transform -1 0 16688 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1670092720
transform 1 0 224 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1670092720
transform -1 0 16688 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1670092720
transform 1 0 224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1670092720
transform -1 0 16688 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1670092720
transform 1 0 224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1670092720
transform -1 0 16688 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1670092720
transform 1 0 224 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1670092720
transform -1 0 16688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1670092720
transform 1 0 224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1670092720
transform -1 0 16688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1670092720
transform 1 0 224 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1670092720
transform -1 0 16688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1670092720
transform 1 0 224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1670092720
transform -1 0 16688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1670092720
transform 1 0 224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1670092720
transform -1 0 16688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1670092720
transform 1 0 224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1670092720
transform -1 0 16688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1670092720
transform 1 0 224 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1670092720
transform -1 0 16688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1670092720
transform 1 0 224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1670092720
transform -1 0 16688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_24 $PDK_ROOT/$PDK/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1670092720
transform 1 0 4144 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_25
timestamp 1670092720
transform 1 0 8064 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_26
timestamp 1670092720
transform 1 0 11984 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_27
timestamp 1670092720
transform 1 0 15904 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_28
timestamp 1670092720
transform 1 0 8176 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_29
timestamp 1670092720
transform 1 0 16128 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_30
timestamp 1670092720
transform 1 0 4144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_31
timestamp 1670092720
transform 1 0 12096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_32
timestamp 1670092720
transform 1 0 8176 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_33
timestamp 1670092720
transform 1 0 16128 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_34
timestamp 1670092720
transform 1 0 4144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_35
timestamp 1670092720
transform 1 0 12096 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_36
timestamp 1670092720
transform 1 0 8176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_37
timestamp 1670092720
transform 1 0 16128 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_38
timestamp 1670092720
transform 1 0 4144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_39
timestamp 1670092720
transform 1 0 12096 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_40
timestamp 1670092720
transform 1 0 8176 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_41
timestamp 1670092720
transform 1 0 16128 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_42
timestamp 1670092720
transform 1 0 4144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_43
timestamp 1670092720
transform 1 0 12096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_44
timestamp 1670092720
transform 1 0 8176 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_45
timestamp 1670092720
transform 1 0 16128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_46
timestamp 1670092720
transform 1 0 4144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_47
timestamp 1670092720
transform 1 0 12096 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_48
timestamp 1670092720
transform 1 0 4144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_49
timestamp 1670092720
transform 1 0 8064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_50
timestamp 1670092720
transform 1 0 11984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_51
timestamp 1670092720
transform 1 0 15904 0 -1 10976
box -86 -86 310 870
<< labels >>
flabel metal4 s 2122 1508 2442 11036 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 6238 1508 6558 11036 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 10354 1508 10674 11036 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 14470 1508 14790 11036 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 4180 1508 4500 11036 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 8296 1508 8616 11036 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 12412 1508 12732 11036 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 16528 1508 16848 11036 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal2 s 560 0 672 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[0]
port 2 nsew signal input
flabel metal2 s 5040 0 5152 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[10]
port 3 nsew signal input
flabel metal2 s 5488 0 5600 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[11]
port 4 nsew signal input
flabel metal2 s 5936 0 6048 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[12]
port 5 nsew signal input
flabel metal2 s 6384 0 6496 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[13]
port 6 nsew signal input
flabel metal2 s 6832 0 6944 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[14]
port 7 nsew signal input
flabel metal2 s 7280 0 7392 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[15]
port 8 nsew signal input
flabel metal2 s 7728 0 7840 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[16]
port 9 nsew signal input
flabel metal2 s 8176 0 8288 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[17]
port 10 nsew signal input
flabel metal2 s 1008 0 1120 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[1]
port 11 nsew signal input
flabel metal2 s 1456 0 1568 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[2]
port 12 nsew signal input
flabel metal2 s 1904 0 2016 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[3]
port 13 nsew signal input
flabel metal2 s 2352 0 2464 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[4]
port 14 nsew signal input
flabel metal2 s 2800 0 2912 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[5]
port 15 nsew signal input
flabel metal2 s 3248 0 3360 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[6]
port 16 nsew signal input
flabel metal2 s 3696 0 3808 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[7]
port 17 nsew signal input
flabel metal2 s 4144 0 4256 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[8]
port 18 nsew signal input
flabel metal2 s 4592 0 4704 800 0 FreeSans 448 90 0 0 mgmt_gpio_in[9]
port 19 nsew signal input
flabel metal2 s 560 12200 672 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[0]
port 20 nsew signal tristate
flabel metal2 s 5040 12200 5152 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[10]
port 21 nsew signal tristate
flabel metal2 s 5488 12200 5600 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[11]
port 22 nsew signal tristate
flabel metal2 s 5936 12200 6048 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[12]
port 23 nsew signal tristate
flabel metal2 s 6384 12200 6496 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[13]
port 24 nsew signal tristate
flabel metal2 s 6832 12200 6944 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[14]
port 25 nsew signal tristate
flabel metal2 s 7280 12200 7392 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[15]
port 26 nsew signal tristate
flabel metal2 s 7728 12200 7840 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[16]
port 27 nsew signal tristate
flabel metal2 s 8176 12200 8288 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[17]
port 28 nsew signal tristate
flabel metal2 s 1008 12200 1120 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[1]
port 29 nsew signal tristate
flabel metal2 s 1456 12200 1568 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[2]
port 30 nsew signal tristate
flabel metal2 s 1904 12200 2016 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[3]
port 31 nsew signal tristate
flabel metal2 s 2352 12200 2464 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[4]
port 32 nsew signal tristate
flabel metal2 s 2800 12200 2912 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[5]
port 33 nsew signal tristate
flabel metal2 s 3248 12200 3360 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[6]
port 34 nsew signal tristate
flabel metal2 s 3696 12200 3808 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[7]
port 35 nsew signal tristate
flabel metal2 s 4144 12200 4256 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[8]
port 36 nsew signal tristate
flabel metal2 s 4592 12200 4704 13000 0 FreeSans 448 90 0 0 mgmt_gpio_in_buf[9]
port 37 nsew signal tristate
flabel metal3 s 0 2128 800 2240 0 FreeSans 448 0 0 0 mgmt_gpio_oeb[0]
port 38 nsew signal input
flabel metal3 s 0 6384 800 6496 0 FreeSans 448 0 0 0 mgmt_gpio_oeb[1]
port 39 nsew signal input
flabel metal3 s 0 10640 800 10752 0 FreeSans 448 0 0 0 mgmt_gpio_oeb[2]
port 40 nsew signal input
flabel metal3 s 16200 2128 17000 2240 0 FreeSans 448 0 0 0 mgmt_gpio_oeb_buf[0]
port 41 nsew signal tristate
flabel metal3 s 16200 6384 17000 6496 0 FreeSans 448 0 0 0 mgmt_gpio_oeb_buf[1]
port 42 nsew signal tristate
flabel metal3 s 16200 10640 17000 10752 0 FreeSans 448 0 0 0 mgmt_gpio_oeb_buf[2]
port 43 nsew signal tristate
flabel metal2 s 8624 12200 8736 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[0]
port 44 nsew signal input
flabel metal2 s 13104 12200 13216 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[10]
port 45 nsew signal input
flabel metal2 s 13552 12200 13664 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[11]
port 46 nsew signal input
flabel metal2 s 14000 12200 14112 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[12]
port 47 nsew signal input
flabel metal2 s 14448 12200 14560 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[13]
port 48 nsew signal input
flabel metal2 s 14896 12200 15008 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[14]
port 49 nsew signal input
flabel metal2 s 15344 12200 15456 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[15]
port 50 nsew signal input
flabel metal2 s 15792 12200 15904 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[16]
port 51 nsew signal input
flabel metal2 s 16240 12200 16352 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[17]
port 52 nsew signal input
flabel metal2 s 9072 12200 9184 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[1]
port 53 nsew signal input
flabel metal2 s 9520 12200 9632 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[2]
port 54 nsew signal input
flabel metal2 s 9968 12200 10080 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[3]
port 55 nsew signal input
flabel metal2 s 10416 12200 10528 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[4]
port 56 nsew signal input
flabel metal2 s 10864 12200 10976 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[5]
port 57 nsew signal input
flabel metal2 s 11312 12200 11424 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[6]
port 58 nsew signal input
flabel metal2 s 11760 12200 11872 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[7]
port 59 nsew signal input
flabel metal2 s 12208 12200 12320 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[8]
port 60 nsew signal input
flabel metal2 s 12656 12200 12768 13000 0 FreeSans 448 90 0 0 mgmt_gpio_out[9]
port 61 nsew signal input
flabel metal2 s 8624 0 8736 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[0]
port 62 nsew signal tristate
flabel metal2 s 13104 0 13216 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[10]
port 63 nsew signal tristate
flabel metal2 s 13552 0 13664 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[11]
port 64 nsew signal tristate
flabel metal2 s 14000 0 14112 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[12]
port 65 nsew signal tristate
flabel metal2 s 14448 0 14560 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[13]
port 66 nsew signal tristate
flabel metal2 s 14896 0 15008 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[14]
port 67 nsew signal tristate
flabel metal2 s 15344 0 15456 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[15]
port 68 nsew signal tristate
flabel metal2 s 15792 0 15904 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[16]
port 69 nsew signal tristate
flabel metal2 s 16240 0 16352 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[17]
port 70 nsew signal tristate
flabel metal2 s 9072 0 9184 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[1]
port 71 nsew signal tristate
flabel metal2 s 9520 0 9632 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[2]
port 72 nsew signal tristate
flabel metal2 s 9968 0 10080 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[3]
port 73 nsew signal tristate
flabel metal2 s 10416 0 10528 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[4]
port 74 nsew signal tristate
flabel metal2 s 10864 0 10976 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[5]
port 75 nsew signal tristate
flabel metal2 s 11312 0 11424 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[6]
port 76 nsew signal tristate
flabel metal2 s 11760 0 11872 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[7]
port 77 nsew signal tristate
flabel metal2 s 12208 0 12320 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[8]
port 78 nsew signal tristate
flabel metal2 s 12656 0 12768 800 0 FreeSans 448 90 0 0 mgmt_gpio_out_buf[9]
port 79 nsew signal tristate
rlabel metal1 8456 10192 8456 10192 0 VDD
rlabel via1 8536 10976 8536 10976 0 VSS
rlabel metal3 1680 8232 1680 8232 0 mgmt_gpio_in[0]
rlabel metal2 6776 1904 6776 1904 0 mgmt_gpio_in[10]
rlabel metal2 6776 3472 6776 3472 0 mgmt_gpio_in[11]
rlabel metal2 7000 4032 7000 4032 0 mgmt_gpio_in[12]
rlabel metal2 7448 2408 7448 2408 0 mgmt_gpio_in[13]
rlabel metal2 6888 4578 6888 4578 0 mgmt_gpio_in[14]
rlabel metal2 7224 2520 7224 2520 0 mgmt_gpio_in[15]
rlabel metal2 7784 4046 7784 4046 0 mgmt_gpio_in[16]
rlabel metal2 8232 3374 8232 3374 0 mgmt_gpio_in[17]
rlabel metal2 2744 7168 2744 7168 0 mgmt_gpio_in[1]
rlabel metal2 1512 2478 1512 2478 0 mgmt_gpio_in[2]
rlabel metal2 2968 8736 2968 8736 0 mgmt_gpio_in[3]
rlabel metal2 2408 1470 2408 1470 0 mgmt_gpio_in[4]
rlabel metal2 3976 3864 3976 3864 0 mgmt_gpio_in[5]
rlabel metal2 3360 3528 3360 3528 0 mgmt_gpio_in[6]
rlabel metal3 4256 5880 4256 5880 0 mgmt_gpio_in[7]
rlabel metal3 2856 1960 2856 1960 0 mgmt_gpio_in[8]
rlabel metal2 4872 2744 4872 2744 0 mgmt_gpio_in[9]
rlabel metal2 952 8372 952 8372 0 mgmt_gpio_in_buf[0]
rlabel metal2 5096 7154 5096 7154 0 mgmt_gpio_in_buf[10]
rlabel metal2 5544 7938 5544 7938 0 mgmt_gpio_in_buf[11]
rlabel metal2 5992 8218 5992 8218 0 mgmt_gpio_in_buf[12]
rlabel metal2 6608 3752 6608 3752 0 mgmt_gpio_in_buf[13]
rlabel metal2 6888 11354 6888 11354 0 mgmt_gpio_in_buf[14]
rlabel metal2 6552 9072 6552 9072 0 mgmt_gpio_in_buf[15]
rlabel metal2 7112 9968 7112 9968 0 mgmt_gpio_in_buf[16]
rlabel metal2 8232 9506 8232 9506 0 mgmt_gpio_in_buf[17]
rlabel metal2 1064 9786 1064 9786 0 mgmt_gpio_in_buf[1]
rlabel metal2 1512 11466 1512 11466 0 mgmt_gpio_in_buf[2]
rlabel metal2 1960 10570 1960 10570 0 mgmt_gpio_in_buf[3]
rlabel metal2 2520 10304 2520 10304 0 mgmt_gpio_in_buf[4]
rlabel metal2 2856 8218 2856 8218 0 mgmt_gpio_in_buf[5]
rlabel metal2 2912 3640 2912 3640 0 mgmt_gpio_in_buf[6]
rlabel metal2 3696 10696 3696 10696 0 mgmt_gpio_in_buf[7]
rlabel metal3 3640 5096 3640 5096 0 mgmt_gpio_in_buf[8]
rlabel metal3 3640 5544 3640 5544 0 mgmt_gpio_in_buf[9]
rlabel metal2 8680 2464 8680 2464 0 mgmt_gpio_oeb[0]
rlabel metal3 854 6440 854 6440 0 mgmt_gpio_oeb[1]
rlabel metal2 12488 9800 12488 9800 0 mgmt_gpio_oeb[2]
rlabel metal2 11032 2408 11032 2408 0 mgmt_gpio_oeb_buf[0]
rlabel metal2 15064 6216 15064 6216 0 mgmt_gpio_oeb_buf[1]
rlabel metal2 14392 10304 14392 10304 0 mgmt_gpio_oeb_buf[2]
rlabel metal3 9184 8232 9184 8232 0 mgmt_gpio_out[0]
rlabel metal2 11704 2128 11704 2128 0 mgmt_gpio_out[10]
rlabel metal2 14504 7616 14504 7616 0 mgmt_gpio_out[11]
rlabel metal2 15512 5600 15512 5600 0 mgmt_gpio_out[12]
rlabel metal2 15176 10864 15176 10864 0 mgmt_gpio_out[13]
rlabel metal2 15624 5880 15624 5880 0 mgmt_gpio_out[14]
rlabel metal2 16072 9968 16072 9968 0 mgmt_gpio_out[15]
rlabel metal3 14280 5880 14280 5880 0 mgmt_gpio_out[16]
rlabel metal2 16240 8232 16240 8232 0 mgmt_gpio_out[17]
rlabel metal2 10584 10864 10584 10864 0 mgmt_gpio_out[1]
rlabel metal2 10808 9856 10808 9856 0 mgmt_gpio_out[2]
rlabel metal3 10528 9016 10528 9016 0 mgmt_gpio_out[3]
rlabel metal3 10976 5208 10976 5208 0 mgmt_gpio_out[4]
rlabel metal2 11312 5208 11312 5208 0 mgmt_gpio_out[5]
rlabel metal2 13832 4760 13832 4760 0 mgmt_gpio_out[6]
rlabel metal2 15288 3136 15288 3136 0 mgmt_gpio_out[7]
rlabel metal3 13496 3528 13496 3528 0 mgmt_gpio_out[8]
rlabel metal2 14616 4592 14616 4592 0 mgmt_gpio_out[9]
rlabel metal2 8680 1358 8680 1358 0 mgmt_gpio_out_buf[0]
rlabel metal2 13160 1414 13160 1414 0 mgmt_gpio_out_buf[10]
rlabel metal2 13608 4046 13608 4046 0 mgmt_gpio_out_buf[11]
rlabel metal2 14056 3766 14056 3766 0 mgmt_gpio_out_buf[12]
rlabel metal2 14504 1246 14504 1246 0 mgmt_gpio_out_buf[13]
rlabel metal2 14952 2982 14952 2982 0 mgmt_gpio_out_buf[14]
rlabel metal3 15064 8904 15064 8904 0 mgmt_gpio_out_buf[15]
rlabel metal2 15848 1750 15848 1750 0 mgmt_gpio_out_buf[16]
rlabel metal2 16296 3094 16296 3094 0 mgmt_gpio_out_buf[17]
rlabel metal2 9128 5614 9128 5614 0 mgmt_gpio_out_buf[1]
rlabel metal2 9576 5222 9576 5222 0 mgmt_gpio_out_buf[2]
rlabel metal2 10024 1974 10024 1974 0 mgmt_gpio_out_buf[3]
rlabel metal2 10472 1414 10472 1414 0 mgmt_gpio_out_buf[4]
rlabel metal2 10920 2198 10920 2198 0 mgmt_gpio_out_buf[5]
rlabel metal2 11368 1694 11368 1694 0 mgmt_gpio_out_buf[6]
rlabel metal2 11816 1246 11816 1246 0 mgmt_gpio_out_buf[7]
rlabel metal2 12264 2198 12264 2198 0 mgmt_gpio_out_buf[8]
rlabel metal2 12712 1078 12712 1078 0 mgmt_gpio_out_buf[9]
<< properties >>
string FIXED_BBOX 0 0 17000 13000
<< end >>
