magic
tech gf180mcuC
magscale 1 10
timestamp 1638586901
<< metal4 >>
rect -746 93 9893 373
<< metal5 >>
rect 5226 10173 5460 10266
tri 4620 10080 4713 10173 se
rect 4713 10080 5460 10173
tri 4526 9893 4620 9986 se
rect 4620 9893 5460 10080
tri 3753 9800 3846 9893 se
rect 3846 9800 4853 9893
rect 3753 9753 4853 9800
tri 3660 9613 3753 9706 se
rect 3753 9660 4760 9753
tri 4760 9660 4853 9753 nw
rect 3753 9613 3966 9660
tri 3966 9613 4013 9660 nw
rect 3360 9473 3966 9613
rect 5226 9566 5460 9893
rect 5226 9520 6440 9566
rect 3360 9380 3873 9473
tri 3873 9380 3966 9473 nw
tri 4853 9426 4946 9520 se
rect 4946 9426 6440 9520
tri 4340 9380 4386 9426 se
rect 4386 9380 6440 9426
tri 3920 8960 4340 9380 se
rect 4340 9333 6440 9380
rect 4340 9053 6253 9333
tri 6253 9240 6346 9333 nw
rect 4340 8960 6160 9053
tri 6160 8960 6253 9053 nw
tri 3826 8586 3920 8680 se
rect 3920 8586 6160 8960
rect 3826 8400 6160 8586
tri 6160 8400 6253 8493 sw
rect 1866 7746 2100 8213
rect 3826 8026 6253 8400
tri 3826 7933 3920 8026 ne
rect 3920 7933 6253 8026
tri 6253 7933 6440 8120 sw
rect 3920 7840 4853 7933
tri 4853 7840 4946 7933 nw
rect 5226 7840 6440 7933
rect 3920 7746 4475 7840
rect 1586 7466 2333 7746
tri 1586 7373 1680 7466 ne
rect 1680 7186 2240 7466
tri 2240 7373 2333 7466 nw
tri 3920 7404 4262 7746 ne
rect 4262 7404 4475 7746
tri 4475 7695 4620 7840 nw
rect 5226 7326 5506 7840
tri 5973 7653 6160 7840 ne
rect 6160 7653 6440 7840
tri 9053 7746 9333 8026 se
rect 9333 7746 9546 8026
tri 8773 7466 9053 7746 se
rect 5226 7280 7093 7326
tri 4853 7186 4946 7280 se
rect 4946 7186 7093 7280
rect 1866 6953 2100 7186
rect 4106 7093 7093 7186
tri 4060 6954 4106 7000 se
rect 4106 6954 6626 7093
rect 1866 6906 2893 6953
tri 4013 6906 4060 6953 se
rect 4060 6906 6626 6954
tri 6626 6906 6813 7093 nw
tri 1120 6813 1213 6906 se
rect 1213 6813 2893 6906
rect 560 6720 2893 6813
tri 93 6160 560 6626 se
rect 560 6253 2520 6720
tri 2520 6626 2613 6720 nw
tri 3640 6626 3920 6906 se
rect 3920 6720 6626 6906
rect 3920 6626 6346 6720
rect 560 6160 2426 6253
tri 2426 6160 2520 6253 nw
tri 3173 6160 3640 6626 se
rect 3640 6160 6346 6626
tri 6346 6440 6626 6720 nw
rect 7606 6673 7840 7000
tri 8120 6813 8773 7466 se
rect 8773 7280 9053 7466
tri 9053 7373 9426 7746 nw
rect 8773 7000 8960 7280
tri 8960 7186 9053 7280 nw
rect 8773 6813 8866 7000
tri 8866 6906 8960 7000 nw
tri 8073 6673 8120 6720 se
rect 8120 6673 8866 6813
rect 7606 6533 8866 6673
tri 0 5786 93 5880 se
rect 93 5786 2426 6160
rect 0 5413 2426 5786
tri 2800 5693 3173 6066 se
rect 3173 5693 6253 6160
tri 6253 6066 6346 6160 nw
tri 7513 6160 7606 6253 se
rect 7606 6160 8773 6533
tri 8773 6440 8866 6533 nw
tri 7466 6066 7513 6113 se
rect 7513 6066 8773 6160
tri 2426 5413 2520 5506 sw
rect 0 4946 2520 5413
tri 0 4853 93 4946 ne
rect 93 4573 2520 4946
rect -653 4386 -373 4433
tri -373 4386 -326 4433 sw
rect -653 4293 -280 4386
tri -280 4293 -186 4386 sw
tri 93 4293 373 4573 ne
rect 373 4480 2520 4573
tri 2753 5273 2800 5320 se
rect 2800 5273 6253 5693
rect 2753 4573 6253 5273
tri 6906 5413 7466 5973 se
rect 7466 5413 8680 6066
tri 8680 5973 8773 6066 nw
tri 6720 5040 6906 5226 se
rect 6906 5040 8680 5413
tri 6580 4853 6720 4993 se
rect 6720 4853 8680 5040
tri 6486 4573 6580 4666 se
rect 6580 4573 8680 4853
rect 2753 4480 8680 4573
tri 8680 4480 8773 4573 sw
rect 373 4386 1213 4480
tri 1213 4386 1306 4480 nw
tri 1586 4386 1680 4480 ne
rect 1680 4386 8773 4480
rect 373 4293 933 4386
rect -653 4200 -93 4293
tri -466 4080 -346 4200 ne
rect -346 4106 -93 4200
tri -93 4106 93 4293 sw
rect 466 4106 933 4293
tri 933 4200 1120 4386 nw
rect 1866 4293 8773 4386
rect -346 4080 186 4106
tri -253 3893 -66 4080 ne
rect -66 4060 186 4080
tri 186 4060 233 4106 sw
rect 466 4060 886 4106
tri 886 4060 933 4106 nw
rect -66 3893 886 4060
tri 26 3826 93 3893 ne
rect 93 3826 886 3893
tri 186 3733 280 3826 ne
rect 280 3733 1440 3826
tri 373 3640 466 3733 ne
rect 466 3640 1440 3733
tri 1440 3640 1626 3826 sw
rect 1866 3640 2146 4293
tri 2386 4200 2480 4293 ne
rect 2480 4200 8773 4293
tri 2520 4013 2706 4200 ne
rect 2706 4013 8773 4200
rect 466 3453 2146 3640
rect 2706 3920 7000 4013
tri 7000 3920 7093 4013 nw
rect 2706 3826 6720 3920
tri 6720 3826 6813 3920 nw
tri 2706 3453 3080 3826 ne
rect 3080 3480 6720 3826
tri 6720 3480 6906 3666 sw
rect 3080 3453 6906 3480
rect 653 3360 2146 3453
tri 2146 3360 2240 3453 sw
rect 3080 3360 4760 3453
tri 4760 3360 4853 3453 nw
tri 5133 3360 5226 3453 ne
rect 5226 3360 6906 3453
tri 653 3266 746 3360 ne
rect 746 3266 2426 3360
tri 2426 3266 2520 3360 sw
tri 933 2706 1493 3266 ne
rect 1493 2520 2800 3266
rect 3080 3173 4013 3360
tri 4013 3266 4106 3360 nw
tri 3080 2893 3360 3173 ne
rect 3360 2893 3733 3173
tri 3733 2893 4013 3173 nw
rect 5320 3173 6906 3360
tri 2800 2520 3173 2893 sw
tri 3360 2800 3453 2893 ne
rect 3453 2520 3733 2893
tri 1400 2333 1493 2426 se
rect 1493 2333 3733 2520
rect 1400 2240 3733 2333
tri 3733 2240 4013 2520 sw
rect 1400 2146 4200 2240
tri 4200 2146 4293 2240 sw
rect 1400 2053 4573 2146
tri 4573 2053 4666 2146 sw
rect 5320 2053 5693 3173
tri 5973 3080 6066 3173 ne
rect 6066 3080 6906 3173
tri 6906 3080 7186 3360 sw
tri 6440 2893 6626 3080 ne
rect 6626 2986 7186 3080
rect 7560 2986 7840 4013
tri 8120 3920 8213 4013 ne
rect 8213 3920 8773 4013
tri 8773 3920 8960 4106 sw
tri 8373 3546 8746 3920 ne
rect 8746 3546 8960 3920
tri 8306 3080 8493 3266 se
rect 8493 3173 9333 3266
tri 9333 3173 9426 3266 sw
rect 8493 3080 9426 3173
tri 8120 2986 8213 3080 se
rect 8213 2986 9426 3080
rect 6626 2940 9426 2986
rect 6626 2893 9333 2940
tri 6906 2706 7093 2893 ne
rect 7093 2706 9333 2893
rect 7093 2473 9893 2706
rect 7093 2426 9426 2473
tri 6440 2053 6813 2426 se
rect 6813 2333 9426 2426
rect 6813 2053 9333 2333
tri 9333 2240 9426 2333 nw
rect 1400 1866 9333 2053
rect 1400 1773 3966 1866
tri 1400 1680 1493 1773 ne
rect 1493 1586 3966 1773
rect 4200 1773 9333 1866
rect 4200 1586 4526 1773
rect 1493 1493 4526 1586
rect 4760 1680 9146 1773
tri 9146 1680 9240 1773 nw
rect 4760 1493 5133 1680
rect 1493 1400 5133 1493
rect 5366 1400 5693 1680
rect 5926 1400 6253 1680
rect 6486 1400 9146 1680
rect 1493 1306 9146 1400
tri 1493 1213 1586 1306 ne
rect 1586 1026 9053 1306
tri 9053 1213 9146 1306 nw
tri 1586 933 1680 1026 ne
rect 1680 840 8773 1026
tri 1680 560 1960 840 ne
rect 1960 466 8773 840
tri 8773 746 9053 1026 nw
tri 1960 373 2053 466 ne
rect 2053 373 8773 466
<< fillblock >>
rect -1680 7093 -1493 7280
rect -840 6906 10000 10373
rect -1306 6533 10000 6906
rect -840 0 10000 6533
<< end >>
