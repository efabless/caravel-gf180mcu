magic
tech gf180mcuD
magscale 1 10
timestamp 1655304105
<< metal1 >>
rect -90 227 -38 240
rect -90 -99 -38 -86
<< via1 >>
rect -90 -86 -38 227
<< metal2 >>
rect -92 227 -36 239
rect -92 -86 -90 227
rect -38 -86 -36 227
rect -92 -99 -36 -86
<< end >>
