magic
tech gf180mcuC
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 0 576 108 756
rect 216 576 324 756
rect 0 504 324 576
rect 36 432 288 504
rect 72 324 252 432
rect 36 252 288 324
rect 0 180 324 252
rect 0 0 108 180
rect 216 0 324 180
<< properties >>
string FIXED_BBOX 0 -216 432 756
<< end >>
