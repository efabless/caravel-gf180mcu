magic
tech gf180mcuD
magscale 1 10
timestamp 1655304105
<< pwell >>
rect -334 -532 334 532
<< mvnmos >>
rect -70 -276 70 324
<< mvndiff >>
rect -158 311 -70 324
rect -158 -263 -145 311
rect -99 -263 -70 311
rect -158 -276 -70 -263
rect 70 311 158 324
rect 70 -263 99 311
rect 145 -263 158 311
rect 70 -276 158 -263
<< mvndiffc >>
rect -145 -263 -99 311
rect 99 -263 145 311
<< mvpsubdiff >>
rect -302 487 302 500
rect -302 441 -186 487
rect 186 441 302 487
rect -302 428 302 441
rect -302 384 -230 428
rect -302 -384 -289 384
rect -243 -384 -230 384
rect 230 384 302 428
rect -302 -428 -230 -384
rect 230 -384 243 384
rect 289 -384 302 384
rect 230 -428 302 -384
rect -302 -500 302 -428
<< mvpsubdiffcont >>
rect -186 441 186 487
rect -289 -384 -243 384
rect 243 -384 289 384
<< polysilicon >>
rect -70 324 70 368
rect -70 -309 70 -276
rect -70 -355 -57 -309
rect 57 -355 70 -309
rect -70 -368 70 -355
<< polycontact >>
rect -57 -355 57 -309
<< metal1 >>
rect -289 441 -186 487
rect 186 441 289 487
rect -289 384 -243 441
rect 243 384 289 441
rect -145 311 -99 322
rect -145 -274 -99 -263
rect 99 311 145 322
rect 99 -274 145 -263
rect -68 -355 -57 -309
rect 57 -355 68 -309
rect -289 -441 -243 -384
rect 243 -441 289 -384
rect -289 -487 289 -441
<< properties >>
string FIXED_BBOX -266 -464 266 464
string gencell nmos_6p0
string library gf180mcu
string parameters w 3.0 l 0.7 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.6 wmin 0.3 full_metal 1 compatible {nmos_3p3 nmos_6p0 nmos_6p0_nat}
<< end >>
