* NGSPICE file created from gpio_control_block.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1 D RN SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlya_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlya_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

.subckt gpio_control_block VDD VSS gpio_defaults[0] gpio_defaults[1] gpio_defaults[2]
+ gpio_defaults[3] gpio_defaults[4] gpio_defaults[5] gpio_defaults[6] gpio_defaults[7]
+ gpio_defaults[8] gpio_defaults[9] mgmt_gpio_in mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_drive_sel[0]
+ pad_gpio_drive_sel[1] pad_gpio_in pad_gpio_inen pad_gpio_out pad_gpio_outen pad_gpio_pulldown_sel
+ pad_gpio_pullup_sel pad_gpio_schmitt_sel pad_gpio_slew_sel resetn resetn_out serial_clock
+ serial_clock_out serial_data_in serial_data_out serial_load serial_load_out user_gpio_in
+ user_gpio_oeb user_gpio_out zero
XANTENNA__074__I resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_062_ _056_/Z gpio_defaults[1] _063_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_045_ _091_/Q mgmt_gpio_oeb _046_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_114_ serial_load serial_load_out VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__092__CLK serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_101 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__109__RN resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_061_ _060_/Z gpio_defaults[0] _061_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_044_ _092_/Q _050_/B1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_113_ serial_clock serial_clock_out VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__062__A2 gpio_defaults[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__071__A2 gpio_defaults[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_102 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_060_ _077_/I _060_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_112_ resetn resetn_out VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_103 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__052__I0 user_gpio_out VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_111_ pad_gpio_in mgmt_gpio_in VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__095__CLK serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_104 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__052__I1 mgmt_gpio_out VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__110__CLK serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__065__A2 gpio_defaults[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_110_ _110_/D resetn serial_clock _110_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_105 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__100__CLK serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__102__RN resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__098__CLK serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_099_ _109_/D _086_/Z _087_/ZN serial_load pad_gpio_pullup_sel VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1
XFILLER_31_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_37_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__113__I serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__068__A2 gpio_defaults[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_098_ _110_/Q _083_/Z _084_/ZN serial_load pad_gpio_drive_sel[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1
XANTENNA__103__CLK serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_097_ _110_/D _080_/Z _081_/ZN serial_load pad_gpio_drive_sel[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1
XFILLER_1_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__105__RN resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_096_ _106_/D _076_/Z _078_/ZN serial_load pad_gpio_schmitt_sel VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1
XFILLER_1_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_079_ _074_/Z gpio_defaults[8] _080_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__106__CLK serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_095_ _107_/D _072_/Z _073_/ZN serial_load pad_gpio_slew_sel VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1
XFILLER_24_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__056__I resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_078_ _077_/Z gpio_defaults[4] _078_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__059__I resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_094_ _105_/D _069_/Z _070_/ZN serial_load _094_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1
XFILLER_10_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_077_ _077_/I _077_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__108__RN resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__091__CLK serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_093_ _104_/D _066_/Z _067_/ZN serial_load pad_gpio_inen VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1
XFILLER_24_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__061__A2 gpio_defaults[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__070__A2 gpio_defaults[3] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_076_ _076_/I _076_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_90 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_059_ resetn _077_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__109__CLK serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_092_ _103_/D _063_/Z _064_/ZN serial_load _092_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1
XTAP_91 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_058_ _058_/I _058_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_075_ _074_/Z gpio_defaults[4] _076_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_19_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_091_ _102_/D _058_/Z _061_/ZN serial_load _091_/Q VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1
XANTENNA__094__CLK serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_074_ resetn _074_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_92 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_057_ _056_/Z gpio_defaults[0] _058_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_32_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_21_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_109_ _109_/D resetn serial_clock _110_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__064__A2 gpio_defaults[1] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__073__A2 gpio_defaults[5] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_93 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__082__A2 gpio_defaults[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_090_ _077_/Z gpio_defaults[6] _090_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_056_ resetn _056_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_073_ _060_/Z gpio_defaults[5] _073_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_108_ _108_/D resetn serial_clock _109_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_072_ _072_/I _072_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_94 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_055_ _055_/I serial_data_out VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__101__RN resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__110__RN resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_107_ _107_/D resetn serial_clock _108_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__097__CLK serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_071_ _056_/Z gpio_defaults[5] _072_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_95 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_84 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_106_ _106_/D resetn serial_clock _107_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_054_ one _054_/A2 _055_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__085__A2 gpio_defaults[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__067__A2 gpio_defaults[2] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_070_ _060_/Z gpio_defaults[3] _070_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_96 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__111__I pad_gpio_in VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_85 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__102__CLK serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_80 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_053_ _053_/I pad_gpio_out VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_105_ _105_/D resetn serial_clock _106_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__114__I serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_81 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_97 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_86 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__104__RN resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_104_ _104_/D resetn serial_clock _105_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_052_ user_gpio_out mgmt_gpio_out _091_/Q _053_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_98 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_87 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_21_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_051_ _051_/I pad_gpio_outen VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_103_ _103_/D resetn serial_clock _104_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__088__A2 gpio_defaults[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__079__A2 gpio_defaults[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_83 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_99 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__105__CLK serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_88 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_102_ _102_/D resetn serial_clock _103_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_32_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_050_ _050_/A1 _050_/A2 _050_/B1 _050_/B2 _051_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_40_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_89 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_2_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__107__RN resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_101_ serial_data_in resetn serial_clock _102_/D VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_22_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_74 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_100_ _108_/D _089_/Z _090_/ZN serial_load pad_gpio_pulldown_sel VDD VSS gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1
XFILLER_0_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__108__CLK serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__101__D serial_data_in VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xconst_source_zero zero VDD VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_75 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_17_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xdata_delay_1 _110_/Q data_delay_2/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlya_2
XPHY_76 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__093__CLK serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_089_ _089_/I _089_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xdata_delay_2 data_delay_2/I _054_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__dlya_2
XANTENNA__081__A2 gpio_defaults[8] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__090__A2 gpio_defaults[6] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_77 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__045__A2 mgmt_gpio_oeb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_088_ _074_/Z gpio_defaults[6] _089_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_33_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_087_ _077_/Z gpio_defaults[7] _087_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__096__CLK serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_79 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_086_ _086_/I _086_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_069_ _069_/I _069_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__084__A2 gpio_defaults[9] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__057__A2 gpio_defaults[0] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__075__A2 gpio_defaults[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__101__CLK serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_085_ _074_/Z gpio_defaults[7] _086_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_068_ _056_/Z gpio_defaults[3] _069_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__112__I resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__103__RN resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_067_ _060_/Z gpio_defaults[2] _067_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__099__CLK serial_load VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_084_ _077_/Z gpio_defaults[9] _084_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__115__I pad_gpio_in VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_083_ _083_/I _083_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_066_ _066_/I _066_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_049_ _094_/Q _050_/B2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__078__A2 gpio_defaults[4] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__087__A2 gpio_defaults[7] VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__104__CLK serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_065_ _056_/Z gpio_defaults[2] _066_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_082_ _074_/Z gpio_defaults[9] _083_/I VDD VSS gf180mcu_fd_sc_mcu7t5v0__or2_1
X_048_ _048_/A1 _091_/Q _050_/A2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__106__RN resetn VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__047__I user_gpio_oeb VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_081_ _077_/Z gpio_defaults[8] _081_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_064_ _060_/Z gpio_defaults[1] _064_/ZN VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xconst_source_one one VDD VSS gf180mcu_fd_sc_mcu7t5v0__tieh
X_047_ user_gpio_oeb _048_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_063_ _063_/I _063_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_080_ _080_/I _080_/Z VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
X_046_ _050_/B1 _046_/A2 _050_/A1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_115_ pad_gpio_in user_gpio_in VDD VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__107__CLK serial_clock VDD VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_100 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

