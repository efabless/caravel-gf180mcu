magic
tech gf180mcuC
magscale 1 5
timestamp 1668824049
<< obsm1 >>
rect 672 463 51296 76145
<< metal2 >>
rect 840 77600 896 78000
rect 1568 77600 1624 78000
rect 2296 77600 2352 78000
rect 3024 77600 3080 78000
rect 3752 77600 3808 78000
rect 4480 77600 4536 78000
rect 5208 77600 5264 78000
rect 5936 77600 5992 78000
rect 6664 77600 6720 78000
rect 7392 77600 7448 78000
rect 8120 77600 8176 78000
rect 8848 77600 8904 78000
rect 9576 77600 9632 78000
rect 10304 77600 10360 78000
rect 11032 77600 11088 78000
rect 11760 77600 11816 78000
rect 12488 77600 12544 78000
rect 13216 77600 13272 78000
rect 13944 77600 14000 78000
rect 14672 77600 14728 78000
rect 15400 77600 15456 78000
rect 16128 77600 16184 78000
rect 16856 77600 16912 78000
rect 17584 77600 17640 78000
rect 18312 77600 18368 78000
rect 19040 77600 19096 78000
rect 19768 77600 19824 78000
rect 20496 77600 20552 78000
rect 21224 77600 21280 78000
rect 21952 77600 22008 78000
rect 22680 77600 22736 78000
rect 23408 77600 23464 78000
rect 24136 77600 24192 78000
rect 24864 77600 24920 78000
rect 25592 77600 25648 78000
rect 26320 77600 26376 78000
rect 27048 77600 27104 78000
rect 27776 77600 27832 78000
rect 28504 77600 28560 78000
rect 29232 77600 29288 78000
rect 29960 77600 30016 78000
rect 30688 77600 30744 78000
rect 31416 77600 31472 78000
rect 32144 77600 32200 78000
rect 32872 77600 32928 78000
rect 33600 77600 33656 78000
rect 34328 77600 34384 78000
rect 35056 77600 35112 78000
rect 35784 77600 35840 78000
rect 36512 77600 36568 78000
rect 37240 77600 37296 78000
rect 37968 77600 38024 78000
rect 38696 77600 38752 78000
rect 39424 77600 39480 78000
rect 40152 77600 40208 78000
rect 40880 77600 40936 78000
rect 41608 77600 41664 78000
rect 42336 77600 42392 78000
rect 43064 77600 43120 78000
rect 43792 77600 43848 78000
rect 44520 77600 44576 78000
rect 45248 77600 45304 78000
rect 45976 77600 46032 78000
rect 46704 77600 46760 78000
rect 47432 77600 47488 78000
rect 48160 77600 48216 78000
rect 48888 77600 48944 78000
rect 49616 77600 49672 78000
rect 50344 77600 50400 78000
rect 51072 77600 51128 78000
rect 1008 0 1064 400
rect 1568 0 1624 400
rect 2128 0 2184 400
rect 2688 0 2744 400
rect 3248 0 3304 400
rect 3808 0 3864 400
rect 4368 0 4424 400
rect 4928 0 4984 400
rect 5488 0 5544 400
rect 6048 0 6104 400
rect 6608 0 6664 400
rect 7168 0 7224 400
rect 7728 0 7784 400
rect 8288 0 8344 400
rect 8848 0 8904 400
rect 9408 0 9464 400
rect 9968 0 10024 400
rect 10528 0 10584 400
rect 11088 0 11144 400
rect 11648 0 11704 400
rect 12208 0 12264 400
rect 12768 0 12824 400
rect 13328 0 13384 400
rect 13888 0 13944 400
rect 14448 0 14504 400
rect 15008 0 15064 400
rect 15568 0 15624 400
rect 16128 0 16184 400
rect 16688 0 16744 400
rect 17248 0 17304 400
rect 17808 0 17864 400
rect 18368 0 18424 400
rect 18928 0 18984 400
rect 19488 0 19544 400
rect 20048 0 20104 400
rect 20608 0 20664 400
rect 21168 0 21224 400
rect 21728 0 21784 400
rect 22288 0 22344 400
rect 22848 0 22904 400
rect 23408 0 23464 400
rect 23968 0 24024 400
rect 24528 0 24584 400
rect 25088 0 25144 400
rect 25648 0 25704 400
rect 26208 0 26264 400
rect 26768 0 26824 400
rect 27328 0 27384 400
rect 27888 0 27944 400
rect 28448 0 28504 400
rect 29008 0 29064 400
rect 29568 0 29624 400
rect 30128 0 30184 400
rect 30688 0 30744 400
rect 31248 0 31304 400
rect 31808 0 31864 400
rect 32368 0 32424 400
rect 32928 0 32984 400
rect 33488 0 33544 400
rect 34048 0 34104 400
rect 34608 0 34664 400
rect 35168 0 35224 400
rect 35728 0 35784 400
rect 36288 0 36344 400
rect 36848 0 36904 400
rect 37408 0 37464 400
rect 37968 0 38024 400
rect 38528 0 38584 400
rect 39088 0 39144 400
rect 39648 0 39704 400
rect 40208 0 40264 400
rect 40768 0 40824 400
rect 41328 0 41384 400
rect 41888 0 41944 400
rect 42448 0 42504 400
rect 43008 0 43064 400
rect 43568 0 43624 400
rect 44128 0 44184 400
rect 44688 0 44744 400
rect 45248 0 45304 400
rect 45808 0 45864 400
rect 46368 0 46424 400
rect 46928 0 46984 400
rect 47488 0 47544 400
rect 48048 0 48104 400
rect 48608 0 48664 400
rect 49168 0 49224 400
rect 49728 0 49784 400
rect 50288 0 50344 400
rect 50848 0 50904 400
<< obsm2 >>
rect 574 77570 810 77658
rect 926 77570 1538 77658
rect 1654 77570 2266 77658
rect 2382 77570 2994 77658
rect 3110 77570 3722 77658
rect 3838 77570 4450 77658
rect 4566 77570 5178 77658
rect 5294 77570 5906 77658
rect 6022 77570 6634 77658
rect 6750 77570 7362 77658
rect 7478 77570 8090 77658
rect 8206 77570 8818 77658
rect 8934 77570 9546 77658
rect 9662 77570 10274 77658
rect 10390 77570 11002 77658
rect 11118 77570 11730 77658
rect 11846 77570 12458 77658
rect 12574 77570 13186 77658
rect 13302 77570 13914 77658
rect 14030 77570 14642 77658
rect 14758 77570 15370 77658
rect 15486 77570 16098 77658
rect 16214 77570 16826 77658
rect 16942 77570 17554 77658
rect 17670 77570 18282 77658
rect 18398 77570 19010 77658
rect 19126 77570 19738 77658
rect 19854 77570 20466 77658
rect 20582 77570 21194 77658
rect 21310 77570 21922 77658
rect 22038 77570 22650 77658
rect 22766 77570 23378 77658
rect 23494 77570 24106 77658
rect 24222 77570 24834 77658
rect 24950 77570 25562 77658
rect 25678 77570 26290 77658
rect 26406 77570 27018 77658
rect 27134 77570 27746 77658
rect 27862 77570 28474 77658
rect 28590 77570 29202 77658
rect 29318 77570 29930 77658
rect 30046 77570 30658 77658
rect 30774 77570 31386 77658
rect 31502 77570 32114 77658
rect 32230 77570 32842 77658
rect 32958 77570 33570 77658
rect 33686 77570 34298 77658
rect 34414 77570 35026 77658
rect 35142 77570 35754 77658
rect 35870 77570 36482 77658
rect 36598 77570 37210 77658
rect 37326 77570 37938 77658
rect 38054 77570 38666 77658
rect 38782 77570 39394 77658
rect 39510 77570 40122 77658
rect 40238 77570 40850 77658
rect 40966 77570 41578 77658
rect 41694 77570 42306 77658
rect 42422 77570 43034 77658
rect 43150 77570 43762 77658
rect 43878 77570 44490 77658
rect 44606 77570 45218 77658
rect 45334 77570 45946 77658
rect 46062 77570 46674 77658
rect 46790 77570 47402 77658
rect 47518 77570 48130 77658
rect 48246 77570 48858 77658
rect 48974 77570 49586 77658
rect 49702 77570 50314 77658
rect 50430 77570 51042 77658
rect 51158 77570 51786 77658
rect 574 430 51786 77570
rect 574 350 978 430
rect 1094 350 1538 430
rect 1654 350 2098 430
rect 2214 350 2658 430
rect 2774 350 3218 430
rect 3334 350 3778 430
rect 3894 350 4338 430
rect 4454 350 4898 430
rect 5014 350 5458 430
rect 5574 350 6018 430
rect 6134 350 6578 430
rect 6694 350 7138 430
rect 7254 350 7698 430
rect 7814 350 8258 430
rect 8374 350 8818 430
rect 8934 350 9378 430
rect 9494 350 9938 430
rect 10054 350 10498 430
rect 10614 350 11058 430
rect 11174 350 11618 430
rect 11734 350 12178 430
rect 12294 350 12738 430
rect 12854 350 13298 430
rect 13414 350 13858 430
rect 13974 350 14418 430
rect 14534 350 14978 430
rect 15094 350 15538 430
rect 15654 350 16098 430
rect 16214 350 16658 430
rect 16774 350 17218 430
rect 17334 350 17778 430
rect 17894 350 18338 430
rect 18454 350 18898 430
rect 19014 350 19458 430
rect 19574 350 20018 430
rect 20134 350 20578 430
rect 20694 350 21138 430
rect 21254 350 21698 430
rect 21814 350 22258 430
rect 22374 350 22818 430
rect 22934 350 23378 430
rect 23494 350 23938 430
rect 24054 350 24498 430
rect 24614 350 25058 430
rect 25174 350 25618 430
rect 25734 350 26178 430
rect 26294 350 26738 430
rect 26854 350 27298 430
rect 27414 350 27858 430
rect 27974 350 28418 430
rect 28534 350 28978 430
rect 29094 350 29538 430
rect 29654 350 30098 430
rect 30214 350 30658 430
rect 30774 350 31218 430
rect 31334 350 31778 430
rect 31894 350 32338 430
rect 32454 350 32898 430
rect 33014 350 33458 430
rect 33574 350 34018 430
rect 34134 350 34578 430
rect 34694 350 35138 430
rect 35254 350 35698 430
rect 35814 350 36258 430
rect 36374 350 36818 430
rect 36934 350 37378 430
rect 37494 350 37938 430
rect 38054 350 38498 430
rect 38614 350 39058 430
rect 39174 350 39618 430
rect 39734 350 40178 430
rect 40294 350 40738 430
rect 40854 350 41298 430
rect 41414 350 41858 430
rect 41974 350 42418 430
rect 42534 350 42978 430
rect 43094 350 43538 430
rect 43654 350 44098 430
rect 44214 350 44658 430
rect 44774 350 45218 430
rect 45334 350 45778 430
rect 45894 350 46338 430
rect 46454 350 46898 430
rect 47014 350 47458 430
rect 47574 350 48018 430
rect 48134 350 48578 430
rect 48694 350 49138 430
rect 49254 350 49698 430
rect 49814 350 50258 430
rect 50374 350 50818 430
rect 50934 350 51786 430
<< metal3 >>
rect 51600 76608 52000 76664
rect 0 75600 400 75656
rect 51600 75432 52000 75488
rect 0 74984 400 75040
rect 0 74368 400 74424
rect 51600 74256 52000 74312
rect 0 73752 400 73808
rect 0 73136 400 73192
rect 51600 73080 52000 73136
rect 0 72520 400 72576
rect 0 71904 400 71960
rect 51600 71904 52000 71960
rect 0 71288 400 71344
rect 0 70672 400 70728
rect 51600 70728 52000 70784
rect 0 70056 400 70112
rect 51600 69552 52000 69608
rect 0 69440 400 69496
rect 0 68824 400 68880
rect 51600 68376 52000 68432
rect 0 68208 400 68264
rect 0 67592 400 67648
rect 51600 67200 52000 67256
rect 0 66976 400 67032
rect 0 66360 400 66416
rect 51600 66024 52000 66080
rect 0 65744 400 65800
rect 0 65128 400 65184
rect 51600 64848 52000 64904
rect 0 64512 400 64568
rect 0 63896 400 63952
rect 51600 63672 52000 63728
rect 0 63280 400 63336
rect 0 62664 400 62720
rect 51600 62496 52000 62552
rect 0 62048 400 62104
rect 0 61432 400 61488
rect 51600 61320 52000 61376
rect 0 60816 400 60872
rect 0 60200 400 60256
rect 51600 60144 52000 60200
rect 0 59584 400 59640
rect 0 58968 400 59024
rect 51600 58968 52000 59024
rect 0 58352 400 58408
rect 0 57736 400 57792
rect 51600 57792 52000 57848
rect 0 57120 400 57176
rect 51600 56616 52000 56672
rect 0 56504 400 56560
rect 0 55888 400 55944
rect 51600 55440 52000 55496
rect 0 55272 400 55328
rect 0 54656 400 54712
rect 51600 54264 52000 54320
rect 0 54040 400 54096
rect 0 53424 400 53480
rect 51600 53088 52000 53144
rect 0 52808 400 52864
rect 0 52192 400 52248
rect 51600 51912 52000 51968
rect 0 51576 400 51632
rect 0 50960 400 51016
rect 51600 50736 52000 50792
rect 0 50344 400 50400
rect 0 49728 400 49784
rect 51600 49560 52000 49616
rect 0 49112 400 49168
rect 0 48496 400 48552
rect 51600 48384 52000 48440
rect 0 47880 400 47936
rect 0 47264 400 47320
rect 51600 47208 52000 47264
rect 0 46648 400 46704
rect 0 46032 400 46088
rect 51600 46032 52000 46088
rect 0 45416 400 45472
rect 0 44800 400 44856
rect 51600 44856 52000 44912
rect 0 44184 400 44240
rect 51600 43680 52000 43736
rect 0 43568 400 43624
rect 0 42952 400 43008
rect 51600 42504 52000 42560
rect 0 42336 400 42392
rect 0 41720 400 41776
rect 51600 41328 52000 41384
rect 0 41104 400 41160
rect 0 40488 400 40544
rect 51600 40152 52000 40208
rect 0 39872 400 39928
rect 0 39256 400 39312
rect 51600 38976 52000 39032
rect 0 38640 400 38696
rect 0 38024 400 38080
rect 51600 37800 52000 37856
rect 0 37408 400 37464
rect 0 36792 400 36848
rect 51600 36624 52000 36680
rect 0 36176 400 36232
rect 0 35560 400 35616
rect 51600 35448 52000 35504
rect 0 34944 400 35000
rect 0 34328 400 34384
rect 51600 34272 52000 34328
rect 0 33712 400 33768
rect 0 33096 400 33152
rect 51600 33096 52000 33152
rect 0 32480 400 32536
rect 0 31864 400 31920
rect 51600 31920 52000 31976
rect 0 31248 400 31304
rect 51600 30744 52000 30800
rect 0 30632 400 30688
rect 0 30016 400 30072
rect 51600 29568 52000 29624
rect 0 29400 400 29456
rect 0 28784 400 28840
rect 51600 28392 52000 28448
rect 0 28168 400 28224
rect 0 27552 400 27608
rect 51600 27216 52000 27272
rect 0 26936 400 26992
rect 0 26320 400 26376
rect 51600 26040 52000 26096
rect 0 25704 400 25760
rect 0 25088 400 25144
rect 51600 24864 52000 24920
rect 0 24472 400 24528
rect 0 23856 400 23912
rect 51600 23688 52000 23744
rect 0 23240 400 23296
rect 0 22624 400 22680
rect 51600 22512 52000 22568
rect 0 22008 400 22064
rect 0 21392 400 21448
rect 51600 21336 52000 21392
rect 0 20776 400 20832
rect 0 20160 400 20216
rect 51600 20160 52000 20216
rect 0 19544 400 19600
rect 0 18928 400 18984
rect 51600 18984 52000 19040
rect 0 18312 400 18368
rect 51600 17808 52000 17864
rect 0 17696 400 17752
rect 0 17080 400 17136
rect 51600 16632 52000 16688
rect 0 16464 400 16520
rect 0 15848 400 15904
rect 51600 15456 52000 15512
rect 0 15232 400 15288
rect 0 14616 400 14672
rect 51600 14280 52000 14336
rect 0 14000 400 14056
rect 0 13384 400 13440
rect 51600 13104 52000 13160
rect 0 12768 400 12824
rect 0 12152 400 12208
rect 51600 11928 52000 11984
rect 0 11536 400 11592
rect 0 10920 400 10976
rect 51600 10752 52000 10808
rect 0 10304 400 10360
rect 0 9688 400 9744
rect 51600 9576 52000 9632
rect 0 9072 400 9128
rect 0 8456 400 8512
rect 51600 8400 52000 8456
rect 0 7840 400 7896
rect 0 7224 400 7280
rect 51600 7224 52000 7280
rect 0 6608 400 6664
rect 0 5992 400 6048
rect 51600 6048 52000 6104
rect 0 5376 400 5432
rect 51600 4872 52000 4928
rect 0 4760 400 4816
rect 0 4144 400 4200
rect 51600 3696 52000 3752
rect 0 3528 400 3584
rect 0 2912 400 2968
rect 51600 2520 52000 2576
rect 0 2296 400 2352
rect 51600 1344 52000 1400
<< obsm3 >>
rect 400 76578 51570 76650
rect 400 75686 51791 76578
rect 430 75570 51791 75686
rect 400 75518 51791 75570
rect 400 75402 51570 75518
rect 400 75070 51791 75402
rect 430 74954 51791 75070
rect 400 74454 51791 74954
rect 430 74342 51791 74454
rect 430 74338 51570 74342
rect 400 74226 51570 74338
rect 400 73838 51791 74226
rect 430 73722 51791 73838
rect 400 73222 51791 73722
rect 430 73166 51791 73222
rect 430 73106 51570 73166
rect 400 73050 51570 73106
rect 400 72606 51791 73050
rect 430 72490 51791 72606
rect 400 71990 51791 72490
rect 430 71874 51570 71990
rect 400 71374 51791 71874
rect 430 71258 51791 71374
rect 400 70814 51791 71258
rect 400 70758 51570 70814
rect 430 70698 51570 70758
rect 430 70642 51791 70698
rect 400 70142 51791 70642
rect 430 70026 51791 70142
rect 400 69638 51791 70026
rect 400 69526 51570 69638
rect 430 69522 51570 69526
rect 430 69410 51791 69522
rect 400 68910 51791 69410
rect 430 68794 51791 68910
rect 400 68462 51791 68794
rect 400 68346 51570 68462
rect 400 68294 51791 68346
rect 430 68178 51791 68294
rect 400 67678 51791 68178
rect 430 67562 51791 67678
rect 400 67286 51791 67562
rect 400 67170 51570 67286
rect 400 67062 51791 67170
rect 430 66946 51791 67062
rect 400 66446 51791 66946
rect 430 66330 51791 66446
rect 400 66110 51791 66330
rect 400 65994 51570 66110
rect 400 65830 51791 65994
rect 430 65714 51791 65830
rect 400 65214 51791 65714
rect 430 65098 51791 65214
rect 400 64934 51791 65098
rect 400 64818 51570 64934
rect 400 64598 51791 64818
rect 430 64482 51791 64598
rect 400 63982 51791 64482
rect 430 63866 51791 63982
rect 400 63758 51791 63866
rect 400 63642 51570 63758
rect 400 63366 51791 63642
rect 430 63250 51791 63366
rect 400 62750 51791 63250
rect 430 62634 51791 62750
rect 400 62582 51791 62634
rect 400 62466 51570 62582
rect 400 62134 51791 62466
rect 430 62018 51791 62134
rect 400 61518 51791 62018
rect 430 61406 51791 61518
rect 430 61402 51570 61406
rect 400 61290 51570 61402
rect 400 60902 51791 61290
rect 430 60786 51791 60902
rect 400 60286 51791 60786
rect 430 60230 51791 60286
rect 430 60170 51570 60230
rect 400 60114 51570 60170
rect 400 59670 51791 60114
rect 430 59554 51791 59670
rect 400 59054 51791 59554
rect 430 58938 51570 59054
rect 400 58438 51791 58938
rect 430 58322 51791 58438
rect 400 57878 51791 58322
rect 400 57822 51570 57878
rect 430 57762 51570 57822
rect 430 57706 51791 57762
rect 400 57206 51791 57706
rect 430 57090 51791 57206
rect 400 56702 51791 57090
rect 400 56590 51570 56702
rect 430 56586 51570 56590
rect 430 56474 51791 56586
rect 400 55974 51791 56474
rect 430 55858 51791 55974
rect 400 55526 51791 55858
rect 400 55410 51570 55526
rect 400 55358 51791 55410
rect 430 55242 51791 55358
rect 400 54742 51791 55242
rect 430 54626 51791 54742
rect 400 54350 51791 54626
rect 400 54234 51570 54350
rect 400 54126 51791 54234
rect 430 54010 51791 54126
rect 400 53510 51791 54010
rect 430 53394 51791 53510
rect 400 53174 51791 53394
rect 400 53058 51570 53174
rect 400 52894 51791 53058
rect 430 52778 51791 52894
rect 400 52278 51791 52778
rect 430 52162 51791 52278
rect 400 51998 51791 52162
rect 400 51882 51570 51998
rect 400 51662 51791 51882
rect 430 51546 51791 51662
rect 400 51046 51791 51546
rect 430 50930 51791 51046
rect 400 50822 51791 50930
rect 400 50706 51570 50822
rect 400 50430 51791 50706
rect 430 50314 51791 50430
rect 400 49814 51791 50314
rect 430 49698 51791 49814
rect 400 49646 51791 49698
rect 400 49530 51570 49646
rect 400 49198 51791 49530
rect 430 49082 51791 49198
rect 400 48582 51791 49082
rect 430 48470 51791 48582
rect 430 48466 51570 48470
rect 400 48354 51570 48466
rect 400 47966 51791 48354
rect 430 47850 51791 47966
rect 400 47350 51791 47850
rect 430 47294 51791 47350
rect 430 47234 51570 47294
rect 400 47178 51570 47234
rect 400 46734 51791 47178
rect 430 46618 51791 46734
rect 400 46118 51791 46618
rect 430 46002 51570 46118
rect 400 45502 51791 46002
rect 430 45386 51791 45502
rect 400 44942 51791 45386
rect 400 44886 51570 44942
rect 430 44826 51570 44886
rect 430 44770 51791 44826
rect 400 44270 51791 44770
rect 430 44154 51791 44270
rect 400 43766 51791 44154
rect 400 43654 51570 43766
rect 430 43650 51570 43654
rect 430 43538 51791 43650
rect 400 43038 51791 43538
rect 430 42922 51791 43038
rect 400 42590 51791 42922
rect 400 42474 51570 42590
rect 400 42422 51791 42474
rect 430 42306 51791 42422
rect 400 41806 51791 42306
rect 430 41690 51791 41806
rect 400 41414 51791 41690
rect 400 41298 51570 41414
rect 400 41190 51791 41298
rect 430 41074 51791 41190
rect 400 40574 51791 41074
rect 430 40458 51791 40574
rect 400 40238 51791 40458
rect 400 40122 51570 40238
rect 400 39958 51791 40122
rect 430 39842 51791 39958
rect 400 39342 51791 39842
rect 430 39226 51791 39342
rect 400 39062 51791 39226
rect 400 38946 51570 39062
rect 400 38726 51791 38946
rect 430 38610 51791 38726
rect 400 38110 51791 38610
rect 430 37994 51791 38110
rect 400 37886 51791 37994
rect 400 37770 51570 37886
rect 400 37494 51791 37770
rect 430 37378 51791 37494
rect 400 36878 51791 37378
rect 430 36762 51791 36878
rect 400 36710 51791 36762
rect 400 36594 51570 36710
rect 400 36262 51791 36594
rect 430 36146 51791 36262
rect 400 35646 51791 36146
rect 430 35534 51791 35646
rect 430 35530 51570 35534
rect 400 35418 51570 35530
rect 400 35030 51791 35418
rect 430 34914 51791 35030
rect 400 34414 51791 34914
rect 430 34358 51791 34414
rect 430 34298 51570 34358
rect 400 34242 51570 34298
rect 400 33798 51791 34242
rect 430 33682 51791 33798
rect 400 33182 51791 33682
rect 430 33066 51570 33182
rect 400 32566 51791 33066
rect 430 32450 51791 32566
rect 400 32006 51791 32450
rect 400 31950 51570 32006
rect 430 31890 51570 31950
rect 430 31834 51791 31890
rect 400 31334 51791 31834
rect 430 31218 51791 31334
rect 400 30830 51791 31218
rect 400 30718 51570 30830
rect 430 30714 51570 30718
rect 430 30602 51791 30714
rect 400 30102 51791 30602
rect 430 29986 51791 30102
rect 400 29654 51791 29986
rect 400 29538 51570 29654
rect 400 29486 51791 29538
rect 430 29370 51791 29486
rect 400 28870 51791 29370
rect 430 28754 51791 28870
rect 400 28478 51791 28754
rect 400 28362 51570 28478
rect 400 28254 51791 28362
rect 430 28138 51791 28254
rect 400 27638 51791 28138
rect 430 27522 51791 27638
rect 400 27302 51791 27522
rect 400 27186 51570 27302
rect 400 27022 51791 27186
rect 430 26906 51791 27022
rect 400 26406 51791 26906
rect 430 26290 51791 26406
rect 400 26126 51791 26290
rect 400 26010 51570 26126
rect 400 25790 51791 26010
rect 430 25674 51791 25790
rect 400 25174 51791 25674
rect 430 25058 51791 25174
rect 400 24950 51791 25058
rect 400 24834 51570 24950
rect 400 24558 51791 24834
rect 430 24442 51791 24558
rect 400 23942 51791 24442
rect 430 23826 51791 23942
rect 400 23774 51791 23826
rect 400 23658 51570 23774
rect 400 23326 51791 23658
rect 430 23210 51791 23326
rect 400 22710 51791 23210
rect 430 22598 51791 22710
rect 430 22594 51570 22598
rect 400 22482 51570 22594
rect 400 22094 51791 22482
rect 430 21978 51791 22094
rect 400 21478 51791 21978
rect 430 21422 51791 21478
rect 430 21362 51570 21422
rect 400 21306 51570 21362
rect 400 20862 51791 21306
rect 430 20746 51791 20862
rect 400 20246 51791 20746
rect 430 20130 51570 20246
rect 400 19630 51791 20130
rect 430 19514 51791 19630
rect 400 19070 51791 19514
rect 400 19014 51570 19070
rect 430 18954 51570 19014
rect 430 18898 51791 18954
rect 400 18398 51791 18898
rect 430 18282 51791 18398
rect 400 17894 51791 18282
rect 400 17782 51570 17894
rect 430 17778 51570 17782
rect 430 17666 51791 17778
rect 400 17166 51791 17666
rect 430 17050 51791 17166
rect 400 16718 51791 17050
rect 400 16602 51570 16718
rect 400 16550 51791 16602
rect 430 16434 51791 16550
rect 400 15934 51791 16434
rect 430 15818 51791 15934
rect 400 15542 51791 15818
rect 400 15426 51570 15542
rect 400 15318 51791 15426
rect 430 15202 51791 15318
rect 400 14702 51791 15202
rect 430 14586 51791 14702
rect 400 14366 51791 14586
rect 400 14250 51570 14366
rect 400 14086 51791 14250
rect 430 13970 51791 14086
rect 400 13470 51791 13970
rect 430 13354 51791 13470
rect 400 13190 51791 13354
rect 400 13074 51570 13190
rect 400 12854 51791 13074
rect 430 12738 51791 12854
rect 400 12238 51791 12738
rect 430 12122 51791 12238
rect 400 12014 51791 12122
rect 400 11898 51570 12014
rect 400 11622 51791 11898
rect 430 11506 51791 11622
rect 400 11006 51791 11506
rect 430 10890 51791 11006
rect 400 10838 51791 10890
rect 400 10722 51570 10838
rect 400 10390 51791 10722
rect 430 10274 51791 10390
rect 400 9774 51791 10274
rect 430 9662 51791 9774
rect 430 9658 51570 9662
rect 400 9546 51570 9658
rect 400 9158 51791 9546
rect 430 9042 51791 9158
rect 400 8542 51791 9042
rect 430 8486 51791 8542
rect 430 8426 51570 8486
rect 400 8370 51570 8426
rect 400 7926 51791 8370
rect 430 7810 51791 7926
rect 400 7310 51791 7810
rect 430 7194 51570 7310
rect 400 6694 51791 7194
rect 430 6578 51791 6694
rect 400 6134 51791 6578
rect 400 6078 51570 6134
rect 430 6018 51570 6078
rect 430 5962 51791 6018
rect 400 5462 51791 5962
rect 430 5346 51791 5462
rect 400 4958 51791 5346
rect 400 4846 51570 4958
rect 430 4842 51570 4846
rect 430 4730 51791 4842
rect 400 4230 51791 4730
rect 430 4114 51791 4230
rect 400 3782 51791 4114
rect 400 3666 51570 3782
rect 400 3614 51791 3666
rect 430 3498 51791 3614
rect 400 2998 51791 3498
rect 430 2882 51791 2998
rect 400 2606 51791 2882
rect 400 2490 51570 2606
rect 400 2382 51791 2490
rect 430 2266 51791 2382
rect 400 1430 51791 2266
rect 400 1314 51570 1430
rect 400 854 51791 1314
<< metal4 >>
rect -418 478 -258 77138
rect -88 808 72 76808
rect 2224 478 2384 77138
rect 2554 478 2714 77138
rect 9904 478 10064 77138
rect 10234 478 10394 77138
rect 17584 478 17744 77138
rect 17914 478 18074 77138
rect 25264 478 25424 77138
rect 25594 478 25754 77138
rect 32944 478 33104 77138
rect 33274 478 33434 77138
rect 40624 478 40784 77138
rect 40954 478 41114 77138
rect 48304 478 48464 77138
rect 48634 478 48794 77138
rect 51896 808 52056 76808
rect 52226 478 52386 77138
<< obsm4 >>
rect 518 1353 2194 76375
rect 2414 1353 2524 76375
rect 2744 1353 9874 76375
rect 10094 1353 10204 76375
rect 10424 1353 17554 76375
rect 17774 1353 17884 76375
rect 18104 1353 25234 76375
rect 25454 1353 25564 76375
rect 25784 1353 32914 76375
rect 33134 1353 33244 76375
rect 33464 1353 40594 76375
rect 40814 1353 40924 76375
rect 41144 1353 48274 76375
rect 48494 1353 48604 76375
rect 48824 1353 51058 76375
<< metal5 >>
rect -418 76978 52386 77138
rect -88 76648 52056 76808
rect -418 73509 52386 73669
rect -418 69599 52386 69759
rect -418 65689 52386 65849
rect -418 61779 52386 61939
rect -418 57869 52386 58029
rect -418 53959 52386 54119
rect -418 50049 52386 50209
rect -418 46139 52386 46299
rect -418 42229 52386 42389
rect -418 38319 52386 38479
rect -418 34409 52386 34569
rect -418 30499 52386 30659
rect -418 26589 52386 26749
rect -418 22679 52386 22839
rect -418 18769 52386 18929
rect -418 14859 52386 15019
rect -418 10949 52386 11109
rect -418 7039 52386 7199
rect -418 3129 52386 3289
rect -88 808 52056 968
rect -418 478 52386 638
<< obsm5 >>
rect 566 73719 51066 75930
rect 566 69809 51066 73459
rect 566 65899 51066 69549
rect 566 61989 51066 65639
rect 566 58079 51066 61729
rect 566 54169 51066 57819
rect 566 50259 51066 53909
rect 566 46349 51066 49999
rect 566 42439 51066 46089
rect 566 38529 51066 42179
rect 566 34619 51066 38269
rect 566 30709 51066 34359
rect 566 26799 51066 30449
rect 566 22889 51066 26539
rect 566 18979 51066 22629
rect 566 15069 51066 18719
rect 566 11159 51066 14809
rect 566 7249 51066 10899
rect 566 3339 51066 6989
rect 566 1686 51066 3079
<< labels >>
rlabel metal4 s -88 808 72 76808 4 VDD
port 1 nsew power bidirectional
rlabel metal5 s -88 808 52056 968 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -88 76648 52056 76808 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 51896 808 52056 76808 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 2224 478 2384 77138 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 9904 478 10064 77138 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 17584 478 17744 77138 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 25264 478 25424 77138 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 32944 478 33104 77138 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 40624 478 40784 77138 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 48304 478 48464 77138 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 3129 52386 3289 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 10949 52386 11109 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 18769 52386 18929 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 26589 52386 26749 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 34409 52386 34569 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 42229 52386 42389 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 50049 52386 50209 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 57869 52386 58029 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 65689 52386 65849 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s -418 73509 52386 73669 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s -418 478 -258 77138 4 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 478 52386 638 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 76978 52386 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 52226 478 52386 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 2554 478 2714 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 10234 478 10394 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 17914 478 18074 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 25594 478 25754 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 33274 478 33434 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 40954 478 41114 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 48634 478 48794 77138 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 7039 52386 7199 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 14859 52386 15019 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 22679 52386 22839 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 30499 52386 30659 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 38319 52386 38479 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 46139 52386 46299 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 53959 52386 54119 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 61779 52386 61939 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s -418 69599 52386 69759 6 VSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 2296 400 2352 6 debug_in
port 3 nsew signal output
rlabel metal3 s 0 2912 400 2968 6 debug_mode
port 4 nsew signal input
rlabel metal3 s 0 3528 400 3584 6 debug_oeb
port 5 nsew signal input
rlabel metal3 s 0 4144 400 4200 6 debug_out
port 6 nsew signal input
rlabel metal3 s 0 5376 400 5432 6 irq[0]
port 7 nsew signal output
rlabel metal3 s 0 5992 400 6048 6 irq[1]
port 8 nsew signal output
rlabel metal3 s 0 6608 400 6664 6 irq[2]
port 9 nsew signal output
rlabel metal2 s 32928 0 32984 400 6 mask_rev_in[0]
port 10 nsew signal input
rlabel metal2 s 38528 0 38584 400 6 mask_rev_in[10]
port 11 nsew signal input
rlabel metal2 s 39088 0 39144 400 6 mask_rev_in[11]
port 12 nsew signal input
rlabel metal2 s 39648 0 39704 400 6 mask_rev_in[12]
port 13 nsew signal input
rlabel metal2 s 40208 0 40264 400 6 mask_rev_in[13]
port 14 nsew signal input
rlabel metal2 s 40768 0 40824 400 6 mask_rev_in[14]
port 15 nsew signal input
rlabel metal2 s 41328 0 41384 400 6 mask_rev_in[15]
port 16 nsew signal input
rlabel metal2 s 41888 0 41944 400 6 mask_rev_in[16]
port 17 nsew signal input
rlabel metal2 s 42448 0 42504 400 6 mask_rev_in[17]
port 18 nsew signal input
rlabel metal2 s 43008 0 43064 400 6 mask_rev_in[18]
port 19 nsew signal input
rlabel metal2 s 43568 0 43624 400 6 mask_rev_in[19]
port 20 nsew signal input
rlabel metal2 s 33488 0 33544 400 6 mask_rev_in[1]
port 21 nsew signal input
rlabel metal2 s 44128 0 44184 400 6 mask_rev_in[20]
port 22 nsew signal input
rlabel metal2 s 44688 0 44744 400 6 mask_rev_in[21]
port 23 nsew signal input
rlabel metal2 s 45248 0 45304 400 6 mask_rev_in[22]
port 24 nsew signal input
rlabel metal2 s 45808 0 45864 400 6 mask_rev_in[23]
port 25 nsew signal input
rlabel metal2 s 46368 0 46424 400 6 mask_rev_in[24]
port 26 nsew signal input
rlabel metal2 s 46928 0 46984 400 6 mask_rev_in[25]
port 27 nsew signal input
rlabel metal2 s 47488 0 47544 400 6 mask_rev_in[26]
port 28 nsew signal input
rlabel metal2 s 48048 0 48104 400 6 mask_rev_in[27]
port 29 nsew signal input
rlabel metal2 s 48608 0 48664 400 6 mask_rev_in[28]
port 30 nsew signal input
rlabel metal2 s 49168 0 49224 400 6 mask_rev_in[29]
port 31 nsew signal input
rlabel metal2 s 34048 0 34104 400 6 mask_rev_in[2]
port 32 nsew signal input
rlabel metal2 s 49728 0 49784 400 6 mask_rev_in[30]
port 33 nsew signal input
rlabel metal2 s 50288 0 50344 400 6 mask_rev_in[31]
port 34 nsew signal input
rlabel metal2 s 34608 0 34664 400 6 mask_rev_in[3]
port 35 nsew signal input
rlabel metal2 s 35168 0 35224 400 6 mask_rev_in[4]
port 36 nsew signal input
rlabel metal2 s 35728 0 35784 400 6 mask_rev_in[5]
port 37 nsew signal input
rlabel metal2 s 36288 0 36344 400 6 mask_rev_in[6]
port 38 nsew signal input
rlabel metal2 s 36848 0 36904 400 6 mask_rev_in[7]
port 39 nsew signal input
rlabel metal2 s 37408 0 37464 400 6 mask_rev_in[8]
port 40 nsew signal input
rlabel metal2 s 37968 0 38024 400 6 mask_rev_in[9]
port 41 nsew signal input
rlabel metal3 s 51600 7224 52000 7280 6 mgmt_gpio_in[0]
port 42 nsew signal input
rlabel metal3 s 51600 42504 52000 42560 6 mgmt_gpio_in[10]
port 43 nsew signal input
rlabel metal3 s 51600 46032 52000 46088 6 mgmt_gpio_in[11]
port 44 nsew signal input
rlabel metal3 s 51600 49560 52000 49616 6 mgmt_gpio_in[12]
port 45 nsew signal input
rlabel metal3 s 51600 53088 52000 53144 6 mgmt_gpio_in[13]
port 46 nsew signal input
rlabel metal3 s 51600 56616 52000 56672 6 mgmt_gpio_in[14]
port 47 nsew signal input
rlabel metal3 s 51600 60144 52000 60200 6 mgmt_gpio_in[15]
port 48 nsew signal input
rlabel metal3 s 51600 63672 52000 63728 6 mgmt_gpio_in[16]
port 49 nsew signal input
rlabel metal3 s 51600 67200 52000 67256 6 mgmt_gpio_in[17]
port 50 nsew signal input
rlabel metal3 s 51600 70728 52000 70784 6 mgmt_gpio_in[18]
port 51 nsew signal input
rlabel metal3 s 51600 74256 52000 74312 6 mgmt_gpio_in[19]
port 52 nsew signal input
rlabel metal3 s 51600 10752 52000 10808 6 mgmt_gpio_in[1]
port 53 nsew signal input
rlabel metal3 s 0 42952 400 43008 6 mgmt_gpio_in[20]
port 54 nsew signal input
rlabel metal3 s 0 44800 400 44856 6 mgmt_gpio_in[21]
port 55 nsew signal input
rlabel metal3 s 0 46648 400 46704 6 mgmt_gpio_in[22]
port 56 nsew signal input
rlabel metal3 s 0 48496 400 48552 6 mgmt_gpio_in[23]
port 57 nsew signal input
rlabel metal3 s 0 50344 400 50400 6 mgmt_gpio_in[24]
port 58 nsew signal input
rlabel metal3 s 0 52192 400 52248 6 mgmt_gpio_in[25]
port 59 nsew signal input
rlabel metal3 s 0 54040 400 54096 6 mgmt_gpio_in[26]
port 60 nsew signal input
rlabel metal3 s 0 55888 400 55944 6 mgmt_gpio_in[27]
port 61 nsew signal input
rlabel metal3 s 0 57736 400 57792 6 mgmt_gpio_in[28]
port 62 nsew signal input
rlabel metal3 s 0 59584 400 59640 6 mgmt_gpio_in[29]
port 63 nsew signal input
rlabel metal3 s 51600 14280 52000 14336 6 mgmt_gpio_in[2]
port 64 nsew signal input
rlabel metal3 s 0 61432 400 61488 6 mgmt_gpio_in[30]
port 65 nsew signal input
rlabel metal3 s 0 63280 400 63336 6 mgmt_gpio_in[31]
port 66 nsew signal input
rlabel metal3 s 0 65128 400 65184 6 mgmt_gpio_in[32]
port 67 nsew signal input
rlabel metal3 s 0 66976 400 67032 6 mgmt_gpio_in[33]
port 68 nsew signal input
rlabel metal3 s 0 68824 400 68880 6 mgmt_gpio_in[34]
port 69 nsew signal input
rlabel metal3 s 0 70672 400 70728 6 mgmt_gpio_in[35]
port 70 nsew signal input
rlabel metal3 s 0 72520 400 72576 6 mgmt_gpio_in[36]
port 71 nsew signal input
rlabel metal3 s 0 74368 400 74424 6 mgmt_gpio_in[37]
port 72 nsew signal input
rlabel metal3 s 51600 17808 52000 17864 6 mgmt_gpio_in[3]
port 73 nsew signal input
rlabel metal3 s 51600 21336 52000 21392 6 mgmt_gpio_in[4]
port 74 nsew signal input
rlabel metal3 s 51600 24864 52000 24920 6 mgmt_gpio_in[5]
port 75 nsew signal input
rlabel metal3 s 51600 28392 52000 28448 6 mgmt_gpio_in[6]
port 76 nsew signal input
rlabel metal3 s 51600 31920 52000 31976 6 mgmt_gpio_in[7]
port 77 nsew signal input
rlabel metal3 s 51600 35448 52000 35504 6 mgmt_gpio_in[8]
port 78 nsew signal input
rlabel metal3 s 51600 38976 52000 39032 6 mgmt_gpio_in[9]
port 79 nsew signal input
rlabel metal3 s 51600 8400 52000 8456 6 mgmt_gpio_oeb[0]
port 80 nsew signal output
rlabel metal3 s 51600 43680 52000 43736 6 mgmt_gpio_oeb[10]
port 81 nsew signal output
rlabel metal3 s 51600 47208 52000 47264 6 mgmt_gpio_oeb[11]
port 82 nsew signal output
rlabel metal3 s 51600 50736 52000 50792 6 mgmt_gpio_oeb[12]
port 83 nsew signal output
rlabel metal3 s 51600 54264 52000 54320 6 mgmt_gpio_oeb[13]
port 84 nsew signal output
rlabel metal3 s 51600 57792 52000 57848 6 mgmt_gpio_oeb[14]
port 85 nsew signal output
rlabel metal3 s 51600 61320 52000 61376 6 mgmt_gpio_oeb[15]
port 86 nsew signal output
rlabel metal3 s 51600 64848 52000 64904 6 mgmt_gpio_oeb[16]
port 87 nsew signal output
rlabel metal3 s 51600 68376 52000 68432 6 mgmt_gpio_oeb[17]
port 88 nsew signal output
rlabel metal3 s 51600 71904 52000 71960 6 mgmt_gpio_oeb[18]
port 89 nsew signal output
rlabel metal3 s 51600 75432 52000 75488 6 mgmt_gpio_oeb[19]
port 90 nsew signal output
rlabel metal3 s 51600 11928 52000 11984 6 mgmt_gpio_oeb[1]
port 91 nsew signal output
rlabel metal3 s 0 43568 400 43624 6 mgmt_gpio_oeb[20]
port 92 nsew signal output
rlabel metal3 s 0 45416 400 45472 6 mgmt_gpio_oeb[21]
port 93 nsew signal output
rlabel metal3 s 0 47264 400 47320 6 mgmt_gpio_oeb[22]
port 94 nsew signal output
rlabel metal3 s 0 49112 400 49168 6 mgmt_gpio_oeb[23]
port 95 nsew signal output
rlabel metal3 s 0 50960 400 51016 6 mgmt_gpio_oeb[24]
port 96 nsew signal output
rlabel metal3 s 0 52808 400 52864 6 mgmt_gpio_oeb[25]
port 97 nsew signal output
rlabel metal3 s 0 54656 400 54712 6 mgmt_gpio_oeb[26]
port 98 nsew signal output
rlabel metal3 s 0 56504 400 56560 6 mgmt_gpio_oeb[27]
port 99 nsew signal output
rlabel metal3 s 0 58352 400 58408 6 mgmt_gpio_oeb[28]
port 100 nsew signal output
rlabel metal3 s 0 60200 400 60256 6 mgmt_gpio_oeb[29]
port 101 nsew signal output
rlabel metal3 s 51600 15456 52000 15512 6 mgmt_gpio_oeb[2]
port 102 nsew signal output
rlabel metal3 s 0 62048 400 62104 6 mgmt_gpio_oeb[30]
port 103 nsew signal output
rlabel metal3 s 0 63896 400 63952 6 mgmt_gpio_oeb[31]
port 104 nsew signal output
rlabel metal3 s 0 65744 400 65800 6 mgmt_gpio_oeb[32]
port 105 nsew signal output
rlabel metal3 s 0 67592 400 67648 6 mgmt_gpio_oeb[33]
port 106 nsew signal output
rlabel metal3 s 0 69440 400 69496 6 mgmt_gpio_oeb[34]
port 107 nsew signal output
rlabel metal3 s 0 71288 400 71344 6 mgmt_gpio_oeb[35]
port 108 nsew signal output
rlabel metal3 s 0 73136 400 73192 6 mgmt_gpio_oeb[36]
port 109 nsew signal output
rlabel metal3 s 0 74984 400 75040 6 mgmt_gpio_oeb[37]
port 110 nsew signal output
rlabel metal3 s 51600 18984 52000 19040 6 mgmt_gpio_oeb[3]
port 111 nsew signal output
rlabel metal3 s 51600 22512 52000 22568 6 mgmt_gpio_oeb[4]
port 112 nsew signal output
rlabel metal3 s 51600 26040 52000 26096 6 mgmt_gpio_oeb[5]
port 113 nsew signal output
rlabel metal3 s 51600 29568 52000 29624 6 mgmt_gpio_oeb[6]
port 114 nsew signal output
rlabel metal3 s 51600 33096 52000 33152 6 mgmt_gpio_oeb[7]
port 115 nsew signal output
rlabel metal3 s 51600 36624 52000 36680 6 mgmt_gpio_oeb[8]
port 116 nsew signal output
rlabel metal3 s 51600 40152 52000 40208 6 mgmt_gpio_oeb[9]
port 117 nsew signal output
rlabel metal3 s 51600 9576 52000 9632 6 mgmt_gpio_out[0]
port 118 nsew signal output
rlabel metal3 s 51600 44856 52000 44912 6 mgmt_gpio_out[10]
port 119 nsew signal output
rlabel metal3 s 51600 48384 52000 48440 6 mgmt_gpio_out[11]
port 120 nsew signal output
rlabel metal3 s 51600 51912 52000 51968 6 mgmt_gpio_out[12]
port 121 nsew signal output
rlabel metal3 s 51600 55440 52000 55496 6 mgmt_gpio_out[13]
port 122 nsew signal output
rlabel metal3 s 51600 58968 52000 59024 6 mgmt_gpio_out[14]
port 123 nsew signal output
rlabel metal3 s 51600 62496 52000 62552 6 mgmt_gpio_out[15]
port 124 nsew signal output
rlabel metal3 s 51600 66024 52000 66080 6 mgmt_gpio_out[16]
port 125 nsew signal output
rlabel metal3 s 51600 69552 52000 69608 6 mgmt_gpio_out[17]
port 126 nsew signal output
rlabel metal3 s 51600 73080 52000 73136 6 mgmt_gpio_out[18]
port 127 nsew signal output
rlabel metal3 s 51600 76608 52000 76664 6 mgmt_gpio_out[19]
port 128 nsew signal output
rlabel metal3 s 51600 13104 52000 13160 6 mgmt_gpio_out[1]
port 129 nsew signal output
rlabel metal3 s 0 44184 400 44240 6 mgmt_gpio_out[20]
port 130 nsew signal output
rlabel metal3 s 0 46032 400 46088 6 mgmt_gpio_out[21]
port 131 nsew signal output
rlabel metal3 s 0 47880 400 47936 6 mgmt_gpio_out[22]
port 132 nsew signal output
rlabel metal3 s 0 49728 400 49784 6 mgmt_gpio_out[23]
port 133 nsew signal output
rlabel metal3 s 0 51576 400 51632 6 mgmt_gpio_out[24]
port 134 nsew signal output
rlabel metal3 s 0 53424 400 53480 6 mgmt_gpio_out[25]
port 135 nsew signal output
rlabel metal3 s 0 55272 400 55328 6 mgmt_gpio_out[26]
port 136 nsew signal output
rlabel metal3 s 0 57120 400 57176 6 mgmt_gpio_out[27]
port 137 nsew signal output
rlabel metal3 s 0 58968 400 59024 6 mgmt_gpio_out[28]
port 138 nsew signal output
rlabel metal3 s 0 60816 400 60872 6 mgmt_gpio_out[29]
port 139 nsew signal output
rlabel metal3 s 51600 16632 52000 16688 6 mgmt_gpio_out[2]
port 140 nsew signal output
rlabel metal3 s 0 62664 400 62720 6 mgmt_gpio_out[30]
port 141 nsew signal output
rlabel metal3 s 0 64512 400 64568 6 mgmt_gpio_out[31]
port 142 nsew signal output
rlabel metal3 s 0 66360 400 66416 6 mgmt_gpio_out[32]
port 143 nsew signal output
rlabel metal3 s 0 68208 400 68264 6 mgmt_gpio_out[33]
port 144 nsew signal output
rlabel metal3 s 0 70056 400 70112 6 mgmt_gpio_out[34]
port 145 nsew signal output
rlabel metal3 s 0 71904 400 71960 6 mgmt_gpio_out[35]
port 146 nsew signal output
rlabel metal3 s 0 73752 400 73808 6 mgmt_gpio_out[36]
port 147 nsew signal output
rlabel metal3 s 0 75600 400 75656 6 mgmt_gpio_out[37]
port 148 nsew signal output
rlabel metal3 s 51600 20160 52000 20216 6 mgmt_gpio_out[3]
port 149 nsew signal output
rlabel metal3 s 51600 23688 52000 23744 6 mgmt_gpio_out[4]
port 150 nsew signal output
rlabel metal3 s 51600 27216 52000 27272 6 mgmt_gpio_out[5]
port 151 nsew signal output
rlabel metal3 s 51600 30744 52000 30800 6 mgmt_gpio_out[6]
port 152 nsew signal output
rlabel metal3 s 51600 34272 52000 34328 6 mgmt_gpio_out[7]
port 153 nsew signal output
rlabel metal3 s 51600 37800 52000 37856 6 mgmt_gpio_out[8]
port 154 nsew signal output
rlabel metal3 s 51600 41328 52000 41384 6 mgmt_gpio_out[9]
port 155 nsew signal output
rlabel metal2 s 1568 0 1624 400 6 pad_flash_clk
port 156 nsew signal output
rlabel metal2 s 2128 0 2184 400 6 pad_flash_clk_oe
port 157 nsew signal output
rlabel metal2 s 2688 0 2744 400 6 pad_flash_csb
port 158 nsew signal output
rlabel metal2 s 3248 0 3304 400 6 pad_flash_csb_oe
port 159 nsew signal output
rlabel metal2 s 3808 0 3864 400 6 pad_flash_io0_di
port 160 nsew signal input
rlabel metal2 s 4368 0 4424 400 6 pad_flash_io0_do
port 161 nsew signal output
rlabel metal2 s 4928 0 4984 400 6 pad_flash_io0_ie
port 162 nsew signal output
rlabel metal2 s 5488 0 5544 400 6 pad_flash_io0_oe
port 163 nsew signal output
rlabel metal2 s 6048 0 6104 400 6 pad_flash_io1_di
port 164 nsew signal input
rlabel metal2 s 6608 0 6664 400 6 pad_flash_io1_do
port 165 nsew signal output
rlabel metal2 s 7168 0 7224 400 6 pad_flash_io1_ie
port 166 nsew signal output
rlabel metal2 s 7728 0 7784 400 6 pad_flash_io1_oe
port 167 nsew signal output
rlabel metal2 s 15008 0 15064 400 6 pll90_sel[0]
port 168 nsew signal output
rlabel metal2 s 15568 0 15624 400 6 pll90_sel[1]
port 169 nsew signal output
rlabel metal2 s 16128 0 16184 400 6 pll90_sel[2]
port 170 nsew signal output
rlabel metal2 s 31248 0 31304 400 6 pll_bypass
port 171 nsew signal output
rlabel metal2 s 9968 0 10024 400 6 pll_dco_ena
port 172 nsew signal output
rlabel metal2 s 10528 0 10584 400 6 pll_div[0]
port 173 nsew signal output
rlabel metal2 s 11088 0 11144 400 6 pll_div[1]
port 174 nsew signal output
rlabel metal2 s 11648 0 11704 400 6 pll_div[2]
port 175 nsew signal output
rlabel metal2 s 12208 0 12264 400 6 pll_div[3]
port 176 nsew signal output
rlabel metal2 s 12768 0 12824 400 6 pll_div[4]
port 177 nsew signal output
rlabel metal2 s 9408 0 9464 400 6 pll_ena
port 178 nsew signal output
rlabel metal2 s 13328 0 13384 400 6 pll_sel[0]
port 179 nsew signal output
rlabel metal2 s 13888 0 13944 400 6 pll_sel[1]
port 180 nsew signal output
rlabel metal2 s 14448 0 14504 400 6 pll_sel[2]
port 181 nsew signal output
rlabel metal2 s 16688 0 16744 400 6 pll_trim[0]
port 182 nsew signal output
rlabel metal2 s 22288 0 22344 400 6 pll_trim[10]
port 183 nsew signal output
rlabel metal2 s 22848 0 22904 400 6 pll_trim[11]
port 184 nsew signal output
rlabel metal2 s 23408 0 23464 400 6 pll_trim[12]
port 185 nsew signal output
rlabel metal2 s 23968 0 24024 400 6 pll_trim[13]
port 186 nsew signal output
rlabel metal2 s 24528 0 24584 400 6 pll_trim[14]
port 187 nsew signal output
rlabel metal2 s 25088 0 25144 400 6 pll_trim[15]
port 188 nsew signal output
rlabel metal2 s 25648 0 25704 400 6 pll_trim[16]
port 189 nsew signal output
rlabel metal2 s 26208 0 26264 400 6 pll_trim[17]
port 190 nsew signal output
rlabel metal2 s 26768 0 26824 400 6 pll_trim[18]
port 191 nsew signal output
rlabel metal2 s 27328 0 27384 400 6 pll_trim[19]
port 192 nsew signal output
rlabel metal2 s 17248 0 17304 400 6 pll_trim[1]
port 193 nsew signal output
rlabel metal2 s 27888 0 27944 400 6 pll_trim[20]
port 194 nsew signal output
rlabel metal2 s 28448 0 28504 400 6 pll_trim[21]
port 195 nsew signal output
rlabel metal2 s 29008 0 29064 400 6 pll_trim[22]
port 196 nsew signal output
rlabel metal2 s 29568 0 29624 400 6 pll_trim[23]
port 197 nsew signal output
rlabel metal2 s 30128 0 30184 400 6 pll_trim[24]
port 198 nsew signal output
rlabel metal2 s 30688 0 30744 400 6 pll_trim[25]
port 199 nsew signal output
rlabel metal2 s 17808 0 17864 400 6 pll_trim[2]
port 200 nsew signal output
rlabel metal2 s 18368 0 18424 400 6 pll_trim[3]
port 201 nsew signal output
rlabel metal2 s 18928 0 18984 400 6 pll_trim[4]
port 202 nsew signal output
rlabel metal2 s 19488 0 19544 400 6 pll_trim[5]
port 203 nsew signal output
rlabel metal2 s 20048 0 20104 400 6 pll_trim[6]
port 204 nsew signal output
rlabel metal2 s 20608 0 20664 400 6 pll_trim[7]
port 205 nsew signal output
rlabel metal2 s 21168 0 21224 400 6 pll_trim[8]
port 206 nsew signal output
rlabel metal2 s 21728 0 21784 400 6 pll_trim[9]
port 207 nsew signal output
rlabel metal2 s 8288 0 8344 400 6 porb
port 208 nsew signal input
rlabel metal2 s 50848 0 50904 400 6 pwr_ctrl_out
port 209 nsew signal output
rlabel metal3 s 0 11536 400 11592 6 qspi_enabled
port 210 nsew signal input
rlabel metal2 s 8848 0 8904 400 6 reset
port 211 nsew signal output
rlabel metal3 s 0 10920 400 10976 6 ser_rx
port 212 nsew signal output
rlabel metal3 s 0 10304 400 10360 6 ser_tx
port 213 nsew signal input
rlabel metal3 s 51600 1344 52000 1400 6 serial_clock
port 214 nsew signal output
rlabel metal3 s 51600 4872 52000 4928 6 serial_data_1
port 215 nsew signal output
rlabel metal3 s 51600 6048 52000 6104 6 serial_data_2
port 216 nsew signal output
rlabel metal3 s 51600 3696 52000 3752 6 serial_load
port 217 nsew signal output
rlabel metal3 s 51600 2520 52000 2576 6 serial_resetn
port 218 nsew signal output
rlabel metal3 s 0 9072 400 9128 6 spi_csb
port 219 nsew signal input
rlabel metal3 s 0 12768 400 12824 6 spi_enabled
port 220 nsew signal input
rlabel metal3 s 0 8456 400 8512 6 spi_sck
port 221 nsew signal input
rlabel metal3 s 0 9688 400 9744 6 spi_sdi
port 222 nsew signal output
rlabel metal3 s 0 7840 400 7896 6 spi_sdo
port 223 nsew signal input
rlabel metal3 s 0 7224 400 7280 6 spi_sdoenb
port 224 nsew signal input
rlabel metal3 s 0 34328 400 34384 6 spimemio_flash_clk
port 225 nsew signal input
rlabel metal3 s 0 34944 400 35000 6 spimemio_flash_csb
port 226 nsew signal input
rlabel metal3 s 0 35560 400 35616 6 spimemio_flash_io0_di
port 227 nsew signal output
rlabel metal3 s 0 36176 400 36232 6 spimemio_flash_io0_do
port 228 nsew signal input
rlabel metal3 s 0 36792 400 36848 6 spimemio_flash_io0_oeb
port 229 nsew signal input
rlabel metal3 s 0 37408 400 37464 6 spimemio_flash_io1_di
port 230 nsew signal output
rlabel metal3 s 0 38024 400 38080 6 spimemio_flash_io1_do
port 231 nsew signal input
rlabel metal3 s 0 38640 400 38696 6 spimemio_flash_io1_oeb
port 232 nsew signal input
rlabel metal3 s 0 39256 400 39312 6 spimemio_flash_io2_di
port 233 nsew signal output
rlabel metal3 s 0 39872 400 39928 6 spimemio_flash_io2_do
port 234 nsew signal input
rlabel metal3 s 0 40488 400 40544 6 spimemio_flash_io2_oeb
port 235 nsew signal input
rlabel metal3 s 0 41104 400 41160 6 spimemio_flash_io3_di
port 236 nsew signal output
rlabel metal3 s 0 41720 400 41776 6 spimemio_flash_io3_do
port 237 nsew signal input
rlabel metal3 s 0 42336 400 42392 6 spimemio_flash_io3_oeb
port 238 nsew signal input
rlabel metal3 s 0 4760 400 4816 6 trap
port 239 nsew signal input
rlabel metal3 s 0 12152 400 12208 6 uart_enabled
port 240 nsew signal input
rlabel metal2 s 1008 0 1064 400 6 user_clock
port 241 nsew signal input
rlabel metal3 s 0 13384 400 13440 6 wb_ack_o
port 242 nsew signal output
rlabel metal2 s 840 77600 896 78000 6 wb_adr_i[0]
port 243 nsew signal input
rlabel metal2 s 8120 77600 8176 78000 6 wb_adr_i[10]
port 244 nsew signal input
rlabel metal2 s 8848 77600 8904 78000 6 wb_adr_i[11]
port 245 nsew signal input
rlabel metal2 s 9576 77600 9632 78000 6 wb_adr_i[12]
port 246 nsew signal input
rlabel metal2 s 10304 77600 10360 78000 6 wb_adr_i[13]
port 247 nsew signal input
rlabel metal2 s 11032 77600 11088 78000 6 wb_adr_i[14]
port 248 nsew signal input
rlabel metal2 s 11760 77600 11816 78000 6 wb_adr_i[15]
port 249 nsew signal input
rlabel metal2 s 12488 77600 12544 78000 6 wb_adr_i[16]
port 250 nsew signal input
rlabel metal2 s 13216 77600 13272 78000 6 wb_adr_i[17]
port 251 nsew signal input
rlabel metal2 s 13944 77600 14000 78000 6 wb_adr_i[18]
port 252 nsew signal input
rlabel metal2 s 14672 77600 14728 78000 6 wb_adr_i[19]
port 253 nsew signal input
rlabel metal2 s 1568 77600 1624 78000 6 wb_adr_i[1]
port 254 nsew signal input
rlabel metal2 s 15400 77600 15456 78000 6 wb_adr_i[20]
port 255 nsew signal input
rlabel metal2 s 16128 77600 16184 78000 6 wb_adr_i[21]
port 256 nsew signal input
rlabel metal2 s 16856 77600 16912 78000 6 wb_adr_i[22]
port 257 nsew signal input
rlabel metal2 s 17584 77600 17640 78000 6 wb_adr_i[23]
port 258 nsew signal input
rlabel metal2 s 18312 77600 18368 78000 6 wb_adr_i[24]
port 259 nsew signal input
rlabel metal2 s 19040 77600 19096 78000 6 wb_adr_i[25]
port 260 nsew signal input
rlabel metal2 s 19768 77600 19824 78000 6 wb_adr_i[26]
port 261 nsew signal input
rlabel metal2 s 20496 77600 20552 78000 6 wb_adr_i[27]
port 262 nsew signal input
rlabel metal2 s 21224 77600 21280 78000 6 wb_adr_i[28]
port 263 nsew signal input
rlabel metal2 s 21952 77600 22008 78000 6 wb_adr_i[29]
port 264 nsew signal input
rlabel metal2 s 2296 77600 2352 78000 6 wb_adr_i[2]
port 265 nsew signal input
rlabel metal2 s 22680 77600 22736 78000 6 wb_adr_i[30]
port 266 nsew signal input
rlabel metal2 s 23408 77600 23464 78000 6 wb_adr_i[31]
port 267 nsew signal input
rlabel metal2 s 3024 77600 3080 78000 6 wb_adr_i[3]
port 268 nsew signal input
rlabel metal2 s 3752 77600 3808 78000 6 wb_adr_i[4]
port 269 nsew signal input
rlabel metal2 s 4480 77600 4536 78000 6 wb_adr_i[5]
port 270 nsew signal input
rlabel metal2 s 5208 77600 5264 78000 6 wb_adr_i[6]
port 271 nsew signal input
rlabel metal2 s 5936 77600 5992 78000 6 wb_adr_i[7]
port 272 nsew signal input
rlabel metal2 s 6664 77600 6720 78000 6 wb_adr_i[8]
port 273 nsew signal input
rlabel metal2 s 7392 77600 7448 78000 6 wb_adr_i[9]
port 274 nsew signal input
rlabel metal2 s 31808 0 31864 400 6 wb_clk_i
port 275 nsew signal input
rlabel metal2 s 51072 77600 51128 78000 6 wb_cyc_i
port 276 nsew signal input
rlabel metal2 s 24136 77600 24192 78000 6 wb_dat_i[0]
port 277 nsew signal input
rlabel metal2 s 31416 77600 31472 78000 6 wb_dat_i[10]
port 278 nsew signal input
rlabel metal2 s 32144 77600 32200 78000 6 wb_dat_i[11]
port 279 nsew signal input
rlabel metal2 s 32872 77600 32928 78000 6 wb_dat_i[12]
port 280 nsew signal input
rlabel metal2 s 33600 77600 33656 78000 6 wb_dat_i[13]
port 281 nsew signal input
rlabel metal2 s 34328 77600 34384 78000 6 wb_dat_i[14]
port 282 nsew signal input
rlabel metal2 s 35056 77600 35112 78000 6 wb_dat_i[15]
port 283 nsew signal input
rlabel metal2 s 35784 77600 35840 78000 6 wb_dat_i[16]
port 284 nsew signal input
rlabel metal2 s 36512 77600 36568 78000 6 wb_dat_i[17]
port 285 nsew signal input
rlabel metal2 s 37240 77600 37296 78000 6 wb_dat_i[18]
port 286 nsew signal input
rlabel metal2 s 37968 77600 38024 78000 6 wb_dat_i[19]
port 287 nsew signal input
rlabel metal2 s 24864 77600 24920 78000 6 wb_dat_i[1]
port 288 nsew signal input
rlabel metal2 s 38696 77600 38752 78000 6 wb_dat_i[20]
port 289 nsew signal input
rlabel metal2 s 39424 77600 39480 78000 6 wb_dat_i[21]
port 290 nsew signal input
rlabel metal2 s 40152 77600 40208 78000 6 wb_dat_i[22]
port 291 nsew signal input
rlabel metal2 s 40880 77600 40936 78000 6 wb_dat_i[23]
port 292 nsew signal input
rlabel metal2 s 41608 77600 41664 78000 6 wb_dat_i[24]
port 293 nsew signal input
rlabel metal2 s 42336 77600 42392 78000 6 wb_dat_i[25]
port 294 nsew signal input
rlabel metal2 s 43064 77600 43120 78000 6 wb_dat_i[26]
port 295 nsew signal input
rlabel metal2 s 43792 77600 43848 78000 6 wb_dat_i[27]
port 296 nsew signal input
rlabel metal2 s 44520 77600 44576 78000 6 wb_dat_i[28]
port 297 nsew signal input
rlabel metal2 s 45248 77600 45304 78000 6 wb_dat_i[29]
port 298 nsew signal input
rlabel metal2 s 25592 77600 25648 78000 6 wb_dat_i[2]
port 299 nsew signal input
rlabel metal2 s 45976 77600 46032 78000 6 wb_dat_i[30]
port 300 nsew signal input
rlabel metal2 s 46704 77600 46760 78000 6 wb_dat_i[31]
port 301 nsew signal input
rlabel metal2 s 26320 77600 26376 78000 6 wb_dat_i[3]
port 302 nsew signal input
rlabel metal2 s 27048 77600 27104 78000 6 wb_dat_i[4]
port 303 nsew signal input
rlabel metal2 s 27776 77600 27832 78000 6 wb_dat_i[5]
port 304 nsew signal input
rlabel metal2 s 28504 77600 28560 78000 6 wb_dat_i[6]
port 305 nsew signal input
rlabel metal2 s 29232 77600 29288 78000 6 wb_dat_i[7]
port 306 nsew signal input
rlabel metal2 s 29960 77600 30016 78000 6 wb_dat_i[8]
port 307 nsew signal input
rlabel metal2 s 30688 77600 30744 78000 6 wb_dat_i[9]
port 308 nsew signal input
rlabel metal3 s 0 14616 400 14672 6 wb_dat_o[0]
port 309 nsew signal output
rlabel metal3 s 0 20776 400 20832 6 wb_dat_o[10]
port 310 nsew signal output
rlabel metal3 s 0 21392 400 21448 6 wb_dat_o[11]
port 311 nsew signal output
rlabel metal3 s 0 22008 400 22064 6 wb_dat_o[12]
port 312 nsew signal output
rlabel metal3 s 0 22624 400 22680 6 wb_dat_o[13]
port 313 nsew signal output
rlabel metal3 s 0 23240 400 23296 6 wb_dat_o[14]
port 314 nsew signal output
rlabel metal3 s 0 23856 400 23912 6 wb_dat_o[15]
port 315 nsew signal output
rlabel metal3 s 0 24472 400 24528 6 wb_dat_o[16]
port 316 nsew signal output
rlabel metal3 s 0 25088 400 25144 6 wb_dat_o[17]
port 317 nsew signal output
rlabel metal3 s 0 25704 400 25760 6 wb_dat_o[18]
port 318 nsew signal output
rlabel metal3 s 0 26320 400 26376 6 wb_dat_o[19]
port 319 nsew signal output
rlabel metal3 s 0 15232 400 15288 6 wb_dat_o[1]
port 320 nsew signal output
rlabel metal3 s 0 26936 400 26992 6 wb_dat_o[20]
port 321 nsew signal output
rlabel metal3 s 0 27552 400 27608 6 wb_dat_o[21]
port 322 nsew signal output
rlabel metal3 s 0 28168 400 28224 6 wb_dat_o[22]
port 323 nsew signal output
rlabel metal3 s 0 28784 400 28840 6 wb_dat_o[23]
port 324 nsew signal output
rlabel metal3 s 0 29400 400 29456 6 wb_dat_o[24]
port 325 nsew signal output
rlabel metal3 s 0 30016 400 30072 6 wb_dat_o[25]
port 326 nsew signal output
rlabel metal3 s 0 30632 400 30688 6 wb_dat_o[26]
port 327 nsew signal output
rlabel metal3 s 0 31248 400 31304 6 wb_dat_o[27]
port 328 nsew signal output
rlabel metal3 s 0 31864 400 31920 6 wb_dat_o[28]
port 329 nsew signal output
rlabel metal3 s 0 32480 400 32536 6 wb_dat_o[29]
port 330 nsew signal output
rlabel metal3 s 0 15848 400 15904 6 wb_dat_o[2]
port 331 nsew signal output
rlabel metal3 s 0 33096 400 33152 6 wb_dat_o[30]
port 332 nsew signal output
rlabel metal3 s 0 33712 400 33768 6 wb_dat_o[31]
port 333 nsew signal output
rlabel metal3 s 0 16464 400 16520 6 wb_dat_o[3]
port 334 nsew signal output
rlabel metal3 s 0 17080 400 17136 6 wb_dat_o[4]
port 335 nsew signal output
rlabel metal3 s 0 17696 400 17752 6 wb_dat_o[5]
port 336 nsew signal output
rlabel metal3 s 0 18312 400 18368 6 wb_dat_o[6]
port 337 nsew signal output
rlabel metal3 s 0 18928 400 18984 6 wb_dat_o[7]
port 338 nsew signal output
rlabel metal3 s 0 19544 400 19600 6 wb_dat_o[8]
port 339 nsew signal output
rlabel metal3 s 0 20160 400 20216 6 wb_dat_o[9]
port 340 nsew signal output
rlabel metal2 s 32368 0 32424 400 6 wb_rstn_i
port 341 nsew signal input
rlabel metal2 s 47432 77600 47488 78000 6 wb_sel_i[0]
port 342 nsew signal input
rlabel metal2 s 48160 77600 48216 78000 6 wb_sel_i[1]
port 343 nsew signal input
rlabel metal2 s 48888 77600 48944 78000 6 wb_sel_i[2]
port 344 nsew signal input
rlabel metal2 s 49616 77600 49672 78000 6 wb_sel_i[3]
port 345 nsew signal input
rlabel metal3 s 0 14000 400 14056 6 wb_stb_i
port 346 nsew signal input
rlabel metal2 s 50344 77600 50400 78000 6 wb_we_i
port 347 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 52000 78000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12831154
string GDS_FILE /home/hosni/GF180/EF/caravel-gf180mcu/openlane/housekeeping/runs/RUN_2022.11.19_02.10.22/results/signoff/housekeeping.magic.gds
string GDS_START 633868
<< end >>

