magic
tech gf180mcuC
magscale 1 5
timestamp 1654634570
<< metal5 >>
rect 108 540 216 648
rect 0 432 324 540
rect 108 0 216 432
<< properties >>
string FIXED_BBOX 0 -216 432 756
<< end >>
