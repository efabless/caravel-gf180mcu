magic
tech gf180mcuC
magscale 1 10
timestamp 1654652987
<< fillblock >>
rect -429 -1786 18270 2667
rect -429 -6331 7951 -1786
use font_2D  font_2D_0 alpha
timestamp 1654634570
transform 1 0 4768 0 1 -1351
box 0 648 864 864
use font_4A  font_4A_0 alpha
timestamp 1654634570
transform 1 0 -158 0 1 -6007
box 0 0 648 1512
use font_4B  font_4B_0 alpha
timestamp 1654634570
transform 1 0 5905 0 1 -3592
box 0 0 648 1512
use font_6C  font_6C_0 alpha
timestamp 1654634570
transform 1 0 5138 0 1 776
box 0 0 216 1512
use font_6C  font_6C_1
timestamp 1654634570
transform 1 0 3478 0 1 -1341
box 0 0 216 1512
use font_6C  font_6C_2
timestamp 1654634570
transform 1 0 6691 0 1 -1356
box 0 0 216 1512
use font_6C  font_6C_3
timestamp 1654634570
transform 1 0 9723 0 1 -1366
box 0 0 216 1512
use font_6C  font_6C_4
timestamp 1654634570
transform 1 0 14500 0 1 782
box 0 0 216 1512
use font_6E  font_6E_0 alpha
timestamp 1654634570
transform 1 0 2528 0 1 -3583
box 0 0 648 1080
use font_6E  font_6E_1
timestamp 1654634570
transform 1 0 1564 0 1 -6016
box 0 0 648 1080
use font_6E  font_6E_2
timestamp 1654634570
transform 1 0 13176 0 1 -1348
box 0 0 648 1080
use font_6F  font_6F_0 alpha
timestamp 1654634570
transform 1 0 879 0 1 -1313
box 0 0 648 1080
use font_6F  font_6F_1
timestamp 1654634570
transform 1 0 1730 0 1 -1323
box 0 0 648 1080
use font_6F  font_6F_2
timestamp 1654634570
transform 1 0 -55 0 1 -3555
box 0 0 648 1080
use font_6F  font_6F_3
timestamp 1654634570
transform 1 0 7131 0 1 -1366
box 0 0 648 1080
use font_6F  font_6F_4
timestamp 1654634570
transform 1 0 11473 0 1 -1339
box 0 0 648 1080
use font_28  font_28_0 alpha
timestamp 1654634570
transform 1 0 8140 0 1 800
box 0 0 432 1512
use font_29  font_29_0 alpha
timestamp 1654634570
transform 1 0 9640 0 1 782
box 0 0 432 1512
use font_30  font_30_0 alpha
timestamp 1654634570
transform 1 0 4923 0 1 -5999
box 0 0 648 1512
use font_32  font_32_0 alpha
timestamp 1654634570
transform 1 0 4053 0 1 -6008
box 0 0 648 1512
use font_32  font_32_1
timestamp 1654634570
transform 1 0 5803 0 1 -6007
box 0 0 648 1512
use font_32  font_32_2
timestamp 1654634570
transform 1 0 6691 0 1 -5999
box 0 0 648 1512
use font_43  font_43_0 alpha
timestamp 1654634570
transform 1 0 -46 0 1 785
box 0 0 648 1512
use font_44  font_44_0 alpha
timestamp 1654634570
transform 1 0 5045 0 1 -3592
box 0 0 648 1512
use font_45  font_45_0 alpha
timestamp 1654634570
transform 1 0 11030 0 1 782
box 0 0 648 1512
use font_46  font_46_0 alpha
timestamp 1654634570
transform 1 0 6907 0 1 794
box 0 0 648 1512
use font_46  font_46_1
timestamp 1654634570
transform 1 0 10621 0 1 -1375
box 0 0 648 1512
use font_47  font_47_0 alpha
timestamp 1654634570
transform 1 0 6027 0 1 794
box 0 0 648 1512
use font_47  font_47_1
timestamp 1654634570
transform 1 0 39 0 1 -1330
box 0 0 648 1512
use font_47  font_47_2
timestamp 1654634570
transform 1 0 5831 0 1 -1330
box 0 0 648 1512
use font_50  font_50_0 alpha
timestamp 1654634570
transform 1 0 4184 0 1 -3574
box 0 0 648 1512
use font_61  font_61_0 alpha
timestamp 1654634570
transform 1 0 806 0 1 776
box 0 0 648 1080
use font_61  font_61_1
timestamp 1654634570
transform 1 0 2537 0 1 776
box 0 0 648 1080
use font_61  font_61_2
timestamp 1654634570
transform 1 0 8853 0 1 -1347
box 0 0 648 1080
use font_61  font_61_3
timestamp 1654634570
transform 1 0 12760 0 1 772
box 0 0 648 1080
use font_62  font_62_0 alpha
timestamp 1654634570
transform 1 0 7992 0 1 -1347
box 0 0 648 1512
use font_62  font_62_1
timestamp 1654634570
transform 1 0 13630 0 1 782
box 0 0 648 1512
use font_63  font_63_0 alpha
timestamp 1654634570
transform 1 0 8780 0 1 970
box 0 0 648 1080
use font_64  font_64_0 alpha
timestamp 1654634570
transform 1 0 14055 0 1 -1330
box 0 0 648 1512
use font_65  font_65_0 alpha
timestamp 1654634570
transform 1 0 4277 0 1 794
box 0 0 648 1080
use font_65  font_65_1
timestamp 1654634570
transform 1 0 3918 0 1 -1341
box 0 0 648 1080
use font_65  font_65_2
timestamp 1654634570
transform 1 0 16432 0 1 -1339
box 0 0 648 1080
use font_65  font_65_3
timestamp 1654634570
transform 1 0 1676 0 1 -3564
box 0 0 648 1080
use font_65  font_65_4
timestamp 1654634570
transform 1 0 2425 0 1 -6008
box 0 0 648 1080
use font_65  font_65_5
timestamp 1654634570
transform 1 0 14930 0 1 782
box 0 0 648 1080
use font_66  font_66_0 alpha
timestamp 1654634570
transform 1 0 11890 0 1 782
box 0 0 648 1512
use font_67  font_67_0 alpha
timestamp 1654634570
transform 1 0 2609 0 1 -1332
box 0 -432 648 1080
use font_69  font_69_0 alpha
timestamp 1654634570
transform 1 0 15777 0 1 -1330
box 0 0 432 1512
use font_70  font_70_0 alpha
timestamp 1654634570
transform 1 0 806 0 1 -3546
box 0 -432 648 1080
use font_72  font_72_0 alpha
timestamp 1654634570
transform 1 0 1667 0 1 776
box 0 0 648 1080
use font_72  font_72_1
timestamp 1654634570
transform 1 0 14916 0 1 -1339
box 0 0 648 1080
use font_73  font_73_0 alpha
timestamp 1654634570
transform 1 0 17302 0 1 -1330
box 0 0 648 1080
use font_73  font_73_1
timestamp 1654634570
transform 1 0 15800 0 1 790
box 0 0 648 1080
use font_73  font_73_2
timestamp 1654634570
transform 1 0 16660 0 1 790
box 0 0 648 1080
use font_75  font_75_0 alpha
timestamp 1654634570
transform 1 0 703 0 1 -6016
box 0 0 648 1080
use font_75  font_75_1
timestamp 1654634570
transform 1 0 12334 0 1 -1330
box 0 0 648 1080
use font_76  font_76_0 alpha
timestamp 1654634570
transform 1 0 3445 0 1 776
box 0 0 648 1080
<< end >>
