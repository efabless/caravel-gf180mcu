* Simple POR testbench

.include /usr/share/pdk/gf180mcuC/libs.ref/gf180mcu_pr/spice/design.hspice
.lib /usr/share/pdk/gf180mcuC/libs.ref/gf180mcu_pr/spice/sm141064.hspice typical
.lib /usr/share/pdk/gf180mcuC/libs.ref/gf180mcu_pr/spice/sm141064.hspice res_typical
.include simple_por.spice

V0 VDD 0 5
V1 In 0 PWL(0 0 100u 5 200u 5 300u 0)

X0 VDD 0 In Out schmitt_inverter

.control
tran 500n 350u
plot V(In) V(Out)
.endc
