magic
tech gf180mcuC
magscale 1 5
timestamp 1668623287
<< fillblock >>
rect 0 0 25330 6045
use alpha_0  alphaX_0 hexdigits
timestamp 1654634570
transform 1 0 22665 0 1 700
box 0 0 1944 4536
use alpha_0  alphaX_1
timestamp 1654634570
transform 1 0 19480 0 1 700
box 0 0 1944 4536
use alpha_0  alphaX_2
timestamp 1654634570
transform 1 0 16355 0 1 700
box 0 0 1944 4536
use alpha_0  alphaX_3
timestamp 1654634570
transform 1 0 13230 0 1 700
box 0 0 1944 4536
use alpha_0  alphaX_4
timestamp 1654634570
transform 1 0 10105 0 1 700
box 0 0 1944 4536
use alpha_0  alphaX_5
timestamp 1654634570
transform 1 0 6980 0 1 700
box 0 0 1944 4536
use alpha_0  alphaX_6
timestamp 1654634570
transform 1 0 3855 0 1 700
box 0 0 1944 4536
use alpha_0  alphaX_7
timestamp 1654634570
transform 1 0 730 0 1 700
box 0 0 1944 4536
<< end >>
