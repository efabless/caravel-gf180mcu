VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel
  CLASS BLOCK ;
  FOREIGN caravel ;
  ORIGIN 0.000 0.000 ;
  SIZE 3890.000 BY 5100.000 ;
  PIN clock
    PORT
      LAYER Metal5 ;
        RECT 1082.500 2.000 1142.500 62.000 ;
    END
  END clock
  PIN flash_clk
    PORT
      LAYER Metal5 ;
        RECT 1907.500 2.000 1967.500 62.000 ;
    END
  END flash_clk
  PIN flash_csb
    PORT
      LAYER Metal5 ;
        RECT 1632.500 2.000 1692.500 62.000 ;
    END
  END flash_csb
  PIN flash_io0
    PORT
      LAYER Metal5 ;
        RECT 2182.500 2.000 2242.500 62.000 ;
    END
  END flash_io0
  PIN flash_io1
    PORT
      LAYER Metal5 ;
        RECT 2457.500 2.000 2517.500 62.000 ;
    END
  END flash_io1
  PIN gpio
    PORT
      LAYER Metal5 ;
        RECT 2732.500 2.000 2792.500 62.000 ;
    END
  END gpio
  PIN mprj_io[0]
    PORT
      LAYER Metal5 ;
        RECT 3818.000 452.500 3878.000 512.500 ;
    END
  END mprj_io[0]
  PIN mprj_io[10]
    PORT
      LAYER Metal5 ;
        RECT 3818.000 3247.500 3878.000 3307.500 ;
    END
  END mprj_io[10]
  PIN mprj_io[11]
    PORT
      LAYER Metal5 ;
        RECT 3818.000 3462.500 3878.000 3522.500 ;
    END
  END mprj_io[11]
  PIN mprj_io[12]
    PORT
      LAYER Metal5 ;
        RECT 3818.000 3677.500 3878.000 3737.500 ;
    END
  END mprj_io[12]
  PIN mprj_io[13]
    PORT
      LAYER Metal5 ;
        RECT 3818.000 4107.500 3878.000 4167.500 ;
    END
  END mprj_io[13]
  PIN mprj_io[14]
    PORT
      LAYER Metal5 ;
        RECT 3818.000 4537.500 3878.000 4597.500 ;
    END
  END mprj_io[14]
  PIN mprj_io[15]
    PORT
      LAYER Metal5 ;
        RECT 3277.500 5008.000 3337.500 5068.000 ;
    END
  END mprj_io[15]
  PIN mprj_io[16]
    PORT
      LAYER Metal5 ;
        RECT 2727.500 5008.000 2787.500 5068.000 ;
    END
  END mprj_io[16]
  PIN mprj_io[17]
    PORT
      LAYER Metal5 ;
        RECT 2452.500 5008.000 2512.500 5068.000 ;
    END
  END mprj_io[17]
  PIN mprj_io[18]
    PORT
      LAYER Metal5 ;
        RECT 2177.500 5008.000 2237.500 5068.000 ;
    END
  END mprj_io[18]
  PIN mprj_io[19]
    PORT
      LAYER Metal5 ;
        RECT 1627.500 5008.000 1687.500 5068.000 ;
    END
  END mprj_io[19]
  PIN mprj_io[1]
    PORT
      LAYER Metal5 ;
        RECT 3818.000 667.500 3878.000 727.500 ;
    END
  END mprj_io[1]
  PIN mprj_io[20]
    PORT
      LAYER Metal5 ;
        RECT 1352.500 5008.000 1412.500 5068.000 ;
    END
  END mprj_io[20]
  PIN mprj_io[21]
    PORT
      LAYER Metal5 ;
        RECT 1077.500 5008.000 1137.500 5068.000 ;
    END
  END mprj_io[21]
  PIN mprj_io[22]
    PORT
      LAYER Metal5 ;
        RECT 802.500 5008.000 862.500 5068.000 ;
    END
  END mprj_io[22]
  PIN mprj_io[23]
    PORT
      LAYER Metal5 ;
        RECT 527.500 5008.000 587.500 5068.000 ;
    END
  END mprj_io[23]
  PIN mprj_io[24]
    PORT
      LAYER Metal5 ;
        RECT 2.000 4532.500 62.000 4592.500 ;
    END
  END mprj_io[24]
  PIN mprj_io[25]
    PORT
      LAYER Metal5 ;
        RECT 2.000 3712.500 62.000 3772.500 ;
    END
  END mprj_io[25]
  PIN mprj_io[26]
    PORT
      LAYER Metal5 ;
        RECT 2.000 3507.500 62.000 3567.500 ;
    END
  END mprj_io[26]
  PIN mprj_io[27]
    PORT
      LAYER Metal5 ;
        RECT 2.000 3302.500 62.000 3362.500 ;
    END
  END mprj_io[27]
  PIN mprj_io[28]
    PORT
      LAYER Metal5 ;
        RECT 2.000 3097.500 62.000 3157.500 ;
    END
  END mprj_io[28]
  PIN mprj_io[29]
    PORT
      LAYER Metal5 ;
        RECT 2.000 2892.500 62.000 2952.500 ;
    END
  END mprj_io[29]
  PIN mprj_io[2]
    PORT
      LAYER Metal5 ;
        RECT 3818.000 882.500 3878.000 942.500 ;
    END
  END mprj_io[2]
  PIN mprj_io[30]
    PORT
      LAYER Metal5 ;
        RECT 2.000 2687.500 62.000 2747.500 ;
    END
  END mprj_io[30]
  PIN mprj_io[31]
    PORT
      LAYER Metal5 ;
        RECT 2.000 2482.500 62.000 2542.500 ;
    END
  END mprj_io[31]
  PIN mprj_io[32]
    PORT
      LAYER Metal5 ;
        RECT 2.000 1867.500 62.000 1927.500 ;
    END
  END mprj_io[32]
  PIN mprj_io[33]
    PORT
      LAYER Metal5 ;
        RECT 2.000 1662.500 62.000 1722.500 ;
    END
  END mprj_io[33]
  PIN mprj_io[34]
    PORT
      LAYER Metal5 ;
        RECT 2.000 1457.500 62.000 1517.500 ;
    END
  END mprj_io[34]
  PIN mprj_io[35]
    PORT
      LAYER Metal5 ;
        RECT 2.000 1252.500 62.000 1312.500 ;
    END
  END mprj_io[35]
  PIN mprj_io[36]
    PORT
      LAYER Metal5 ;
        RECT 2.000 1047.500 62.000 1107.500 ;
    END
  END mprj_io[36]
  PIN mprj_io[37]
    PORT
      LAYER Metal5 ;
        RECT 2.000 842.500 62.000 902.500 ;
    END
  END mprj_io[37]
  PIN mprj_io[3]
    PORT
      LAYER Metal5 ;
        RECT 3818.000 1097.500 3878.000 1157.500 ;
    END
  END mprj_io[3]
  PIN mprj_io[4]
    PORT
      LAYER Metal5 ;
        RECT 3818.000 1312.500 3878.000 1372.500 ;
    END
  END mprj_io[4]
  PIN mprj_io[5]
    PORT
      LAYER Metal5 ;
        RECT 3818.000 1527.500 3878.000 1587.500 ;
    END
  END mprj_io[5]
  PIN mprj_io[6]
    PORT
      LAYER Metal5 ;
        RECT 3818.000 1742.500 3878.000 1802.500 ;
    END
  END mprj_io[6]
  PIN mprj_io[7]
    PORT
      LAYER Metal5 ;
        RECT 3818.000 2602.500 3878.000 2662.500 ;
    END
  END mprj_io[7]
  PIN mprj_io[8]
    PORT
      LAYER Metal5 ;
        RECT 3818.000 2817.500 3878.000 2877.500 ;
    END
  END mprj_io[8]
  PIN mprj_io[9]
    PORT
      LAYER Metal5 ;
        RECT 3818.000 3032.500 3878.000 3092.500 ;
    END
  END mprj_io[9]
  PIN resetb
    PORT
      LAYER Metal5 ;
        RECT 807.500 2.000 867.500 62.000 ;
    END
  END resetb
  PIN vdd
    PORT
      LAYER Metal5 ;
        RECT 3818.000 2387.500 3878.000 2447.500 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3818.000 3892.500 3878.000 3952.500 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3818.000 4322.500 3878.000 4382.500 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3282.500 2.000 3342.500 62.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.000 4327.500 62.000 4387.500 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.000 4122.500 62.000 4182.500 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.000 2277.500 62.000 2337.500 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.000 637.500 62.000 697.500 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.000 432.500 62.000 492.500 ;
    END
  END vdd
  PIN vss
    PORT
      LAYER Metal5 ;
        RECT 3002.500 5008.000 3062.500 5068.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1902.500 5008.000 1962.500 5068.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3818.000 1957.500 3878.000 2017.500 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3818.000 2172.500 3878.000 2232.500 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 532.500 2.000 592.500 62.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 1357.500 2.000 1417.500 62.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 3007.500 2.000 3067.500 62.000 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.000 3917.500 62.000 3977.500 ;
    END
    PORT
      LAYER Metal5 ;
        RECT 2.000 2072.500 62.000 2132.500 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 65.540 65.540 3814.460 5004.460 ;
      LAYER Metal2 ;
        RECT 0.000 0.000 3880.000 5070.000 ;
      LAYER Metal3 ;
        RECT 0.000 0.000 3880.000 5070.000 ;
      LAYER Metal4 ;
        RECT 0.000 0.000 3880.000 5070.000 ;
      LAYER Metal5 ;
        RECT 0.000 5068.500 3880.000 5070.000 ;
        RECT 0.000 5007.500 527.000 5068.500 ;
        RECT 588.000 5007.500 802.000 5068.500 ;
        RECT 863.000 5007.500 1077.000 5068.500 ;
        RECT 1138.000 5007.500 1352.000 5068.500 ;
        RECT 1413.000 5007.500 1627.000 5068.500 ;
        RECT 1688.000 5007.500 1902.000 5068.500 ;
        RECT 1963.000 5007.500 2177.000 5068.500 ;
        RECT 2238.000 5007.500 2452.000 5068.500 ;
        RECT 2513.000 5007.500 2727.000 5068.500 ;
        RECT 2788.000 5007.500 3002.000 5068.500 ;
        RECT 3063.000 5007.500 3277.000 5068.500 ;
        RECT 3338.000 5007.500 3880.000 5068.500 ;
        RECT 0.000 4598.000 3880.000 5007.500 ;
        RECT 0.000 4593.000 3817.500 4598.000 ;
        RECT 0.000 4532.000 1.500 4593.000 ;
        RECT 62.500 4537.000 3817.500 4593.000 ;
        RECT 3878.500 4537.000 3880.000 4598.000 ;
        RECT 62.500 4532.000 3880.000 4537.000 ;
        RECT 0.000 4388.000 3880.000 4532.000 ;
        RECT 0.000 4327.000 1.500 4388.000 ;
        RECT 62.500 4383.000 3880.000 4388.000 ;
        RECT 62.500 4327.000 3817.500 4383.000 ;
        RECT 0.000 4322.000 3817.500 4327.000 ;
        RECT 3878.500 4322.000 3880.000 4383.000 ;
        RECT 0.000 4183.000 3880.000 4322.000 ;
        RECT 0.000 4122.000 1.500 4183.000 ;
        RECT 62.500 4168.000 3880.000 4183.000 ;
        RECT 62.500 4122.000 3817.500 4168.000 ;
        RECT 0.000 4107.000 3817.500 4122.000 ;
        RECT 3878.500 4107.000 3880.000 4168.000 ;
        RECT 0.000 3978.000 3880.000 4107.000 ;
        RECT 0.000 3917.000 1.500 3978.000 ;
        RECT 62.500 3953.000 3880.000 3978.000 ;
        RECT 62.500 3917.000 3817.500 3953.000 ;
        RECT 0.000 3892.000 3817.500 3917.000 ;
        RECT 3878.500 3892.000 3880.000 3953.000 ;
        RECT 0.000 3773.000 3880.000 3892.000 ;
        RECT 0.000 3712.000 1.500 3773.000 ;
        RECT 62.500 3738.000 3880.000 3773.000 ;
        RECT 62.500 3712.000 3817.500 3738.000 ;
        RECT 0.000 3677.000 3817.500 3712.000 ;
        RECT 3878.500 3677.000 3880.000 3738.000 ;
        RECT 0.000 3568.000 3880.000 3677.000 ;
        RECT 0.000 3507.000 1.500 3568.000 ;
        RECT 62.500 3523.000 3880.000 3568.000 ;
        RECT 62.500 3507.000 3817.500 3523.000 ;
        RECT 0.000 3462.000 3817.500 3507.000 ;
        RECT 3878.500 3462.000 3880.000 3523.000 ;
        RECT 0.000 3363.000 3880.000 3462.000 ;
        RECT 0.000 3302.000 1.500 3363.000 ;
        RECT 62.500 3308.000 3880.000 3363.000 ;
        RECT 62.500 3302.000 3817.500 3308.000 ;
        RECT 0.000 3247.000 3817.500 3302.000 ;
        RECT 3878.500 3247.000 3880.000 3308.000 ;
        RECT 0.000 3158.000 3880.000 3247.000 ;
        RECT 0.000 3097.000 1.500 3158.000 ;
        RECT 62.500 3097.000 3880.000 3158.000 ;
        RECT 0.000 3093.000 3880.000 3097.000 ;
        RECT 0.000 3032.000 3817.500 3093.000 ;
        RECT 3878.500 3032.000 3880.000 3093.000 ;
        RECT 0.000 2953.000 3880.000 3032.000 ;
        RECT 0.000 2892.000 1.500 2953.000 ;
        RECT 62.500 2892.000 3880.000 2953.000 ;
        RECT 0.000 2878.000 3880.000 2892.000 ;
        RECT 0.000 2817.000 3817.500 2878.000 ;
        RECT 3878.500 2817.000 3880.000 2878.000 ;
        RECT 0.000 2748.000 3880.000 2817.000 ;
        RECT 0.000 2687.000 1.500 2748.000 ;
        RECT 62.500 2687.000 3880.000 2748.000 ;
        RECT 0.000 2663.000 3880.000 2687.000 ;
        RECT 0.000 2602.000 3817.500 2663.000 ;
        RECT 3878.500 2602.000 3880.000 2663.000 ;
        RECT 0.000 2543.000 3880.000 2602.000 ;
        RECT 0.000 2482.000 1.500 2543.000 ;
        RECT 62.500 2482.000 3880.000 2543.000 ;
        RECT 0.000 2448.000 3880.000 2482.000 ;
        RECT 0.000 2387.000 3817.500 2448.000 ;
        RECT 3878.500 2387.000 3880.000 2448.000 ;
        RECT 0.000 2338.000 3880.000 2387.000 ;
        RECT 0.000 2277.000 1.500 2338.000 ;
        RECT 62.500 2277.000 3880.000 2338.000 ;
        RECT 0.000 2233.000 3880.000 2277.000 ;
        RECT 0.000 2172.000 3817.500 2233.000 ;
        RECT 3878.500 2172.000 3880.000 2233.000 ;
        RECT 0.000 2133.000 3880.000 2172.000 ;
        RECT 0.000 2072.000 1.500 2133.000 ;
        RECT 62.500 2072.000 3880.000 2133.000 ;
        RECT 0.000 2018.000 3880.000 2072.000 ;
        RECT 0.000 1957.000 3817.500 2018.000 ;
        RECT 3878.500 1957.000 3880.000 2018.000 ;
        RECT 0.000 1928.000 3880.000 1957.000 ;
        RECT 0.000 1867.000 1.500 1928.000 ;
        RECT 62.500 1867.000 3880.000 1928.000 ;
        RECT 0.000 1803.000 3880.000 1867.000 ;
        RECT 0.000 1742.000 3817.500 1803.000 ;
        RECT 3878.500 1742.000 3880.000 1803.000 ;
        RECT 0.000 1723.000 3880.000 1742.000 ;
        RECT 0.000 1662.000 1.500 1723.000 ;
        RECT 62.500 1662.000 3880.000 1723.000 ;
        RECT 0.000 1588.000 3880.000 1662.000 ;
        RECT 0.000 1527.000 3817.500 1588.000 ;
        RECT 3878.500 1527.000 3880.000 1588.000 ;
        RECT 0.000 1518.000 3880.000 1527.000 ;
        RECT 0.000 1457.000 1.500 1518.000 ;
        RECT 62.500 1457.000 3880.000 1518.000 ;
        RECT 0.000 1373.000 3880.000 1457.000 ;
        RECT 0.000 1313.000 3817.500 1373.000 ;
        RECT 0.000 1252.000 1.500 1313.000 ;
        RECT 62.500 1312.000 3817.500 1313.000 ;
        RECT 3878.500 1312.000 3880.000 1373.000 ;
        RECT 62.500 1252.000 3880.000 1312.000 ;
        RECT 0.000 1158.000 3880.000 1252.000 ;
        RECT 0.000 1108.000 3817.500 1158.000 ;
        RECT 0.000 1047.000 1.500 1108.000 ;
        RECT 62.500 1097.000 3817.500 1108.000 ;
        RECT 3878.500 1097.000 3880.000 1158.000 ;
        RECT 62.500 1047.000 3880.000 1097.000 ;
        RECT 0.000 943.000 3880.000 1047.000 ;
        RECT 0.000 903.000 3817.500 943.000 ;
        RECT 0.000 842.000 1.500 903.000 ;
        RECT 62.500 882.000 3817.500 903.000 ;
        RECT 3878.500 882.000 3880.000 943.000 ;
        RECT 62.500 842.000 3880.000 882.000 ;
        RECT 0.000 728.000 3880.000 842.000 ;
        RECT 0.000 698.000 3817.500 728.000 ;
        RECT 0.000 637.000 1.500 698.000 ;
        RECT 62.500 667.000 3817.500 698.000 ;
        RECT 3878.500 667.000 3880.000 728.000 ;
        RECT 62.500 637.000 3880.000 667.000 ;
        RECT 0.000 513.000 3880.000 637.000 ;
        RECT 0.000 493.000 3817.500 513.000 ;
        RECT 0.000 432.000 1.500 493.000 ;
        RECT 62.500 452.000 3817.500 493.000 ;
        RECT 3878.500 452.000 3880.000 513.000 ;
        RECT 62.500 432.000 3880.000 452.000 ;
        RECT 0.000 62.500 3880.000 432.000 ;
        RECT 0.000 1.500 532.000 62.500 ;
        RECT 593.000 1.500 807.000 62.500 ;
        RECT 868.000 1.500 1082.000 62.500 ;
        RECT 1143.000 1.500 1357.000 62.500 ;
        RECT 1418.000 1.500 1632.000 62.500 ;
        RECT 1693.000 1.500 1907.000 62.500 ;
        RECT 1968.000 1.500 2182.000 62.500 ;
        RECT 2243.000 1.500 2457.000 62.500 ;
        RECT 2518.000 1.500 2732.000 62.500 ;
        RECT 2793.000 1.500 3007.000 62.500 ;
        RECT 3068.000 1.500 3282.000 62.500 ;
        RECT 3343.000 1.500 3880.000 62.500 ;
        RECT 0.000 0.000 3880.000 1.500 ;
  END
END caravel
END LIBRARY

