* Simple POR testbench (No. 2:  Running at slow VDD ramp (but not too slow))

.include /usr/share/pdk/gf180mcuC/libs.tech/ngspice/design.ngspice
.lib /usr/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice typical
.lib /usr/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /usr/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.ngspice mimcap_typical
.include simple_por.spice

* Very slow ramp up and down.  Ramp is about half the POR delay time.
* The POR should behave correctly for any power supply ramp up to around
* this risetime.
V0 VDD 0 PWL(0 0 1u 0 20m 5 80m 5 100m 0)

X0 VDD 0 PORB POR simple_por

.control
tran 1u 101m
plot V(VDD) V(POR) V(PORB)
.endc
