magic
tech gf180mcuD
magscale 1 10
timestamp 1655304105
<< error_p >>
rect -48 -255 -37 -209
<< nwell >>
rect -368 -486 378 486
<< mvpmos >>
rect -50 -176 60 224
<< mvpdiff >>
rect -138 211 -50 224
rect -138 -163 -125 211
rect -79 -163 -50 211
rect -138 -176 -50 -163
rect 60 211 148 224
rect 60 -163 89 211
rect 135 -163 148 211
rect 60 -176 148 -163
<< mvpdiffc >>
rect -125 -163 -79 211
rect 89 -163 135 211
<< mvnsubdiff >>
rect -282 387 292 400
rect -282 341 -166 387
rect 166 341 292 387
rect -282 328 292 341
rect -282 284 -210 328
rect -282 -284 -269 284
rect -223 -284 -210 284
rect 220 284 292 328
rect -282 -328 -210 -284
rect 220 -284 233 284
rect 279 -284 292 284
rect 220 -328 292 -284
rect -282 -400 292 -328
<< mvnsubdiffcont >>
rect -166 341 166 387
rect -269 -284 -223 284
rect 233 -284 279 284
<< polysilicon >>
rect -50 224 60 268
rect -50 -209 60 -176
rect -50 -255 -37 -209
rect 47 -255 60 -209
rect -50 -268 60 -255
<< polycontact >>
rect -37 -255 47 -209
<< metal1 >>
rect -269 341 -166 387
rect 166 341 279 387
rect -269 284 -223 341
rect 233 284 279 341
rect -125 211 -79 222
rect -125 -174 -79 -163
rect 89 211 135 222
rect 89 -174 135 -163
rect -48 -255 -37 -209
rect 47 -255 58 -209
rect -269 -341 -223 -284
rect 233 -341 279 -284
rect -269 -387 279 -341
<< properties >>
string FIXED_BBOX -246 -364 246 364
string gencell pmos_6p0
string library gf180mcu
string parameters w 2.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.5 wmin 0.3 full_metal 1 compatible {pmos_3p3 pmos_6p0}
<< end >>
