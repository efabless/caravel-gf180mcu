* NGSPICE file created from caravel.ext - technology: gf180mcuC

* Black-box entry subcircuit for gpio_control_block abstract view
.subckt gpio_control_block VDD VSS gpio_defaults[0] gpio_defaults[1] gpio_defaults[2]
+ gpio_defaults[3] gpio_defaults[4] gpio_defaults[5] gpio_defaults[6] gpio_defaults[7]
+ gpio_defaults[8] gpio_defaults[9] mgmt_gpio_in mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_drive_sel[0]
+ pad_gpio_drive_sel[1] pad_gpio_in pad_gpio_inen pad_gpio_out pad_gpio_outen pad_gpio_pulldown_sel
+ pad_gpio_pullup_sel pad_gpio_schmitt_sel pad_gpio_slew_sel resetn resetn_out serial_clock
+ serial_clock_out serial_data_in serial_data_out serial_load serial_load_out user_gpio_in
+ user_gpio_oeb user_gpio_out zero
.ends

* Black-box entry subcircuit for gpio_defaults_block abstract view
.subckt gpio_defaults_block gpio_defaults[0] gpio_defaults[1] gpio_defaults[2] gpio_defaults[3]
+ gpio_defaults[4] gpio_defaults[5] gpio_defaults[6] gpio_defaults[7] gpio_defaults[8]
+ gpio_defaults[9] VDD VSS
.ends

* Black-box entry subcircuit for digital_pll abstract view
.subckt digital_pll VDD VSS clockp[0] clockp[1] dco div[0] div[1] div[2] div[3] div[4]
+ enable ext_trim[0] ext_trim[10] ext_trim[11] ext_trim[12] ext_trim[13] ext_trim[14]
+ ext_trim[15] ext_trim[16] ext_trim[17] ext_trim[18] ext_trim[19] ext_trim[1] ext_trim[20]
+ ext_trim[21] ext_trim[22] ext_trim[23] ext_trim[24] ext_trim[25] ext_trim[2] ext_trim[3]
+ ext_trim[4] ext_trim[5] ext_trim[6] ext_trim[7] ext_trim[8] ext_trim[9] osc resetb
.ends

* Black-box entry subcircuit for GF_NI_FILL10 abstract view
.subckt GF_NI_FILL10 DVDD DVSS VDD VSS
.ends

* Black-box entry subcircuit for GF_NI_IN_S abstract view
.subckt GF_NI_IN_S DVDD DVSS PAD PD PU VDD VSS Y
.ends

* Black-box entry subcircuit for GF_NI_DVSS abstract view
.subckt GF_NI_DVSS DVDD DVSS VDD
.ends

* Black-box entry subcircuit for GF_NI_DVDD abstract view
.subckt GF_NI_DVDD DVDD DVSS VSS
.ends

* Black-box entry subcircuit for GF_NI_FILL5 abstract view
.subckt GF_NI_FILL5 DVDD DVSS VDD VSS
.ends

* Black-box entry subcircuit for GF_NI_BI_T abstract view
.subckt GF_NI_BI_T A CS DVDD DVSS IE OE PAD PD PDRV0 PDRV1 PU SL VDD VSS Y
.ends

* Black-box entry subcircuit for GF_NI_IN_C abstract view
.subckt GF_NI_IN_C DVDD DVSS PAD PD PU VDD VSS Y
.ends

* Black-box entry subcircuit for GF_NI_COR abstract view
.subckt GF_NI_COR DVDD DVSS VDD VSS
.ends

.subckt chip_io clock clock_core flash_clk flash_clk_core flash_clk_oe_core flash_csb
+ flash_csb_core flash_csb_oe_core flash_io0 flash_io0_di_core flash_io0_do_core flash_io0_ie_core
+ flash_io0_oe_core flash_io1 flash_io1_di_core flash_io1_do_core flash_io1_ie_core
+ flash_io1_oe_core gpio gpio_drive_select_core[0] gpio_drive_select_core[1] gpio_in_core
+ gpio_inen_core gpio_out_core gpio_outen_core gpio_pd_select gpio_pu_select gpio_schmitt_select
+ gpio_slew_select mprj_io[0] mprj_io[10] mprj_io[11] mprj_io[12] mprj_io[13] mprj_io[14]
+ mprj_io[15] mprj_io[16] mprj_io[17] mprj_io[18] mprj_io[19] mprj_io[1] mprj_io[20]
+ mprj_io[21] mprj_io[22] mprj_io[23] mprj_io[24] mprj_io[25] mprj_io[26] mprj_io[27]
+ mprj_io[28] mprj_io[29] mprj_io[2] mprj_io[30] mprj_io[31] mprj_io[32] mprj_io[33]
+ mprj_io[34] mprj_io[35] mprj_io[36] mprj_io[37] mprj_io[3] mprj_io[4] mprj_io[5]
+ mprj_io[6] mprj_io[7] mprj_io[8] mprj_io[9] mprj_io_drive_sel[0] mprj_io_drive_sel[10]
+ mprj_io_drive_sel[11] mprj_io_drive_sel[12] mprj_io_drive_sel[13] mprj_io_drive_sel[14]
+ mprj_io_drive_sel[15] mprj_io_drive_sel[16] mprj_io_drive_sel[17] mprj_io_drive_sel[18]
+ mprj_io_drive_sel[19] mprj_io_drive_sel[1] mprj_io_drive_sel[20] mprj_io_drive_sel[21]
+ mprj_io_drive_sel[22] mprj_io_drive_sel[23] mprj_io_drive_sel[24] mprj_io_drive_sel[25]
+ mprj_io_drive_sel[26] mprj_io_drive_sel[27] mprj_io_drive_sel[28] mprj_io_drive_sel[29]
+ mprj_io_drive_sel[2] mprj_io_drive_sel[30] mprj_io_drive_sel[31] mprj_io_drive_sel[32]
+ mprj_io_drive_sel[33] mprj_io_drive_sel[34] mprj_io_drive_sel[35] mprj_io_drive_sel[36]
+ mprj_io_drive_sel[37] mprj_io_drive_sel[38] mprj_io_drive_sel[39] mprj_io_drive_sel[3]
+ mprj_io_drive_sel[40] mprj_io_drive_sel[41] mprj_io_drive_sel[42] mprj_io_drive_sel[43]
+ mprj_io_drive_sel[44] mprj_io_drive_sel[45] mprj_io_drive_sel[46] mprj_io_drive_sel[47]
+ mprj_io_drive_sel[48] mprj_io_drive_sel[49] mprj_io_drive_sel[4] mprj_io_drive_sel[51]
+ mprj_io_drive_sel[525] mprj_io_drive_sel[52] mprj_io_drive_sel[53] mprj_io_drive_sel[54]
+ mprj_io_drive_sel[55] mprj_io_drive_sel[56] mprj_io_drive_sel[57] mprj_io_drive_sel[58]
+ mprj_io_drive_sel[59] mprj_io_drive_sel[5] mprj_io_drive_sel[61] mprj_io_drive_sel[62]
+ mprj_io_drive_sel[63] mprj_io_drive_sel[64] mprj_io_drive_sel[65] mprj_io_drive_sel[66]
+ mprj_io_drive_sel[67] mprj_io_drive_sel[68] mprj_io_drive_sel[69] mprj_io_drive_sel[6]
+ mprj_io_drive_sel[70] mprj_io_drive_sel[71] mprj_io_drive_sel[72] mprj_io_drive_sel[73]
+ mprj_io_drive_sel[74] mprj_io_drive_sel[75] mprj_io_drive_sel[7] mprj_io_drive_sel[8]
+ mprj_io_drive_sel[9] mprj_io_in[0] mprj_io_in[10] mprj_io_in[11] mprj_io_in[12]
+ mprj_io_in[13] mprj_io_in[14] mprj_io_in[15] mprj_io_in[16] mprj_io_in[17] mprj_io_in[18]
+ mprj_io_in[19] mprj_io_in[1] mprj_io_in[20] mprj_io_in[21] mprj_io_in[22] mprj_io_in[23]
+ mprj_io_in[24] mprj_io_in[25] mprj_io_in[26] mprj_io_in[27] mprj_io_in[28] mprj_io_in[29]
+ mprj_io_in[2] mprj_io_in[30] mprj_io_in[31] mprj_io_in[32] mprj_io_in[33] mprj_io_in[34]
+ mprj_io_in[35] mprj_io_in[36] mprj_io_in[37] mprj_io_in[3] mprj_io_in[4] mprj_io_in[5]
+ mprj_io_in[6] mprj_io_in[7] mprj_io_in[8] mprj_io_in[9] mprj_io_inen[0] mprj_io_inen[10]
+ mprj_io_inen[11] mprj_io_inen[12] mprj_io_inen[13] mprj_io_inen[14] mprj_io_inen[15]
+ mprj_io_inen[16] mprj_io_inen[17] mprj_io_inen[18] mprj_io_inen[19] mprj_io_inen[1]
+ mprj_io_inen[20] mprj_io_inen[21] mprj_io_inen[22] mprj_io_inen[23] mprj_io_inen[24]
+ mprj_io_inen[25] mprj_io_inen[26] mprj_io_inen[27] mprj_io_inen[28] mprj_io_inen[29]
+ mprj_io_inen[2] mprj_io_inen[30] mprj_io_inen[31] mprj_io_inen[32] mprj_io_inen[33]
+ mprj_io_inen[34] mprj_io_inen[35] mprj_io_inen[36] mprj_io_inen[37] mprj_io_inen[3]
+ mprj_io_inen[4] mprj_io_inen[5] mprj_io_inen[6] mprj_io_inen[7] mprj_io_inen[8]
+ mprj_io_inen[9] mprj_io_out[0] mprj_io_out[10] mprj_io_out[11] mprj_io_out[12] mprj_io_out[13]
+ mprj_io_out[14] mprj_io_out[15] mprj_io_out[16] mprj_io_out[17] mprj_io_out[18]
+ mprj_io_out[19] mprj_io_out[1] mprj_io_out[20] mprj_io_out[21] mprj_io_out[22] mprj_io_out[23]
+ mprj_io_out[24] mprj_io_out[25] mprj_io_out[26] mprj_io_out[27] mprj_io_out[28]
+ mprj_io_out[29] mprj_io_out[2] mprj_io_out[30] mprj_io_out[31] mprj_io_out[32] mprj_io_out[33]
+ mprj_io_out[34] mprj_io_out[35] mprj_io_out[36] mprj_io_out[37] mprj_io_out[3] mprj_io_out[4]
+ mprj_io_out[5] mprj_io_out[6] mprj_io_out[7] mprj_io_out[8] mprj_io_out[9] mprj_io_outen[0]
+ mprj_io_outen[10] mprj_io_outen[11] mprj_io_outen[12] mprj_io_outen[13] mprj_io_outen[14]
+ mprj_io_outen[15] mprj_io_outen[16] mprj_io_outen[17] mprj_io_outen[18] mprj_io_outen[19]
+ mprj_io_outen[1] mprj_io_outen[20] mprj_io_outen[21] mprj_io_outen[22] mprj_io_outen[23]
+ mprj_io_outen[24] mprj_io_outen[25] mprj_io_outen[26] mprj_io_outen[27] mprj_io_outen[28]
+ mprj_io_outen[29] mprj_io_outen[2] mprj_io_outen[30] mprj_io_outen[31] mprj_io_outen[32]
+ mprj_io_outen[33] mprj_io_outen[34] mprj_io_outen[35] mprj_io_outen[36] mprj_io_outen[37]
+ mprj_io_outen[3] mprj_io_outen[4] mprj_io_outen[5] mprj_io_outen[6] mprj_io_outen[7]
+ mprj_io_outen[8] mprj_io_outen[9] mprj_io_pd_select[0] mprj_io_pd_select[10] mprj_io_pd_select[11]
+ mprj_io_pd_select[12] mprj_io_pd_select[13] mprj_io_pd_select[14] mprj_io_pd_select[15]
+ mprj_io_pd_select[16] mprj_io_pd_select[17] mprj_io_pd_select[18] mprj_io_pd_select[19]
+ mprj_io_pd_select[1] mprj_io_pd_select[20] mprj_io_pd_select[21] mprj_io_pd_select[22]
+ mprj_io_pd_select[23] mprj_io_pd_select[24] mprj_io_pd_select[25] mprj_io_pd_select[26]
+ mprj_io_pd_select[27] mprj_io_pd_select[28] mprj_io_pd_select[29] mprj_io_pd_select[2]
+ mprj_io_pd_select[30] mprj_io_pd_select[31] mprj_io_pd_select[32] mprj_io_pd_select[33]
+ mprj_io_pd_select[34] mprj_io_pd_select[35] mprj_io_pd_select[36] mprj_io_pd_select[37]
+ mprj_io_pd_select[3] mprj_io_pd_select[4] mprj_io_pd_select[5] mprj_io_pd_select[6]
+ mprj_io_pd_select[7] mprj_io_pd_select[8] mprj_io_pd_select[9] mprj_io_pu_select[0]
+ mprj_io_pu_select[10] mprj_io_pu_select[11] mprj_io_pu_select[12] mprj_io_pu_select[13]
+ mprj_io_pu_select[14] mprj_io_pu_select[15] mprj_io_pu_select[16] mprj_io_pu_select[17]
+ mprj_io_pu_select[18] mprj_io_pu_select[19] mprj_io_pu_select[1] mprj_io_pu_select[20]
+ mprj_io_pu_select[21] mprj_io_pu_select[22] mprj_io_pu_select[23] mprj_io_pu_select[24]
+ mprj_io_pu_select[25] mprj_io_pu_select[26] mprj_io_pu_select[27] mprj_io_pu_select[28]
+ mprj_io_pu_select[29] mprj_io_pu_select[2] mprj_io_pu_select[30] mprj_io_pu_select[31]
+ mprj_io_pu_select[32] mprj_io_pu_select[33] mprj_io_pu_select[34] mprj_io_pu_select[35]
+ mprj_io_pu_select[36] mprj_io_pu_select[37] mprj_io_pu_select[3] mprj_io_pu_select[4]
+ mprj_io_pu_select[5] mprj_io_pu_select[6] mprj_io_pu_select[7] mprj_io_pu_select[8]
+ mprj_io_pu_select[9] mprj_io_schmitt_select[0] mprj_io_schmitt_select[10] mprj_io_schmitt_select[11]
+ mprj_io_schmitt_select[12] mprj_io_schmitt_select[13] mprj_io_schmitt_select[14]
+ mprj_io_schmitt_select[15] mprj_io_schmitt_select[16] mprj_io_schmitt_select[17]
+ mprj_io_schmitt_select[18] mprj_io_schmitt_select[19] mprj_io_schmitt_select[1]
+ mprj_io_schmitt_select[20] mprj_io_schmitt_select[21] mprj_io_schmitt_select[22]
+ mprj_io_schmitt_select[23] mprj_io_schmitt_select[24] mprj_io_schmitt_select[25]
+ mprj_io_schmitt_select[26] mprj_io_schmitt_select[27] mprj_io_schmitt_select[28]
+ mprj_io_schmitt_select[29] mprj_io_schmitt_select[2] mprj_io_schmitt_select[30]
+ mprj_io_schmitt_select[31] mprj_io_schmitt_select[32] mprj_io_schmitt_select[33]
+ mprj_io_schmitt_select[34] mprj_io_schmitt_select[35] mprj_io_schmitt_select[36]
+ mprj_io_schmitt_select[37] mprj_io_schmitt_select[3] mprj_io_schmitt_select[4] mprj_io_schmitt_select[5]
+ mprj_io_schmitt_select[6] mprj_io_schmitt_select[7] mprj_io_schmitt_select[8] mprj_io_schmitt_select[9]
+ mprj_io_slew_select[0] mprj_io_slew_select[10] mprj_io_slew_select[11] mprj_io_slew_select[12]
+ mprj_io_slew_select[13] mprj_io_slew_select[14] mprj_io_slew_select[15] mprj_io_slew_select[16]
+ mprj_io_slew_select[17] mprj_io_slew_select[18] mprj_io_slew_select[19] mprj_io_slew_select[1]
+ mprj_io_slew_select[20] mprj_io_slew_select[21] mprj_io_slew_select[22] mprj_io_slew_select[23]
+ mprj_io_slew_select[24] mprj_io_slew_select[25] mprj_io_slew_select[26] mprj_io_slew_select[27]
+ mprj_io_slew_select[28] mprj_io_slew_select[29] mprj_io_slew_select[2] mprj_io_slew_select[30]
+ mprj_io_slew_select[31] mprj_io_slew_select[32] mprj_io_slew_select[33] mprj_io_slew_select[34]
+ mprj_io_slew_select[35] mprj_io_slew_select[36] mprj_io_slew_select[37] mprj_io_slew_select[3]
+ mprj_io_slew_select[4] mprj_io_slew_select[5] mprj_io_slew_select[6] mprj_io_slew_select[7]
+ mprj_io_slew_select[8] mprj_io_slew_select[9] resetb resetb_core vdd vss GF_NI_COR_3/VSS
+ GF_NI_COR_3/VDD
XGF_NI_FILL10_513 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_524 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_535 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_546 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_557 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_568 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_579 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_502 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_94 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_83 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_72 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_61 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_50 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_398 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_387 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_376 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_365 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_354 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_343 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_332 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_321 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_310 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_140 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_151 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_162 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_173 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_184 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_195 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_909 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_706 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_717 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_728 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_739 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_514 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_525 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_536 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_547 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_558 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_569 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_503 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_95 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_84 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_73 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_62 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_51 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_40 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_399 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_388 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_377 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_366 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_355 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_344 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_333 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_322 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_311 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_300 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_130 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_141 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_152 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_163 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_174 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_185 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_196 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_707 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_718 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_729 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_515 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_526 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_537 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_504 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_548 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_559 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_96 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_85 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_74 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_63 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_52 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_41 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_30 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_389 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_378 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_367 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_356 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_345 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_334 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_323 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_312 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_301 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_890 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_120 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_131 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_142 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_153 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_164 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_175 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_186 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_197 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_708 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_719 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_516 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_527 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_538 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_549 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_505 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_97 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_86 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_75 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_64 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_53 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_42 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_31 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_20 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_379 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_368 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_357 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_346 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_335 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_324 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_313 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_302 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_880 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_891 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_110 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_121 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_132 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_143 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_154 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_165 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_176 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_187 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_198 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_709 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_517 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_528 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_539 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_506 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_87 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_65 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_76 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_54 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_43 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_32 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_21 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_10 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_98 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_303 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_369 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_358 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_347 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_336 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_325 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_314 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_870 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_881 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_892 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_IN_S_0 GF_NI_COR_3/VDD GF_NI_COR_3/VSS resetb GF_NI_IN_S_0/PD GF_NI_IN_S_0/PU
+ GF_NI_COR_3/VDD GF_NI_COR_3/VSS resetb_core GF_NI_IN_S
XGF_NI_FILL10_100 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_111 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_122 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_133 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_144 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_155 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_166 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_177 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_188 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_199 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_DVSS_0 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_DVSS
XGF_NI_FILL10_518 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_529 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_507 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_44 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_33 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_22 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_11 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_66 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_77 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_55 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_88 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_99 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_359 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_348 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_337 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_326 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_315 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_304 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_860 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_882 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_893 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_871 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_101 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_112 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_123 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_134 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_145 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_156 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_167 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_178 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_690 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_189 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_DVSS_1 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_DVSS
XGF_NI_FILL10_519 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_508 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_67 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_45 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_56 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_34 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_23 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_12 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_78 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_89 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_349 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_338 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_327 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_316 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_305 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_850 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_861 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_872 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_883 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_894 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_102 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_113 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_124 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_135 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_146 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_157 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_168 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_179 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_680 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_691 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_DVSS_2 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_DVSS
XGF_NI_FILL10_509 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_68 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_46 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_57 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_35 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_24 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_13 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_79 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_339 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_328 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_317 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_306 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_840 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_851 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_862 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_873 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_884 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_895 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_DVDD_0 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VSS GF_NI_DVDD
XGF_NI_FILL10_103 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_114 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_125 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_136 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_147 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_158 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_169 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_670 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_681 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_692 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL5_0 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL5
XGF_NI_DVSS_3 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_DVSS
XGF_NI_FILL10_69 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_58 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_47 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_36 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_25 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_14 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_329 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_318 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_307 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_830 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_841 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_852 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_863 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_874 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_885 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_896 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_DVDD_1 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VSS GF_NI_DVDD
XGF_NI_FILL10_104 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_115 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_126 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_137 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_148 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_159 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_660 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_671 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_682 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_693 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL5_1 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL5
XGF_NI_FILL10_490 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_DVSS_4 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_DVSS
XGF_NI_FILL10_59 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_48 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_37 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_26 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_15 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_319 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_308 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_820 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_831 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_842 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_853 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_864 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_875 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_DVDD_2 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VSS GF_NI_DVDD
XGF_NI_FILL10_897 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_886 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_105 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_116 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_127 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_138 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_149 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_650 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_661 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_672 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_683 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_694 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL5_2 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL5
XGF_NI_FILL10_491 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_480 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_0 flash_csb_core GF_NI_BI_T_0/CS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_BI_T_0/IE
+ flash_csb_oe_core flash_csb GF_NI_BI_T_0/PD GF_NI_BI_T_0/PDRV0 GF_NI_BI_T_0/PDRV1
+ GF_NI_BI_T_0/PU GF_NI_BI_T_0/SL GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_BI_T_0/Y GF_NI_BI_T
XGF_NI_DVSS_5 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_DVSS
XGF_NI_FILL10_49 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_38 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_27 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_16 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_309 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_810 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_821 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_832 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_843 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_854 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_865 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_876 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_887 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_898 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_DVDD_3 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VSS GF_NI_DVDD
XGF_NI_FILL10_106 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_117 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_128 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_139 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_640 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_651 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_662 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_673 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_684 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_695 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_492 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_481 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_470 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_1 flash_clk_core GF_NI_BI_T_1/CS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_BI_T_1/IE
+ flash_clk_oe_core flash_clk GF_NI_BI_T_1/PD GF_NI_BI_T_1/PDRV0 GF_NI_BI_T_1/PDRV1
+ GF_NI_BI_T_1/PU GF_NI_BI_T_1/SL GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_BI_T_1/Y GF_NI_BI_T
XGF_NI_DVSS_6 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_DVSS
XGF_NI_FILL10_39 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_28 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_17 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_811 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_822 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_833 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_844 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_855 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_866 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_877 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_888 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_899 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_800 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_DVDD_4 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VSS GF_NI_DVDD
XGF_NI_FILL10_630 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_107 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_118 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_129 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_641 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_652 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_663 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_674 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_685 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_696 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_493 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_482 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_471 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_460 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_2 flash_io0_do_core GF_NI_BI_T_2/CS GF_NI_COR_3/VDD GF_NI_COR_3/VSS flash_io0_ie_core
+ flash_io0_oe_core flash_io0 GF_NI_BI_T_2/PD GF_NI_BI_T_2/PDRV0 GF_NI_BI_T_2/PDRV1
+ GF_NI_BI_T_2/PU GF_NI_BI_T_2/SL GF_NI_COR_3/VDD GF_NI_COR_3/VSS flash_io0_di_core
+ GF_NI_BI_T
XGF_NI_FILL10_290 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_29 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_18 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_801 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_812 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_823 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_834 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_845 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_867 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_878 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_889 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_856 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_DVDD_5 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VSS GF_NI_DVDD
XGF_NI_FILL10_108 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_119 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_620 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_631 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_642 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_653 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_664 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_675 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_686 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_697 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_494 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_483 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_472 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_461 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_450 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_3 flash_io1_do_core GF_NI_BI_T_3/CS GF_NI_COR_3/VDD GF_NI_COR_3/VSS flash_io1_ie_core
+ flash_io1_oe_core flash_io1 GF_NI_BI_T_3/PD GF_NI_BI_T_3/PDRV0 GF_NI_BI_T_3/PDRV1
+ GF_NI_BI_T_3/PU GF_NI_BI_T_3/SL GF_NI_COR_3/VDD GF_NI_COR_3/VSS flash_io1_di_core
+ GF_NI_BI_T
XGF_NI_DVSS_8 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_DVSS
XGF_NI_FILL10_280 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_291 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_19 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_802 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_813 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_824 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_835 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_846 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_857 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_868 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_879 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_109 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_610 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_621 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_632 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_643 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_654 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_665 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_676 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_687 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_698 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_495 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_484 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_473 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_462 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_451 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_440 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_4 gpio_out_core gpio_schmitt_select GF_NI_COR_3/VDD GF_NI_COR_3/VSS gpio_inen_core
+ gpio_outen_core gpio gpio_pd_select gpio_drive_select_core[0] gpio_drive_select_core[1]
+ gpio_pu_select gpio_slew_select GF_NI_COR_3/VDD GF_NI_COR_3/VSS gpio_in_core GF_NI_BI_T
XGF_NI_DVSS_9 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_DVSS
XGF_NI_FILL10_292 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_270 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_281 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1040 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_803 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_814 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_825 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_836 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_858 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_869 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_847 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_DVDD_7 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VSS GF_NI_DVDD
XGF_NI_FILL10_600 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_611 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_622 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_633 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_644 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_655 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_666 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_677 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_688 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_699 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_496 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_485 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_474 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_463 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_452 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_441 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_430 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_5 mprj_io_out[0] mprj_io_schmitt_select[0] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[0] mprj_io_outen[0] mprj_io[0] mprj_io_pd_select[0] mprj_io_drive_sel[0]
+ mprj_io_drive_sel[1] mprj_io_pu_select[0] mprj_io_slew_select[0] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[0] GF_NI_BI_T
XGF_NI_FILL10_260 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_271 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_282 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_293 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1041 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1030 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_DVDD_8 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VSS GF_NI_DVDD
XGF_NI_FILL10_804 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_815 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_826 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_837 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_848 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_859 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_601 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_612 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_623 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_634 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_645 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_656 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_667 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_678 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_689 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_497 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_486 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_475 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_464 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_453 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_442 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_431 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_420 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_6 mprj_io_out[1] mprj_io_schmitt_select[1] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[1] mprj_io_outen[1] mprj_io[1] mprj_io_pd_select[1] mprj_io_drive_sel[2]
+ mprj_io_drive_sel[3] mprj_io_pu_select[1] mprj_io_slew_select[1] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[1] GF_NI_BI_T
XGF_NI_FILL10_294 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1042 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_250 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1031 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1020 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_261 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_272 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_283 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_805 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_816 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_838 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_849 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_827 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_DVDD_9 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VSS GF_NI_DVDD
XGF_NI_FILL10_602 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_613 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_624 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_635 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_646 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_657 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_668 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_679 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_498 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_487 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_476 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_465 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_454 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_443 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_432 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_421 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_410 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_7 mprj_io_out[2] mprj_io_schmitt_select[2] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[2] mprj_io_outen[2] mprj_io[2] mprj_io_pd_select[2] mprj_io_drive_sel[5]
+ mprj_io_drive_sel[4] mprj_io_pu_select[2] mprj_io_slew_select[2] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[2] GF_NI_BI_T
XGF_NI_FILL10_295 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_240 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_251 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1010 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_262 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_273 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_284 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_0 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_1043 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1032 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1021 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_806 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_817 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_828 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_839 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_603 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_614 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_625 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_636 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_647 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_658 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_669 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_499 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_488 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_477 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_466 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_455 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_444 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_433 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_422 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_411 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_400 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_8 mprj_io_out[3] mprj_io_schmitt_select[3] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[3] mprj_io_outen[3] mprj_io[3] mprj_io_pd_select[3] mprj_io_drive_sel[7]
+ mprj_io_drive_sel[6] mprj_io_pu_select[3] mprj_io_slew_select[3] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[3] GF_NI_BI_T
XGF_NI_FILL10_296 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_230 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_241 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_252 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_263 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_274 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_285 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_1044 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1033 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1022 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1011 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1000 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_807 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_829 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_818 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_604 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_615 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_626 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_637 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_648 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_659 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_412 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_401 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_489 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_478 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_467 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_456 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_445 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_434 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_423 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_9 mprj_io_out[4] mprj_io_schmitt_select[4] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[4] mprj_io_outen[4] mprj_io[4] mprj_io_pd_select[4] mprj_io_drive_sel[9]
+ mprj_io_drive_sel[8] mprj_io_pu_select[4] mprj_io_slew_select[4] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[4] GF_NI_BI_T
XGF_NI_FILL10_990 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_297 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_220 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_231 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_242 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_253 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_264 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_275 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_286 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_2 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_1045 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1034 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1001 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_808 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_819 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_605 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_616 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_627 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_638 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_649 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_479 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_468 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_457 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_446 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_435 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_424 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_413 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_402 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_980 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_991 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_210 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_221 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_232 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_243 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_254 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_265 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_276 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_287 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_298 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_3 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_1046 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1035 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1024 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1013 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1002 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_809 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_606 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_617 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_628 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_639 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_469 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_458 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_447 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_436 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_425 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_414 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_403 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_970 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_981 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_992 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_40 mprj_io_out[33] mprj_io_schmitt_select[33] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[33] mprj_io_outen[33] mprj_io[33] mprj_io_pd_select[33] mprj_io_drive_sel[66]
+ mprj_io_drive_sel[67] mprj_io_pu_select[33] mprj_io_slew_select[33] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[33] GF_NI_BI_T
XGF_NI_FILL10_299 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1047 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_200 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_211 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_222 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_233 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_244 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_255 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1036 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1025 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1014 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_266 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_277 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1003 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_288 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_4 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_607 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_618 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_629 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_459 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_448 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_437 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_426 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_415 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_404 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_960 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_971 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_982 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_993 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_30 mprj_io_out[28] mprj_io_schmitt_select[28] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[28] mprj_io_outen[28] mprj_io[28] mprj_io_pd_select[28] mprj_io_drive_sel[56]
+ mprj_io_drive_sel[57] mprj_io_pu_select[28] mprj_io_slew_select[28] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[28] GF_NI_BI_T
XGF_NI_BI_T_41 mprj_io_out[34] mprj_io_schmitt_select[34] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[34] mprj_io_outen[34] mprj_io[34] mprj_io_pd_select[34] mprj_io_drive_sel[68]
+ mprj_io_drive_sel[69] mprj_io_pu_select[34] mprj_io_slew_select[34] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[34] GF_NI_BI_T
XGF_NI_FILL10_289 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_201 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_212 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_223 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_234 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_245 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_256 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1026 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1015 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_267 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_278 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1004 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_790 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_5 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_608 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_619 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_449 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_438 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_427 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_416 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_405 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_950 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_961 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_972 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_983 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_994 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_20 mprj_io_out[13] mprj_io_schmitt_select[13] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[13] mprj_io_outen[13] mprj_io[12] mprj_io_pd_select[13] mprj_io_drive_sel[26]
+ mprj_io_drive_sel[27] mprj_io_pu_select[13] mprj_io_slew_select[13] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[13] GF_NI_BI_T
XGF_NI_BI_T_31 mprj_io_out[29] mprj_io_schmitt_select[29] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[29] mprj_io_outen[29] mprj_io[29] mprj_io_pd_select[29] mprj_io_drive_sel[58]
+ mprj_io_drive_sel[59] mprj_io_pu_select[29] mprj_io_slew_select[29] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[29] GF_NI_BI_T
XGF_NI_BI_T_42 mprj_io_out[36] mprj_io_schmitt_select[36] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[36] mprj_io_outen[36] mprj_io[36] mprj_io_pd_select[36] mprj_io_drive_sel[72]
+ mprj_io_drive_sel[73] mprj_io_pu_select[36] mprj_io_slew_select[36] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[36] GF_NI_BI_T
XGF_NI_FILL10_202 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_213 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_224 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_235 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_246 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_257 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_268 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_279 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_780 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_791 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_6 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_1038 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1027 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1016 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1005 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_609 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_428 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_417 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_406 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_439 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_940 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_951 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_962 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_973 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_21 mprj_io_out[20] mprj_io_schmitt_select[20] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[20] mprj_io_outen[20] mprj_io[20] mprj_io_pd_select[20] mprj_io_drive_sel[40]
+ mprj_io_drive_sel[41] mprj_io_pu_select[20] mprj_io_slew_select[20] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[20] GF_NI_BI_T
XGF_NI_BI_T_32 mprj_io_out[30] mprj_io_schmitt_select[30] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[30] mprj_io_outen[30] mprj_io[30] mprj_io_pd_select[30] mprj_io_drive_sel[63]
+ mprj_io_drive_sel[61] mprj_io_pu_select[30] mprj_io_slew_select[30] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[30] GF_NI_BI_T
XGF_NI_BI_T_10 mprj_io_out[5] mprj_io_schmitt_select[5] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[5] mprj_io_outen[5] mprj_io[5] mprj_io_pd_select[5] mprj_io_drive_sel[11]
+ mprj_io_drive_sel[10] mprj_io_pu_select[5] mprj_io_slew_select[5] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[5] GF_NI_BI_T
XGF_NI_FILL10_995 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_203 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_214 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_225 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_236 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_247 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_258 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_269 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_770 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_781 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_792 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_7 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_1039 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1028 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1017 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1006 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_429 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_418 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_407 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_22 mprj_io_out[12] mprj_io_schmitt_select[12] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[12] mprj_io_outen[12] mprj_io[13] mprj_io_pd_select[12] mprj_io_drive_sel[25]
+ mprj_io_drive_sel[24] mprj_io_pu_select[12] mprj_io_slew_select[12] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[12] GF_NI_BI_T
XGF_NI_BI_T_33 mprj_io_out[25] mprj_io_schmitt_select[25] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[25] mprj_io_outen[25] mprj_io[25] mprj_io_pd_select[25] mprj_io_drive_sel[525]
+ mprj_io_drive_sel[51] mprj_io_pu_select[25] mprj_io_slew_select[25] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[25] GF_NI_BI_T
XGF_NI_FILL10_930 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_941 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_952 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_963 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_11 mprj_io_out[6] mprj_io_schmitt_select[6] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[6] mprj_io_outen[6] mprj_io[6] mprj_io_pd_select[6] mprj_io_drive_sel[13]
+ mprj_io_drive_sel[12] mprj_io_pu_select[6] mprj_io_slew_select[6] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[6] GF_NI_BI_T
XGF_NI_FILL10_974 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_985 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_996 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_204 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_215 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_226 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_237 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_259 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_248 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_760 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_771 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_782 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_793 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_8 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_1029 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1018 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1007 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_590 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_419 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_408 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_920 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_931 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_942 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_953 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_964 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_975 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_997 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_986 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_12 mprj_io_out[18] mprj_io_schmitt_select[18] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[18] mprj_io_outen[18] mprj_io[18] mprj_io_pd_select[18] mprj_io_drive_sel[36]
+ mprj_io_drive_sel[37] mprj_io_pu_select[18] mprj_io_slew_select[18] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[18] GF_NI_BI_T
XGF_NI_BI_T_23 mprj_io_out[21] mprj_io_schmitt_select[21] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[21] mprj_io_outen[21] mprj_io[21] mprj_io_pd_select[21] mprj_io_drive_sel[42]
+ mprj_io_drive_sel[43] mprj_io_pu_select[21] mprj_io_slew_select[21] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[21] GF_NI_BI_T
XGF_NI_BI_T_34 mprj_io_out[26] mprj_io_schmitt_select[26] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[26] mprj_io_outen[26] mprj_io[26] mprj_io_pd_select[26] mprj_io_drive_sel[52]
+ mprj_io_drive_sel[53] mprj_io_pu_select[26] mprj_io_slew_select[26] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[26] GF_NI_BI_T
XGF_NI_FILL10_750 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_205 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_216 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_227 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_238 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_249 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1019 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1008 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_772 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_783 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_794 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_9 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_761 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_580 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_591 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_409 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_910 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_921 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_932 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_943 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_965 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_976 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_987 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_13 mprj_io_out[22] mprj_io_schmitt_select[22] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[22] mprj_io_outen[22] mprj_io[22] mprj_io_pd_select[22] mprj_io_drive_sel[44]
+ mprj_io_drive_sel[45] mprj_io_pu_select[22] mprj_io_slew_select[22] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[22] GF_NI_BI_T
XGF_NI_BI_T_24 mprj_io_out[14] mprj_io_schmitt_select[14] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[14] mprj_io_outen[14] mprj_io[14] mprj_io_pd_select[14] mprj_io_drive_sel[28]
+ mprj_io_drive_sel[29] mprj_io_pu_select[14] mprj_io_slew_select[14] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[14] GF_NI_BI_T
XGF_NI_BI_T_35 mprj_io_out[27] mprj_io_schmitt_select[27] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[27] mprj_io_outen[27] mprj_io[27] mprj_io_pd_select[27] mprj_io_drive_sel[54]
+ mprj_io_drive_sel[55] mprj_io_pu_select[27] mprj_io_slew_select[27] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[27] GF_NI_BI_T
XGF_NI_FILL10_206 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_217 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_228 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_239 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_1009 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_740 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_751 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_762 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_784 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_795 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_773 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_570 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_581 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_592 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_900 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_911 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_922 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_933 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_944 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_955 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_966 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_977 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_999 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_988 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_25 mprj_io_out[15] mprj_io_schmitt_select[15] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[15] mprj_io_outen[15] mprj_io[15] mprj_io_pd_select[15] mprj_io_drive_sel[30]
+ mprj_io_drive_sel[31] mprj_io_pu_select[15] mprj_io_slew_select[15] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[15] GF_NI_BI_T
XGF_NI_BI_T_14 mprj_io_out[19] mprj_io_schmitt_select[19] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[19] mprj_io_outen[19] mprj_io[19] mprj_io_pd_select[19] mprj_io_drive_sel[38]
+ mprj_io_drive_sel[39] mprj_io_pu_select[19] mprj_io_slew_select[19] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[19] GF_NI_BI_T
XGF_NI_BI_T_36 mprj_io_out[31] mprj_io_schmitt_select[31] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[31] mprj_io_outen[31] mprj_io[31] mprj_io_pd_select[31] mprj_io_drive_sel[62]
+ mprj_io_drive_sel[63] mprj_io_pu_select[31] mprj_io_slew_select[31] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[31] GF_NI_BI_T
XGF_NI_FILL10_207 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_218 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_229 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_730 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_741 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_752 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_763 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_774 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_796 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_785 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_560 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_571 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_582 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_593 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_390 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_912 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_923 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_934 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_945 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_956 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_967 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_978 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_901 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_989 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_26 mprj_io_out[16] mprj_io_schmitt_select[16] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[16] mprj_io_outen[16] mprj_io[16] mprj_io_pd_select[16] mprj_io_drive_sel[32]
+ mprj_io_drive_sel[33] mprj_io_pu_select[16] mprj_io_slew_select[16] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[16] GF_NI_BI_T
XGF_NI_BI_T_15 mprj_io_out[7] mprj_io_schmitt_select[7] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[7] mprj_io_outen[7] mprj_io[7] mprj_io_pd_select[7] mprj_io_drive_sel[15]
+ mprj_io_drive_sel[14] mprj_io_pu_select[7] mprj_io_slew_select[7] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[7] GF_NI_BI_T
XGF_NI_BI_T_37 mprj_io_out[37] mprj_io_schmitt_select[37] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[37] mprj_io_outen[37] mprj_io[37] mprj_io_pd_select[37] mprj_io_drive_sel[74]
+ mprj_io_drive_sel[75] mprj_io_pu_select[37] mprj_io_slew_select[37] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[37] GF_NI_BI_T
XGF_NI_FILL10_208 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_219 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_720 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_731 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_742 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_753 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_764 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_775 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_786 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_797 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_550 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_561 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_572 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_583 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_594 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_391 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_380 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_27 mprj_io_out[17] mprj_io_schmitt_select[17] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[17] mprj_io_outen[17] mprj_io[17] mprj_io_pd_select[17] mprj_io_drive_sel[34]
+ mprj_io_drive_sel[35] mprj_io_pu_select[17] mprj_io_slew_select[17] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[17] GF_NI_BI_T
XGF_NI_BI_T_16 mprj_io_out[8] mprj_io_schmitt_select[8] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[8] mprj_io_outen[8] mprj_io[8] mprj_io_pd_select[8] mprj_io_drive_sel[17]
+ mprj_io_drive_sel[16] mprj_io_pu_select[8] mprj_io_slew_select[8] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[8] GF_NI_BI_T
XGF_NI_FILL10_902 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_913 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_924 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_935 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_946 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_957 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_968 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_979 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_38 mprj_io_out[35] mprj_io_schmitt_select[35] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[35] mprj_io_outen[35] mprj_io[35] mprj_io_pd_select[35] mprj_io_drive_sel[70]
+ mprj_io_drive_sel[71] mprj_io_pu_select[35] mprj_io_slew_select[35] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[35] GF_NI_BI_T
XGF_NI_IN_C_0 GF_NI_COR_3/VDD GF_NI_COR_3/VSS clock GF_NI_IN_C_0/PD GF_NI_IN_C_0/PU
+ GF_NI_COR_3/VDD GF_NI_COR_3/VSS clock_core GF_NI_IN_C
XGF_NI_FILL10_209 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_710 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_721 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_732 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_743 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_754 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_765 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_776 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_787 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_798 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_540 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_551 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_562 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_573 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_584 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_595 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_392 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_381 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_370 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_COR_0 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR
XGF_NI_FILL10_903 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_914 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_936 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_947 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_958 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_925 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_28 mprj_io_out[23] mprj_io_schmitt_select[23] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[23] mprj_io_outen[23] mprj_io[23] mprj_io_pd_select[23] mprj_io_drive_sel[46]
+ mprj_io_drive_sel[47] mprj_io_pu_select[23] mprj_io_slew_select[23] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[23] GF_NI_BI_T
XGF_NI_BI_T_17 mprj_io_out[9] mprj_io_schmitt_select[9] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[9] mprj_io_outen[9] mprj_io[9] mprj_io_pd_select[9] mprj_io_drive_sel[19]
+ mprj_io_drive_sel[18] mprj_io_pu_select[9] mprj_io_slew_select[9] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[9] GF_NI_BI_T
XGF_NI_BI_T_39 mprj_io_out[32] mprj_io_schmitt_select[32] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[32] mprj_io_outen[32] mprj_io[32] mprj_io_pd_select[32] mprj_io_drive_sel[64]
+ mprj_io_drive_sel[65] mprj_io_pu_select[32] mprj_io_slew_select[32] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[32] GF_NI_BI_T
XGF_NI_FILL10_700 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_711 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_722 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_733 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_744 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_755 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_766 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_777 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_788 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_799 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_530 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_541 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_552 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_563 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_574 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_585 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_596 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_393 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_382 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_371 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_360 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_COR_1 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR
XGF_NI_FILL10_190 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_904 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_915 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_926 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_937 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_948 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_959 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_29 mprj_io_out[24] mprj_io_schmitt_select[24] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[24] mprj_io_outen[24] mprj_io[24] mprj_io_pd_select[24] mprj_io_drive_sel[48]
+ mprj_io_drive_sel[49] mprj_io_pu_select[24] mprj_io_slew_select[24] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[24] GF_NI_BI_T
XGF_NI_BI_T_18 mprj_io_out[10] mprj_io_schmitt_select[10] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[10] mprj_io_outen[10] mprj_io[10] mprj_io_pd_select[10] mprj_io_drive_sel[21]
+ mprj_io_drive_sel[20] mprj_io_pu_select[10] mprj_io_slew_select[10] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[10] GF_NI_BI_T
XGF_NI_FILL10_701 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_712 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_723 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_734 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_745 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_756 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_767 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_778 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_789 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_520 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_531 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_553 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_542 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_564 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_575 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_586 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_597 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_90 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_COR_2 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR
XGF_NI_FILL10_394 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_383 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_372 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_361 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_350 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_180 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_191 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_905 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_927 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_938 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_949 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_916 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_BI_T_19 mprj_io_out[11] mprj_io_schmitt_select[11] GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ mprj_io_inen[11] mprj_io_outen[11] mprj_io[11] mprj_io_pd_select[11] mprj_io_drive_sel[23]
+ mprj_io_drive_sel[22] mprj_io_pu_select[11] mprj_io_slew_select[11] GF_NI_COR_3/VDD
+ GF_NI_COR_3/VSS mprj_io_in[11] GF_NI_BI_T
XGF_NI_FILL10_702 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_713 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_724 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_735 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_746 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_757 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_768 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_779 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_521 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_510 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_532 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_543 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_554 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_565 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_576 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_587 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_598 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_80 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_91 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_COR_3 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR
XGF_NI_FILL10_395 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_384 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_373 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_362 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_351 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_340 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_170 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_181 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_192 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_906 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_917 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_928 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_703 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_714 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_725 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_736 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_747 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_758 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_769 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_522 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_533 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_544 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_555 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_566 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_577 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_588 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_599 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_511 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_500 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_81 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_70 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_92 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_396 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_385 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_374 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_363 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_352 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_341 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_330 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_160 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_171 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_182 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_193 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_907 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_918 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_929 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_704 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_715 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_726 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_737 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_748 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_759 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_523 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_534 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_545 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_556 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_567 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_578 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_589 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_512 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_501 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_82 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_71 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_60 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_93 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_FILL10
XGF_NI_FILL10_397 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_386 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_375 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_364 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_353 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_342 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_331 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_320 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_150 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_161 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_172 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_183 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_194 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_908 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_919 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_705 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_716 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_727 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_738 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
XGF_NI_FILL10_749 GF_NI_COR_3/VDD GF_NI_COR_3/VSS GF_NI_COR_3/VDD GF_NI_COR_3/VSS
+ GF_NI_FILL10
.ends

* Black-box entry subcircuit for mgmt_core_wrapper abstract view
.subckt mgmt_core_wrapper VDD VSS core_clk core_rstn debug_in debug_mode debug_oeb
+ debug_out flash_clk flash_csb flash_io0_di flash_io0_do flash_io0_oeb flash_io1_di
+ flash_io1_do flash_io1_oeb flash_io2_di flash_io2_do flash_io2_oeb flash_io3_di
+ flash_io3_do flash_io3_oeb gpio_in_pad gpio_inenb_pad gpio_mode0_pad gpio_mode1_pad
+ gpio_out_pad gpio_outenb_pad hk_ack_i hk_cyc_o hk_dat_i[0] hk_dat_i[10] hk_dat_i[11]
+ hk_dat_i[12] hk_dat_i[13] hk_dat_i[14] hk_dat_i[15] hk_dat_i[16] hk_dat_i[17] hk_dat_i[18]
+ hk_dat_i[19] hk_dat_i[1] hk_dat_i[20] hk_dat_i[21] hk_dat_i[22] hk_dat_i[23] hk_dat_i[24]
+ hk_dat_i[25] hk_dat_i[26] hk_dat_i[27] hk_dat_i[28] hk_dat_i[29] hk_dat_i[2] hk_dat_i[30]
+ hk_dat_i[31] hk_dat_i[3] hk_dat_i[4] hk_dat_i[5] hk_dat_i[6] hk_dat_i[7] hk_dat_i[8]
+ hk_dat_i[9] hk_stb_o irq[0] irq[1] irq[2] irq[3] irq[4] irq[5] la_iena[0] la_iena[10]
+ la_iena[11] la_iena[12] la_iena[13] la_iena[14] la_iena[15] la_iena[16] la_iena[17]
+ la_iena[18] la_iena[19] la_iena[1] la_iena[20] la_iena[21] la_iena[22] la_iena[23]
+ la_iena[24] la_iena[25] la_iena[26] la_iena[27] la_iena[28] la_iena[29] la_iena[2]
+ la_iena[30] la_iena[31] la_iena[32] la_iena[33] la_iena[34] la_iena[35] la_iena[36]
+ la_iena[37] la_iena[38] la_iena[39] la_iena[3] la_iena[40] la_iena[41] la_iena[42]
+ la_iena[43] la_iena[44] la_iena[45] la_iena[46] la_iena[47] la_iena[48] la_iena[49]
+ la_iena[4] la_iena[50] la_iena[51] la_iena[52] la_iena[53] la_iena[54] la_iena[55]
+ la_iena[56] la_iena[57] la_iena[58] la_iena[59] la_iena[5] la_iena[60] la_iena[61]
+ la_iena[62] la_iena[63] la_iena[6] la_iena[7] la_iena[8] la_iena[9] la_input[0]
+ la_input[10] la_input[11] la_input[12] la_input[13] la_input[14] la_input[15] la_input[16]
+ la_input[17] la_input[18] la_input[19] la_input[1] la_input[20] la_input[21] la_input[22]
+ la_input[23] la_input[24] la_input[25] la_input[26] la_input[27] la_input[28] la_input[29]
+ la_input[2] la_input[30] la_input[31] la_input[32] la_input[33] la_input[34] la_input[35]
+ la_input[36] la_input[37] la_input[38] la_input[39] la_input[3] la_input[40] la_input[41]
+ la_input[42] la_input[43] la_input[44] la_input[45] la_input[46] la_input[47] la_input[48]
+ la_input[49] la_input[4] la_input[50] la_input[51] la_input[52] la_input[53] la_input[54]
+ la_input[55] la_input[56] la_input[57] la_input[58] la_input[59] la_input[5] la_input[60]
+ la_input[61] la_input[62] la_input[63] la_input[6] la_input[7] la_input[8] la_input[9]
+ la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15]
+ la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21]
+ la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28]
+ la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34]
+ la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40]
+ la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47]
+ la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53]
+ la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5]
+ la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7] la_oenb[8]
+ la_oenb[9] la_output[0] la_output[10] la_output[11] la_output[12] la_output[13]
+ la_output[14] la_output[15] la_output[16] la_output[17] la_output[18] la_output[19]
+ la_output[1] la_output[20] la_output[21] la_output[22] la_output[23] la_output[24]
+ la_output[25] la_output[26] la_output[27] la_output[28] la_output[29] la_output[2]
+ la_output[30] la_output[31] la_output[32] la_output[33] la_output[34] la_output[35]
+ la_output[36] la_output[37] la_output[38] la_output[39] la_output[3] la_output[40]
+ la_output[41] la_output[42] la_output[43] la_output[44] la_output[45] la_output[46]
+ la_output[47] la_output[48] la_output[49] la_output[4] la_output[50] la_output[51]
+ la_output[52] la_output[53] la_output[54] la_output[55] la_output[56] la_output[57]
+ la_output[58] la_output[59] la_output[5] la_output[60] la_output[61] la_output[62]
+ la_output[63] la_output[6] la_output[7] la_output[8] la_output[9] mprj_ack_i mprj_adr_o[0]
+ mprj_adr_o[10] mprj_adr_o[11] mprj_adr_o[12] mprj_adr_o[13] mprj_adr_o[14] mprj_adr_o[15]
+ mprj_adr_o[16] mprj_adr_o[17] mprj_adr_o[18] mprj_adr_o[19] mprj_adr_o[1] mprj_adr_o[20]
+ mprj_adr_o[21] mprj_adr_o[22] mprj_adr_o[23] mprj_adr_o[24] mprj_adr_o[25] mprj_adr_o[26]
+ mprj_adr_o[27] mprj_adr_o[28] mprj_adr_o[29] mprj_adr_o[2] mprj_adr_o[30] mprj_adr_o[31]
+ mprj_adr_o[3] mprj_adr_o[4] mprj_adr_o[5] mprj_adr_o[6] mprj_adr_o[7] mprj_adr_o[8]
+ mprj_adr_o[9] mprj_cyc_o mprj_dat_i[0] mprj_dat_i[10] mprj_dat_i[11] mprj_dat_i[12]
+ mprj_dat_i[13] mprj_dat_i[14] mprj_dat_i[15] mprj_dat_i[16] mprj_dat_i[17] mprj_dat_i[18]
+ mprj_dat_i[19] mprj_dat_i[1] mprj_dat_i[20] mprj_dat_i[21] mprj_dat_i[22] mprj_dat_i[23]
+ mprj_dat_i[24] mprj_dat_i[25] mprj_dat_i[26] mprj_dat_i[27] mprj_dat_i[28] mprj_dat_i[29]
+ mprj_dat_i[2] mprj_dat_i[30] mprj_dat_i[31] mprj_dat_i[3] mprj_dat_i[4] mprj_dat_i[5]
+ mprj_dat_i[6] mprj_dat_i[7] mprj_dat_i[8] mprj_dat_i[9] mprj_dat_o[0] mprj_dat_o[10]
+ mprj_dat_o[11] mprj_dat_o[12] mprj_dat_o[13] mprj_dat_o[14] mprj_dat_o[15] mprj_dat_o[16]
+ mprj_dat_o[17] mprj_dat_o[18] mprj_dat_o[19] mprj_dat_o[1] mprj_dat_o[20] mprj_dat_o[21]
+ mprj_dat_o[22] mprj_dat_o[23] mprj_dat_o[24] mprj_dat_o[25] mprj_dat_o[26] mprj_dat_o[27]
+ mprj_dat_o[28] mprj_dat_o[29] mprj_dat_o[2] mprj_dat_o[30] mprj_dat_o[31] mprj_dat_o[3]
+ mprj_dat_o[4] mprj_dat_o[5] mprj_dat_o[6] mprj_dat_o[7] mprj_dat_o[8] mprj_dat_o[9]
+ mprj_sel_o[0] mprj_sel_o[1] mprj_sel_o[2] mprj_sel_o[3] mprj_stb_o mprj_wb_iena
+ mprj_we_o qspi_enabled ser_rx ser_tx spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb trap uart_enabled user_irq_ena[0] user_irq_ena[1] user_irq_ena[2]
.ends

* Black-box entry subcircuit for simple_por abstract view
.subckt simple_por vdd vss porb por
.ends

* Black-box entry subcircuit for caravel_clocking abstract view
.subckt caravel_clocking VDD VSS core_clk ext_clk ext_clk_sel ext_reset pll_clk pll_clk90
+ resetb resetb_sync sel2[0] sel2[1] sel2[2] sel[0] sel[1] sel[2] user_clk
.ends

* Black-box entry subcircuit for spare_logic_block abstract view
.subckt spare_logic_block VDD VSS spare_xfq[0] spare_xfq[1] spare_xi[0] spare_xi[1]
+ spare_xi[2] spare_xi[3] spare_xib spare_xmx[0] spare_xmx[1] spare_xna[0] spare_xna[1]
+ spare_xno[0] spare_xno[1] spare_xz[0] spare_xz[10] spare_xz[11] spare_xz[12] spare_xz[13]
+ spare_xz[14] spare_xz[15] spare_xz[16] spare_xz[17] spare_xz[18] spare_xz[19] spare_xz[1]
+ spare_xz[20] spare_xz[21] spare_xz[22] spare_xz[23] spare_xz[24] spare_xz[25] spare_xz[26]
+ spare_xz[27] spare_xz[28] spare_xz[29] spare_xz[2] spare_xz[30] spare_xz[3] spare_xz[4]
+ spare_xz[5] spare_xz[6] spare_xz[7] spare_xz[8] spare_xz[9]
.ends

* Black-box entry subcircuit for user_id_programming abstract view
.subckt user_id_programming mask_rev[0] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[13]
+ mask_rev[14] mask_rev[15] mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[1]
+ mask_rev[20] mask_rev[21] mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26]
+ mask_rev[27] mask_rev[28] mask_rev[29] mask_rev[2] mask_rev[30] mask_rev[31] mask_rev[3]
+ mask_rev[4] mask_rev[5] mask_rev[6] mask_rev[7] mask_rev[8] mask_rev[9] VDD VSS
.ends

* Black-box entry subcircuit for mgmt_protect abstract view
.subckt mgmt_protect VDD VSS caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0]
+ la_data_in_core[10] la_data_in_core[11] la_data_in_core[12] la_data_in_core[13]
+ la_data_in_core[14] la_data_in_core[15] la_data_in_core[16] la_data_in_core[17]
+ la_data_in_core[18] la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21]
+ la_data_in_core[22] la_data_in_core[23] la_data_in_core[24] la_data_in_core[25]
+ la_data_in_core[26] la_data_in_core[27] la_data_in_core[28] la_data_in_core[29]
+ la_data_in_core[2] la_data_in_core[30] la_data_in_core[31] la_data_in_core[32] la_data_in_core[33]
+ la_data_in_core[34] la_data_in_core[35] la_data_in_core[36] la_data_in_core[37]
+ la_data_in_core[38] la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41]
+ la_data_in_core[42] la_data_in_core[43] la_data_in_core[44] la_data_in_core[45]
+ la_data_in_core[46] la_data_in_core[47] la_data_in_core[48] la_data_in_core[49]
+ la_data_in_core[4] la_data_in_core[50] la_data_in_core[51] la_data_in_core[52] la_data_in_core[53]
+ la_data_in_core[54] la_data_in_core[55] la_data_in_core[56] la_data_in_core[57]
+ la_data_in_core[58] la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61]
+ la_data_in_core[62] la_data_in_core[63] la_data_in_core[6] la_data_in_core[7] la_data_in_core[8]
+ la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[10] la_data_in_mprj[11] la_data_in_mprj[12]
+ la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15] la_data_in_mprj[16]
+ la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19] la_data_in_mprj[1] la_data_in_mprj[20]
+ la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23] la_data_in_mprj[24]
+ la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27] la_data_in_mprj[28]
+ la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31] la_data_in_mprj[32]
+ la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35] la_data_in_mprj[36]
+ la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39] la_data_in_mprj[3] la_data_in_mprj[40]
+ la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43] la_data_in_mprj[44]
+ la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47] la_data_in_mprj[48]
+ la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51] la_data_in_mprj[52]
+ la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55] la_data_in_mprj[56]
+ la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59] la_data_in_mprj[5] la_data_in_mprj[60]
+ la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63] la_data_in_mprj[6] la_data_in_mprj[7]
+ la_data_in_mprj[8] la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[10] la_data_out_core[11]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[6] la_data_out_core[7] la_data_out_core[8]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[10] la_data_out_mprj[11]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[6] la_data_out_mprj[7] la_data_out_mprj[8]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[10] la_iena_mprj[11] la_iena_mprj[12]
+ la_iena_mprj[13] la_iena_mprj[14] la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17]
+ la_iena_mprj[18] la_iena_mprj[19] la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21]
+ la_iena_mprj[22] la_iena_mprj[23] la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26]
+ la_iena_mprj[27] la_iena_mprj[28] la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30]
+ la_iena_mprj[31] la_iena_mprj[32] la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35]
+ la_iena_mprj[36] la_iena_mprj[37] la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3]
+ la_iena_mprj[40] la_iena_mprj[41] la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44]
+ la_iena_mprj[45] la_iena_mprj[46] la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49]
+ la_iena_mprj[4] la_iena_mprj[50] la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53]
+ la_iena_mprj[54] la_iena_mprj[55] la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58]
+ la_iena_mprj[59] la_iena_mprj[5] la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62]
+ la_iena_mprj[63] la_iena_mprj[6] la_iena_mprj[7] la_iena_mprj[8] la_iena_mprj[9]
+ la_oenb_core[0] la_oenb_core[10] la_oenb_core[11] la_oenb_core[12] la_oenb_core[13]
+ la_oenb_core[14] la_oenb_core[15] la_oenb_core[16] la_oenb_core[17] la_oenb_core[18]
+ la_oenb_core[19] la_oenb_core[1] la_oenb_core[20] la_oenb_core[21] la_oenb_core[22]
+ la_oenb_core[23] la_oenb_core[24] la_oenb_core[25] la_oenb_core[26] la_oenb_core[27]
+ la_oenb_core[28] la_oenb_core[29] la_oenb_core[2] la_oenb_core[30] la_oenb_core[31]
+ la_oenb_core[32] la_oenb_core[33] la_oenb_core[34] la_oenb_core[35] la_oenb_core[36]
+ la_oenb_core[37] la_oenb_core[38] la_oenb_core[39] la_oenb_core[3] la_oenb_core[40]
+ la_oenb_core[41] la_oenb_core[42] la_oenb_core[43] la_oenb_core[44] la_oenb_core[45]
+ la_oenb_core[46] la_oenb_core[47] la_oenb_core[48] la_oenb_core[49] la_oenb_core[4]
+ la_oenb_core[50] la_oenb_core[51] la_oenb_core[52] la_oenb_core[53] la_oenb_core[54]
+ la_oenb_core[55] la_oenb_core[56] la_oenb_core[57] la_oenb_core[58] la_oenb_core[59]
+ la_oenb_core[5] la_oenb_core[60] la_oenb_core[61] la_oenb_core[62] la_oenb_core[63]
+ la_oenb_core[6] la_oenb_core[7] la_oenb_core[8] la_oenb_core[9] la_oenb_mprj[0]
+ la_oenb_mprj[10] la_oenb_mprj[11] la_oenb_mprj[12] la_oenb_mprj[13] la_oenb_mprj[14]
+ la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18] la_oenb_mprj[19]
+ la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22] la_oenb_mprj[23]
+ la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27] la_oenb_mprj[28]
+ la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31] la_oenb_mprj[32]
+ la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36] la_oenb_mprj[37]
+ la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40] la_oenb_mprj[41]
+ la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45] la_oenb_mprj[46]
+ la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4] la_oenb_mprj[50]
+ la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54] la_oenb_mprj[55]
+ la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59] la_oenb_mprj[5]
+ la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63] la_oenb_mprj[6]
+ la_oenb_mprj[7] la_oenb_mprj[8] la_oenb_mprj[9] mprj_ack_i_core mprj_ack_i_user
+ mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11] mprj_adr_o_core[12] mprj_adr_o_core[13]
+ mprj_adr_o_core[14] mprj_adr_o_core[15] mprj_adr_o_core[16] mprj_adr_o_core[17]
+ mprj_adr_o_core[18] mprj_adr_o_core[19] mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21]
+ mprj_adr_o_core[22] mprj_adr_o_core[23] mprj_adr_o_core[24] mprj_adr_o_core[25]
+ mprj_adr_o_core[26] mprj_adr_o_core[27] mprj_adr_o_core[28] mprj_adr_o_core[29]
+ mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31] mprj_adr_o_core[3] mprj_adr_o_core[4]
+ mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7] mprj_adr_o_core[8] mprj_adr_o_core[9]
+ mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11] mprj_adr_o_user[12] mprj_adr_o_user[13]
+ mprj_adr_o_user[14] mprj_adr_o_user[15] mprj_adr_o_user[16] mprj_adr_o_user[17]
+ mprj_adr_o_user[18] mprj_adr_o_user[19] mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21]
+ mprj_adr_o_user[22] mprj_adr_o_user[23] mprj_adr_o_user[24] mprj_adr_o_user[25]
+ mprj_adr_o_user[26] mprj_adr_o_user[27] mprj_adr_o_user[28] mprj_adr_o_user[29]
+ mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31] mprj_adr_o_user[3] mprj_adr_o_user[4]
+ mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7] mprj_adr_o_user[8] mprj_adr_o_user[9]
+ mprj_cyc_o_core mprj_cyc_o_user mprj_dat_i_core[0] mprj_dat_i_core[10] mprj_dat_i_core[11]
+ mprj_dat_i_core[12] mprj_dat_i_core[13] mprj_dat_i_core[14] mprj_dat_i_core[15]
+ mprj_dat_i_core[16] mprj_dat_i_core[17] mprj_dat_i_core[18] mprj_dat_i_core[19]
+ mprj_dat_i_core[1] mprj_dat_i_core[20] mprj_dat_i_core[21] mprj_dat_i_core[22] mprj_dat_i_core[23]
+ mprj_dat_i_core[24] mprj_dat_i_core[25] mprj_dat_i_core[26] mprj_dat_i_core[27]
+ mprj_dat_i_core[28] mprj_dat_i_core[29] mprj_dat_i_core[2] mprj_dat_i_core[30] mprj_dat_i_core[31]
+ mprj_dat_i_core[3] mprj_dat_i_core[4] mprj_dat_i_core[5] mprj_dat_i_core[6] mprj_dat_i_core[7]
+ mprj_dat_i_core[8] mprj_dat_i_core[9] mprj_dat_i_user[0] mprj_dat_i_user[10] mprj_dat_i_user[11]
+ mprj_dat_i_user[12] mprj_dat_i_user[13] mprj_dat_i_user[14] mprj_dat_i_user[15]
+ mprj_dat_i_user[16] mprj_dat_i_user[17] mprj_dat_i_user[18] mprj_dat_i_user[19]
+ mprj_dat_i_user[1] mprj_dat_i_user[20] mprj_dat_i_user[21] mprj_dat_i_user[22] mprj_dat_i_user[23]
+ mprj_dat_i_user[24] mprj_dat_i_user[25] mprj_dat_i_user[26] mprj_dat_i_user[27]
+ mprj_dat_i_user[28] mprj_dat_i_user[29] mprj_dat_i_user[2] mprj_dat_i_user[30] mprj_dat_i_user[31]
+ mprj_dat_i_user[3] mprj_dat_i_user[4] mprj_dat_i_user[5] mprj_dat_i_user[6] mprj_dat_i_user[7]
+ mprj_dat_i_user[8] mprj_dat_i_user[9] mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11]
+ mprj_dat_o_core[12] mprj_dat_o_core[13] mprj_dat_o_core[14] mprj_dat_o_core[15]
+ mprj_dat_o_core[16] mprj_dat_o_core[17] mprj_dat_o_core[18] mprj_dat_o_core[19]
+ mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21] mprj_dat_o_core[22] mprj_dat_o_core[23]
+ mprj_dat_o_core[24] mprj_dat_o_core[25] mprj_dat_o_core[26] mprj_dat_o_core[27]
+ mprj_dat_o_core[28] mprj_dat_o_core[29] mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31]
+ mprj_dat_o_core[3] mprj_dat_o_core[4] mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7]
+ mprj_dat_o_core[8] mprj_dat_o_core[9] mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11]
+ mprj_dat_o_user[12] mprj_dat_o_user[13] mprj_dat_o_user[14] mprj_dat_o_user[15]
+ mprj_dat_o_user[16] mprj_dat_o_user[17] mprj_dat_o_user[18] mprj_dat_o_user[19]
+ mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21] mprj_dat_o_user[22] mprj_dat_o_user[23]
+ mprj_dat_o_user[24] mprj_dat_o_user[25] mprj_dat_o_user[26] mprj_dat_o_user[27]
+ mprj_dat_o_user[28] mprj_dat_o_user[29] mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31]
+ mprj_dat_o_user[3] mprj_dat_o_user[4] mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7]
+ mprj_dat_o_user[8] mprj_dat_o_user[9] mprj_iena_wb mprj_sel_o_core[0] mprj_sel_o_core[1]
+ mprj_sel_o_core[2] mprj_sel_o_core[3] mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2]
+ mprj_sel_o_user[3] mprj_stb_o_core mprj_stb_o_user mprj_we_o_core mprj_we_o_user
+ user_clock user_clock2 user_irq[0] user_irq[1] user_irq[2] user_irq_core[0] user_irq_core[1]
+ user_irq_core[2] user_irq_ena[0] user_irq_ena[1] user_irq_ena[2] user_reset
.ends

* Black-box entry subcircuit for gpio_defaults_block_009 abstract view
.subckt gpio_defaults_block_009 gpio_defaults[0] gpio_defaults[1] gpio_defaults[2]
+ gpio_defaults[3] gpio_defaults[4] gpio_defaults[5] gpio_defaults[6] gpio_defaults[7]
+ gpio_defaults[8] gpio_defaults[9] VDD VSS
.ends

* Black-box entry subcircuit for gpio_defaults_block_007 abstract view
.subckt gpio_defaults_block_007 gpio_defaults[0] gpio_defaults[1] gpio_defaults[2]
+ gpio_defaults[3] gpio_defaults[4] gpio_defaults[5] gpio_defaults[6] gpio_defaults[7]
+ gpio_defaults[8] gpio_defaults[9] VDD VSS
.ends

* Black-box entry subcircuit for user_project_wrapper abstract view
.subckt user_project_wrapper io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
.ends

* Black-box entry subcircuit for housekeeping abstract view
.subckt housekeeping VDD VSS debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oe
+ pad_flash_csb pad_flash_csb_oe pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ie
+ pad_flash_io0_oe pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ie pad_flash_io1_oe
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out qspi_enabled reset
+ ser_rx ser_tx serial_clock serial_data_1 serial_data_2 serial_load serial_resetn
+ spi_csb spi_enabled spi_sck spi_sdi spi_sdo spi_sdoenb spimemio_flash_clk spimemio_flash_csb
+ spimemio_flash_io0_di spimemio_flash_io0_do spimemio_flash_io0_oeb spimemio_flash_io1_di
+ spimemio_flash_io1_do spimemio_flash_io1_oeb spimemio_flash_io2_di spimemio_flash_io2_do
+ spimemio_flash_io2_oeb spimemio_flash_io3_di spimemio_flash_io3_do spimemio_flash_io3_oeb
+ trap uart_enabled user_clock wb_ack_o wb_adr_i[0] wb_adr_i[10] wb_adr_i[11] wb_adr_i[12]
+ wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17] wb_adr_i[18] wb_adr_i[19]
+ wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23] wb_adr_i[24] wb_adr_i[25]
+ wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2] wb_adr_i[30] wb_adr_i[31]
+ wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7] wb_adr_i[8] wb_adr_i[9]
+ wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11] wb_dat_i[12] wb_dat_i[13]
+ wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18] wb_dat_i[19] wb_dat_i[1]
+ wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24] wb_dat_i[25] wb_dat_i[26]
+ wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30] wb_dat_i[31] wb_dat_i[3]
+ wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8] wb_dat_i[9] wb_dat_o[0]
+ wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14] wb_dat_o[15] wb_dat_o[16]
+ wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20] wb_dat_o[21] wb_dat_o[22]
+ wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27] wb_dat_o[28] wb_dat_o[29]
+ wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4] wb_dat_o[5] wb_dat_o[6]
+ wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0] wb_sel_i[1] wb_sel_i[2]
+ wb_sel_i[3] wb_stb_i wb_we_i
.ends

.subckt caravel clock flash_clk flash_csb flash_io0 flash_io1 gpio mprj_io[0] mprj_io[10]
+ mprj_io[11] mprj_io[12] mprj_io[13] mprj_io[14] mprj_io[15] mprj_io[16] mprj_io[17]
+ mprj_io[18] mprj_io[19] mprj_io[1] mprj_io[20] mprj_io[21] mprj_io[22] mprj_io[23]
+ mprj_io[24] mprj_io[25] mprj_io[26] mprj_io[27] mprj_io[28] mprj_io[29] mprj_io[2]
+ mprj_io[30] mprj_io[31] mprj_io[32] mprj_io[33] mprj_io[34] mprj_io[35] mprj_io[36]
+ mprj_io[37] mprj_io[3] mprj_io[4] mprj_io[5] mprj_io[6] mprj_io[7] mprj_io[8] mprj_io[9]
+ resetb vdd vss
Xgpio_control_in_2\[0\] soc/VDD soc/VSS gpio_defaults_block_6/gpio_defaults[0] gpio_defaults_block_6/gpio_defaults[1]
+ gpio_defaults_block_6/gpio_defaults[2] gpio_defaults_block_6/gpio_defaults[3] gpio_defaults_block_6/gpio_defaults[4]
+ gpio_defaults_block_6/gpio_defaults[5] gpio_defaults_block_6/gpio_defaults[6] gpio_defaults_block_6/gpio_defaults[7]
+ gpio_defaults_block_6/gpio_defaults[8] gpio_defaults_block_6/gpio_defaults[9] housekeeping/mgmt_gpio_in[19]
+ gpio_control_in_2\[0\]/zero housekeeping/mgmt_gpio_out[19] gpio_control_in_2\[0\]/one
+ padframe/mprj_io_drive_sel[38] padframe/mprj_io_drive_sel[39] padframe/mprj_io_in[19]
+ padframe/mprj_io_inen[19] padframe/mprj_io_out[19] padframe/mprj_io_outen[19] padframe/mprj_io_pd_select[19]
+ padframe/mprj_io_pu_select[19] padframe/mprj_io_schmitt_select[19] padframe/mprj_io_slew_select[19]
+ gpio_control_in_2\[0\]/resetn gpio_control_in_2\[0\]/resetn_out gpio_control_in_2\[0\]/serial_clock
+ gpio_control_in_2\[0\]/serial_clock_out gpio_control_in_2\[0\]/serial_data_in gpio_control_in_2\[0\]/serial_data_out
+ gpio_control_in_2\[0\]/serial_load gpio_control_in_2\[0\]/serial_load_out mprj/io_in[19]
+ mprj/io_oeb[19] mprj/io_out[19] gpio_control_in_2\[0\]/zero gpio_control_block
Xgpio_defaults_block_11 gpio_defaults_block_11/gpio_defaults[0] gpio_defaults_block_11/gpio_defaults[1]
+ gpio_defaults_block_11/gpio_defaults[2] gpio_defaults_block_11/gpio_defaults[3]
+ gpio_defaults_block_11/gpio_defaults[4] gpio_defaults_block_11/gpio_defaults[5]
+ gpio_defaults_block_11/gpio_defaults[6] gpio_defaults_block_11/gpio_defaults[7]
+ gpio_defaults_block_11/gpio_defaults[8] gpio_defaults_block_11/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_22 gpio_defaults_block_22/gpio_defaults[0] gpio_defaults_block_22/gpio_defaults[1]
+ gpio_defaults_block_22/gpio_defaults[2] gpio_defaults_block_22/gpio_defaults[3]
+ gpio_defaults_block_22/gpio_defaults[4] gpio_defaults_block_22/gpio_defaults[5]
+ gpio_defaults_block_22/gpio_defaults[6] gpio_defaults_block_22/gpio_defaults[7]
+ gpio_defaults_block_22/gpio_defaults[8] gpio_defaults_block_22/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_in_1\[6\] soc/VDD soc/VSS gpio_defaults_block_1/gpio_defaults[0] gpio_defaults_block_1/gpio_defaults[1]
+ gpio_defaults_block_1/gpio_defaults[2] gpio_defaults_block_1/gpio_defaults[3] gpio_defaults_block_1/gpio_defaults[4]
+ gpio_defaults_block_1/gpio_defaults[5] gpio_defaults_block_1/gpio_defaults[6] gpio_defaults_block_1/gpio_defaults[7]
+ gpio_defaults_block_1/gpio_defaults[8] gpio_defaults_block_1/gpio_defaults[9] housekeeping/mgmt_gpio_in[14]
+ gpio_control_in_1\[6\]/zero housekeeping/mgmt_gpio_out[14] gpio_control_in_1\[6\]/one
+ padframe/mprj_io_drive_sel[28] padframe/mprj_io_drive_sel[29] padframe/mprj_io_in[14]
+ padframe/mprj_io_inen[14] padframe/mprj_io_out[14] padframe/mprj_io_outen[14] padframe/mprj_io_pd_select[14]
+ padframe/mprj_io_pu_select[14] padframe/mprj_io_schmitt_select[14] padframe/mprj_io_slew_select[14]
+ gpio_control_in_1\[6\]/resetn gpio_control_in_1\[7\]/resetn gpio_control_in_1\[6\]/serial_clock
+ gpio_control_in_1\[7\]/serial_clock gpio_control_in_1\[6\]/serial_data_in gpio_control_in_1\[7\]/serial_data_in
+ gpio_control_in_1\[6\]/serial_load gpio_control_in_1\[7\]/serial_load mprj/io_in[14]
+ mprj/io_oeb[14] mprj/io_out[14] gpio_control_in_1\[6\]/zero gpio_control_block
Xgpio_defaults_block_12 gpio_defaults_block_12/gpio_defaults[0] gpio_defaults_block_12/gpio_defaults[1]
+ gpio_defaults_block_12/gpio_defaults[2] gpio_defaults_block_12/gpio_defaults[3]
+ gpio_defaults_block_12/gpio_defaults[4] gpio_defaults_block_12/gpio_defaults[5]
+ gpio_defaults_block_12/gpio_defaults[6] gpio_defaults_block_12/gpio_defaults[7]
+ gpio_defaults_block_12/gpio_defaults[8] gpio_defaults_block_12/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_23 gpio_defaults_block_23/gpio_defaults[0] gpio_defaults_block_23/gpio_defaults[1]
+ gpio_defaults_block_23/gpio_defaults[2] gpio_defaults_block_23/gpio_defaults[3]
+ gpio_defaults_block_23/gpio_defaults[4] gpio_defaults_block_23/gpio_defaults[5]
+ gpio_defaults_block_23/gpio_defaults[6] gpio_defaults_block_23/gpio_defaults[7]
+ gpio_defaults_block_23/gpio_defaults[8] gpio_defaults_block_23/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xpll soc/VDD soc/VSS pll/clockp[0] pll/clockp[1] pll/dco pll/div[0] pll/div[1] pll/div[2]
+ pll/div[3] pll/div[4] pll/enable pll/ext_trim[0] pll/ext_trim[10] pll/ext_trim[11]
+ pll/ext_trim[12] pll/ext_trim[13] pll/ext_trim[14] pll/ext_trim[15] pll/ext_trim[16]
+ pll/ext_trim[17] pll/ext_trim[18] pll/ext_trim[19] pll/ext_trim[1] pll/ext_trim[20]
+ pll/ext_trim[21] pll/ext_trim[22] pll/ext_trim[23] pll/ext_trim[24] pll/ext_trim[25]
+ pll/ext_trim[2] pll/ext_trim[3] pll/ext_trim[4] pll/ext_trim[5] pll/ext_trim[6]
+ pll/ext_trim[7] pll/ext_trim[8] pll/ext_trim[9] pll/osc pll/resetb digital_pll
Xpadframe clock pll/osc flash_clk padframe/flash_clk_core padframe/flash_clk_oe_core
+ flash_csb padframe/flash_csb_core padframe/flash_csb_oe_core flash_io0 padframe/flash_io0_di_core
+ padframe/flash_io0_do_core padframe/flash_io0_ie_core padframe/flash_io0_oe_core
+ flash_io1 padframe/flash_io1_di_core padframe/flash_io1_do_core padframe/flash_io1_ie_core
+ padframe/flash_io1_oe_core gpio soc/gpio_mode0_pad soc/gpio_mode1_pad soc/gpio_in_pad
+ soc/gpio_inenb_pad soc/gpio_out_pad soc/gpio_outenb_pad padframe/gpio_pd_select
+ padframe/gpio_pu_select padframe/gpio_schmitt_select padframe/gpio_slew_select mprj_io[0]
+ mprj_io[10] mprj_io[11] mprj_io[12] mprj_io[13] mprj_io[14] mprj_io[15] mprj_io[16]
+ mprj_io[17] mprj_io[18] mprj_io[19] mprj_io[1] mprj_io[20] mprj_io[21] mprj_io[22]
+ mprj_io[23] mprj_io[24] mprj_io[25] mprj_io[26] mprj_io[27] mprj_io[28] mprj_io[29]
+ mprj_io[2] mprj_io[30] mprj_io[31] mprj_io[32] mprj_io[33] mprj_io[34] mprj_io[35]
+ mprj_io[36] mprj_io[37] mprj_io[3] mprj_io[4] mprj_io[5] mprj_io[6] mprj_io[7] mprj_io[8]
+ mprj_io[9] padframe/mprj_io_drive_sel[0] padframe/mprj_io_drive_sel[10] padframe/mprj_io_drive_sel[11]
+ padframe/mprj_io_drive_sel[12] padframe/mprj_io_drive_sel[13] padframe/mprj_io_drive_sel[14]
+ padframe/mprj_io_drive_sel[15] padframe/mprj_io_drive_sel[16] padframe/mprj_io_drive_sel[17]
+ padframe/mprj_io_drive_sel[18] padframe/mprj_io_drive_sel[19] padframe/mprj_io_drive_sel[1]
+ padframe/mprj_io_drive_sel[20] padframe/mprj_io_drive_sel[21] padframe/mprj_io_drive_sel[22]
+ padframe/mprj_io_drive_sel[23] padframe/mprj_io_drive_sel[24] padframe/mprj_io_drive_sel[25]
+ padframe/mprj_io_drive_sel[26] padframe/mprj_io_drive_sel[27] padframe/mprj_io_drive_sel[28]
+ padframe/mprj_io_drive_sel[29] padframe/mprj_io_drive_sel[2] padframe/mprj_io_drive_sel[30]
+ padframe/mprj_io_drive_sel[31] padframe/mprj_io_drive_sel[32] padframe/mprj_io_drive_sel[33]
+ padframe/mprj_io_drive_sel[34] padframe/mprj_io_drive_sel[35] padframe/mprj_io_drive_sel[36]
+ padframe/mprj_io_drive_sel[37] padframe/mprj_io_drive_sel[38] padframe/mprj_io_drive_sel[39]
+ padframe/mprj_io_drive_sel[3] padframe/mprj_io_drive_sel[40] padframe/mprj_io_drive_sel[41]
+ padframe/mprj_io_drive_sel[42] padframe/mprj_io_drive_sel[43] padframe/mprj_io_drive_sel[44]
+ padframe/mprj_io_drive_sel[45] padframe/mprj_io_drive_sel[46] padframe/mprj_io_drive_sel[47]
+ padframe/mprj_io_drive_sel[48] padframe/mprj_io_drive_sel[49] padframe/mprj_io_drive_sel[4]
+ padframe/mprj_io_drive_sel[51] padframe/mprj_io_drive_sel[525] padframe/mprj_io_drive_sel[52]
+ padframe/mprj_io_drive_sel[53] padframe/mprj_io_drive_sel[54] padframe/mprj_io_drive_sel[55]
+ padframe/mprj_io_drive_sel[56] padframe/mprj_io_drive_sel[57] padframe/mprj_io_drive_sel[58]
+ padframe/mprj_io_drive_sel[59] padframe/mprj_io_drive_sel[5] padframe/mprj_io_drive_sel[61]
+ padframe/mprj_io_drive_sel[62] padframe/mprj_io_drive_sel[63] padframe/mprj_io_drive_sel[64]
+ padframe/mprj_io_drive_sel[65] padframe/mprj_io_drive_sel[66] padframe/mprj_io_drive_sel[67]
+ padframe/mprj_io_drive_sel[68] padframe/mprj_io_drive_sel[69] padframe/mprj_io_drive_sel[6]
+ padframe/mprj_io_drive_sel[70] padframe/mprj_io_drive_sel[71] padframe/mprj_io_drive_sel[72]
+ padframe/mprj_io_drive_sel[73] padframe/mprj_io_drive_sel[74] padframe/mprj_io_drive_sel[75]
+ padframe/mprj_io_drive_sel[7] padframe/mprj_io_drive_sel[8] padframe/mprj_io_drive_sel[9]
+ padframe/mprj_io_in[0] padframe/mprj_io_in[10] padframe/mprj_io_in[11] padframe/mprj_io_in[12]
+ padframe/mprj_io_in[13] padframe/mprj_io_in[14] padframe/mprj_io_in[15] padframe/mprj_io_in[16]
+ padframe/mprj_io_in[17] padframe/mprj_io_in[18] padframe/mprj_io_in[19] padframe/mprj_io_in[1]
+ padframe/mprj_io_in[20] padframe/mprj_io_in[21] padframe/mprj_io_in[22] padframe/mprj_io_in[23]
+ padframe/mprj_io_in[24] padframe/mprj_io_in[25] padframe/mprj_io_in[26] padframe/mprj_io_in[27]
+ padframe/mprj_io_in[28] padframe/mprj_io_in[29] padframe/mprj_io_in[2] padframe/mprj_io_in[30]
+ padframe/mprj_io_in[31] padframe/mprj_io_in[32] padframe/mprj_io_in[33] padframe/mprj_io_in[34]
+ padframe/mprj_io_in[35] padframe/mprj_io_in[36] padframe/mprj_io_in[37] padframe/mprj_io_in[3]
+ padframe/mprj_io_in[4] padframe/mprj_io_in[5] padframe/mprj_io_in[6] padframe/mprj_io_in[7]
+ padframe/mprj_io_in[8] padframe/mprj_io_in[9] padframe/mprj_io_inen[0] padframe/mprj_io_inen[10]
+ padframe/mprj_io_inen[11] padframe/mprj_io_inen[12] padframe/mprj_io_inen[13] padframe/mprj_io_inen[14]
+ padframe/mprj_io_inen[15] padframe/mprj_io_inen[16] padframe/mprj_io_inen[17] padframe/mprj_io_inen[18]
+ padframe/mprj_io_inen[19] padframe/mprj_io_inen[1] padframe/mprj_io_inen[20] padframe/mprj_io_inen[21]
+ padframe/mprj_io_inen[22] padframe/mprj_io_inen[23] padframe/mprj_io_inen[24] padframe/mprj_io_inen[25]
+ padframe/mprj_io_inen[26] padframe/mprj_io_inen[27] padframe/mprj_io_inen[28] padframe/mprj_io_inen[29]
+ padframe/mprj_io_inen[2] padframe/mprj_io_inen[30] padframe/mprj_io_inen[31] padframe/mprj_io_inen[32]
+ padframe/mprj_io_inen[33] padframe/mprj_io_inen[34] padframe/mprj_io_inen[35] padframe/mprj_io_inen[36]
+ padframe/mprj_io_inen[37] padframe/mprj_io_inen[3] padframe/mprj_io_inen[4] padframe/mprj_io_inen[5]
+ padframe/mprj_io_inen[6] padframe/mprj_io_inen[7] padframe/mprj_io_inen[8] padframe/mprj_io_inen[9]
+ padframe/mprj_io_out[0] padframe/mprj_io_out[10] padframe/mprj_io_out[11] padframe/mprj_io_out[12]
+ padframe/mprj_io_out[13] padframe/mprj_io_out[14] padframe/mprj_io_out[15] padframe/mprj_io_out[16]
+ padframe/mprj_io_out[17] padframe/mprj_io_out[18] padframe/mprj_io_out[19] padframe/mprj_io_out[1]
+ padframe/mprj_io_out[20] padframe/mprj_io_out[21] padframe/mprj_io_out[22] padframe/mprj_io_out[23]
+ padframe/mprj_io_out[24] padframe/mprj_io_out[25] padframe/mprj_io_out[26] padframe/mprj_io_out[27]
+ padframe/mprj_io_out[28] padframe/mprj_io_out[29] padframe/mprj_io_out[2] padframe/mprj_io_out[30]
+ padframe/mprj_io_out[31] padframe/mprj_io_out[32] padframe/mprj_io_out[33] padframe/mprj_io_out[34]
+ padframe/mprj_io_out[35] padframe/mprj_io_out[36] padframe/mprj_io_out[37] padframe/mprj_io_out[3]
+ padframe/mprj_io_out[4] padframe/mprj_io_out[5] padframe/mprj_io_out[6] padframe/mprj_io_out[7]
+ padframe/mprj_io_out[8] padframe/mprj_io_out[9] padframe/mprj_io_outen[0] padframe/mprj_io_outen[10]
+ padframe/mprj_io_outen[11] padframe/mprj_io_outen[12] padframe/mprj_io_outen[13]
+ padframe/mprj_io_outen[14] padframe/mprj_io_outen[15] padframe/mprj_io_outen[16]
+ padframe/mprj_io_outen[17] padframe/mprj_io_outen[18] padframe/mprj_io_outen[19]
+ padframe/mprj_io_outen[1] padframe/mprj_io_outen[20] padframe/mprj_io_outen[21]
+ padframe/mprj_io_outen[22] padframe/mprj_io_outen[23] padframe/mprj_io_outen[24]
+ padframe/mprj_io_outen[25] padframe/mprj_io_outen[26] padframe/mprj_io_outen[27]
+ padframe/mprj_io_outen[28] padframe/mprj_io_outen[29] padframe/mprj_io_outen[2]
+ padframe/mprj_io_outen[30] padframe/mprj_io_outen[31] padframe/mprj_io_outen[32]
+ padframe/mprj_io_outen[33] padframe/mprj_io_outen[34] padframe/mprj_io_outen[35]
+ padframe/mprj_io_outen[36] padframe/mprj_io_outen[37] padframe/mprj_io_outen[3]
+ padframe/mprj_io_outen[4] padframe/mprj_io_outen[5] padframe/mprj_io_outen[6] padframe/mprj_io_outen[7]
+ padframe/mprj_io_outen[8] padframe/mprj_io_outen[9] padframe/mprj_io_pd_select[0]
+ padframe/mprj_io_pd_select[10] padframe/mprj_io_pd_select[11] padframe/mprj_io_pd_select[12]
+ padframe/mprj_io_pd_select[13] padframe/mprj_io_pd_select[14] padframe/mprj_io_pd_select[15]
+ padframe/mprj_io_pd_select[16] padframe/mprj_io_pd_select[17] padframe/mprj_io_pd_select[18]
+ padframe/mprj_io_pd_select[19] padframe/mprj_io_pd_select[1] padframe/mprj_io_pd_select[20]
+ padframe/mprj_io_pd_select[21] padframe/mprj_io_pd_select[22] padframe/mprj_io_pd_select[23]
+ padframe/mprj_io_pd_select[24] padframe/mprj_io_pd_select[25] padframe/mprj_io_pd_select[26]
+ padframe/mprj_io_pd_select[27] padframe/mprj_io_pd_select[28] padframe/mprj_io_pd_select[29]
+ padframe/mprj_io_pd_select[2] padframe/mprj_io_pd_select[30] padframe/mprj_io_pd_select[31]
+ padframe/mprj_io_pd_select[32] padframe/mprj_io_pd_select[33] padframe/mprj_io_pd_select[34]
+ padframe/mprj_io_pd_select[35] padframe/mprj_io_pd_select[36] padframe/mprj_io_pd_select[37]
+ padframe/mprj_io_pd_select[3] padframe/mprj_io_pd_select[4] padframe/mprj_io_pd_select[5]
+ padframe/mprj_io_pd_select[6] padframe/mprj_io_pd_select[7] padframe/mprj_io_pd_select[8]
+ padframe/mprj_io_pd_select[9] padframe/mprj_io_pu_select[0] padframe/mprj_io_pu_select[10]
+ padframe/mprj_io_pu_select[11] padframe/mprj_io_pu_select[12] padframe/mprj_io_pu_select[13]
+ padframe/mprj_io_pu_select[14] padframe/mprj_io_pu_select[15] padframe/mprj_io_pu_select[16]
+ padframe/mprj_io_pu_select[17] padframe/mprj_io_pu_select[18] padframe/mprj_io_pu_select[19]
+ padframe/mprj_io_pu_select[1] padframe/mprj_io_pu_select[20] padframe/mprj_io_pu_select[21]
+ padframe/mprj_io_pu_select[22] padframe/mprj_io_pu_select[23] padframe/mprj_io_pu_select[24]
+ padframe/mprj_io_pu_select[25] padframe/mprj_io_pu_select[26] padframe/mprj_io_pu_select[27]
+ padframe/mprj_io_pu_select[28] padframe/mprj_io_pu_select[29] padframe/mprj_io_pu_select[2]
+ padframe/mprj_io_pu_select[30] padframe/mprj_io_pu_select[31] padframe/mprj_io_pu_select[32]
+ padframe/mprj_io_pu_select[33] padframe/mprj_io_pu_select[34] padframe/mprj_io_pu_select[35]
+ padframe/mprj_io_pu_select[36] padframe/mprj_io_pu_select[37] padframe/mprj_io_pu_select[3]
+ padframe/mprj_io_pu_select[4] padframe/mprj_io_pu_select[5] padframe/mprj_io_pu_select[6]
+ padframe/mprj_io_pu_select[7] padframe/mprj_io_pu_select[8] padframe/mprj_io_pu_select[9]
+ padframe/mprj_io_schmitt_select[0] padframe/mprj_io_schmitt_select[10] padframe/mprj_io_schmitt_select[11]
+ padframe/mprj_io_schmitt_select[12] padframe/mprj_io_schmitt_select[13] padframe/mprj_io_schmitt_select[14]
+ padframe/mprj_io_schmitt_select[15] padframe/mprj_io_schmitt_select[16] padframe/mprj_io_schmitt_select[17]
+ padframe/mprj_io_schmitt_select[18] padframe/mprj_io_schmitt_select[19] padframe/mprj_io_schmitt_select[1]
+ padframe/mprj_io_schmitt_select[20] padframe/mprj_io_schmitt_select[21] padframe/mprj_io_schmitt_select[22]
+ padframe/mprj_io_schmitt_select[23] padframe/mprj_io_schmitt_select[24] padframe/mprj_io_schmitt_select[25]
+ padframe/mprj_io_schmitt_select[26] padframe/mprj_io_schmitt_select[27] padframe/mprj_io_schmitt_select[28]
+ padframe/mprj_io_schmitt_select[29] padframe/mprj_io_schmitt_select[2] padframe/mprj_io_schmitt_select[30]
+ padframe/mprj_io_schmitt_select[31] padframe/mprj_io_schmitt_select[32] padframe/mprj_io_schmitt_select[33]
+ padframe/mprj_io_schmitt_select[34] padframe/mprj_io_schmitt_select[35] padframe/mprj_io_schmitt_select[36]
+ padframe/mprj_io_schmitt_select[37] padframe/mprj_io_schmitt_select[3] padframe/mprj_io_schmitt_select[4]
+ padframe/mprj_io_schmitt_select[5] padframe/mprj_io_schmitt_select[6] padframe/mprj_io_schmitt_select[7]
+ padframe/mprj_io_schmitt_select[8] padframe/mprj_io_schmitt_select[9] padframe/mprj_io_slew_select[0]
+ padframe/mprj_io_slew_select[10] padframe/mprj_io_slew_select[11] padframe/mprj_io_slew_select[12]
+ padframe/mprj_io_slew_select[13] padframe/mprj_io_slew_select[14] padframe/mprj_io_slew_select[15]
+ padframe/mprj_io_slew_select[16] padframe/mprj_io_slew_select[17] padframe/mprj_io_slew_select[18]
+ padframe/mprj_io_slew_select[19] padframe/mprj_io_slew_select[1] padframe/mprj_io_slew_select[20]
+ padframe/mprj_io_slew_select[21] padframe/mprj_io_slew_select[22] padframe/mprj_io_slew_select[23]
+ padframe/mprj_io_slew_select[24] padframe/mprj_io_slew_select[25] padframe/mprj_io_slew_select[26]
+ padframe/mprj_io_slew_select[27] padframe/mprj_io_slew_select[28] padframe/mprj_io_slew_select[29]
+ padframe/mprj_io_slew_select[2] padframe/mprj_io_slew_select[30] padframe/mprj_io_slew_select[31]
+ padframe/mprj_io_slew_select[32] padframe/mprj_io_slew_select[33] padframe/mprj_io_slew_select[34]
+ padframe/mprj_io_slew_select[35] padframe/mprj_io_slew_select[36] padframe/mprj_io_slew_select[37]
+ padframe/mprj_io_slew_select[3] padframe/mprj_io_slew_select[4] padframe/mprj_io_slew_select[5]
+ padframe/mprj_io_slew_select[6] padframe/mprj_io_slew_select[7] padframe/mprj_io_slew_select[8]
+ padframe/mprj_io_slew_select[9] resetb pll/resetb vdd vss soc/VSS soc/VDD chip_io
Xgpio_defaults_block_13 gpio_defaults_block_13/gpio_defaults[0] gpio_defaults_block_13/gpio_defaults[1]
+ gpio_defaults_block_13/gpio_defaults[2] gpio_defaults_block_13/gpio_defaults[3]
+ gpio_defaults_block_13/gpio_defaults[4] gpio_defaults_block_13/gpio_defaults[5]
+ gpio_defaults_block_13/gpio_defaults[6] gpio_defaults_block_13/gpio_defaults[7]
+ gpio_defaults_block_13/gpio_defaults[8] gpio_defaults_block_13/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_24 gpio_defaults_block_24/gpio_defaults[0] gpio_defaults_block_24/gpio_defaults[1]
+ gpio_defaults_block_24/gpio_defaults[2] gpio_defaults_block_24/gpio_defaults[3]
+ gpio_defaults_block_24/gpio_defaults[4] gpio_defaults_block_24/gpio_defaults[5]
+ gpio_defaults_block_24/gpio_defaults[6] gpio_defaults_block_24/gpio_defaults[7]
+ gpio_defaults_block_24/gpio_defaults[8] gpio_defaults_block_24/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_in_2\[14\] soc/VDD soc/VSS gpio_defaults_block_27/gpio_defaults[0] gpio_defaults_block_27/gpio_defaults[1]
+ gpio_defaults_block_27/gpio_defaults[2] gpio_defaults_block_27/gpio_defaults[3]
+ gpio_defaults_block_27/gpio_defaults[4] gpio_defaults_block_27/gpio_defaults[5]
+ gpio_defaults_block_27/gpio_defaults[6] gpio_defaults_block_27/gpio_defaults[7]
+ gpio_defaults_block_27/gpio_defaults[8] gpio_defaults_block_27/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[33] gpio_control_in_2\[14\]/zero housekeeping/mgmt_gpio_out[33]
+ gpio_control_in_2\[14\]/one padframe/mprj_io_drive_sel[66] padframe/mprj_io_drive_sel[67]
+ padframe/mprj_io_in[33] padframe/mprj_io_inen[33] padframe/mprj_io_out[33] padframe/mprj_io_outen[33]
+ padframe/mprj_io_pd_select[33] padframe/mprj_io_pu_select[33] padframe/mprj_io_schmitt_select[33]
+ padframe/mprj_io_slew_select[33] gpio_control_in_2\[14\]/resetn gpio_control_in_2\[13\]/resetn
+ gpio_control_in_2\[14\]/serial_clock gpio_control_in_2\[13\]/serial_clock gpio_control_in_2\[14\]/serial_data_in
+ gpio_control_in_2\[13\]/serial_data_in gpio_control_in_2\[14\]/serial_load gpio_control_in_2\[13\]/serial_load
+ mprj/io_in[33] mprj/io_oeb[33] mprj/io_out[33] gpio_control_in_2\[14\]/zero gpio_control_block
Xgpio_control_in_1a\[3\] soc/VDD soc/VSS gpio_defaults_block_28/gpio_defaults[0] gpio_defaults_block_28/gpio_defaults[1]
+ gpio_defaults_block_28/gpio_defaults[2] gpio_defaults_block_28/gpio_defaults[3]
+ gpio_defaults_block_28/gpio_defaults[4] gpio_defaults_block_28/gpio_defaults[5]
+ gpio_defaults_block_28/gpio_defaults[6] gpio_defaults_block_28/gpio_defaults[7]
+ gpio_defaults_block_28/gpio_defaults[8] gpio_defaults_block_28/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[5] gpio_control_in_1a\[3\]/zero housekeeping/mgmt_gpio_out[5]
+ gpio_control_in_1a\[3\]/one padframe/mprj_io_drive_sel[11] padframe/mprj_io_drive_sel[10]
+ padframe/mprj_io_in[5] padframe/mprj_io_inen[5] padframe/mprj_io_out[5] padframe/mprj_io_outen[5]
+ padframe/mprj_io_pd_select[5] padframe/mprj_io_pu_select[5] padframe/mprj_io_schmitt_select[5]
+ padframe/mprj_io_slew_select[5] gpio_control_in_1a\[3\]/resetn gpio_control_in_1a\[4\]/resetn
+ gpio_control_in_1a\[3\]/serial_clock gpio_control_in_1a\[4\]/serial_clock gpio_control_in_1a\[3\]/serial_data_in
+ gpio_control_in_1a\[4\]/serial_data_in gpio_control_in_1a\[3\]/serial_load gpio_control_in_1a\[4\]/serial_load
+ mprj/io_in[5] mprj/io_oeb[5] mprj/io_out[5] gpio_control_in_1a\[3\]/zero gpio_control_block
Xgpio_control_bidir_2\[0\] soc/VDD soc/VSS gpio_defaults_block_30/gpio_defaults[0]
+ gpio_defaults_block_30/gpio_defaults[1] gpio_defaults_block_30/gpio_defaults[2]
+ gpio_defaults_block_30/gpio_defaults[3] gpio_defaults_block_30/gpio_defaults[4]
+ gpio_defaults_block_30/gpio_defaults[5] gpio_defaults_block_30/gpio_defaults[6]
+ gpio_defaults_block_30/gpio_defaults[7] gpio_defaults_block_30/gpio_defaults[8]
+ gpio_defaults_block_30/gpio_defaults[9] housekeeping/mgmt_gpio_in[35] housekeeping/mgmt_gpio_oeb[35]
+ housekeeping/mgmt_gpio_out[35] gpio_control_bidir_2\[0\]/one padframe/mprj_io_drive_sel[70]
+ padframe/mprj_io_drive_sel[71] padframe/mprj_io_in[35] padframe/mprj_io_inen[35]
+ padframe/mprj_io_out[35] padframe/mprj_io_outen[35] padframe/mprj_io_pd_select[35]
+ padframe/mprj_io_pu_select[35] padframe/mprj_io_schmitt_select[35] padframe/mprj_io_slew_select[35]
+ gpio_control_bidir_2\[0\]/resetn gpio_control_in_2\[15\]/resetn gpio_control_bidir_2\[0\]/serial_clock
+ gpio_control_in_2\[15\]/serial_clock gpio_control_bidir_2\[0\]/serial_data_in gpio_control_in_2\[15\]/serial_data_in
+ gpio_control_bidir_2\[0\]/serial_load gpio_control_in_2\[15\]/serial_load mprj/io_in[35]
+ mprj/io_oeb[35] mprj/io_out[35] gpio_control_bidir_2\[0\]/zero gpio_control_block
Xsoc soc/VDD soc/VSS soc/core_clk soc/core_rstn soc/debug_in soc/debug_mode soc/debug_oeb
+ soc/debug_out soc/flash_clk soc/flash_csb soc/flash_io0_di soc/flash_io0_do soc/flash_io0_oeb
+ soc/flash_io1_di soc/flash_io1_do soc/flash_io1_oeb soc/flash_io2_di soc/flash_io2_do
+ soc/flash_io2_oeb soc/flash_io3_di soc/flash_io3_do soc/flash_io3_oeb soc/gpio_in_pad
+ soc/gpio_inenb_pad soc/gpio_mode0_pad soc/gpio_mode1_pad soc/gpio_out_pad soc/gpio_outenb_pad
+ soc/hk_ack_i soc/hk_cyc_o soc/hk_dat_i[0] soc/hk_dat_i[10] soc/hk_dat_i[11] soc/hk_dat_i[12]
+ soc/hk_dat_i[13] soc/hk_dat_i[14] soc/hk_dat_i[15] soc/hk_dat_i[16] soc/hk_dat_i[17]
+ soc/hk_dat_i[18] soc/hk_dat_i[19] soc/hk_dat_i[1] soc/hk_dat_i[20] soc/hk_dat_i[21]
+ soc/hk_dat_i[22] soc/hk_dat_i[23] soc/hk_dat_i[24] soc/hk_dat_i[25] soc/hk_dat_i[26]
+ soc/hk_dat_i[27] soc/hk_dat_i[28] soc/hk_dat_i[29] soc/hk_dat_i[2] soc/hk_dat_i[30]
+ soc/hk_dat_i[31] soc/hk_dat_i[3] soc/hk_dat_i[4] soc/hk_dat_i[5] soc/hk_dat_i[6]
+ soc/hk_dat_i[7] soc/hk_dat_i[8] soc/hk_dat_i[9] soc/hk_stb_o soc/irq[0] soc/irq[1]
+ soc/irq[2] soc/irq[3] soc/irq[4] soc/irq[5] soc/la_iena[0] soc/la_iena[10] soc/la_iena[11]
+ soc/la_iena[12] soc/la_iena[13] soc/la_iena[14] soc/la_iena[15] soc/la_iena[16]
+ soc/la_iena[17] soc/la_iena[18] soc/la_iena[19] soc/la_iena[1] soc/la_iena[20] soc/la_iena[21]
+ soc/la_iena[22] soc/la_iena[23] soc/la_iena[24] soc/la_iena[25] soc/la_iena[26]
+ soc/la_iena[27] soc/la_iena[28] soc/la_iena[29] soc/la_iena[2] soc/la_iena[30] soc/la_iena[31]
+ soc/la_iena[32] soc/la_iena[33] soc/la_iena[34] soc/la_iena[35] soc/la_iena[36]
+ soc/la_iena[37] soc/la_iena[38] soc/la_iena[39] soc/la_iena[3] soc/la_iena[40] soc/la_iena[41]
+ soc/la_iena[42] soc/la_iena[43] soc/la_iena[44] soc/la_iena[45] soc/la_iena[46]
+ soc/la_iena[47] soc/la_iena[48] soc/la_iena[49] soc/la_iena[4] soc/la_iena[50] soc/la_iena[51]
+ soc/la_iena[52] soc/la_iena[53] soc/la_iena[54] soc/la_iena[55] soc/la_iena[56]
+ soc/la_iena[57] soc/la_iena[58] soc/la_iena[59] soc/la_iena[5] soc/la_iena[60] soc/la_iena[61]
+ soc/la_iena[62] soc/la_iena[63] soc/la_iena[6] soc/la_iena[7] soc/la_iena[8] soc/la_iena[9]
+ soc/la_input[0] soc/la_input[10] soc/la_input[11] soc/la_input[12] soc/la_input[13]
+ soc/la_input[14] soc/la_input[15] soc/la_input[16] soc/la_input[17] soc/la_input[18]
+ soc/la_input[19] soc/la_input[1] soc/la_input[20] soc/la_input[21] soc/la_input[22]
+ soc/la_input[23] soc/la_input[24] soc/la_input[25] soc/la_input[26] soc/la_input[27]
+ soc/la_input[28] soc/la_input[29] soc/la_input[2] soc/la_input[30] soc/la_input[31]
+ soc/la_input[32] soc/la_input[33] soc/la_input[34] soc/la_input[35] soc/la_input[36]
+ soc/la_input[37] soc/la_input[38] soc/la_input[39] soc/la_input[3] soc/la_input[40]
+ soc/la_input[41] soc/la_input[42] soc/la_input[43] soc/la_input[44] soc/la_input[45]
+ soc/la_input[46] soc/la_input[47] soc/la_input[48] soc/la_input[49] soc/la_input[4]
+ soc/la_input[50] soc/la_input[51] soc/la_input[52] soc/la_input[53] soc/la_input[54]
+ soc/la_input[55] soc/la_input[56] soc/la_input[57] soc/la_input[58] soc/la_input[59]
+ soc/la_input[5] soc/la_input[60] soc/la_input[61] soc/la_input[62] soc/la_input[63]
+ soc/la_input[6] soc/la_input[7] soc/la_input[8] soc/la_input[9] soc/la_oenb[0] soc/la_oenb[10]
+ soc/la_oenb[11] soc/la_oenb[12] soc/la_oenb[13] soc/la_oenb[14] soc/la_oenb[15]
+ soc/la_oenb[16] soc/la_oenb[17] soc/la_oenb[18] soc/la_oenb[19] soc/la_oenb[1] soc/la_oenb[20]
+ soc/la_oenb[21] soc/la_oenb[22] soc/la_oenb[23] soc/la_oenb[24] soc/la_oenb[25]
+ soc/la_oenb[26] soc/la_oenb[27] soc/la_oenb[28] soc/la_oenb[29] soc/la_oenb[2] soc/la_oenb[30]
+ soc/la_oenb[31] soc/la_oenb[32] soc/la_oenb[33] soc/la_oenb[34] soc/la_oenb[35]
+ soc/la_oenb[36] soc/la_oenb[37] soc/la_oenb[38] soc/la_oenb[39] soc/la_oenb[3] soc/la_oenb[40]
+ soc/la_oenb[41] soc/la_oenb[42] soc/la_oenb[43] soc/la_oenb[44] soc/la_oenb[45]
+ soc/la_oenb[46] soc/la_oenb[47] soc/la_oenb[48] soc/la_oenb[49] soc/la_oenb[4] soc/la_oenb[50]
+ soc/la_oenb[51] soc/la_oenb[52] soc/la_oenb[53] soc/la_oenb[54] soc/la_oenb[55]
+ soc/la_oenb[56] soc/la_oenb[57] soc/la_oenb[58] soc/la_oenb[59] soc/la_oenb[5] soc/la_oenb[60]
+ soc/la_oenb[61] soc/la_oenb[62] soc/la_oenb[63] soc/la_oenb[6] soc/la_oenb[7] soc/la_oenb[8]
+ soc/la_oenb[9] soc/la_output[0] soc/la_output[10] soc/la_output[11] soc/la_output[12]
+ soc/la_output[13] soc/la_output[14] soc/la_output[15] soc/la_output[16] soc/la_output[17]
+ soc/la_output[18] soc/la_output[19] soc/la_output[1] soc/la_output[20] soc/la_output[21]
+ soc/la_output[22] soc/la_output[23] soc/la_output[24] soc/la_output[25] soc/la_output[26]
+ soc/la_output[27] soc/la_output[28] soc/la_output[29] soc/la_output[2] soc/la_output[30]
+ soc/la_output[31] soc/la_output[32] soc/la_output[33] soc/la_output[34] soc/la_output[35]
+ soc/la_output[36] soc/la_output[37] soc/la_output[38] soc/la_output[39] soc/la_output[3]
+ soc/la_output[40] soc/la_output[41] soc/la_output[42] soc/la_output[43] soc/la_output[44]
+ soc/la_output[45] soc/la_output[46] soc/la_output[47] soc/la_output[48] soc/la_output[49]
+ soc/la_output[4] soc/la_output[50] soc/la_output[51] soc/la_output[52] soc/la_output[53]
+ soc/la_output[54] soc/la_output[55] soc/la_output[56] soc/la_output[57] soc/la_output[58]
+ soc/la_output[59] soc/la_output[5] soc/la_output[60] soc/la_output[61] soc/la_output[62]
+ soc/la_output[63] soc/la_output[6] soc/la_output[7] soc/la_output[8] soc/la_output[9]
+ soc/mprj_ack_i soc/mprj_adr_o[0] soc/mprj_adr_o[10] soc/mprj_adr_o[11] soc/mprj_adr_o[12]
+ soc/mprj_adr_o[13] soc/mprj_adr_o[14] soc/mprj_adr_o[15] soc/mprj_adr_o[16] soc/mprj_adr_o[17]
+ soc/mprj_adr_o[18] soc/mprj_adr_o[19] soc/mprj_adr_o[1] soc/mprj_adr_o[20] soc/mprj_adr_o[21]
+ soc/mprj_adr_o[22] soc/mprj_adr_o[23] soc/mprj_adr_o[24] soc/mprj_adr_o[25] soc/mprj_adr_o[26]
+ soc/mprj_adr_o[27] soc/mprj_adr_o[28] soc/mprj_adr_o[29] soc/mprj_adr_o[2] soc/mprj_adr_o[30]
+ soc/mprj_adr_o[31] soc/mprj_adr_o[3] soc/mprj_adr_o[4] soc/mprj_adr_o[5] soc/mprj_adr_o[6]
+ soc/mprj_adr_o[7] soc/mprj_adr_o[8] soc/mprj_adr_o[9] soc/mprj_cyc_o soc/mprj_dat_i[0]
+ soc/mprj_dat_i[10] soc/mprj_dat_i[11] soc/mprj_dat_i[12] soc/mprj_dat_i[13] soc/mprj_dat_i[14]
+ soc/mprj_dat_i[15] soc/mprj_dat_i[16] soc/mprj_dat_i[17] soc/mprj_dat_i[18] soc/mprj_dat_i[19]
+ soc/mprj_dat_i[1] soc/mprj_dat_i[20] soc/mprj_dat_i[21] soc/mprj_dat_i[22] soc/mprj_dat_i[23]
+ soc/mprj_dat_i[24] soc/mprj_dat_i[25] soc/mprj_dat_i[26] soc/mprj_dat_i[27] soc/mprj_dat_i[28]
+ soc/mprj_dat_i[29] soc/mprj_dat_i[2] soc/mprj_dat_i[30] soc/mprj_dat_i[31] soc/mprj_dat_i[3]
+ soc/mprj_dat_i[4] soc/mprj_dat_i[5] soc/mprj_dat_i[6] soc/mprj_dat_i[7] soc/mprj_dat_i[8]
+ soc/mprj_dat_i[9] soc/mprj_dat_o[0] soc/mprj_dat_o[10] soc/mprj_dat_o[11] soc/mprj_dat_o[12]
+ soc/mprj_dat_o[13] soc/mprj_dat_o[14] soc/mprj_dat_o[15] soc/mprj_dat_o[16] soc/mprj_dat_o[17]
+ soc/mprj_dat_o[18] soc/mprj_dat_o[19] soc/mprj_dat_o[1] soc/mprj_dat_o[20] soc/mprj_dat_o[21]
+ soc/mprj_dat_o[22] soc/mprj_dat_o[23] soc/mprj_dat_o[24] soc/mprj_dat_o[25] soc/mprj_dat_o[26]
+ soc/mprj_dat_o[27] soc/mprj_dat_o[28] soc/mprj_dat_o[29] soc/mprj_dat_o[2] soc/mprj_dat_o[30]
+ soc/mprj_dat_o[31] soc/mprj_dat_o[3] soc/mprj_dat_o[4] soc/mprj_dat_o[5] soc/mprj_dat_o[6]
+ soc/mprj_dat_o[7] soc/mprj_dat_o[8] soc/mprj_dat_o[9] soc/mprj_sel_o[0] soc/mprj_sel_o[1]
+ soc/mprj_sel_o[2] soc/mprj_sel_o[3] soc/mprj_stb_o soc/mprj_wb_iena soc/mprj_we_o
+ soc/qspi_enabled soc/ser_rx soc/ser_tx soc/spi_csb soc/spi_enabled soc/spi_sck soc/spi_sdi
+ soc/spi_sdo soc/spi_sdoenb soc/trap soc/uart_enabled soc/user_irq_ena[0] soc/user_irq_ena[1]
+ soc/user_irq_ena[2] mgmt_core_wrapper
Xgpio_defaults_block_14 gpio_defaults_block_14/gpio_defaults[0] gpio_defaults_block_14/gpio_defaults[1]
+ gpio_defaults_block_14/gpio_defaults[2] gpio_defaults_block_14/gpio_defaults[3]
+ gpio_defaults_block_14/gpio_defaults[4] gpio_defaults_block_14/gpio_defaults[5]
+ gpio_defaults_block_14/gpio_defaults[6] gpio_defaults_block_14/gpio_defaults[7]
+ gpio_defaults_block_14/gpio_defaults[8] gpio_defaults_block_14/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_in_2\[9\] soc/VDD soc/VSS gpio_defaults_block_18/gpio_defaults[0] gpio_defaults_block_18/gpio_defaults[1]
+ gpio_defaults_block_18/gpio_defaults[2] gpio_defaults_block_18/gpio_defaults[3]
+ gpio_defaults_block_18/gpio_defaults[4] gpio_defaults_block_18/gpio_defaults[5]
+ gpio_defaults_block_18/gpio_defaults[6] gpio_defaults_block_18/gpio_defaults[7]
+ gpio_defaults_block_18/gpio_defaults[8] gpio_defaults_block_18/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[28] gpio_control_in_2\[9\]/zero housekeeping/mgmt_gpio_out[28]
+ gpio_control_in_2\[9\]/one padframe/mprj_io_drive_sel[56] padframe/mprj_io_drive_sel[57]
+ padframe/mprj_io_in[28] padframe/mprj_io_inen[28] padframe/mprj_io_out[28] padframe/mprj_io_outen[28]
+ padframe/mprj_io_pd_select[28] padframe/mprj_io_pu_select[28] padframe/mprj_io_schmitt_select[28]
+ padframe/mprj_io_slew_select[28] gpio_control_in_2\[9\]/resetn gpio_control_in_2\[8\]/resetn
+ gpio_control_in_2\[9\]/serial_clock gpio_control_in_2\[8\]/serial_clock gpio_control_in_2\[9\]/serial_data_in
+ gpio_control_in_2\[8\]/serial_data_in gpio_control_in_2\[9\]/serial_load gpio_control_in_2\[8\]/serial_load
+ mprj/io_in[28] mprj/io_oeb[28] mprj/io_out[28] gpio_control_in_2\[9\]/zero gpio_control_block
Xgpio_defaults_block_25 gpio_defaults_block_25/gpio_defaults[0] gpio_defaults_block_25/gpio_defaults[1]
+ gpio_defaults_block_25/gpio_defaults[2] gpio_defaults_block_25/gpio_defaults[3]
+ gpio_defaults_block_25/gpio_defaults[4] gpio_defaults_block_25/gpio_defaults[5]
+ gpio_defaults_block_25/gpio_defaults[6] gpio_defaults_block_25/gpio_defaults[7]
+ gpio_defaults_block_25/gpio_defaults[8] gpio_defaults_block_25/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xsimple_por_0 soc/VDD soc/VSS simple_por_0/porb simple_por_0/por simple_por
Xgpio_control_in_1\[4\] soc/VDD soc/VSS gpio_defaults_block_11/gpio_defaults[0] gpio_defaults_block_11/gpio_defaults[1]
+ gpio_defaults_block_11/gpio_defaults[2] gpio_defaults_block_11/gpio_defaults[3]
+ gpio_defaults_block_11/gpio_defaults[4] gpio_defaults_block_11/gpio_defaults[5]
+ gpio_defaults_block_11/gpio_defaults[6] gpio_defaults_block_11/gpio_defaults[7]
+ gpio_defaults_block_11/gpio_defaults[8] gpio_defaults_block_11/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[12] gpio_control_in_1\[4\]/zero housekeeping/mgmt_gpio_out[12]
+ gpio_control_in_1\[4\]/one padframe/mprj_io_drive_sel[25] padframe/mprj_io_drive_sel[24]
+ padframe/mprj_io_in[12] padframe/mprj_io_inen[12] padframe/mprj_io_out[12] padframe/mprj_io_outen[12]
+ padframe/mprj_io_pd_select[12] padframe/mprj_io_pu_select[12] padframe/mprj_io_schmitt_select[12]
+ padframe/mprj_io_slew_select[12] gpio_control_in_1\[4\]/resetn gpio_control_in_1\[5\]/resetn
+ gpio_control_in_1\[4\]/serial_clock gpio_control_in_1\[5\]/serial_clock gpio_control_in_1\[4\]/serial_data_in
+ gpio_control_in_1\[5\]/serial_data_in gpio_control_in_1\[4\]/serial_load gpio_control_in_1\[5\]/serial_load
+ mprj/io_in[12] mprj/io_oeb[12] mprj/io_out[12] gpio_control_in_1\[4\]/zero gpio_control_block
Xgpio_defaults_block_15 gpio_defaults_block_15/gpio_defaults[0] gpio_defaults_block_15/gpio_defaults[1]
+ gpio_defaults_block_15/gpio_defaults[2] gpio_defaults_block_15/gpio_defaults[3]
+ gpio_defaults_block_15/gpio_defaults[4] gpio_defaults_block_15/gpio_defaults[5]
+ gpio_defaults_block_15/gpio_defaults[6] gpio_defaults_block_15/gpio_defaults[7]
+ gpio_defaults_block_15/gpio_defaults[8] gpio_defaults_block_15/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_26 gpio_defaults_block_26/gpio_defaults[0] gpio_defaults_block_26/gpio_defaults[1]
+ gpio_defaults_block_26/gpio_defaults[2] gpio_defaults_block_26/gpio_defaults[3]
+ gpio_defaults_block_26/gpio_defaults[4] gpio_defaults_block_26/gpio_defaults[5]
+ gpio_defaults_block_26/gpio_defaults[6] gpio_defaults_block_26/gpio_defaults[7]
+ gpio_defaults_block_26/gpio_defaults[8] gpio_defaults_block_26/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_16 gpio_defaults_block_16/gpio_defaults[0] gpio_defaults_block_16/gpio_defaults[1]
+ gpio_defaults_block_16/gpio_defaults[2] gpio_defaults_block_16/gpio_defaults[3]
+ gpio_defaults_block_16/gpio_defaults[4] gpio_defaults_block_16/gpio_defaults[5]
+ gpio_defaults_block_16/gpio_defaults[6] gpio_defaults_block_16/gpio_defaults[7]
+ gpio_defaults_block_16/gpio_defaults[8] gpio_defaults_block_16/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_in_2\[12\] soc/VDD soc/VSS gpio_defaults_block_22/gpio_defaults[0] gpio_defaults_block_22/gpio_defaults[1]
+ gpio_defaults_block_22/gpio_defaults[2] gpio_defaults_block_22/gpio_defaults[3]
+ gpio_defaults_block_22/gpio_defaults[4] gpio_defaults_block_22/gpio_defaults[5]
+ gpio_defaults_block_22/gpio_defaults[6] gpio_defaults_block_22/gpio_defaults[7]
+ gpio_defaults_block_22/gpio_defaults[8] gpio_defaults_block_22/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[31] gpio_control_in_2\[12\]/zero housekeeping/mgmt_gpio_out[31]
+ gpio_control_in_2\[12\]/one padframe/mprj_io_drive_sel[62] padframe/mprj_io_drive_sel[63]
+ padframe/mprj_io_in[31] padframe/mprj_io_inen[31] padframe/mprj_io_out[31] padframe/mprj_io_outen[31]
+ padframe/mprj_io_pd_select[31] padframe/mprj_io_pu_select[31] padframe/mprj_io_schmitt_select[31]
+ padframe/mprj_io_slew_select[31] gpio_control_in_2\[12\]/resetn gpio_control_in_2\[11\]/resetn
+ gpio_control_in_2\[12\]/serial_clock gpio_control_in_2\[11\]/serial_clock gpio_control_in_2\[12\]/serial_data_in
+ gpio_control_in_2\[11\]/serial_data_in gpio_control_in_2\[12\]/serial_load gpio_control_in_2\[11\]/serial_load
+ mprj/io_in[31] mprj/io_oeb[31] mprj/io_out[31] gpio_control_in_2\[12\]/zero gpio_control_block
Xgpio_defaults_block_27 gpio_defaults_block_27/gpio_defaults[0] gpio_defaults_block_27/gpio_defaults[1]
+ gpio_defaults_block_27/gpio_defaults[2] gpio_defaults_block_27/gpio_defaults[3]
+ gpio_defaults_block_27/gpio_defaults[4] gpio_defaults_block_27/gpio_defaults[5]
+ gpio_defaults_block_27/gpio_defaults[6] gpio_defaults_block_27/gpio_defaults[7]
+ gpio_defaults_block_27/gpio_defaults[8] gpio_defaults_block_27/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_in_1a\[1\] soc/VDD soc/VSS gpio_control_in_1a\[1\]/gpio_defaults[0]
+ gpio_control_in_1a\[1\]/gpio_defaults[1] gpio_control_in_1a\[1\]/gpio_defaults[2]
+ gpio_control_in_1a\[1\]/gpio_defaults[3] gpio_control_in_1a\[1\]/gpio_defaults[4]
+ gpio_control_in_1a\[1\]/gpio_defaults[5] gpio_control_in_1a\[1\]/gpio_defaults[6]
+ gpio_control_in_1a\[1\]/gpio_defaults[7] gpio_control_in_1a\[1\]/gpio_defaults[8]
+ gpio_control_in_1a\[1\]/gpio_defaults[9] housekeeping/mgmt_gpio_in[3] gpio_control_in_1a\[1\]/zero
+ housekeeping/mgmt_gpio_out[3] gpio_control_in_1a\[1\]/one padframe/mprj_io_drive_sel[7]
+ padframe/mprj_io_drive_sel[6] padframe/mprj_io_in[3] padframe/mprj_io_inen[3] padframe/mprj_io_out[3]
+ padframe/mprj_io_outen[3] padframe/mprj_io_pd_select[3] padframe/mprj_io_pu_select[3]
+ padframe/mprj_io_schmitt_select[3] padframe/mprj_io_slew_select[3] gpio_control_in_1a\[1\]/resetn
+ gpio_control_in_1a\[2\]/resetn gpio_control_in_1a\[1\]/serial_clock gpio_control_in_1a\[2\]/serial_clock
+ gpio_control_in_1a\[1\]/serial_data_in gpio_control_in_1a\[2\]/serial_data_in gpio_control_in_1a\[1\]/serial_load
+ gpio_control_in_1a\[2\]/serial_load mprj/io_in[3] mprj/io_oeb[3] mprj/io_out[3]
+ gpio_control_in_1a\[1\]/zero gpio_control_block
Xclock_ctrl soc/VDD soc/VSS soc/core_clk pll/osc clock_ctrl/ext_clk_sel housekeeping/reset
+ pll/clockp[1] pll/clockp[0] pll/resetb soc/core_rstn clock_ctrl/sel2[0] clock_ctrl/sel2[1]
+ clock_ctrl/sel2[2] clock_ctrl/sel[0] clock_ctrl/sel[1] clock_ctrl/sel[2] clock_ctrl/user_clk
+ caravel_clocking
Xgpio_control_in_2\[7\] soc/VDD soc/VSS gpio_defaults_block_13/gpio_defaults[0] gpio_defaults_block_13/gpio_defaults[1]
+ gpio_defaults_block_13/gpio_defaults[2] gpio_defaults_block_13/gpio_defaults[3]
+ gpio_defaults_block_13/gpio_defaults[4] gpio_defaults_block_13/gpio_defaults[5]
+ gpio_defaults_block_13/gpio_defaults[6] gpio_defaults_block_13/gpio_defaults[7]
+ gpio_defaults_block_13/gpio_defaults[8] gpio_defaults_block_13/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[26] gpio_control_in_2\[7\]/zero housekeeping/mgmt_gpio_out[26]
+ gpio_control_in_2\[7\]/one padframe/mprj_io_drive_sel[52] padframe/mprj_io_drive_sel[53]
+ padframe/mprj_io_in[26] padframe/mprj_io_inen[26] padframe/mprj_io_out[26] padframe/mprj_io_outen[26]
+ padframe/mprj_io_pd_select[26] padframe/mprj_io_pu_select[26] padframe/mprj_io_schmitt_select[26]
+ padframe/mprj_io_slew_select[26] gpio_control_in_2\[7\]/resetn gpio_control_in_2\[6\]/resetn
+ gpio_control_in_2\[7\]/serial_clock gpio_control_in_2\[6\]/serial_clock gpio_control_in_2\[7\]/serial_data_in
+ gpio_control_in_2\[6\]/serial_data_in gpio_control_in_2\[7\]/serial_load gpio_control_in_2\[6\]/serial_load
+ mprj/io_in[26] mprj/io_oeb[26] mprj/io_out[26] gpio_control_in_2\[7\]/zero gpio_control_block
Xgpio_defaults_block_17 gpio_defaults_block_17/gpio_defaults[0] gpio_defaults_block_17/gpio_defaults[1]
+ gpio_defaults_block_17/gpio_defaults[2] gpio_defaults_block_17/gpio_defaults[3]
+ gpio_defaults_block_17/gpio_defaults[4] gpio_defaults_block_17/gpio_defaults[5]
+ gpio_defaults_block_17/gpio_defaults[6] gpio_defaults_block_17/gpio_defaults[7]
+ gpio_defaults_block_17/gpio_defaults[8] gpio_defaults_block_17/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_28 gpio_defaults_block_28/gpio_defaults[0] gpio_defaults_block_28/gpio_defaults[1]
+ gpio_defaults_block_28/gpio_defaults[2] gpio_defaults_block_28/gpio_defaults[3]
+ gpio_defaults_block_28/gpio_defaults[4] gpio_defaults_block_28/gpio_defaults[5]
+ gpio_defaults_block_28/gpio_defaults[6] gpio_defaults_block_28/gpio_defaults[7]
+ gpio_defaults_block_28/gpio_defaults[8] gpio_defaults_block_28/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_in_1\[2\] soc/VDD soc/VSS gpio_defaults_block_16/gpio_defaults[0] gpio_defaults_block_16/gpio_defaults[1]
+ gpio_defaults_block_16/gpio_defaults[2] gpio_defaults_block_16/gpio_defaults[3]
+ gpio_defaults_block_16/gpio_defaults[4] gpio_defaults_block_16/gpio_defaults[5]
+ gpio_defaults_block_16/gpio_defaults[6] gpio_defaults_block_16/gpio_defaults[7]
+ gpio_defaults_block_16/gpio_defaults[8] gpio_defaults_block_16/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[10] gpio_control_in_1\[2\]/zero housekeeping/mgmt_gpio_out[10]
+ gpio_control_in_1\[2\]/one padframe/mprj_io_drive_sel[21] padframe/mprj_io_drive_sel[20]
+ padframe/mprj_io_in[10] padframe/mprj_io_inen[10] padframe/mprj_io_out[10] padframe/mprj_io_outen[10]
+ padframe/mprj_io_pd_select[10] padframe/mprj_io_pu_select[10] padframe/mprj_io_schmitt_select[10]
+ padframe/mprj_io_slew_select[10] gpio_control_in_1\[2\]/resetn gpio_control_in_1\[3\]/resetn
+ gpio_control_in_1\[2\]/serial_clock gpio_control_in_1\[3\]/serial_clock gpio_control_in_1\[2\]/serial_data_in
+ gpio_control_in_1\[3\]/serial_data_in gpio_control_in_1\[2\]/serial_load gpio_control_in_1\[3\]/serial_load
+ mprj/io_in[10] mprj/io_oeb[10] mprj/io_out[10] gpio_control_in_1\[2\]/zero gpio_control_block
Xgpio_defaults_block_18 gpio_defaults_block_18/gpio_defaults[0] gpio_defaults_block_18/gpio_defaults[1]
+ gpio_defaults_block_18/gpio_defaults[2] gpio_defaults_block_18/gpio_defaults[3]
+ gpio_defaults_block_18/gpio_defaults[4] gpio_defaults_block_18/gpio_defaults[5]
+ gpio_defaults_block_18/gpio_defaults[6] gpio_defaults_block_18/gpio_defaults[7]
+ gpio_defaults_block_18/gpio_defaults[8] gpio_defaults_block_18/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_19 gpio_defaults_block_19/gpio_defaults[0] gpio_defaults_block_19/gpio_defaults[1]
+ gpio_defaults_block_19/gpio_defaults[2] gpio_defaults_block_19/gpio_defaults[3]
+ gpio_defaults_block_19/gpio_defaults[4] gpio_defaults_block_19/gpio_defaults[5]
+ gpio_defaults_block_19/gpio_defaults[6] gpio_defaults_block_19/gpio_defaults[7]
+ gpio_defaults_block_19/gpio_defaults[8] gpio_defaults_block_19/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_29 gpio_defaults_block_29/gpio_defaults[0] gpio_defaults_block_29/gpio_defaults[1]
+ gpio_defaults_block_29/gpio_defaults[2] gpio_defaults_block_29/gpio_defaults[3]
+ gpio_defaults_block_29/gpio_defaults[4] gpio_defaults_block_29/gpio_defaults[5]
+ gpio_defaults_block_29/gpio_defaults[6] gpio_defaults_block_29/gpio_defaults[7]
+ gpio_defaults_block_29/gpio_defaults[8] gpio_defaults_block_29/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_in_2\[10\] soc/VDD soc/VSS gpio_defaults_block_17/gpio_defaults[0] gpio_defaults_block_17/gpio_defaults[1]
+ gpio_defaults_block_17/gpio_defaults[2] gpio_defaults_block_17/gpio_defaults[3]
+ gpio_defaults_block_17/gpio_defaults[4] gpio_defaults_block_17/gpio_defaults[5]
+ gpio_defaults_block_17/gpio_defaults[6] gpio_defaults_block_17/gpio_defaults[7]
+ gpio_defaults_block_17/gpio_defaults[8] gpio_defaults_block_17/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[29] gpio_control_in_2\[10\]/zero housekeeping/mgmt_gpio_out[29]
+ gpio_control_in_2\[10\]/one padframe/mprj_io_drive_sel[58] padframe/mprj_io_drive_sel[59]
+ padframe/mprj_io_in[29] padframe/mprj_io_inen[29] padframe/mprj_io_out[29] padframe/mprj_io_outen[29]
+ padframe/mprj_io_pd_select[29] padframe/mprj_io_pu_select[29] padframe/mprj_io_schmitt_select[29]
+ padframe/mprj_io_slew_select[29] gpio_control_in_2\[10\]/resetn gpio_control_in_2\[9\]/resetn
+ gpio_control_in_2\[10\]/serial_clock gpio_control_in_2\[9\]/serial_clock gpio_control_in_2\[10\]/serial_data_in
+ gpio_control_in_2\[9\]/serial_data_in gpio_control_in_2\[10\]/serial_load gpio_control_in_2\[9\]/serial_load
+ mprj/io_in[29] mprj/io_oeb[29] mprj/io_out[29] gpio_control_in_2\[10\]/zero gpio_control_block
Xgpio_defaults_block_0 gpio_defaults_block_0/gpio_defaults[0] gpio_defaults_block_0/gpio_defaults[1]
+ gpio_defaults_block_0/gpio_defaults[2] gpio_defaults_block_0/gpio_defaults[3] gpio_defaults_block_0/gpio_defaults[4]
+ gpio_defaults_block_0/gpio_defaults[5] gpio_defaults_block_0/gpio_defaults[6] gpio_defaults_block_0/gpio_defaults[7]
+ gpio_defaults_block_0/gpio_defaults[8] gpio_defaults_block_0/gpio_defaults[9] gpio_defaults_block_0/VDD
+ gpio_defaults_block_0/VSS gpio_defaults_block
Xgpio_control_in_1\[10\] soc/VDD soc/VSS gpio_defaults_block_4/gpio_defaults[0] gpio_defaults_block_4/gpio_defaults[1]
+ gpio_defaults_block_4/gpio_defaults[2] gpio_defaults_block_4/gpio_defaults[3] gpio_defaults_block_4/gpio_defaults[4]
+ gpio_defaults_block_4/gpio_defaults[5] gpio_defaults_block_4/gpio_defaults[6] gpio_defaults_block_4/gpio_defaults[7]
+ gpio_defaults_block_4/gpio_defaults[8] gpio_defaults_block_4/gpio_defaults[9] housekeeping/mgmt_gpio_in[18]
+ gpio_control_in_1\[10\]/zero housekeeping/mgmt_gpio_out[18] gpio_control_in_1\[10\]/one
+ padframe/mprj_io_drive_sel[36] padframe/mprj_io_drive_sel[37] padframe/mprj_io_in[18]
+ padframe/mprj_io_inen[18] padframe/mprj_io_out[18] padframe/mprj_io_outen[18] padframe/mprj_io_pd_select[18]
+ padframe/mprj_io_pu_select[18] padframe/mprj_io_schmitt_select[18] padframe/mprj_io_slew_select[18]
+ gpio_control_in_1\[10\]/resetn gpio_control_in_1\[10\]/resetn_out gpio_control_in_1\[10\]/serial_clock
+ gpio_control_in_1\[10\]/serial_clock_out gpio_control_in_1\[9\]/serial_data_out
+ gpio_control_in_1\[10\]/serial_data_out gpio_control_in_1\[10\]/serial_load gpio_control_in_1\[10\]/serial_load_out
+ mprj/io_in[18] mprj/io_oeb[18] mprj/io_out[18] gpio_control_in_1\[10\]/zero gpio_control_block
Xgpio_control_in_2\[5\] soc/VDD soc/VSS gpio_defaults_block_10/gpio_defaults[0] gpio_defaults_block_10/gpio_defaults[1]
+ gpio_defaults_block_10/gpio_defaults[2] gpio_defaults_block_10/gpio_defaults[3]
+ gpio_defaults_block_10/gpio_defaults[4] gpio_defaults_block_10/gpio_defaults[5]
+ gpio_defaults_block_10/gpio_defaults[6] gpio_defaults_block_10/gpio_defaults[7]
+ gpio_defaults_block_10/gpio_defaults[8] gpio_defaults_block_10/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[24] gpio_control_in_2\[5\]/zero housekeeping/mgmt_gpio_out[24]
+ gpio_control_in_2\[5\]/one padframe/mprj_io_drive_sel[48] padframe/mprj_io_drive_sel[49]
+ padframe/mprj_io_in[24] padframe/mprj_io_inen[24] padframe/mprj_io_out[24] padframe/mprj_io_outen[24]
+ padframe/mprj_io_pd_select[24] padframe/mprj_io_pu_select[24] padframe/mprj_io_schmitt_select[24]
+ padframe/mprj_io_slew_select[24] gpio_control_in_2\[5\]/resetn gpio_control_in_2\[4\]/resetn
+ gpio_control_in_2\[5\]/serial_clock gpio_control_in_2\[4\]/serial_clock gpio_control_in_2\[5\]/serial_data_in
+ gpio_control_in_2\[4\]/serial_data_in gpio_control_in_2\[5\]/serial_load gpio_control_in_2\[4\]/serial_load
+ mprj/io_in[24] mprj/io_oeb[24] mprj/io_out[24] gpio_control_in_2\[5\]/zero gpio_control_block
Xgpio_control_in_1\[0\] soc/VDD soc/VSS gpio_defaults_block_21/gpio_defaults[0] gpio_defaults_block_21/gpio_defaults[1]
+ gpio_defaults_block_21/gpio_defaults[2] gpio_defaults_block_21/gpio_defaults[3]
+ gpio_defaults_block_21/gpio_defaults[4] gpio_defaults_block_21/gpio_defaults[5]
+ gpio_defaults_block_21/gpio_defaults[6] gpio_defaults_block_21/gpio_defaults[7]
+ gpio_defaults_block_21/gpio_defaults[8] gpio_defaults_block_21/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[8] gpio_control_in_1\[0\]/zero housekeeping/mgmt_gpio_out[8]
+ gpio_control_in_1\[0\]/one padframe/mprj_io_drive_sel[17] padframe/mprj_io_drive_sel[16]
+ padframe/mprj_io_in[8] padframe/mprj_io_inen[8] padframe/mprj_io_out[8] padframe/mprj_io_outen[8]
+ padframe/mprj_io_pd_select[8] padframe/mprj_io_pu_select[8] padframe/mprj_io_schmitt_select[8]
+ padframe/mprj_io_slew_select[8] gpio_control_in_1\[0\]/resetn gpio_control_in_1\[1\]/resetn
+ gpio_control_in_1\[0\]/serial_clock gpio_control_in_1\[1\]/serial_clock gpio_control_in_1\[0\]/serial_data_in
+ gpio_control_in_1\[1\]/serial_data_in gpio_control_in_1\[0\]/serial_load gpio_control_in_1\[1\]/serial_load
+ mprj/io_in[8] mprj/io_oeb[8] mprj/io_out[8] gpio_control_in_1\[0\]/zero gpio_control_block
Xgpio_defaults_block_1 gpio_defaults_block_1/gpio_defaults[0] gpio_defaults_block_1/gpio_defaults[1]
+ gpio_defaults_block_1/gpio_defaults[2] gpio_defaults_block_1/gpio_defaults[3] gpio_defaults_block_1/gpio_defaults[4]
+ gpio_defaults_block_1/gpio_defaults[5] gpio_defaults_block_1/gpio_defaults[6] gpio_defaults_block_1/gpio_defaults[7]
+ gpio_defaults_block_1/gpio_defaults[8] gpio_defaults_block_1/gpio_defaults[9] soc/VDD
+ soc/VSS gpio_defaults_block
Xspare_logic\[3\] soc/VDD soc/VSS spare_logic\[3\]/spare_xfq[0] spare_logic\[3\]/spare_xfq[1]
+ spare_logic\[3\]/spare_xi[0] spare_logic\[3\]/spare_xi[1] spare_logic\[3\]/spare_xi[2]
+ spare_logic\[3\]/spare_xi[3] spare_logic\[3\]/spare_xib spare_logic\[3\]/spare_xmx[0]
+ spare_logic\[3\]/spare_xmx[1] spare_logic\[3\]/spare_xna[0] spare_logic\[3\]/spare_xna[1]
+ spare_logic\[3\]/spare_xno[0] spare_logic\[3\]/spare_xno[1] spare_logic\[3\]/spare_xz[0]
+ spare_logic\[3\]/spare_xz[10] spare_logic\[3\]/spare_xz[11] spare_logic\[3\]/spare_xz[12]
+ spare_logic\[3\]/spare_xz[13] spare_logic\[3\]/spare_xz[14] spare_logic\[3\]/spare_xz[15]
+ spare_logic\[3\]/spare_xz[16] spare_logic\[3\]/spare_xz[17] spare_logic\[3\]/spare_xz[18]
+ spare_logic\[3\]/spare_xz[19] spare_logic\[3\]/spare_xz[1] spare_logic\[3\]/spare_xz[20]
+ spare_logic\[3\]/spare_xz[21] spare_logic\[3\]/spare_xz[22] spare_logic\[3\]/spare_xz[23]
+ spare_logic\[3\]/spare_xz[24] spare_logic\[3\]/spare_xz[25] spare_logic\[3\]/spare_xz[26]
+ spare_logic\[3\]/spare_xz[27] spare_logic\[3\]/spare_xz[28] spare_logic\[3\]/spare_xz[29]
+ spare_logic\[3\]/spare_xz[2] spare_logic\[3\]/spare_xz[30] spare_logic\[3\]/spare_xz[3]
+ spare_logic\[3\]/spare_xz[4] spare_logic\[3\]/spare_xz[5] spare_logic\[3\]/spare_xz[6]
+ spare_logic\[3\]/spare_xz[7] spare_logic\[3\]/spare_xz[8] spare_logic\[3\]/spare_xz[9]
+ spare_logic_block
Xuser_id_value user_id_value/mask_rev[0] user_id_value/mask_rev[10] user_id_value/mask_rev[11]
+ user_id_value/mask_rev[12] user_id_value/mask_rev[13] user_id_value/mask_rev[14]
+ user_id_value/mask_rev[15] user_id_value/mask_rev[16] user_id_value/mask_rev[17]
+ user_id_value/mask_rev[18] user_id_value/mask_rev[19] user_id_value/mask_rev[1]
+ user_id_value/mask_rev[20] user_id_value/mask_rev[21] user_id_value/mask_rev[22]
+ user_id_value/mask_rev[23] user_id_value/mask_rev[24] user_id_value/mask_rev[25]
+ user_id_value/mask_rev[26] user_id_value/mask_rev[27] user_id_value/mask_rev[28]
+ user_id_value/mask_rev[29] user_id_value/mask_rev[2] user_id_value/mask_rev[30]
+ user_id_value/mask_rev[31] user_id_value/mask_rev[3] user_id_value/mask_rev[4] user_id_value/mask_rev[5]
+ user_id_value/mask_rev[6] user_id_value/mask_rev[7] user_id_value/mask_rev[8] user_id_value/mask_rev[9]
+ user_id_value/VDD user_id_value/VSS user_id_programming
Xgpio_defaults_block_2 gpio_defaults_block_2/gpio_defaults[0] gpio_defaults_block_2/gpio_defaults[1]
+ gpio_defaults_block_2/gpio_defaults[2] gpio_defaults_block_2/gpio_defaults[3] gpio_defaults_block_2/gpio_defaults[4]
+ gpio_defaults_block_2/gpio_defaults[5] gpio_defaults_block_2/gpio_defaults[6] gpio_defaults_block_2/gpio_defaults[7]
+ gpio_defaults_block_2/gpio_defaults[8] gpio_defaults_block_2/gpio_defaults[9] gpio_defaults_block_2/VDD
+ gpio_defaults_block_2/VSS gpio_defaults_block
Xgpio_control_in_2\[3\] soc/VDD soc/VSS gpio_defaults_block_9/gpio_defaults[0] gpio_defaults_block_9/gpio_defaults[1]
+ gpio_defaults_block_9/gpio_defaults[2] gpio_defaults_block_9/gpio_defaults[3] gpio_defaults_block_9/gpio_defaults[4]
+ gpio_defaults_block_9/gpio_defaults[5] gpio_defaults_block_9/gpio_defaults[6] gpio_defaults_block_9/gpio_defaults[7]
+ gpio_defaults_block_9/gpio_defaults[8] gpio_defaults_block_9/gpio_defaults[9] housekeeping/mgmt_gpio_in[22]
+ gpio_control_in_2\[3\]/zero housekeeping/mgmt_gpio_out[22] gpio_control_in_2\[3\]/one
+ padframe/mprj_io_drive_sel[44] padframe/mprj_io_drive_sel[45] padframe/mprj_io_in[22]
+ padframe/mprj_io_inen[22] padframe/mprj_io_out[22] padframe/mprj_io_outen[22] padframe/mprj_io_pd_select[22]
+ padframe/mprj_io_pu_select[22] padframe/mprj_io_schmitt_select[22] padframe/mprj_io_slew_select[22]
+ gpio_control_in_2\[3\]/resetn gpio_control_in_2\[2\]/resetn gpio_control_in_2\[3\]/serial_clock
+ gpio_control_in_2\[2\]/serial_clock gpio_control_in_2\[3\]/serial_data_in gpio_control_in_2\[2\]/serial_data_in
+ gpio_control_in_2\[3\]/serial_load gpio_control_in_2\[2\]/serial_load mprj/io_in[22]
+ mprj/io_oeb[22] mprj/io_out[22] gpio_control_in_2\[3\]/zero gpio_control_block
Xgpio_defaults_block_3 gpio_defaults_block_3/gpio_defaults[0] gpio_defaults_block_3/gpio_defaults[1]
+ gpio_defaults_block_3/gpio_defaults[2] gpio_defaults_block_3/gpio_defaults[3] gpio_defaults_block_3/gpio_defaults[4]
+ gpio_defaults_block_3/gpio_defaults[5] gpio_defaults_block_3/gpio_defaults[6] gpio_defaults_block_3/gpio_defaults[7]
+ gpio_defaults_block_3/gpio_defaults[8] gpio_defaults_block_3/gpio_defaults[9] gpio_defaults_block_3/VDD
+ gpio_defaults_block_3/VSS gpio_defaults_block
Xgpio_control_bidir_1\[0\] soc/VDD soc/VSS gpio_defaults_block_009_1/gpio_defaults[0]
+ gpio_defaults_block_009_1/gpio_defaults[1] gpio_defaults_block_009_1/gpio_defaults[2]
+ gpio_defaults_block_009_1/gpio_defaults[3] gpio_defaults_block_009_1/gpio_defaults[4]
+ gpio_defaults_block_009_1/gpio_defaults[5] gpio_defaults_block_009_1/gpio_defaults[6]
+ gpio_defaults_block_009_1/gpio_defaults[7] gpio_defaults_block_009_1/gpio_defaults[8]
+ gpio_defaults_block_009_1/gpio_defaults[9] housekeeping/mgmt_gpio_in[0] housekeeping/mgmt_gpio_oeb[0]
+ housekeeping/mgmt_gpio_out[0] gpio_control_bidir_1\[0\]/one padframe/mprj_io_drive_sel[0]
+ padframe/mprj_io_drive_sel[1] padframe/mprj_io_in[0] padframe/mprj_io_inen[0] padframe/mprj_io_out[0]
+ padframe/mprj_io_outen[0] padframe/mprj_io_pd_select[0] padframe/mprj_io_pu_select[0]
+ padframe/mprj_io_schmitt_select[0] padframe/mprj_io_slew_select[0] housekeeping/serial_resetn
+ gpio_control_bidir_1\[1\]/resetn housekeeping/serial_clock gpio_control_bidir_1\[1\]/serial_clock
+ housekeeping/serial_data_1 gpio_control_bidir_1\[1\]/serial_data_in housekeeping/serial_load
+ gpio_control_bidir_1\[1\]/serial_load mprj/io_in[0] mprj/io_oeb[0] mprj/io_out[0]
+ gpio_control_bidir_1\[0\]/zero gpio_control_block
Xgpio_control_in_1\[9\] soc/VDD soc/VSS gpio_defaults_block_3/gpio_defaults[0] gpio_defaults_block_3/gpio_defaults[1]
+ gpio_defaults_block_3/gpio_defaults[2] gpio_defaults_block_3/gpio_defaults[3] gpio_defaults_block_3/gpio_defaults[4]
+ gpio_defaults_block_3/gpio_defaults[5] gpio_defaults_block_3/gpio_defaults[6] gpio_defaults_block_3/gpio_defaults[7]
+ gpio_defaults_block_3/gpio_defaults[8] gpio_defaults_block_3/gpio_defaults[9] housekeeping/mgmt_gpio_in[17]
+ gpio_control_in_1\[9\]/zero housekeeping/mgmt_gpio_out[17] gpio_control_in_1\[9\]/one
+ padframe/mprj_io_drive_sel[34] padframe/mprj_io_drive_sel[35] padframe/mprj_io_in[17]
+ padframe/mprj_io_inen[17] padframe/mprj_io_out[17] padframe/mprj_io_outen[17] padframe/mprj_io_pd_select[17]
+ padframe/mprj_io_pu_select[17] padframe/mprj_io_schmitt_select[17] padframe/mprj_io_slew_select[17]
+ gpio_control_in_1\[9\]/resetn gpio_control_in_1\[10\]/resetn gpio_control_in_1\[9\]/serial_clock
+ gpio_control_in_1\[10\]/serial_clock gpio_control_in_1\[9\]/serial_data_in gpio_control_in_1\[9\]/serial_data_out
+ gpio_control_in_1\[9\]/serial_load gpio_control_in_1\[10\]/serial_load mprj/io_in[17]
+ mprj/io_oeb[17] mprj/io_out[17] gpio_control_in_1\[9\]/zero gpio_control_block
Xgpio_defaults_block_4 gpio_defaults_block_4/gpio_defaults[0] gpio_defaults_block_4/gpio_defaults[1]
+ gpio_defaults_block_4/gpio_defaults[2] gpio_defaults_block_4/gpio_defaults[3] gpio_defaults_block_4/gpio_defaults[4]
+ gpio_defaults_block_4/gpio_defaults[5] gpio_defaults_block_4/gpio_defaults[6] gpio_defaults_block_4/gpio_defaults[7]
+ gpio_defaults_block_4/gpio_defaults[8] gpio_defaults_block_4/gpio_defaults[9] gpio_defaults_block_4/VDD
+ gpio_defaults_block_4/VSS gpio_defaults_block
Xgpio_defaults_block_5 gpio_defaults_block_5/gpio_defaults[0] gpio_defaults_block_5/gpio_defaults[1]
+ gpio_defaults_block_5/gpio_defaults[2] gpio_defaults_block_5/gpio_defaults[3] gpio_defaults_block_5/gpio_defaults[4]
+ gpio_defaults_block_5/gpio_defaults[5] gpio_defaults_block_5/gpio_defaults[6] gpio_defaults_block_5/gpio_defaults[7]
+ gpio_defaults_block_5/gpio_defaults[8] gpio_defaults_block_5/gpio_defaults[9] gpio_defaults_block_5/VDD
+ gpio_defaults_block_5/VSS gpio_defaults_block
Xspare_logic\[1\] soc/VDD soc/VSS spare_logic\[1\]/spare_xfq[0] spare_logic\[1\]/spare_xfq[1]
+ spare_logic\[1\]/spare_xi[0] spare_logic\[1\]/spare_xi[1] spare_logic\[1\]/spare_xi[2]
+ spare_logic\[1\]/spare_xi[3] spare_logic\[1\]/spare_xib spare_logic\[1\]/spare_xmx[0]
+ spare_logic\[1\]/spare_xmx[1] spare_logic\[1\]/spare_xna[0] spare_logic\[1\]/spare_xna[1]
+ spare_logic\[1\]/spare_xno[0] spare_logic\[1\]/spare_xno[1] spare_logic\[1\]/spare_xz[0]
+ spare_logic\[1\]/spare_xz[10] spare_logic\[1\]/spare_xz[11] spare_logic\[1\]/spare_xz[12]
+ spare_logic\[1\]/spare_xz[13] spare_logic\[1\]/spare_xz[14] spare_logic\[1\]/spare_xz[15]
+ spare_logic\[1\]/spare_xz[16] spare_logic\[1\]/spare_xz[17] spare_logic\[1\]/spare_xz[18]
+ spare_logic\[1\]/spare_xz[19] spare_logic\[1\]/spare_xz[1] spare_logic\[1\]/spare_xz[20]
+ spare_logic\[1\]/spare_xz[21] spare_logic\[1\]/spare_xz[22] spare_logic\[1\]/spare_xz[23]
+ spare_logic\[1\]/spare_xz[24] spare_logic\[1\]/spare_xz[25] spare_logic\[1\]/spare_xz[26]
+ spare_logic\[1\]/spare_xz[27] spare_logic\[1\]/spare_xz[28] spare_logic\[1\]/spare_xz[29]
+ spare_logic\[1\]/spare_xz[2] spare_logic\[1\]/spare_xz[30] spare_logic\[1\]/spare_xz[3]
+ spare_logic\[1\]/spare_xz[4] spare_logic\[1\]/spare_xz[5] spare_logic\[1\]/spare_xz[6]
+ spare_logic\[1\]/spare_xz[7] spare_logic\[1\]/spare_xz[8] spare_logic\[1\]/spare_xz[9]
+ spare_logic_block
Xgpio_defaults_block_6 gpio_defaults_block_6/gpio_defaults[0] gpio_defaults_block_6/gpio_defaults[1]
+ gpio_defaults_block_6/gpio_defaults[2] gpio_defaults_block_6/gpio_defaults[3] gpio_defaults_block_6/gpio_defaults[4]
+ gpio_defaults_block_6/gpio_defaults[5] gpio_defaults_block_6/gpio_defaults[6] gpio_defaults_block_6/gpio_defaults[7]
+ gpio_defaults_block_6/gpio_defaults[8] gpio_defaults_block_6/gpio_defaults[9] gpio_defaults_block_6/VDD
+ gpio_defaults_block_6/VSS gpio_defaults_block
Xgpio_control_in_2\[1\] soc/VDD soc/VSS gpio_defaults_block_5/gpio_defaults[0] gpio_defaults_block_5/gpio_defaults[1]
+ gpio_defaults_block_5/gpio_defaults[2] gpio_defaults_block_5/gpio_defaults[3] gpio_defaults_block_5/gpio_defaults[4]
+ gpio_defaults_block_5/gpio_defaults[5] gpio_defaults_block_5/gpio_defaults[6] gpio_defaults_block_5/gpio_defaults[7]
+ gpio_defaults_block_5/gpio_defaults[8] gpio_defaults_block_5/gpio_defaults[9] housekeeping/mgmt_gpio_in[20]
+ gpio_control_in_2\[1\]/zero housekeeping/mgmt_gpio_out[20] gpio_control_in_2\[1\]/one
+ padframe/mprj_io_drive_sel[40] padframe/mprj_io_drive_sel[41] padframe/mprj_io_in[20]
+ padframe/mprj_io_inen[20] padframe/mprj_io_out[20] padframe/mprj_io_outen[20] padframe/mprj_io_pd_select[20]
+ padframe/mprj_io_pu_select[20] padframe/mprj_io_schmitt_select[20] padframe/mprj_io_slew_select[20]
+ gpio_control_in_2\[1\]/resetn gpio_control_in_2\[0\]/resetn gpio_control_in_2\[1\]/serial_clock
+ gpio_control_in_2\[0\]/serial_clock gpio_control_in_2\[1\]/serial_data_in gpio_control_in_2\[0\]/serial_data_in
+ gpio_control_in_2\[1\]/serial_load gpio_control_in_2\[0\]/serial_load mprj/io_in[20]
+ mprj/io_oeb[20] mprj/io_out[20] gpio_control_in_2\[1\]/zero gpio_control_block
Xgpio_defaults_block_7 gpio_defaults_block_7/gpio_defaults[0] gpio_defaults_block_7/gpio_defaults[1]
+ gpio_defaults_block_7/gpio_defaults[2] gpio_defaults_block_7/gpio_defaults[3] gpio_defaults_block_7/gpio_defaults[4]
+ gpio_defaults_block_7/gpio_defaults[5] gpio_defaults_block_7/gpio_defaults[6] gpio_defaults_block_7/gpio_defaults[7]
+ gpio_defaults_block_7/gpio_defaults[8] gpio_defaults_block_7/gpio_defaults[9] gpio_defaults_block_7/VDD
+ gpio_defaults_block_7/VSS gpio_defaults_block
Xgpio_control_in_1\[7\] soc/VDD soc/VSS gpio_defaults_block_0/gpio_defaults[0] gpio_defaults_block_0/gpio_defaults[1]
+ gpio_defaults_block_0/gpio_defaults[2] gpio_defaults_block_0/gpio_defaults[3] gpio_defaults_block_0/gpio_defaults[4]
+ gpio_defaults_block_0/gpio_defaults[5] gpio_defaults_block_0/gpio_defaults[6] gpio_defaults_block_0/gpio_defaults[7]
+ gpio_defaults_block_0/gpio_defaults[8] gpio_defaults_block_0/gpio_defaults[9] housekeeping/mgmt_gpio_in[15]
+ gpio_control_in_1\[7\]/zero housekeeping/mgmt_gpio_out[15] gpio_control_in_1\[7\]/one
+ padframe/mprj_io_drive_sel[30] padframe/mprj_io_drive_sel[31] padframe/mprj_io_in[15]
+ padframe/mprj_io_inen[15] padframe/mprj_io_out[15] padframe/mprj_io_outen[15] padframe/mprj_io_pd_select[15]
+ padframe/mprj_io_pu_select[15] padframe/mprj_io_schmitt_select[15] padframe/mprj_io_slew_select[15]
+ gpio_control_in_1\[7\]/resetn gpio_control_in_1\[8\]/resetn gpio_control_in_1\[7\]/serial_clock
+ gpio_control_in_1\[8\]/serial_clock gpio_control_in_1\[7\]/serial_data_in gpio_control_in_1\[8\]/serial_data_in
+ gpio_control_in_1\[7\]/serial_load gpio_control_in_1\[8\]/serial_load mprj/io_in[15]
+ mprj/io_oeb[15] mprj/io_out[15] gpio_control_in_1\[7\]/zero gpio_control_block
Xgpio_defaults_block_8 gpio_defaults_block_8/gpio_defaults[0] gpio_defaults_block_8/gpio_defaults[1]
+ gpio_defaults_block_8/gpio_defaults[2] gpio_defaults_block_8/gpio_defaults[3] gpio_defaults_block_8/gpio_defaults[4]
+ gpio_defaults_block_8/gpio_defaults[5] gpio_defaults_block_8/gpio_defaults[6] gpio_defaults_block_8/gpio_defaults[7]
+ gpio_defaults_block_8/gpio_defaults[8] gpio_defaults_block_8/gpio_defaults[9] gpio_defaults_block_8/VDD
+ gpio_defaults_block_8/VSS gpio_defaults_block
Xgpio_control_in_1a\[4\] soc/VDD soc/VSS gpio_defaults_block_26/gpio_defaults[0] gpio_defaults_block_26/gpio_defaults[1]
+ gpio_defaults_block_26/gpio_defaults[2] gpio_defaults_block_26/gpio_defaults[3]
+ gpio_defaults_block_26/gpio_defaults[4] gpio_defaults_block_26/gpio_defaults[5]
+ gpio_defaults_block_26/gpio_defaults[6] gpio_defaults_block_26/gpio_defaults[7]
+ gpio_defaults_block_26/gpio_defaults[8] gpio_defaults_block_26/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[6] gpio_control_in_1a\[4\]/zero housekeeping/mgmt_gpio_out[6]
+ gpio_control_in_1a\[4\]/one padframe/mprj_io_drive_sel[13] padframe/mprj_io_drive_sel[12]
+ padframe/mprj_io_in[6] padframe/mprj_io_inen[6] padframe/mprj_io_out[6] padframe/mprj_io_outen[6]
+ padframe/mprj_io_pd_select[6] padframe/mprj_io_pu_select[6] padframe/mprj_io_schmitt_select[6]
+ padframe/mprj_io_slew_select[6] gpio_control_in_1a\[4\]/resetn gpio_control_in_1a\[5\]/resetn
+ gpio_control_in_1a\[4\]/serial_clock gpio_control_in_1a\[5\]/serial_clock gpio_control_in_1a\[4\]/serial_data_in
+ gpio_control_in_1a\[5\]/serial_data_in gpio_control_in_1a\[4\]/serial_load gpio_control_in_1a\[5\]/serial_load
+ mprj/io_in[6] mprj/io_oeb[6] mprj/io_out[6] gpio_control_in_1a\[4\]/zero gpio_control_block
Xmgmt_buffers soc/VDD soc/VSS soc/core_clk clock_ctrl/user_clk soc/core_rstn mprj/la_data_in[0]
+ mprj/la_data_in[10] mprj/la_data_in[11] mprj/la_data_in[12] mprj/la_data_in[13]
+ mprj/la_data_in[14] mprj/la_data_in[15] mprj/la_data_in[16] mprj/la_data_in[17]
+ mprj/la_data_in[18] mprj/la_data_in[19] mprj/la_data_in[1] mprj/la_data_in[20] mprj/la_data_in[21]
+ mprj/la_data_in[22] mprj/la_data_in[23] mprj/la_data_in[24] mprj/la_data_in[25]
+ mprj/la_data_in[26] mprj/la_data_in[27] mprj/la_data_in[28] mprj/la_data_in[29]
+ mprj/la_data_in[2] mprj/la_data_in[30] mprj/la_data_in[31] mprj/la_data_in[32] mprj/la_data_in[33]
+ mprj/la_data_in[34] mprj/la_data_in[35] mprj/la_data_in[36] mprj/la_data_in[37]
+ mprj/la_data_in[38] mprj/la_data_in[39] mprj/la_data_in[3] mprj/la_data_in[40] mprj/la_data_in[41]
+ mprj/la_data_in[42] mprj/la_data_in[43] mprj/la_data_in[44] mprj/la_data_in[45]
+ mprj/la_data_in[46] mprj/la_data_in[47] mprj/la_data_in[48] mprj/la_data_in[49]
+ mprj/la_data_in[4] mprj/la_data_in[50] mprj/la_data_in[51] mprj/la_data_in[52] mprj/la_data_in[53]
+ mprj/la_data_in[54] mprj/la_data_in[55] mprj/la_data_in[56] mprj/la_data_in[57]
+ mprj/la_data_in[58] mprj/la_data_in[59] mprj/la_data_in[5] mprj/la_data_in[60] mprj/la_data_in[61]
+ mprj/la_data_in[62] mprj/la_data_in[63] mprj/la_data_in[6] mprj/la_data_in[7] mprj/la_data_in[8]
+ mprj/la_data_in[9] soc/la_input[0] soc/la_input[10] soc/la_input[11] soc/la_input[12]
+ soc/la_input[13] soc/la_input[14] soc/la_input[15] soc/la_input[16] soc/la_input[17]
+ soc/la_input[18] soc/la_input[19] soc/la_input[1] soc/la_input[20] soc/la_input[21]
+ soc/la_input[22] soc/la_input[23] soc/la_input[24] soc/la_input[25] soc/la_input[26]
+ soc/la_input[27] soc/la_input[28] soc/la_input[29] soc/la_input[2] soc/la_input[30]
+ soc/la_input[31] soc/la_input[32] soc/la_input[33] soc/la_input[34] soc/la_input[35]
+ soc/la_input[36] soc/la_input[37] soc/la_input[38] soc/la_input[39] soc/la_input[3]
+ soc/la_input[40] soc/la_input[41] soc/la_input[42] soc/la_input[43] soc/la_input[44]
+ soc/la_input[45] soc/la_input[46] soc/la_input[47] soc/la_input[48] soc/la_input[49]
+ soc/la_input[4] soc/la_input[50] soc/la_input[51] soc/la_input[52] soc/la_input[53]
+ soc/la_input[54] soc/la_input[55] soc/la_input[56] soc/la_input[57] soc/la_input[58]
+ soc/la_input[59] soc/la_input[5] soc/la_input[60] soc/la_input[61] soc/la_input[62]
+ soc/la_input[63] soc/la_input[6] soc/la_input[7] soc/la_input[8] soc/la_input[9]
+ mprj/la_data_out[0] mprj/la_data_out[10] mprj/la_data_out[11] mprj/la_data_out[12]
+ mprj/la_data_out[13] mprj/la_data_out[14] mprj/la_data_out[15] mprj/la_data_out[16]
+ mprj/la_data_out[17] mprj/la_data_out[18] mprj/la_data_out[19] mprj/la_data_out[1]
+ mprj/la_data_out[20] mprj/la_data_out[21] mprj/la_data_out[22] mprj/la_data_out[23]
+ mprj/la_data_out[24] mprj/la_data_out[25] mprj/la_data_out[26] mprj/la_data_out[27]
+ mprj/la_data_out[28] mprj/la_data_out[29] mprj/la_data_out[2] mprj/la_data_out[30]
+ mprj/la_data_out[31] mprj/la_data_out[32] mprj/la_data_out[33] mprj/la_data_out[34]
+ mprj/la_data_out[35] mprj/la_data_out[36] mprj/la_data_out[37] mprj/la_data_out[38]
+ mprj/la_data_out[39] mprj/la_data_out[3] mprj/la_data_out[40] mprj/la_data_out[41]
+ mprj/la_data_out[42] mprj/la_data_out[43] mprj/la_data_out[44] mprj/la_data_out[45]
+ mprj/la_data_out[46] mprj/la_data_out[47] mprj/la_data_out[48] mprj/la_data_out[49]
+ mprj/la_data_out[4] mprj/la_data_out[50] mprj/la_data_out[51] mprj/la_data_out[52]
+ mprj/la_data_out[53] mprj/la_data_out[54] mprj/la_data_out[55] mprj/la_data_out[56]
+ mprj/la_data_out[57] mprj/la_data_out[58] mprj/la_data_out[59] mprj/la_data_out[5]
+ mprj/la_data_out[60] mprj/la_data_out[61] mprj/la_data_out[62] mprj/la_data_out[63]
+ mprj/la_data_out[6] mprj/la_data_out[7] mprj/la_data_out[8] mprj/la_data_out[9]
+ soc/la_output[0] soc/la_output[10] soc/la_output[11] soc/la_output[12] soc/la_output[13]
+ soc/la_output[14] soc/la_output[15] soc/la_output[16] soc/la_output[17] soc/la_output[18]
+ soc/la_output[19] soc/la_output[1] soc/la_output[20] soc/la_output[21] soc/la_output[22]
+ soc/la_output[23] soc/la_output[24] soc/la_output[25] soc/la_output[26] soc/la_output[27]
+ soc/la_output[28] soc/la_output[29] soc/la_output[2] soc/la_output[30] soc/la_output[31]
+ soc/la_output[32] soc/la_output[33] soc/la_output[34] soc/la_output[35] soc/la_output[36]
+ soc/la_output[37] soc/la_output[38] soc/la_output[39] soc/la_output[3] soc/la_output[40]
+ soc/la_output[41] soc/la_output[42] soc/la_output[43] soc/la_output[44] soc/la_output[45]
+ soc/la_output[46] soc/la_output[47] soc/la_output[48] soc/la_output[49] soc/la_output[4]
+ soc/la_output[50] soc/la_output[51] soc/la_output[52] soc/la_output[53] soc/la_output[54]
+ soc/la_output[55] soc/la_output[56] soc/la_output[57] soc/la_output[58] soc/la_output[59]
+ soc/la_output[5] soc/la_output[60] soc/la_output[61] soc/la_output[62] soc/la_output[63]
+ soc/la_output[6] soc/la_output[7] soc/la_output[8] soc/la_output[9] soc/la_iena[0]
+ soc/la_iena[10] soc/la_iena[11] soc/la_iena[12] soc/la_iena[13] soc/la_iena[14]
+ soc/la_iena[15] soc/la_iena[16] soc/la_iena[17] soc/la_iena[18] soc/la_iena[19]
+ soc/la_iena[1] soc/la_iena[20] soc/la_iena[21] soc/la_iena[22] soc/la_iena[23] soc/la_iena[24]
+ soc/la_iena[25] soc/la_iena[26] soc/la_iena[27] soc/la_iena[28] soc/la_iena[29]
+ soc/la_iena[2] soc/la_iena[30] soc/la_iena[31] soc/la_iena[32] soc/la_iena[33] soc/la_iena[34]
+ soc/la_iena[35] soc/la_iena[36] soc/la_iena[37] soc/la_iena[38] soc/la_iena[39]
+ soc/la_iena[3] soc/la_iena[40] soc/la_iena[41] soc/la_iena[42] soc/la_iena[43] soc/la_iena[44]
+ soc/la_iena[45] soc/la_iena[46] soc/la_iena[47] soc/la_iena[48] soc/la_iena[49]
+ soc/la_iena[4] soc/la_iena[50] soc/la_iena[51] soc/la_iena[52] soc/la_iena[53] soc/la_iena[54]
+ soc/la_iena[55] soc/la_iena[56] soc/la_iena[57] soc/la_iena[58] soc/la_iena[59]
+ soc/la_iena[5] soc/la_iena[60] soc/la_iena[61] soc/la_iena[62] soc/la_iena[63] soc/la_iena[6]
+ soc/la_iena[7] soc/la_iena[8] soc/la_iena[9] mprj/la_oenb[0] mprj/la_oenb[10] mprj/la_oenb[11]
+ mprj/la_oenb[12] mprj/la_oenb[13] mprj/la_oenb[14] mprj/la_oenb[15] mprj/la_oenb[16]
+ mprj/la_oenb[17] mprj/la_oenb[18] mprj/la_oenb[19] mprj/la_oenb[1] mprj/la_oenb[20]
+ mprj/la_oenb[21] mprj/la_oenb[22] mprj/la_oenb[23] mprj/la_oenb[24] mprj/la_oenb[25]
+ mprj/la_oenb[26] mprj/la_oenb[27] mprj/la_oenb[28] mprj/la_oenb[29] mprj/la_oenb[2]
+ mprj/la_oenb[30] mprj/la_oenb[31] mprj/la_oenb[32] mprj/la_oenb[33] mprj/la_oenb[34]
+ mprj/la_oenb[35] mprj/la_oenb[36] mprj/la_oenb[37] mprj/la_oenb[38] mprj/la_oenb[39]
+ mprj/la_oenb[3] mprj/la_oenb[40] mprj/la_oenb[41] mprj/la_oenb[42] mprj/la_oenb[43]
+ mprj/la_oenb[44] mprj/la_oenb[45] mprj/la_oenb[46] mprj/la_oenb[47] mprj/la_oenb[48]
+ mprj/la_oenb[49] mprj/la_oenb[4] mprj/la_oenb[50] mprj/la_oenb[51] mprj/la_oenb[52]
+ mprj/la_oenb[53] mprj/la_oenb[54] mprj/la_oenb[55] mprj/la_oenb[56] mprj/la_oenb[57]
+ mprj/la_oenb[58] mprj/la_oenb[59] mprj/la_oenb[5] mprj/la_oenb[60] mprj/la_oenb[61]
+ mprj/la_oenb[62] mprj/la_oenb[63] mprj/la_oenb[6] mprj/la_oenb[7] mprj/la_oenb[8]
+ mprj/la_oenb[9] soc/la_oenb[0] soc/la_oenb[10] soc/la_oenb[11] soc/la_oenb[12] soc/la_oenb[13]
+ soc/la_oenb[14] soc/la_oenb[15] soc/la_oenb[16] soc/la_oenb[17] soc/la_oenb[18]
+ soc/la_oenb[19] soc/la_oenb[1] soc/la_oenb[20] soc/la_oenb[21] soc/la_oenb[22] soc/la_oenb[23]
+ soc/la_oenb[24] soc/la_oenb[25] soc/la_oenb[26] soc/la_oenb[27] soc/la_oenb[28]
+ soc/la_oenb[29] soc/la_oenb[2] soc/la_oenb[30] soc/la_oenb[31] soc/la_oenb[32] soc/la_oenb[33]
+ soc/la_oenb[34] soc/la_oenb[35] soc/la_oenb[36] soc/la_oenb[37] soc/la_oenb[38]
+ soc/la_oenb[39] soc/la_oenb[3] soc/la_oenb[40] soc/la_oenb[41] soc/la_oenb[42] soc/la_oenb[43]
+ soc/la_oenb[44] soc/la_oenb[45] soc/la_oenb[46] soc/la_oenb[47] soc/la_oenb[48]
+ soc/la_oenb[49] soc/la_oenb[4] soc/la_oenb[50] soc/la_oenb[51] soc/la_oenb[52] soc/la_oenb[53]
+ soc/la_oenb[54] soc/la_oenb[55] soc/la_oenb[56] soc/la_oenb[57] soc/la_oenb[58]
+ soc/la_oenb[59] soc/la_oenb[5] soc/la_oenb[60] soc/la_oenb[61] soc/la_oenb[62] soc/la_oenb[63]
+ soc/la_oenb[6] soc/la_oenb[7] soc/la_oenb[8] soc/la_oenb[9] soc/mprj_ack_i mprj/wbs_ack_o
+ soc/mprj_adr_o[0] soc/mprj_adr_o[10] soc/mprj_adr_o[11] soc/mprj_adr_o[12] soc/mprj_adr_o[13]
+ soc/mprj_adr_o[14] soc/mprj_adr_o[15] soc/mprj_adr_o[16] soc/mprj_adr_o[17] soc/mprj_adr_o[18]
+ soc/mprj_adr_o[19] soc/mprj_adr_o[1] soc/mprj_adr_o[20] soc/mprj_adr_o[21] soc/mprj_adr_o[22]
+ soc/mprj_adr_o[23] soc/mprj_adr_o[24] soc/mprj_adr_o[25] soc/mprj_adr_o[26] soc/mprj_adr_o[27]
+ soc/mprj_adr_o[28] soc/mprj_adr_o[29] soc/mprj_adr_o[2] soc/mprj_adr_o[30] soc/mprj_adr_o[31]
+ soc/mprj_adr_o[3] soc/mprj_adr_o[4] soc/mprj_adr_o[5] soc/mprj_adr_o[6] soc/mprj_adr_o[7]
+ soc/mprj_adr_o[8] soc/mprj_adr_o[9] mprj/wbs_adr_i[0] mprj/wbs_adr_i[10] mprj/wbs_adr_i[11]
+ mprj/wbs_adr_i[12] mprj/wbs_adr_i[13] mprj/wbs_adr_i[14] mprj/wbs_adr_i[15] mprj/wbs_adr_i[16]
+ mprj/wbs_adr_i[17] mprj/wbs_adr_i[18] mprj/wbs_adr_i[19] mprj/wbs_adr_i[1] mprj/wbs_adr_i[20]
+ mprj/wbs_adr_i[21] mprj/wbs_adr_i[22] mprj/wbs_adr_i[23] mprj/wbs_adr_i[24] mprj/wbs_adr_i[25]
+ mprj/wbs_adr_i[26] mprj/wbs_adr_i[27] mprj/wbs_adr_i[28] mprj/wbs_adr_i[29] mprj/wbs_adr_i[2]
+ mprj/wbs_adr_i[30] mprj/wbs_adr_i[31] mprj/wbs_adr_i[3] mprj/wbs_adr_i[4] mprj/wbs_adr_i[5]
+ mprj/wbs_adr_i[6] mprj/wbs_adr_i[7] mprj/wbs_adr_i[8] mprj/wbs_adr_i[9] soc/mprj_cyc_o
+ mprj/wbs_cyc_i soc/mprj_dat_i[0] soc/mprj_dat_i[10] soc/mprj_dat_i[11] soc/mprj_dat_i[12]
+ soc/mprj_dat_i[13] soc/mprj_dat_i[14] soc/mprj_dat_i[15] soc/mprj_dat_i[16] soc/mprj_dat_i[17]
+ soc/mprj_dat_i[18] soc/mprj_dat_i[19] soc/mprj_dat_i[1] soc/mprj_dat_i[20] soc/mprj_dat_i[21]
+ soc/mprj_dat_i[22] soc/mprj_dat_i[23] soc/mprj_dat_i[24] soc/mprj_dat_i[25] soc/mprj_dat_i[26]
+ soc/mprj_dat_i[27] soc/mprj_dat_i[28] soc/mprj_dat_i[29] soc/mprj_dat_i[2] soc/mprj_dat_i[30]
+ soc/mprj_dat_i[31] soc/mprj_dat_i[3] soc/mprj_dat_i[4] soc/mprj_dat_i[5] soc/mprj_dat_i[6]
+ soc/mprj_dat_i[7] soc/mprj_dat_i[8] soc/mprj_dat_i[9] mprj/wbs_dat_o[0] mprj/wbs_dat_o[10]
+ mprj/wbs_dat_o[11] mprj/wbs_dat_o[12] mprj/wbs_dat_o[13] mprj/wbs_dat_o[14] mprj/wbs_dat_o[15]
+ mprj/wbs_dat_o[16] mprj/wbs_dat_o[17] mprj/wbs_dat_o[18] mprj/wbs_dat_o[19] mprj/wbs_dat_o[1]
+ mprj/wbs_dat_o[20] mprj/wbs_dat_o[21] mprj/wbs_dat_o[22] mprj/wbs_dat_o[23] mprj/wbs_dat_o[24]
+ mprj/wbs_dat_o[25] mprj/wbs_dat_o[26] mprj/wbs_dat_o[27] mprj/wbs_dat_o[28] mprj/wbs_dat_o[29]
+ mprj/wbs_dat_o[2] mprj/wbs_dat_o[30] mprj/wbs_dat_o[31] mprj/wbs_dat_o[3] mprj/wbs_dat_o[4]
+ mprj/wbs_dat_o[5] mprj/wbs_dat_o[6] mprj/wbs_dat_o[7] mprj/wbs_dat_o[8] mprj/wbs_dat_o[9]
+ soc/mprj_dat_o[0] soc/mprj_dat_o[10] soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13]
+ soc/mprj_dat_o[14] soc/mprj_dat_o[15] soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18]
+ soc/mprj_dat_o[19] soc/mprj_dat_o[1] soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22]
+ soc/mprj_dat_o[23] soc/mprj_dat_o[24] soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27]
+ soc/mprj_dat_o[28] soc/mprj_dat_o[29] soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31]
+ soc/mprj_dat_o[3] soc/mprj_dat_o[4] soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7]
+ soc/mprj_dat_o[8] soc/mprj_dat_o[9] mprj/wbs_dat_i[0] mprj/wbs_dat_i[10] mprj/wbs_dat_i[11]
+ mprj/wbs_dat_i[12] mprj/wbs_dat_i[13] mprj/wbs_dat_i[14] mprj/wbs_dat_i[15] mprj/wbs_dat_i[16]
+ mprj/wbs_dat_i[17] mprj/wbs_dat_i[18] mprj/wbs_dat_i[19] mprj/wbs_dat_i[1] mprj/wbs_dat_i[20]
+ mprj/wbs_dat_i[21] mprj/wbs_dat_i[22] mprj/wbs_dat_i[23] mprj/wbs_dat_i[24] mprj/wbs_dat_i[25]
+ mprj/wbs_dat_i[26] mprj/wbs_dat_i[27] mprj/wbs_dat_i[28] mprj/wbs_dat_i[29] mprj/wbs_dat_i[2]
+ mprj/wbs_dat_i[30] mprj/wbs_dat_i[31] mprj/wbs_dat_i[3] mprj/wbs_dat_i[4] mprj/wbs_dat_i[5]
+ mprj/wbs_dat_i[6] mprj/wbs_dat_i[7] mprj/wbs_dat_i[8] mprj/wbs_dat_i[9] soc/mprj_wb_iena
+ soc/mprj_sel_o[0] soc/mprj_sel_o[1] soc/mprj_sel_o[2] soc/mprj_sel_o[3] mprj/wbs_sel_i[0]
+ mprj/wbs_sel_i[1] mprj/wbs_sel_i[2] mprj/wbs_sel_i[3] soc/mprj_stb_o mprj/wbs_stb_i
+ soc/mprj_we_o mprj/wbs_we_i mprj/wb_clk_i mprj/user_clock2 soc/irq[0] soc/irq[1]
+ soc/irq[2] mprj/user_irq[0] mprj/user_irq[1] mprj/user_irq[2] soc/user_irq_ena[0]
+ soc/user_irq_ena[1] soc/user_irq_ena[2] mprj/wb_rst_i mgmt_protect
Xgpio_defaults_block_009_0 gpio_defaults_block_009_0/gpio_defaults[0] gpio_defaults_block_009_0/gpio_defaults[1]
+ gpio_defaults_block_009_0/gpio_defaults[2] gpio_defaults_block_009_0/gpio_defaults[3]
+ gpio_defaults_block_009_0/gpio_defaults[4] gpio_defaults_block_009_0/gpio_defaults[5]
+ gpio_defaults_block_009_0/gpio_defaults[6] gpio_defaults_block_009_0/gpio_defaults[7]
+ gpio_defaults_block_009_0/gpio_defaults[8] gpio_defaults_block_009_0/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block_009
Xgpio_defaults_block_009_1 gpio_defaults_block_009_1/gpio_defaults[0] gpio_defaults_block_009_1/gpio_defaults[1]
+ gpio_defaults_block_009_1/gpio_defaults[2] gpio_defaults_block_009_1/gpio_defaults[3]
+ gpio_defaults_block_009_1/gpio_defaults[4] gpio_defaults_block_009_1/gpio_defaults[5]
+ gpio_defaults_block_009_1/gpio_defaults[6] gpio_defaults_block_009_1/gpio_defaults[7]
+ gpio_defaults_block_009_1/gpio_defaults[8] gpio_defaults_block_009_1/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block_009
Xgpio_defaults_block_9 gpio_defaults_block_9/gpio_defaults[0] gpio_defaults_block_9/gpio_defaults[1]
+ gpio_defaults_block_9/gpio_defaults[2] gpio_defaults_block_9/gpio_defaults[3] gpio_defaults_block_9/gpio_defaults[4]
+ gpio_defaults_block_9/gpio_defaults[5] gpio_defaults_block_9/gpio_defaults[6] gpio_defaults_block_9/gpio_defaults[7]
+ gpio_defaults_block_9/gpio_defaults[8] gpio_defaults_block_9/gpio_defaults[9] gpio_defaults_block_9/VDD
+ gpio_defaults_block_9/VSS gpio_defaults_block
Xgpio_control_in_2\[15\] soc/VDD soc/VSS gpio_defaults_block_29/gpio_defaults[0] gpio_defaults_block_29/gpio_defaults[1]
+ gpio_defaults_block_29/gpio_defaults[2] gpio_defaults_block_29/gpio_defaults[3]
+ gpio_defaults_block_29/gpio_defaults[4] gpio_defaults_block_29/gpio_defaults[5]
+ gpio_defaults_block_29/gpio_defaults[6] gpio_defaults_block_29/gpio_defaults[7]
+ gpio_defaults_block_29/gpio_defaults[8] gpio_defaults_block_29/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[34] gpio_control_in_2\[15\]/zero housekeeping/mgmt_gpio_out[34]
+ gpio_control_in_2\[15\]/one padframe/mprj_io_drive_sel[68] padframe/mprj_io_drive_sel[69]
+ padframe/mprj_io_in[34] padframe/mprj_io_inen[34] padframe/mprj_io_out[34] padframe/mprj_io_outen[34]
+ padframe/mprj_io_pd_select[34] padframe/mprj_io_pu_select[34] padframe/mprj_io_schmitt_select[34]
+ padframe/mprj_io_slew_select[34] gpio_control_in_2\[15\]/resetn gpio_control_in_2\[14\]/resetn
+ gpio_control_in_2\[15\]/serial_clock gpio_control_in_2\[14\]/serial_clock gpio_control_in_2\[15\]/serial_data_in
+ gpio_control_in_2\[14\]/serial_data_in gpio_control_in_2\[15\]/serial_load gpio_control_in_2\[14\]/serial_load
+ mprj/io_in[34] mprj/io_oeb[34] mprj/io_out[34] gpio_control_in_2\[15\]/zero gpio_control_block
Xgpio_control_bidir_2\[1\] soc/VDD soc/VSS gpio_defaults_block_31/gpio_defaults[0]
+ gpio_defaults_block_31/gpio_defaults[1] gpio_defaults_block_31/gpio_defaults[2]
+ gpio_defaults_block_31/gpio_defaults[3] gpio_defaults_block_31/gpio_defaults[4]
+ gpio_defaults_block_31/gpio_defaults[5] gpio_defaults_block_31/gpio_defaults[6]
+ gpio_defaults_block_31/gpio_defaults[7] gpio_defaults_block_31/gpio_defaults[8]
+ gpio_defaults_block_31/gpio_defaults[9] housekeeping/mgmt_gpio_in[36] housekeeping/mgmt_gpio_oeb[36]
+ housekeeping/mgmt_gpio_out[36] gpio_control_bidir_2\[1\]/one padframe/mprj_io_drive_sel[72]
+ padframe/mprj_io_drive_sel[73] padframe/mprj_io_in[36] padframe/mprj_io_inen[36]
+ padframe/mprj_io_out[36] padframe/mprj_io_outen[36] padframe/mprj_io_pd_select[36]
+ padframe/mprj_io_pu_select[36] padframe/mprj_io_schmitt_select[36] padframe/mprj_io_slew_select[36]
+ gpio_control_bidir_2\[1\]/resetn gpio_control_bidir_2\[0\]/resetn gpio_control_bidir_2\[1\]/serial_clock
+ gpio_control_bidir_2\[0\]/serial_clock gpio_control_bidir_2\[1\]/serial_data_in
+ gpio_control_bidir_2\[0\]/serial_data_in gpio_control_bidir_2\[1\]/serial_load gpio_control_bidir_2\[0\]/serial_load
+ mprj/io_in[36] mprj/io_oeb[36] mprj/io_out[36] gpio_control_bidir_2\[1\]/zero gpio_control_block
Xgpio_control_in_1\[5\] soc/VDD soc/VSS gpio_defaults_block_12/gpio_defaults[0] gpio_defaults_block_12/gpio_defaults[1]
+ gpio_defaults_block_12/gpio_defaults[2] gpio_defaults_block_12/gpio_defaults[3]
+ gpio_defaults_block_12/gpio_defaults[4] gpio_defaults_block_12/gpio_defaults[5]
+ gpio_defaults_block_12/gpio_defaults[6] gpio_defaults_block_12/gpio_defaults[7]
+ gpio_defaults_block_12/gpio_defaults[8] gpio_defaults_block_12/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[13] gpio_control_in_1\[5\]/zero housekeeping/mgmt_gpio_out[13]
+ gpio_control_in_1\[5\]/one padframe/mprj_io_drive_sel[26] padframe/mprj_io_drive_sel[27]
+ padframe/mprj_io_in[13] padframe/mprj_io_inen[13] padframe/mprj_io_out[13] padframe/mprj_io_outen[13]
+ padframe/mprj_io_pd_select[13] padframe/mprj_io_pu_select[13] padframe/mprj_io_schmitt_select[13]
+ padframe/mprj_io_slew_select[13] gpio_control_in_1\[5\]/resetn gpio_control_in_1\[6\]/resetn
+ gpio_control_in_1\[5\]/serial_clock gpio_control_in_1\[6\]/serial_clock gpio_control_in_1\[5\]/serial_data_in
+ gpio_control_in_1\[6\]/serial_data_in gpio_control_in_1\[5\]/serial_load gpio_control_in_1\[6\]/serial_load
+ mprj/io_in[13] mprj/io_oeb[13] mprj/io_out[13] gpio_control_in_1\[5\]/zero gpio_control_block
Xgpio_defaults_block_007_0 gpio_control_in_1a\[2\]/gpio_defaults[0] gpio_control_in_1a\[2\]/gpio_defaults[1]
+ gpio_control_in_1a\[2\]/gpio_defaults[2] gpio_control_in_1a\[2\]/gpio_defaults[3]
+ gpio_control_in_1a\[2\]/gpio_defaults[4] gpio_control_in_1a\[2\]/gpio_defaults[5]
+ gpio_control_in_1a\[2\]/gpio_defaults[6] gpio_control_in_1a\[2\]/gpio_defaults[7]
+ gpio_control_in_1a\[2\]/gpio_defaults[8] gpio_control_in_1a\[2\]/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block_007
Xgpio_control_in_2\[13\] soc/VDD soc/VSS gpio_defaults_block_25/gpio_defaults[0] gpio_defaults_block_25/gpio_defaults[1]
+ gpio_defaults_block_25/gpio_defaults[2] gpio_defaults_block_25/gpio_defaults[3]
+ gpio_defaults_block_25/gpio_defaults[4] gpio_defaults_block_25/gpio_defaults[5]
+ gpio_defaults_block_25/gpio_defaults[6] gpio_defaults_block_25/gpio_defaults[7]
+ gpio_defaults_block_25/gpio_defaults[8] gpio_defaults_block_25/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[32] gpio_control_in_2\[13\]/zero housekeeping/mgmt_gpio_out[32]
+ gpio_control_in_2\[13\]/one padframe/mprj_io_drive_sel[64] padframe/mprj_io_drive_sel[65]
+ padframe/mprj_io_in[32] padframe/mprj_io_inen[32] padframe/mprj_io_out[32] padframe/mprj_io_outen[32]
+ padframe/mprj_io_pd_select[32] padframe/mprj_io_pu_select[32] padframe/mprj_io_schmitt_select[32]
+ padframe/mprj_io_slew_select[32] gpio_control_in_2\[13\]/resetn gpio_control_in_2\[12\]/resetn
+ gpio_control_in_2\[13\]/serial_clock gpio_control_in_2\[12\]/serial_clock gpio_control_in_2\[13\]/serial_data_in
+ gpio_control_in_2\[12\]/serial_data_in gpio_control_in_2\[13\]/serial_load gpio_control_in_2\[12\]/serial_load
+ mprj/io_in[32] mprj/io_oeb[32] mprj/io_out[32] gpio_control_in_2\[13\]/zero gpio_control_block
Xgpio_control_in_1a\[2\] soc/VDD soc/VSS gpio_control_in_1a\[2\]/gpio_defaults[0]
+ gpio_control_in_1a\[2\]/gpio_defaults[1] gpio_control_in_1a\[2\]/gpio_defaults[2]
+ gpio_control_in_1a\[2\]/gpio_defaults[3] gpio_control_in_1a\[2\]/gpio_defaults[4]
+ gpio_control_in_1a\[2\]/gpio_defaults[5] gpio_control_in_1a\[2\]/gpio_defaults[6]
+ gpio_control_in_1a\[2\]/gpio_defaults[7] gpio_control_in_1a\[2\]/gpio_defaults[8]
+ gpio_control_in_1a\[2\]/gpio_defaults[9] housekeeping/mgmt_gpio_in[4] gpio_control_in_1a\[2\]/zero
+ housekeeping/mgmt_gpio_out[4] gpio_control_in_1a\[2\]/one padframe/mprj_io_drive_sel[9]
+ padframe/mprj_io_drive_sel[8] padframe/mprj_io_in[4] padframe/mprj_io_inen[4] padframe/mprj_io_out[4]
+ padframe/mprj_io_outen[4] padframe/mprj_io_pd_select[4] padframe/mprj_io_pu_select[4]
+ padframe/mprj_io_schmitt_select[4] padframe/mprj_io_slew_select[4] gpio_control_in_1a\[2\]/resetn
+ gpio_control_in_1a\[3\]/resetn gpio_control_in_1a\[2\]/serial_clock gpio_control_in_1a\[3\]/serial_clock
+ gpio_control_in_1a\[2\]/serial_data_in gpio_control_in_1a\[3\]/serial_data_in gpio_control_in_1a\[2\]/serial_load
+ gpio_control_in_1a\[3\]/serial_load mprj/io_in[4] mprj/io_oeb[4] mprj/io_out[4]
+ gpio_control_in_1a\[2\]/zero gpio_control_block
Xgpio_defaults_block_007_1 gpio_control_in_1a\[1\]/gpio_defaults[0] gpio_control_in_1a\[1\]/gpio_defaults[1]
+ gpio_control_in_1a\[1\]/gpio_defaults[2] gpio_control_in_1a\[1\]/gpio_defaults[3]
+ gpio_control_in_1a\[1\]/gpio_defaults[4] gpio_control_in_1a\[1\]/gpio_defaults[5]
+ gpio_control_in_1a\[1\]/gpio_defaults[6] gpio_control_in_1a\[1\]/gpio_defaults[7]
+ gpio_control_in_1a\[1\]/gpio_defaults[8] gpio_control_in_1a\[1\]/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block_007
Xgpio_control_in_2\[8\] soc/VDD soc/VSS gpio_defaults_block_19/gpio_defaults[0] gpio_defaults_block_19/gpio_defaults[1]
+ gpio_defaults_block_19/gpio_defaults[2] gpio_defaults_block_19/gpio_defaults[3]
+ gpio_defaults_block_19/gpio_defaults[4] gpio_defaults_block_19/gpio_defaults[5]
+ gpio_defaults_block_19/gpio_defaults[6] gpio_defaults_block_19/gpio_defaults[7]
+ gpio_defaults_block_19/gpio_defaults[8] gpio_defaults_block_19/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[27] gpio_control_in_2\[8\]/zero housekeeping/mgmt_gpio_out[27]
+ gpio_control_in_2\[8\]/one padframe/mprj_io_drive_sel[54] padframe/mprj_io_drive_sel[55]
+ padframe/mprj_io_in[27] padframe/mprj_io_inen[27] padframe/mprj_io_out[27] padframe/mprj_io_outen[27]
+ padframe/mprj_io_pd_select[27] padframe/mprj_io_pu_select[27] padframe/mprj_io_schmitt_select[27]
+ padframe/mprj_io_slew_select[27] gpio_control_in_2\[8\]/resetn gpio_control_in_2\[7\]/resetn
+ gpio_control_in_2\[8\]/serial_clock gpio_control_in_2\[7\]/serial_clock gpio_control_in_2\[8\]/serial_data_in
+ gpio_control_in_2\[7\]/serial_data_in gpio_control_in_2\[8\]/serial_load gpio_control_in_2\[7\]/serial_load
+ mprj/io_in[27] mprj/io_oeb[27] mprj/io_out[27] gpio_control_in_2\[8\]/zero gpio_control_block
Xgpio_defaults_block_007_2 gpio_control_in_1a\[0\]/gpio_defaults[0] gpio_control_in_1a\[0\]/gpio_defaults[1]
+ gpio_control_in_1a\[0\]/gpio_defaults[2] gpio_control_in_1a\[0\]/gpio_defaults[3]
+ gpio_control_in_1a\[0\]/gpio_defaults[4] gpio_control_in_1a\[0\]/gpio_defaults[5]
+ gpio_control_in_1a\[0\]/gpio_defaults[6] gpio_control_in_1a\[0\]/gpio_defaults[7]
+ gpio_control_in_1a\[0\]/gpio_defaults[8] gpio_control_in_1a\[0\]/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block_007
Xgpio_control_in_1\[3\] soc/VDD soc/VSS gpio_defaults_block_15/gpio_defaults[0] gpio_defaults_block_15/gpio_defaults[1]
+ gpio_defaults_block_15/gpio_defaults[2] gpio_defaults_block_15/gpio_defaults[3]
+ gpio_defaults_block_15/gpio_defaults[4] gpio_defaults_block_15/gpio_defaults[5]
+ gpio_defaults_block_15/gpio_defaults[6] gpio_defaults_block_15/gpio_defaults[7]
+ gpio_defaults_block_15/gpio_defaults[8] gpio_defaults_block_15/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[11] gpio_control_in_1\[3\]/zero housekeeping/mgmt_gpio_out[11]
+ gpio_control_in_1\[3\]/one padframe/mprj_io_drive_sel[23] padframe/mprj_io_drive_sel[22]
+ padframe/mprj_io_in[11] padframe/mprj_io_inen[11] padframe/mprj_io_out[11] padframe/mprj_io_outen[11]
+ padframe/mprj_io_pd_select[11] padframe/mprj_io_pu_select[11] padframe/mprj_io_schmitt_select[11]
+ padframe/mprj_io_slew_select[11] gpio_control_in_1\[3\]/resetn gpio_control_in_1\[4\]/resetn
+ gpio_control_in_1\[3\]/serial_clock gpio_control_in_1\[4\]/serial_clock gpio_control_in_1\[3\]/serial_data_in
+ gpio_control_in_1\[4\]/serial_data_in gpio_control_in_1\[3\]/serial_load gpio_control_in_1\[4\]/serial_load
+ mprj/io_in[11] mprj/io_oeb[11] mprj/io_out[11] gpio_control_in_1\[3\]/zero gpio_control_block
Xgpio_control_in_2\[11\] soc/VDD soc/VSS gpio_defaults_block_23/gpio_defaults[0] gpio_defaults_block_23/gpio_defaults[1]
+ gpio_defaults_block_23/gpio_defaults[2] gpio_defaults_block_23/gpio_defaults[3]
+ gpio_defaults_block_23/gpio_defaults[4] gpio_defaults_block_23/gpio_defaults[5]
+ gpio_defaults_block_23/gpio_defaults[6] gpio_defaults_block_23/gpio_defaults[7]
+ gpio_defaults_block_23/gpio_defaults[8] gpio_defaults_block_23/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[30] gpio_control_in_2\[11\]/zero housekeeping/mgmt_gpio_out[30]
+ gpio_control_in_2\[11\]/one padframe/mprj_io_drive_sel[63] padframe/mprj_io_drive_sel[61]
+ padframe/mprj_io_in[30] padframe/mprj_io_inen[30] padframe/mprj_io_out[30] padframe/mprj_io_outen[30]
+ padframe/mprj_io_pd_select[30] padframe/mprj_io_pu_select[30] padframe/mprj_io_schmitt_select[30]
+ padframe/mprj_io_slew_select[30] gpio_control_in_2\[11\]/resetn gpio_control_in_2\[10\]/resetn
+ gpio_control_in_2\[11\]/serial_clock gpio_control_in_2\[10\]/serial_clock gpio_control_in_2\[11\]/serial_data_in
+ gpio_control_in_2\[10\]/serial_data_in gpio_control_in_2\[11\]/serial_load gpio_control_in_2\[10\]/serial_load
+ mprj/io_in[30] mprj/io_oeb[30] mprj/io_out[30] gpio_control_in_2\[11\]/zero gpio_control_block
Xgpio_control_in_1a\[0\] soc/VDD soc/VSS gpio_control_in_1a\[0\]/gpio_defaults[0]
+ gpio_control_in_1a\[0\]/gpio_defaults[1] gpio_control_in_1a\[0\]/gpio_defaults[2]
+ gpio_control_in_1a\[0\]/gpio_defaults[3] gpio_control_in_1a\[0\]/gpio_defaults[4]
+ gpio_control_in_1a\[0\]/gpio_defaults[5] gpio_control_in_1a\[0\]/gpio_defaults[6]
+ gpio_control_in_1a\[0\]/gpio_defaults[7] gpio_control_in_1a\[0\]/gpio_defaults[8]
+ gpio_control_in_1a\[0\]/gpio_defaults[9] housekeeping/mgmt_gpio_in[2] gpio_control_in_1a\[0\]/zero
+ housekeeping/mgmt_gpio_out[2] gpio_control_in_1a\[0\]/one padframe/mprj_io_drive_sel[5]
+ padframe/mprj_io_drive_sel[4] padframe/mprj_io_in[2] padframe/mprj_io_inen[2] padframe/mprj_io_out[2]
+ padframe/mprj_io_outen[2] padframe/mprj_io_pd_select[2] padframe/mprj_io_pu_select[2]
+ padframe/mprj_io_schmitt_select[2] padframe/mprj_io_slew_select[2] gpio_control_in_1a\[0\]/resetn
+ gpio_control_in_1a\[1\]/resetn gpio_control_in_1a\[0\]/serial_clock gpio_control_in_1a\[1\]/serial_clock
+ gpio_control_in_1a\[0\]/serial_data_in gpio_control_in_1a\[1\]/serial_data_in gpio_control_in_1a\[0\]/serial_load
+ gpio_control_in_1a\[1\]/serial_load mprj/io_in[2] mprj/io_oeb[2] mprj/io_out[2]
+ gpio_control_in_1a\[0\]/zero gpio_control_block
Xgpio_control_in_2\[6\] soc/VDD soc/VSS gpio_defaults_block_14/gpio_defaults[0] gpio_defaults_block_14/gpio_defaults[1]
+ gpio_defaults_block_14/gpio_defaults[2] gpio_defaults_block_14/gpio_defaults[3]
+ gpio_defaults_block_14/gpio_defaults[4] gpio_defaults_block_14/gpio_defaults[5]
+ gpio_defaults_block_14/gpio_defaults[6] gpio_defaults_block_14/gpio_defaults[7]
+ gpio_defaults_block_14/gpio_defaults[8] gpio_defaults_block_14/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[25] gpio_control_in_2\[6\]/zero housekeeping/mgmt_gpio_out[25]
+ gpio_control_in_2\[6\]/one padframe/mprj_io_drive_sel[525] padframe/mprj_io_drive_sel[51]
+ padframe/mprj_io_in[25] padframe/mprj_io_inen[25] padframe/mprj_io_out[25] padframe/mprj_io_outen[25]
+ padframe/mprj_io_pd_select[25] padframe/mprj_io_pu_select[25] padframe/mprj_io_schmitt_select[25]
+ padframe/mprj_io_slew_select[25] gpio_control_in_2\[6\]/resetn gpio_control_in_2\[5\]/resetn
+ gpio_control_in_2\[6\]/serial_clock gpio_control_in_2\[5\]/serial_clock gpio_control_in_2\[6\]/serial_data_in
+ gpio_control_in_2\[5\]/serial_data_in gpio_control_in_2\[6\]/serial_load gpio_control_in_2\[5\]/serial_load
+ mprj/io_in[25] mprj/io_oeb[25] mprj/io_out[25] gpio_control_in_2\[6\]/zero gpio_control_block
Xgpio_control_in_1\[1\] soc/VDD soc/VSS gpio_defaults_block_20/gpio_defaults[0] gpio_defaults_block_20/gpio_defaults[1]
+ gpio_defaults_block_20/gpio_defaults[2] gpio_defaults_block_20/gpio_defaults[3]
+ gpio_defaults_block_20/gpio_defaults[4] gpio_defaults_block_20/gpio_defaults[5]
+ gpio_defaults_block_20/gpio_defaults[6] gpio_defaults_block_20/gpio_defaults[7]
+ gpio_defaults_block_20/gpio_defaults[8] gpio_defaults_block_20/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[9] gpio_control_in_1\[1\]/zero housekeeping/mgmt_gpio_out[9]
+ gpio_control_in_1\[1\]/one padframe/mprj_io_drive_sel[19] padframe/mprj_io_drive_sel[18]
+ padframe/mprj_io_in[9] padframe/mprj_io_inen[9] padframe/mprj_io_out[9] padframe/mprj_io_outen[9]
+ padframe/mprj_io_pd_select[9] padframe/mprj_io_pu_select[9] padframe/mprj_io_schmitt_select[9]
+ padframe/mprj_io_slew_select[9] gpio_control_in_1\[1\]/resetn gpio_control_in_1\[2\]/resetn
+ gpio_control_in_1\[1\]/serial_clock gpio_control_in_1\[2\]/serial_clock gpio_control_in_1\[1\]/serial_data_in
+ gpio_control_in_1\[2\]/serial_data_in gpio_control_in_1\[1\]/serial_load gpio_control_in_1\[2\]/serial_load
+ mprj/io_in[9] mprj/io_oeb[9] mprj/io_out[9] gpio_control_in_1\[1\]/zero gpio_control_block
Xmprj mprj/io_in[0] mprj/io_in[10] mprj/io_in[11] mprj/io_in[12] mprj/io_in[13] mprj/io_in[14]
+ mprj/io_in[15] mprj/io_in[16] mprj/io_in[17] mprj/io_in[18] mprj/io_in[19] mprj/io_in[1]
+ mprj/io_in[20] mprj/io_in[21] mprj/io_in[22] mprj/io_in[23] mprj/io_in[24] mprj/io_in[25]
+ mprj/io_in[26] mprj/io_in[27] mprj/io_in[28] mprj/io_in[29] mprj/io_in[2] mprj/io_in[30]
+ mprj/io_in[31] mprj/io_in[32] mprj/io_in[33] mprj/io_in[34] mprj/io_in[35] mprj/io_in[36]
+ mprj/io_in[37] mprj/io_in[3] mprj/io_in[4] mprj/io_in[5] mprj/io_in[6] mprj/io_in[7]
+ mprj/io_in[8] mprj/io_in[9] mprj/io_oeb[0] mprj/io_oeb[10] mprj/io_oeb[11] mprj/io_oeb[12]
+ mprj/io_oeb[13] mprj/io_oeb[14] mprj/io_oeb[15] mprj/io_oeb[16] mprj/io_oeb[17]
+ mprj/io_oeb[18] mprj/io_oeb[19] mprj/io_oeb[1] mprj/io_oeb[20] mprj/io_oeb[21] mprj/io_oeb[22]
+ mprj/io_oeb[23] mprj/io_oeb[24] mprj/io_oeb[25] mprj/io_oeb[26] mprj/io_oeb[27]
+ mprj/io_oeb[28] mprj/io_oeb[29] mprj/io_oeb[2] mprj/io_oeb[30] mprj/io_oeb[31] mprj/io_oeb[32]
+ mprj/io_oeb[33] mprj/io_oeb[34] mprj/io_oeb[35] mprj/io_oeb[36] mprj/io_oeb[37]
+ mprj/io_oeb[3] mprj/io_oeb[4] mprj/io_oeb[5] mprj/io_oeb[6] mprj/io_oeb[7] mprj/io_oeb[8]
+ mprj/io_oeb[9] mprj/io_out[0] mprj/io_out[10] mprj/io_out[11] mprj/io_out[12] mprj/io_out[13]
+ mprj/io_out[14] mprj/io_out[15] mprj/io_out[16] mprj/io_out[17] mprj/io_out[18]
+ mprj/io_out[19] mprj/io_out[1] mprj/io_out[20] mprj/io_out[21] mprj/io_out[22] mprj/io_out[23]
+ mprj/io_out[24] mprj/io_out[25] mprj/io_out[26] mprj/io_out[27] mprj/io_out[28]
+ mprj/io_out[29] mprj/io_out[2] mprj/io_out[30] mprj/io_out[31] mprj/io_out[32] mprj/io_out[33]
+ mprj/io_out[34] mprj/io_out[35] mprj/io_out[36] mprj/io_out[37] mprj/io_out[3] mprj/io_out[4]
+ mprj/io_out[5] mprj/io_out[6] mprj/io_out[7] mprj/io_out[8] mprj/io_out[9] mprj/la_data_in[0]
+ mprj/la_data_in[10] mprj/la_data_in[11] mprj/la_data_in[12] mprj/la_data_in[13]
+ mprj/la_data_in[14] mprj/la_data_in[15] mprj/la_data_in[16] mprj/la_data_in[17]
+ mprj/la_data_in[18] mprj/la_data_in[19] mprj/la_data_in[1] mprj/la_data_in[20] mprj/la_data_in[21]
+ mprj/la_data_in[22] mprj/la_data_in[23] mprj/la_data_in[24] mprj/la_data_in[25]
+ mprj/la_data_in[26] mprj/la_data_in[27] mprj/la_data_in[28] mprj/la_data_in[29]
+ mprj/la_data_in[2] mprj/la_data_in[30] mprj/la_data_in[31] mprj/la_data_in[32] mprj/la_data_in[33]
+ mprj/la_data_in[34] mprj/la_data_in[35] mprj/la_data_in[36] mprj/la_data_in[37]
+ mprj/la_data_in[38] mprj/la_data_in[39] mprj/la_data_in[3] mprj/la_data_in[40] mprj/la_data_in[41]
+ mprj/la_data_in[42] mprj/la_data_in[43] mprj/la_data_in[44] mprj/la_data_in[45]
+ mprj/la_data_in[46] mprj/la_data_in[47] mprj/la_data_in[48] mprj/la_data_in[49]
+ mprj/la_data_in[4] mprj/la_data_in[50] mprj/la_data_in[51] mprj/la_data_in[52] mprj/la_data_in[53]
+ mprj/la_data_in[54] mprj/la_data_in[55] mprj/la_data_in[56] mprj/la_data_in[57]
+ mprj/la_data_in[58] mprj/la_data_in[59] mprj/la_data_in[5] mprj/la_data_in[60] mprj/la_data_in[61]
+ mprj/la_data_in[62] mprj/la_data_in[63] mprj/la_data_in[6] mprj/la_data_in[7] mprj/la_data_in[8]
+ mprj/la_data_in[9] mprj/la_data_out[0] mprj/la_data_out[10] mprj/la_data_out[11]
+ mprj/la_data_out[12] mprj/la_data_out[13] mprj/la_data_out[14] mprj/la_data_out[15]
+ mprj/la_data_out[16] mprj/la_data_out[17] mprj/la_data_out[18] mprj/la_data_out[19]
+ mprj/la_data_out[1] mprj/la_data_out[20] mprj/la_data_out[21] mprj/la_data_out[22]
+ mprj/la_data_out[23] mprj/la_data_out[24] mprj/la_data_out[25] mprj/la_data_out[26]
+ mprj/la_data_out[27] mprj/la_data_out[28] mprj/la_data_out[29] mprj/la_data_out[2]
+ mprj/la_data_out[30] mprj/la_data_out[31] mprj/la_data_out[32] mprj/la_data_out[33]
+ mprj/la_data_out[34] mprj/la_data_out[35] mprj/la_data_out[36] mprj/la_data_out[37]
+ mprj/la_data_out[38] mprj/la_data_out[39] mprj/la_data_out[3] mprj/la_data_out[40]
+ mprj/la_data_out[41] mprj/la_data_out[42] mprj/la_data_out[43] mprj/la_data_out[44]
+ mprj/la_data_out[45] mprj/la_data_out[46] mprj/la_data_out[47] mprj/la_data_out[48]
+ mprj/la_data_out[49] mprj/la_data_out[4] mprj/la_data_out[50] mprj/la_data_out[51]
+ mprj/la_data_out[52] mprj/la_data_out[53] mprj/la_data_out[54] mprj/la_data_out[55]
+ mprj/la_data_out[56] mprj/la_data_out[57] mprj/la_data_out[58] mprj/la_data_out[59]
+ mprj/la_data_out[5] mprj/la_data_out[60] mprj/la_data_out[61] mprj/la_data_out[62]
+ mprj/la_data_out[63] mprj/la_data_out[6] mprj/la_data_out[7] mprj/la_data_out[8]
+ mprj/la_data_out[9] mprj/la_oenb[0] mprj/la_oenb[10] mprj/la_oenb[11] mprj/la_oenb[12]
+ mprj/la_oenb[13] mprj/la_oenb[14] mprj/la_oenb[15] mprj/la_oenb[16] mprj/la_oenb[17]
+ mprj/la_oenb[18] mprj/la_oenb[19] mprj/la_oenb[1] mprj/la_oenb[20] mprj/la_oenb[21]
+ mprj/la_oenb[22] mprj/la_oenb[23] mprj/la_oenb[24] mprj/la_oenb[25] mprj/la_oenb[26]
+ mprj/la_oenb[27] mprj/la_oenb[28] mprj/la_oenb[29] mprj/la_oenb[2] mprj/la_oenb[30]
+ mprj/la_oenb[31] mprj/la_oenb[32] mprj/la_oenb[33] mprj/la_oenb[34] mprj/la_oenb[35]
+ mprj/la_oenb[36] mprj/la_oenb[37] mprj/la_oenb[38] mprj/la_oenb[39] mprj/la_oenb[3]
+ mprj/la_oenb[40] mprj/la_oenb[41] mprj/la_oenb[42] mprj/la_oenb[43] mprj/la_oenb[44]
+ mprj/la_oenb[45] mprj/la_oenb[46] mprj/la_oenb[47] mprj/la_oenb[48] mprj/la_oenb[49]
+ mprj/la_oenb[4] mprj/la_oenb[50] mprj/la_oenb[51] mprj/la_oenb[52] mprj/la_oenb[53]
+ mprj/la_oenb[54] mprj/la_oenb[55] mprj/la_oenb[56] mprj/la_oenb[57] mprj/la_oenb[58]
+ mprj/la_oenb[59] mprj/la_oenb[5] mprj/la_oenb[60] mprj/la_oenb[61] mprj/la_oenb[62]
+ mprj/la_oenb[63] mprj/la_oenb[6] mprj/la_oenb[7] mprj/la_oenb[8] mprj/la_oenb[9]
+ mprj/user_clock2 mprj/user_irq[0] mprj/user_irq[1] mprj/user_irq[2] soc/VDD soc/VSS
+ mprj/wb_clk_i mprj/wb_rst_i mprj/wbs_ack_o mprj/wbs_adr_i[0] mprj/wbs_adr_i[10]
+ mprj/wbs_adr_i[11] mprj/wbs_adr_i[12] mprj/wbs_adr_i[13] mprj/wbs_adr_i[14] mprj/wbs_adr_i[15]
+ mprj/wbs_adr_i[16] mprj/wbs_adr_i[17] mprj/wbs_adr_i[18] mprj/wbs_adr_i[19] mprj/wbs_adr_i[1]
+ mprj/wbs_adr_i[20] mprj/wbs_adr_i[21] mprj/wbs_adr_i[22] mprj/wbs_adr_i[23] mprj/wbs_adr_i[24]
+ mprj/wbs_adr_i[25] mprj/wbs_adr_i[26] mprj/wbs_adr_i[27] mprj/wbs_adr_i[28] mprj/wbs_adr_i[29]
+ mprj/wbs_adr_i[2] mprj/wbs_adr_i[30] mprj/wbs_adr_i[31] mprj/wbs_adr_i[3] mprj/wbs_adr_i[4]
+ mprj/wbs_adr_i[5] mprj/wbs_adr_i[6] mprj/wbs_adr_i[7] mprj/wbs_adr_i[8] mprj/wbs_adr_i[9]
+ mprj/wbs_cyc_i mprj/wbs_dat_i[0] mprj/wbs_dat_i[10] mprj/wbs_dat_i[11] mprj/wbs_dat_i[12]
+ mprj/wbs_dat_i[13] mprj/wbs_dat_i[14] mprj/wbs_dat_i[15] mprj/wbs_dat_i[16] mprj/wbs_dat_i[17]
+ mprj/wbs_dat_i[18] mprj/wbs_dat_i[19] mprj/wbs_dat_i[1] mprj/wbs_dat_i[20] mprj/wbs_dat_i[21]
+ mprj/wbs_dat_i[22] mprj/wbs_dat_i[23] mprj/wbs_dat_i[24] mprj/wbs_dat_i[25] mprj/wbs_dat_i[26]
+ mprj/wbs_dat_i[27] mprj/wbs_dat_i[28] mprj/wbs_dat_i[29] mprj/wbs_dat_i[2] mprj/wbs_dat_i[30]
+ mprj/wbs_dat_i[31] mprj/wbs_dat_i[3] mprj/wbs_dat_i[4] mprj/wbs_dat_i[5] mprj/wbs_dat_i[6]
+ mprj/wbs_dat_i[7] mprj/wbs_dat_i[8] mprj/wbs_dat_i[9] mprj/wbs_dat_o[0] mprj/wbs_dat_o[10]
+ mprj/wbs_dat_o[11] mprj/wbs_dat_o[12] mprj/wbs_dat_o[13] mprj/wbs_dat_o[14] mprj/wbs_dat_o[15]
+ mprj/wbs_dat_o[16] mprj/wbs_dat_o[17] mprj/wbs_dat_o[18] mprj/wbs_dat_o[19] mprj/wbs_dat_o[1]
+ mprj/wbs_dat_o[20] mprj/wbs_dat_o[21] mprj/wbs_dat_o[22] mprj/wbs_dat_o[23] mprj/wbs_dat_o[24]
+ mprj/wbs_dat_o[25] mprj/wbs_dat_o[26] mprj/wbs_dat_o[27] mprj/wbs_dat_o[28] mprj/wbs_dat_o[29]
+ mprj/wbs_dat_o[2] mprj/wbs_dat_o[30] mprj/wbs_dat_o[31] mprj/wbs_dat_o[3] mprj/wbs_dat_o[4]
+ mprj/wbs_dat_o[5] mprj/wbs_dat_o[6] mprj/wbs_dat_o[7] mprj/wbs_dat_o[8] mprj/wbs_dat_o[9]
+ mprj/wbs_sel_i[0] mprj/wbs_sel_i[1] mprj/wbs_sel_i[2] mprj/wbs_sel_i[3] mprj/wbs_stb_i
+ mprj/wbs_we_i user_project_wrapper
Xgpio_control_in_2\[4\] soc/VDD soc/VSS gpio_defaults_block_8/gpio_defaults[0] gpio_defaults_block_8/gpio_defaults[1]
+ gpio_defaults_block_8/gpio_defaults[2] gpio_defaults_block_8/gpio_defaults[3] gpio_defaults_block_8/gpio_defaults[4]
+ gpio_defaults_block_8/gpio_defaults[5] gpio_defaults_block_8/gpio_defaults[6] gpio_defaults_block_8/gpio_defaults[7]
+ gpio_defaults_block_8/gpio_defaults[8] gpio_defaults_block_8/gpio_defaults[9] housekeeping/mgmt_gpio_in[23]
+ gpio_control_in_2\[4\]/zero housekeeping/mgmt_gpio_out[23] gpio_control_in_2\[4\]/one
+ padframe/mprj_io_drive_sel[46] padframe/mprj_io_drive_sel[47] padframe/mprj_io_in[23]
+ padframe/mprj_io_inen[23] padframe/mprj_io_out[23] padframe/mprj_io_outen[23] padframe/mprj_io_pd_select[23]
+ padframe/mprj_io_pu_select[23] padframe/mprj_io_schmitt_select[23] padframe/mprj_io_slew_select[23]
+ gpio_control_in_2\[4\]/resetn gpio_control_in_2\[3\]/resetn gpio_control_in_2\[4\]/serial_clock
+ gpio_control_in_2\[3\]/serial_clock gpio_control_in_2\[4\]/serial_data_in gpio_control_in_2\[3\]/serial_data_in
+ gpio_control_in_2\[4\]/serial_load gpio_control_in_2\[3\]/serial_load mprj/io_in[23]
+ mprj/io_oeb[23] mprj/io_out[23] gpio_control_in_2\[4\]/zero gpio_control_block
Xgpio_control_bidir_1\[1\] soc/VDD soc/VSS gpio_defaults_block_009_0/gpio_defaults[0]
+ gpio_defaults_block_009_0/gpio_defaults[1] gpio_defaults_block_009_0/gpio_defaults[2]
+ gpio_defaults_block_009_0/gpio_defaults[3] gpio_defaults_block_009_0/gpio_defaults[4]
+ gpio_defaults_block_009_0/gpio_defaults[5] gpio_defaults_block_009_0/gpio_defaults[6]
+ gpio_defaults_block_009_0/gpio_defaults[7] gpio_defaults_block_009_0/gpio_defaults[8]
+ gpio_defaults_block_009_0/gpio_defaults[9] housekeeping/mgmt_gpio_in[1] housekeeping/mgmt_gpio_oeb[1]
+ housekeeping/mgmt_gpio_out[1] gpio_control_bidir_1\[1\]/one padframe/mprj_io_drive_sel[2]
+ padframe/mprj_io_drive_sel[3] padframe/mprj_io_in[1] padframe/mprj_io_inen[1] padframe/mprj_io_out[1]
+ padframe/mprj_io_outen[1] padframe/mprj_io_pd_select[1] padframe/mprj_io_pu_select[1]
+ padframe/mprj_io_schmitt_select[1] padframe/mprj_io_slew_select[1] gpio_control_bidir_1\[1\]/resetn
+ gpio_control_in_1a\[0\]/resetn gpio_control_bidir_1\[1\]/serial_clock gpio_control_in_1a\[0\]/serial_clock
+ gpio_control_bidir_1\[1\]/serial_data_in gpio_control_in_1a\[0\]/serial_data_in
+ gpio_control_bidir_1\[1\]/serial_load gpio_control_in_1a\[0\]/serial_load mprj/io_in[1]
+ mprj/io_oeb[1] mprj/io_out[1] gpio_control_bidir_1\[1\]/zero gpio_control_block
Xspare_logic\[2\] soc/VDD soc/VSS spare_logic\[2\]/spare_xfq[0] spare_logic\[2\]/spare_xfq[1]
+ spare_logic\[2\]/spare_xi[0] spare_logic\[2\]/spare_xi[1] spare_logic\[2\]/spare_xi[2]
+ spare_logic\[2\]/spare_xi[3] spare_logic\[2\]/spare_xib spare_logic\[2\]/spare_xmx[0]
+ spare_logic\[2\]/spare_xmx[1] spare_logic\[2\]/spare_xna[0] spare_logic\[2\]/spare_xna[1]
+ spare_logic\[2\]/spare_xno[0] spare_logic\[2\]/spare_xno[1] spare_logic\[2\]/spare_xz[0]
+ spare_logic\[2\]/spare_xz[10] spare_logic\[2\]/spare_xz[11] spare_logic\[2\]/spare_xz[12]
+ spare_logic\[2\]/spare_xz[13] spare_logic\[2\]/spare_xz[14] spare_logic\[2\]/spare_xz[15]
+ spare_logic\[2\]/spare_xz[16] spare_logic\[2\]/spare_xz[17] spare_logic\[2\]/spare_xz[18]
+ spare_logic\[2\]/spare_xz[19] spare_logic\[2\]/spare_xz[1] spare_logic\[2\]/spare_xz[20]
+ spare_logic\[2\]/spare_xz[21] spare_logic\[2\]/spare_xz[22] spare_logic\[2\]/spare_xz[23]
+ spare_logic\[2\]/spare_xz[24] spare_logic\[2\]/spare_xz[25] spare_logic\[2\]/spare_xz[26]
+ spare_logic\[2\]/spare_xz[27] spare_logic\[2\]/spare_xz[28] spare_logic\[2\]/spare_xz[29]
+ spare_logic\[2\]/spare_xz[2] spare_logic\[2\]/spare_xz[30] spare_logic\[2\]/spare_xz[3]
+ spare_logic\[2\]/spare_xz[4] spare_logic\[2\]/spare_xz[5] spare_logic\[2\]/spare_xz[6]
+ spare_logic\[2\]/spare_xz[7] spare_logic\[2\]/spare_xz[8] spare_logic\[2\]/spare_xz[9]
+ spare_logic_block
Xhousekeeping soc/VDD soc/VSS soc/debug_in soc/debug_mode soc/debug_oeb soc/debug_out
+ soc/irq[3] soc/irq[4] soc/irq[5] user_id_value/mask_rev[0] user_id_value/mask_rev[10]
+ user_id_value/mask_rev[11] user_id_value/mask_rev[12] user_id_value/mask_rev[13]
+ user_id_value/mask_rev[14] user_id_value/mask_rev[15] user_id_value/mask_rev[16]
+ user_id_value/mask_rev[17] user_id_value/mask_rev[18] user_id_value/mask_rev[19]
+ user_id_value/mask_rev[1] user_id_value/mask_rev[20] user_id_value/mask_rev[21]
+ user_id_value/mask_rev[22] user_id_value/mask_rev[23] user_id_value/mask_rev[24]
+ user_id_value/mask_rev[25] user_id_value/mask_rev[26] user_id_value/mask_rev[27]
+ user_id_value/mask_rev[28] user_id_value/mask_rev[29] user_id_value/mask_rev[2]
+ user_id_value/mask_rev[30] user_id_value/mask_rev[31] user_id_value/mask_rev[3]
+ user_id_value/mask_rev[4] user_id_value/mask_rev[5] user_id_value/mask_rev[6] user_id_value/mask_rev[7]
+ user_id_value/mask_rev[8] user_id_value/mask_rev[9] housekeeping/mgmt_gpio_in[0]
+ housekeeping/mgmt_gpio_in[10] housekeeping/mgmt_gpio_in[11] housekeeping/mgmt_gpio_in[12]
+ housekeeping/mgmt_gpio_in[13] housekeeping/mgmt_gpio_in[14] housekeeping/mgmt_gpio_in[15]
+ housekeeping/mgmt_gpio_in[16] housekeeping/mgmt_gpio_in[17] housekeeping/mgmt_gpio_in[18]
+ housekeeping/mgmt_gpio_in[19] housekeeping/mgmt_gpio_in[1] housekeeping/mgmt_gpio_in[20]
+ housekeeping/mgmt_gpio_in[21] housekeeping/mgmt_gpio_in[22] housekeeping/mgmt_gpio_in[23]
+ housekeeping/mgmt_gpio_in[24] housekeeping/mgmt_gpio_in[25] housekeeping/mgmt_gpio_in[26]
+ housekeeping/mgmt_gpio_in[27] housekeeping/mgmt_gpio_in[28] housekeeping/mgmt_gpio_in[29]
+ housekeeping/mgmt_gpio_in[2] housekeeping/mgmt_gpio_in[30] housekeeping/mgmt_gpio_in[31]
+ housekeeping/mgmt_gpio_in[32] housekeeping/mgmt_gpio_in[33] housekeeping/mgmt_gpio_in[34]
+ housekeeping/mgmt_gpio_in[35] housekeeping/mgmt_gpio_in[36] housekeeping/mgmt_gpio_in[37]
+ housekeeping/mgmt_gpio_in[3] housekeeping/mgmt_gpio_in[4] housekeeping/mgmt_gpio_in[5]
+ housekeeping/mgmt_gpio_in[6] housekeeping/mgmt_gpio_in[7] housekeeping/mgmt_gpio_in[8]
+ housekeeping/mgmt_gpio_in[9] housekeeping/mgmt_gpio_oeb[0] housekeeping/mgmt_gpio_oeb[10]
+ housekeeping/mgmt_gpio_oeb[11] housekeeping/mgmt_gpio_oeb[12] housekeeping/mgmt_gpio_oeb[13]
+ housekeeping/mgmt_gpio_oeb[14] housekeeping/mgmt_gpio_oeb[15] housekeeping/mgmt_gpio_oeb[16]
+ housekeeping/mgmt_gpio_oeb[17] housekeeping/mgmt_gpio_oeb[18] housekeeping/mgmt_gpio_oeb[19]
+ housekeeping/mgmt_gpio_oeb[1] housekeeping/mgmt_gpio_oeb[20] housekeeping/mgmt_gpio_oeb[21]
+ housekeeping/mgmt_gpio_oeb[22] housekeeping/mgmt_gpio_oeb[23] housekeeping/mgmt_gpio_oeb[24]
+ housekeeping/mgmt_gpio_oeb[25] housekeeping/mgmt_gpio_oeb[26] housekeeping/mgmt_gpio_oeb[27]
+ housekeeping/mgmt_gpio_oeb[28] housekeeping/mgmt_gpio_oeb[29] housekeeping/mgmt_gpio_oeb[2]
+ housekeeping/mgmt_gpio_oeb[30] housekeeping/mgmt_gpio_oeb[31] housekeeping/mgmt_gpio_oeb[32]
+ housekeeping/mgmt_gpio_oeb[33] housekeeping/mgmt_gpio_oeb[34] housekeeping/mgmt_gpio_oeb[35]
+ housekeeping/mgmt_gpio_oeb[36] housekeeping/mgmt_gpio_oeb[37] housekeeping/mgmt_gpio_oeb[3]
+ housekeeping/mgmt_gpio_oeb[4] housekeeping/mgmt_gpio_oeb[5] housekeeping/mgmt_gpio_oeb[6]
+ housekeeping/mgmt_gpio_oeb[7] housekeeping/mgmt_gpio_oeb[8] housekeeping/mgmt_gpio_oeb[9]
+ housekeeping/mgmt_gpio_out[0] housekeeping/mgmt_gpio_out[10] housekeeping/mgmt_gpio_out[11]
+ housekeeping/mgmt_gpio_out[12] housekeeping/mgmt_gpio_out[13] housekeeping/mgmt_gpio_out[14]
+ housekeeping/mgmt_gpio_out[15] housekeeping/mgmt_gpio_out[16] housekeeping/mgmt_gpio_out[17]
+ housekeeping/mgmt_gpio_out[18] housekeeping/mgmt_gpio_out[19] housekeeping/mgmt_gpio_out[1]
+ housekeeping/mgmt_gpio_out[20] housekeeping/mgmt_gpio_out[21] housekeeping/mgmt_gpio_out[22]
+ housekeeping/mgmt_gpio_out[23] housekeeping/mgmt_gpio_out[24] housekeeping/mgmt_gpio_out[25]
+ housekeeping/mgmt_gpio_out[26] housekeeping/mgmt_gpio_out[27] housekeeping/mgmt_gpio_out[28]
+ housekeeping/mgmt_gpio_out[29] housekeeping/mgmt_gpio_out[2] housekeeping/mgmt_gpio_out[30]
+ housekeeping/mgmt_gpio_out[31] housekeeping/mgmt_gpio_out[32] housekeeping/mgmt_gpio_out[33]
+ housekeeping/mgmt_gpio_out[34] housekeeping/mgmt_gpio_out[35] housekeeping/mgmt_gpio_out[36]
+ housekeeping/mgmt_gpio_out[37] housekeeping/mgmt_gpio_out[3] housekeeping/mgmt_gpio_out[4]
+ housekeeping/mgmt_gpio_out[5] housekeeping/mgmt_gpio_out[6] housekeeping/mgmt_gpio_out[7]
+ housekeeping/mgmt_gpio_out[8] housekeeping/mgmt_gpio_out[9] padframe/flash_clk_core
+ padframe/flash_clk_oe_core padframe/flash_csb_core padframe/flash_csb_oe_core padframe/flash_io0_di_core
+ padframe/flash_io0_do_core padframe/flash_io0_ie_core padframe/flash_io0_oe_core
+ padframe/flash_io1_di_core padframe/flash_io1_do_core padframe/flash_io1_ie_core
+ padframe/flash_io1_oe_core clock_ctrl/sel2[0] clock_ctrl/sel2[1] clock_ctrl/sel2[2]
+ clock_ctrl/ext_clk_sel pll/dco pll/div[0] pll/div[1] pll/div[2] pll/div[3] pll/div[4]
+ pll/enable clock_ctrl/sel[0] clock_ctrl/sel[1] clock_ctrl/sel[2] pll/ext_trim[0]
+ pll/ext_trim[10] pll/ext_trim[11] pll/ext_trim[12] pll/ext_trim[13] pll/ext_trim[14]
+ pll/ext_trim[15] pll/ext_trim[16] pll/ext_trim[17] pll/ext_trim[18] pll/ext_trim[19]
+ pll/ext_trim[1] pll/ext_trim[20] pll/ext_trim[21] pll/ext_trim[22] pll/ext_trim[23]
+ pll/ext_trim[24] pll/ext_trim[25] pll/ext_trim[2] pll/ext_trim[3] pll/ext_trim[4]
+ pll/ext_trim[5] pll/ext_trim[6] pll/ext_trim[7] pll/ext_trim[8] pll/ext_trim[9]
+ simple_por_0/porb housekeeping/pwr_ctrl_out soc/qspi_enabled housekeeping/reset
+ soc/ser_rx soc/ser_tx housekeeping/serial_clock housekeeping/serial_data_1 housekeeping/serial_data_2
+ housekeeping/serial_load housekeeping/serial_resetn soc/spi_csb soc/spi_enabled
+ soc/spi_sck soc/spi_sdi soc/spi_sdo soc/spi_sdoenb soc/flash_clk soc/flash_csb soc/flash_io0_di
+ soc/flash_io0_do soc/flash_io0_oeb soc/flash_io1_di soc/flash_io1_do soc/flash_io1_oeb
+ soc/flash_io2_di soc/flash_io2_do soc/flash_io2_oeb soc/flash_io3_di soc/flash_io3_do
+ soc/flash_io3_oeb soc/trap soc/uart_enabled clock_ctrl/user_clk soc/hk_ack_i soc/mprj_adr_o[0]
+ soc/mprj_adr_o[10] soc/mprj_adr_o[11] soc/mprj_adr_o[12] soc/mprj_adr_o[13] soc/mprj_adr_o[14]
+ soc/mprj_adr_o[15] soc/mprj_adr_o[16] soc/mprj_adr_o[17] soc/mprj_adr_o[18] soc/mprj_adr_o[19]
+ soc/mprj_adr_o[1] soc/mprj_adr_o[20] soc/mprj_adr_o[21] soc/mprj_adr_o[22] soc/mprj_adr_o[23]
+ soc/mprj_adr_o[24] soc/mprj_adr_o[25] soc/mprj_adr_o[26] soc/mprj_adr_o[27] soc/mprj_adr_o[28]
+ soc/mprj_adr_o[29] soc/mprj_adr_o[2] soc/mprj_adr_o[30] soc/mprj_adr_o[31] soc/mprj_adr_o[3]
+ soc/mprj_adr_o[4] soc/mprj_adr_o[5] soc/mprj_adr_o[6] soc/mprj_adr_o[7] soc/mprj_adr_o[8]
+ soc/mprj_adr_o[9] soc/core_clk soc/hk_cyc_o soc/mprj_dat_o[0] soc/mprj_dat_o[10]
+ soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13] soc/mprj_dat_o[14] soc/mprj_dat_o[15]
+ soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18] soc/mprj_dat_o[19] soc/mprj_dat_o[1]
+ soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22] soc/mprj_dat_o[23] soc/mprj_dat_o[24]
+ soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27] soc/mprj_dat_o[28] soc/mprj_dat_o[29]
+ soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31] soc/mprj_dat_o[3] soc/mprj_dat_o[4]
+ soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7] soc/mprj_dat_o[8] soc/mprj_dat_o[9]
+ soc/hk_dat_i[0] soc/hk_dat_i[10] soc/hk_dat_i[11] soc/hk_dat_i[12] soc/hk_dat_i[13]
+ soc/hk_dat_i[14] soc/hk_dat_i[15] soc/hk_dat_i[16] soc/hk_dat_i[17] soc/hk_dat_i[18]
+ soc/hk_dat_i[19] soc/hk_dat_i[1] soc/hk_dat_i[20] soc/hk_dat_i[21] soc/hk_dat_i[22]
+ soc/hk_dat_i[23] soc/hk_dat_i[24] soc/hk_dat_i[25] soc/hk_dat_i[26] soc/hk_dat_i[27]
+ soc/hk_dat_i[28] soc/hk_dat_i[29] soc/hk_dat_i[2] soc/hk_dat_i[30] soc/hk_dat_i[31]
+ soc/hk_dat_i[3] soc/hk_dat_i[4] soc/hk_dat_i[5] soc/hk_dat_i[6] soc/hk_dat_i[7]
+ soc/hk_dat_i[8] soc/hk_dat_i[9] soc/core_rstn soc/mprj_sel_o[0] soc/mprj_sel_o[1]
+ soc/mprj_sel_o[2] soc/mprj_sel_o[3] soc/hk_stb_o soc/mprj_we_o housekeeping
Xgpio_control_in_2\[2\] soc/VDD soc/VSS gpio_defaults_block_7/gpio_defaults[0] gpio_defaults_block_7/gpio_defaults[1]
+ gpio_defaults_block_7/gpio_defaults[2] gpio_defaults_block_7/gpio_defaults[3] gpio_defaults_block_7/gpio_defaults[4]
+ gpio_defaults_block_7/gpio_defaults[5] gpio_defaults_block_7/gpio_defaults[6] gpio_defaults_block_7/gpio_defaults[7]
+ gpio_defaults_block_7/gpio_defaults[8] gpio_defaults_block_7/gpio_defaults[9] housekeeping/mgmt_gpio_in[21]
+ gpio_control_in_2\[2\]/zero housekeeping/mgmt_gpio_out[21] gpio_control_in_2\[2\]/one
+ padframe/mprj_io_drive_sel[42] padframe/mprj_io_drive_sel[43] padframe/mprj_io_in[21]
+ padframe/mprj_io_inen[21] padframe/mprj_io_out[21] padframe/mprj_io_outen[21] padframe/mprj_io_pd_select[21]
+ padframe/mprj_io_pu_select[21] padframe/mprj_io_schmitt_select[21] padframe/mprj_io_slew_select[21]
+ gpio_control_in_2\[2\]/resetn gpio_control_in_2\[1\]/resetn gpio_control_in_2\[2\]/serial_clock
+ gpio_control_in_2\[1\]/serial_clock gpio_control_in_2\[2\]/serial_data_in gpio_control_in_2\[1\]/serial_data_in
+ gpio_control_in_2\[2\]/serial_load gpio_control_in_2\[1\]/serial_load mprj/io_in[21]
+ mprj/io_oeb[21] mprj/io_out[21] gpio_control_in_2\[2\]/zero gpio_control_block
Xgpio_control_in_1\[8\] soc/VDD soc/VSS gpio_defaults_block_2/gpio_defaults[0] gpio_defaults_block_2/gpio_defaults[1]
+ gpio_defaults_block_2/gpio_defaults[2] gpio_defaults_block_2/gpio_defaults[3] gpio_defaults_block_2/gpio_defaults[4]
+ gpio_defaults_block_2/gpio_defaults[5] gpio_defaults_block_2/gpio_defaults[6] gpio_defaults_block_2/gpio_defaults[7]
+ gpio_defaults_block_2/gpio_defaults[8] gpio_defaults_block_2/gpio_defaults[9] housekeeping/mgmt_gpio_in[16]
+ gpio_control_in_1\[8\]/zero housekeeping/mgmt_gpio_out[16] gpio_control_in_1\[8\]/one
+ padframe/mprj_io_drive_sel[32] padframe/mprj_io_drive_sel[33] padframe/mprj_io_in[16]
+ padframe/mprj_io_inen[16] padframe/mprj_io_out[16] padframe/mprj_io_outen[16] padframe/mprj_io_pd_select[16]
+ padframe/mprj_io_pu_select[16] padframe/mprj_io_schmitt_select[16] padframe/mprj_io_slew_select[16]
+ gpio_control_in_1\[8\]/resetn gpio_control_in_1\[9\]/resetn gpio_control_in_1\[8\]/serial_clock
+ gpio_control_in_1\[9\]/serial_clock gpio_control_in_1\[8\]/serial_data_in gpio_control_in_1\[9\]/serial_data_in
+ gpio_control_in_1\[8\]/serial_load gpio_control_in_1\[9\]/serial_load mprj/io_in[16]
+ mprj/io_oeb[16] mprj/io_out[16] gpio_control_in_1\[8\]/zero gpio_control_block
Xspare_logic\[0\] soc/VDD soc/VSS spare_logic\[0\]/spare_xfq[0] spare_logic\[0\]/spare_xfq[1]
+ spare_logic\[0\]/spare_xi[0] spare_logic\[0\]/spare_xi[1] spare_logic\[0\]/spare_xi[2]
+ spare_logic\[0\]/spare_xi[3] spare_logic\[0\]/spare_xib spare_logic\[0\]/spare_xmx[0]
+ spare_logic\[0\]/spare_xmx[1] spare_logic\[0\]/spare_xna[0] spare_logic\[0\]/spare_xna[1]
+ spare_logic\[0\]/spare_xno[0] spare_logic\[0\]/spare_xno[1] spare_logic\[0\]/spare_xz[0]
+ spare_logic\[0\]/spare_xz[10] spare_logic\[0\]/spare_xz[11] spare_logic\[0\]/spare_xz[12]
+ spare_logic\[0\]/spare_xz[13] spare_logic\[0\]/spare_xz[14] spare_logic\[0\]/spare_xz[15]
+ spare_logic\[0\]/spare_xz[16] spare_logic\[0\]/spare_xz[17] spare_logic\[0\]/spare_xz[18]
+ spare_logic\[0\]/spare_xz[19] spare_logic\[0\]/spare_xz[1] spare_logic\[0\]/spare_xz[20]
+ spare_logic\[0\]/spare_xz[21] spare_logic\[0\]/spare_xz[22] spare_logic\[0\]/spare_xz[23]
+ spare_logic\[0\]/spare_xz[24] spare_logic\[0\]/spare_xz[25] spare_logic\[0\]/spare_xz[26]
+ spare_logic\[0\]/spare_xz[27] spare_logic\[0\]/spare_xz[28] spare_logic\[0\]/spare_xz[29]
+ spare_logic\[0\]/spare_xz[2] spare_logic\[0\]/spare_xz[30] spare_logic\[0\]/spare_xz[3]
+ spare_logic\[0\]/spare_xz[4] spare_logic\[0\]/spare_xz[5] spare_logic\[0\]/spare_xz[6]
+ spare_logic\[0\]/spare_xz[7] spare_logic\[0\]/spare_xz[8] spare_logic\[0\]/spare_xz[9]
+ spare_logic_block
Xgpio_defaults_block_30 gpio_defaults_block_30/gpio_defaults[0] gpio_defaults_block_30/gpio_defaults[1]
+ gpio_defaults_block_30/gpio_defaults[2] gpio_defaults_block_30/gpio_defaults[3]
+ gpio_defaults_block_30/gpio_defaults[4] gpio_defaults_block_30/gpio_defaults[5]
+ gpio_defaults_block_30/gpio_defaults[6] gpio_defaults_block_30/gpio_defaults[7]
+ gpio_defaults_block_30/gpio_defaults[8] gpio_defaults_block_30/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_10 gpio_defaults_block_10/gpio_defaults[0] gpio_defaults_block_10/gpio_defaults[1]
+ gpio_defaults_block_10/gpio_defaults[2] gpio_defaults_block_10/gpio_defaults[3]
+ gpio_defaults_block_10/gpio_defaults[4] gpio_defaults_block_10/gpio_defaults[5]
+ gpio_defaults_block_10/gpio_defaults[6] gpio_defaults_block_10/gpio_defaults[7]
+ gpio_defaults_block_10/gpio_defaults[8] gpio_defaults_block_10/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_20 gpio_defaults_block_20/gpio_defaults[0] gpio_defaults_block_20/gpio_defaults[1]
+ gpio_defaults_block_20/gpio_defaults[2] gpio_defaults_block_20/gpio_defaults[3]
+ gpio_defaults_block_20/gpio_defaults[4] gpio_defaults_block_20/gpio_defaults[5]
+ gpio_defaults_block_20/gpio_defaults[6] gpio_defaults_block_20/gpio_defaults[7]
+ gpio_defaults_block_20/gpio_defaults[8] gpio_defaults_block_20/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_21 gpio_defaults_block_21/gpio_defaults[0] gpio_defaults_block_21/gpio_defaults[1]
+ gpio_defaults_block_21/gpio_defaults[2] gpio_defaults_block_21/gpio_defaults[3]
+ gpio_defaults_block_21/gpio_defaults[4] gpio_defaults_block_21/gpio_defaults[5]
+ gpio_defaults_block_21/gpio_defaults[6] gpio_defaults_block_21/gpio_defaults[7]
+ gpio_defaults_block_21/gpio_defaults[8] gpio_defaults_block_21/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_in_1a\[5\] soc/VDD soc/VSS gpio_defaults_block_24/gpio_defaults[0] gpio_defaults_block_24/gpio_defaults[1]
+ gpio_defaults_block_24/gpio_defaults[2] gpio_defaults_block_24/gpio_defaults[3]
+ gpio_defaults_block_24/gpio_defaults[4] gpio_defaults_block_24/gpio_defaults[5]
+ gpio_defaults_block_24/gpio_defaults[6] gpio_defaults_block_24/gpio_defaults[7]
+ gpio_defaults_block_24/gpio_defaults[8] gpio_defaults_block_24/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[7] gpio_control_in_1a\[5\]/zero housekeeping/mgmt_gpio_out[7]
+ gpio_control_in_1a\[5\]/one padframe/mprj_io_drive_sel[15] padframe/mprj_io_drive_sel[14]
+ padframe/mprj_io_in[7] padframe/mprj_io_inen[7] padframe/mprj_io_out[7] padframe/mprj_io_outen[7]
+ padframe/mprj_io_pd_select[7] padframe/mprj_io_pu_select[7] padframe/mprj_io_schmitt_select[7]
+ padframe/mprj_io_slew_select[7] gpio_control_in_1a\[5\]/resetn gpio_control_in_1\[0\]/resetn
+ gpio_control_in_1a\[5\]/serial_clock gpio_control_in_1\[0\]/serial_clock gpio_control_in_1a\[5\]/serial_data_in
+ gpio_control_in_1\[0\]/serial_data_in gpio_control_in_1a\[5\]/serial_load gpio_control_in_1\[0\]/serial_load
+ mprj/io_in[7] mprj/io_oeb[7] mprj/io_out[7] gpio_control_in_1a\[5\]/zero gpio_control_block
Xgpio_defaults_block_31 gpio_defaults_block_31/gpio_defaults[0] gpio_defaults_block_31/gpio_defaults[1]
+ gpio_defaults_block_31/gpio_defaults[2] gpio_defaults_block_31/gpio_defaults[3]
+ gpio_defaults_block_31/gpio_defaults[4] gpio_defaults_block_31/gpio_defaults[5]
+ gpio_defaults_block_31/gpio_defaults[6] gpio_defaults_block_31/gpio_defaults[7]
+ gpio_defaults_block_31/gpio_defaults[8] gpio_defaults_block_31/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_defaults_block_32 gpio_defaults_block_32/gpio_defaults[0] gpio_defaults_block_32/gpio_defaults[1]
+ gpio_defaults_block_32/gpio_defaults[2] gpio_defaults_block_32/gpio_defaults[3]
+ gpio_defaults_block_32/gpio_defaults[4] gpio_defaults_block_32/gpio_defaults[5]
+ gpio_defaults_block_32/gpio_defaults[6] gpio_defaults_block_32/gpio_defaults[7]
+ gpio_defaults_block_32/gpio_defaults[8] gpio_defaults_block_32/gpio_defaults[9]
+ soc/VDD soc/VSS gpio_defaults_block
Xgpio_control_bidir_2\[2\] soc/VDD soc/VSS gpio_defaults_block_32/gpio_defaults[0]
+ gpio_defaults_block_32/gpio_defaults[1] gpio_defaults_block_32/gpio_defaults[2]
+ gpio_defaults_block_32/gpio_defaults[3] gpio_defaults_block_32/gpio_defaults[4]
+ gpio_defaults_block_32/gpio_defaults[5] gpio_defaults_block_32/gpio_defaults[6]
+ gpio_defaults_block_32/gpio_defaults[7] gpio_defaults_block_32/gpio_defaults[8]
+ gpio_defaults_block_32/gpio_defaults[9] housekeeping/mgmt_gpio_in[37] housekeeping/mgmt_gpio_oeb[37]
+ housekeeping/mgmt_gpio_out[37] gpio_control_bidir_2\[2\]/one padframe/mprj_io_drive_sel[74]
+ padframe/mprj_io_drive_sel[75] padframe/mprj_io_in[37] padframe/mprj_io_inen[37]
+ padframe/mprj_io_out[37] padframe/mprj_io_outen[37] padframe/mprj_io_pd_select[37]
+ padframe/mprj_io_pu_select[37] padframe/mprj_io_schmitt_select[37] padframe/mprj_io_slew_select[37]
+ housekeeping/serial_resetn gpio_control_bidir_2\[1\]/resetn housekeeping/serial_clock
+ gpio_control_bidir_2\[1\]/serial_clock housekeeping/serial_data_2 gpio_control_bidir_2\[1\]/serial_data_in
+ housekeeping/serial_load gpio_control_bidir_2\[1\]/serial_load mprj/io_in[37] mprj/io_oeb[37]
+ mprj/io_out[37] gpio_control_bidir_2\[2\]/zero gpio_control_block
.ends

