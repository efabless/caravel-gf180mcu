magic
tech gf180mcuC
magscale 1 10
timestamp 1655473305
<< checkpaint >>
rect -2000 -2000 222000 17000
<< obsm1 >>
rect 74 86 218624 14922
<< metal2 >>
rect 280 14200 392 15000
rect 952 14200 1064 15000
rect 1736 14200 1848 15000
rect 2408 14200 2520 15000
rect 3192 14200 3304 15000
rect 3864 14200 3976 15000
rect 4648 14200 4760 15000
rect 5320 14200 5432 15000
rect 6104 14200 6216 15000
rect 6776 14200 6888 15000
rect 7560 14200 7672 15000
rect 8232 14200 8344 15000
rect 9016 14200 9128 15000
rect 9688 14200 9800 15000
rect 10472 14200 10584 15000
rect 11144 14200 11256 15000
rect 11928 14200 12040 15000
rect 12600 14200 12712 15000
rect 13384 14200 13496 15000
rect 14056 14200 14168 15000
rect 14840 14200 14952 15000
rect 15512 14200 15624 15000
rect 16296 14200 16408 15000
rect 16968 14200 17080 15000
rect 17752 14200 17864 15000
rect 18424 14200 18536 15000
rect 19208 14200 19320 15000
rect 19880 14200 19992 15000
rect 20664 14200 20776 15000
rect 21336 14200 21448 15000
rect 22120 14200 22232 15000
rect 22792 14200 22904 15000
rect 23576 14200 23688 15000
rect 24248 14200 24360 15000
rect 25032 14200 25144 15000
rect 25704 14200 25816 15000
rect 26488 14200 26600 15000
rect 27160 14200 27272 15000
rect 27944 14200 28056 15000
rect 28616 14200 28728 15000
rect 29400 14200 29512 15000
rect 30072 14200 30184 15000
rect 30856 14200 30968 15000
rect 31528 14200 31640 15000
rect 32312 14200 32424 15000
rect 32984 14200 33096 15000
rect 33768 14200 33880 15000
rect 34440 14200 34552 15000
rect 35224 14200 35336 15000
rect 35896 14200 36008 15000
rect 36680 14200 36792 15000
rect 37352 14200 37464 15000
rect 38136 14200 38248 15000
rect 38808 14200 38920 15000
rect 39592 14200 39704 15000
rect 40264 14200 40376 15000
rect 41048 14200 41160 15000
rect 41720 14200 41832 15000
rect 42504 14200 42616 15000
rect 43176 14200 43288 15000
rect 43960 14200 44072 15000
rect 44632 14200 44744 15000
rect 45416 14200 45528 15000
rect 46088 14200 46200 15000
rect 46872 14200 46984 15000
rect 47544 14200 47656 15000
rect 48328 14200 48440 15000
rect 49000 14200 49112 15000
rect 49784 14200 49896 15000
rect 50456 14200 50568 15000
rect 51240 14200 51352 15000
rect 51912 14200 52024 15000
rect 52696 14200 52808 15000
rect 53368 14200 53480 15000
rect 54152 14200 54264 15000
rect 54824 14200 54936 15000
rect 55608 14200 55720 15000
rect 56392 14200 56504 15000
rect 57064 14200 57176 15000
rect 57848 14200 57960 15000
rect 58520 14200 58632 15000
rect 59304 14200 59416 15000
rect 59976 14200 60088 15000
rect 60760 14200 60872 15000
rect 61432 14200 61544 15000
rect 62216 14200 62328 15000
rect 62888 14200 63000 15000
rect 63672 14200 63784 15000
rect 64344 14200 64456 15000
rect 65128 14200 65240 15000
rect 65800 14200 65912 15000
rect 66584 14200 66696 15000
rect 67256 14200 67368 15000
rect 68040 14200 68152 15000
rect 68712 14200 68824 15000
rect 69496 14200 69608 15000
rect 70168 14200 70280 15000
rect 70952 14200 71064 15000
rect 71624 14200 71736 15000
rect 72408 14200 72520 15000
rect 73080 14200 73192 15000
rect 73864 14200 73976 15000
rect 74536 14200 74648 15000
rect 75320 14200 75432 15000
rect 75992 14200 76104 15000
rect 76776 14200 76888 15000
rect 77448 14200 77560 15000
rect 78232 14200 78344 15000
rect 78904 14200 79016 15000
rect 79688 14200 79800 15000
rect 80360 14200 80472 15000
rect 81144 14200 81256 15000
rect 81816 14200 81928 15000
rect 82600 14200 82712 15000
rect 83272 14200 83384 15000
rect 84056 14200 84168 15000
rect 84728 14200 84840 15000
rect 85512 14200 85624 15000
rect 86184 14200 86296 15000
rect 86968 14200 87080 15000
rect 87640 14200 87752 15000
rect 88424 14200 88536 15000
rect 89096 14200 89208 15000
rect 89880 14200 89992 15000
rect 90552 14200 90664 15000
rect 91336 14200 91448 15000
rect 92008 14200 92120 15000
rect 92792 14200 92904 15000
rect 93464 14200 93576 15000
rect 94248 14200 94360 15000
rect 94920 14200 95032 15000
rect 95704 14200 95816 15000
rect 96376 14200 96488 15000
rect 97160 14200 97272 15000
rect 97832 14200 97944 15000
rect 98616 14200 98728 15000
rect 99288 14200 99400 15000
rect 100072 14200 100184 15000
rect 100744 14200 100856 15000
rect 101528 14200 101640 15000
rect 102200 14200 102312 15000
rect 102984 14200 103096 15000
rect 103656 14200 103768 15000
rect 104440 14200 104552 15000
rect 105112 14200 105224 15000
rect 105896 14200 106008 15000
rect 106568 14200 106680 15000
rect 107352 14200 107464 15000
rect 108024 14200 108136 15000
rect 108808 14200 108920 15000
rect 109480 14200 109592 15000
rect 110264 14200 110376 15000
rect 111048 14200 111160 15000
rect 111720 14200 111832 15000
rect 112504 14200 112616 15000
rect 113176 14200 113288 15000
rect 113960 14200 114072 15000
rect 114632 14200 114744 15000
rect 115416 14200 115528 15000
rect 116088 14200 116200 15000
rect 116872 14200 116984 15000
rect 117544 14200 117656 15000
rect 118328 14200 118440 15000
rect 119000 14200 119112 15000
rect 119784 14200 119896 15000
rect 120456 14200 120568 15000
rect 121240 14200 121352 15000
rect 121912 14200 122024 15000
rect 122696 14200 122808 15000
rect 123368 14200 123480 15000
rect 124152 14200 124264 15000
rect 124824 14200 124936 15000
rect 125608 14200 125720 15000
rect 126280 14200 126392 15000
rect 127064 14200 127176 15000
rect 127736 14200 127848 15000
rect 128520 14200 128632 15000
rect 129192 14200 129304 15000
rect 129976 14200 130088 15000
rect 130648 14200 130760 15000
rect 131432 14200 131544 15000
rect 132104 14200 132216 15000
rect 132888 14200 133000 15000
rect 133560 14200 133672 15000
rect 134344 14200 134456 15000
rect 135016 14200 135128 15000
rect 135800 14200 135912 15000
rect 136472 14200 136584 15000
rect 137256 14200 137368 15000
rect 137928 14200 138040 15000
rect 138712 14200 138824 15000
rect 139384 14200 139496 15000
rect 140168 14200 140280 15000
rect 140840 14200 140952 15000
rect 141624 14200 141736 15000
rect 142296 14200 142408 15000
rect 143080 14200 143192 15000
rect 143752 14200 143864 15000
rect 144536 14200 144648 15000
rect 145208 14200 145320 15000
rect 145992 14200 146104 15000
rect 146664 14200 146776 15000
rect 147448 14200 147560 15000
rect 148120 14200 148232 15000
rect 148904 14200 149016 15000
rect 149576 14200 149688 15000
rect 150360 14200 150472 15000
rect 151032 14200 151144 15000
rect 151816 14200 151928 15000
rect 152488 14200 152600 15000
rect 153272 14200 153384 15000
rect 153944 14200 154056 15000
rect 154728 14200 154840 15000
rect 155400 14200 155512 15000
rect 156184 14200 156296 15000
rect 156856 14200 156968 15000
rect 157640 14200 157752 15000
rect 158312 14200 158424 15000
rect 159096 14200 159208 15000
rect 159768 14200 159880 15000
rect 160552 14200 160664 15000
rect 161224 14200 161336 15000
rect 162008 14200 162120 15000
rect 162680 14200 162792 15000
rect 163464 14200 163576 15000
rect 164136 14200 164248 15000
rect 164920 14200 165032 15000
rect 165704 14200 165816 15000
rect 166376 14200 166488 15000
rect 167160 14200 167272 15000
rect 167832 14200 167944 15000
rect 168616 14200 168728 15000
rect 169288 14200 169400 15000
rect 170072 14200 170184 15000
rect 170744 14200 170856 15000
rect 171528 14200 171640 15000
rect 172200 14200 172312 15000
rect 172984 14200 173096 15000
rect 173656 14200 173768 15000
rect 174440 14200 174552 15000
rect 175112 14200 175224 15000
rect 175896 14200 176008 15000
rect 176568 14200 176680 15000
rect 177352 14200 177464 15000
rect 178024 14200 178136 15000
rect 178808 14200 178920 15000
rect 179480 14200 179592 15000
rect 180264 14200 180376 15000
rect 180936 14200 181048 15000
rect 181720 14200 181832 15000
rect 182392 14200 182504 15000
rect 183176 14200 183288 15000
rect 183848 14200 183960 15000
rect 184632 14200 184744 15000
rect 185304 14200 185416 15000
rect 186088 14200 186200 15000
rect 186760 14200 186872 15000
rect 187544 14200 187656 15000
rect 188216 14200 188328 15000
rect 189000 14200 189112 15000
rect 189672 14200 189784 15000
rect 190456 14200 190568 15000
rect 191128 14200 191240 15000
rect 191912 14200 192024 15000
rect 192584 14200 192696 15000
rect 193368 14200 193480 15000
rect 194040 14200 194152 15000
rect 194824 14200 194936 15000
rect 195496 14200 195608 15000
rect 196280 14200 196392 15000
rect 196952 14200 197064 15000
rect 197736 14200 197848 15000
rect 198408 14200 198520 15000
rect 199192 14200 199304 15000
rect 199864 14200 199976 15000
rect 200648 14200 200760 15000
rect 201320 14200 201432 15000
rect 202104 14200 202216 15000
rect 202776 14200 202888 15000
rect 203560 14200 203672 15000
rect 204232 14200 204344 15000
rect 205016 14200 205128 15000
rect 205688 14200 205800 15000
rect 206472 14200 206584 15000
rect 207144 14200 207256 15000
rect 207928 14200 208040 15000
rect 208600 14200 208712 15000
rect 209384 14200 209496 15000
rect 210056 14200 210168 15000
rect 210840 14200 210952 15000
rect 211512 14200 211624 15000
rect 212296 14200 212408 15000
rect 212968 14200 213080 15000
rect 213752 14200 213864 15000
rect 214424 14200 214536 15000
rect 215208 14200 215320 15000
rect 215880 14200 215992 15000
rect 216664 14200 216776 15000
rect 217336 14200 217448 15000
rect 218120 14200 218232 15000
rect 218792 14200 218904 15000
rect 219576 14200 219688 15000
rect 168 0 280 800
rect 728 0 840 800
rect 1288 0 1400 800
rect 1960 0 2072 800
rect 2520 0 2632 800
rect 3192 0 3304 800
rect 3752 0 3864 800
rect 4424 0 4536 800
rect 4984 0 5096 800
rect 5544 0 5656 800
rect 6216 0 6328 800
rect 6776 0 6888 800
rect 7448 0 7560 800
rect 8008 0 8120 800
rect 8680 0 8792 800
rect 9240 0 9352 800
rect 9912 0 10024 800
rect 10472 0 10584 800
rect 11032 0 11144 800
rect 11704 0 11816 800
rect 12264 0 12376 800
rect 12936 0 13048 800
rect 13496 0 13608 800
rect 14168 0 14280 800
rect 14728 0 14840 800
rect 15400 0 15512 800
rect 15960 0 16072 800
rect 16520 0 16632 800
rect 17192 0 17304 800
rect 17752 0 17864 800
rect 18424 0 18536 800
rect 18984 0 19096 800
rect 19656 0 19768 800
rect 20216 0 20328 800
rect 20888 0 21000 800
rect 21448 0 21560 800
rect 22008 0 22120 800
rect 22680 0 22792 800
rect 23240 0 23352 800
rect 23912 0 24024 800
rect 24472 0 24584 800
rect 25144 0 25256 800
rect 25704 0 25816 800
rect 26376 0 26488 800
rect 26936 0 27048 800
rect 27496 0 27608 800
rect 28168 0 28280 800
rect 28728 0 28840 800
rect 29400 0 29512 800
rect 29960 0 30072 800
rect 30632 0 30744 800
rect 31192 0 31304 800
rect 31864 0 31976 800
rect 32424 0 32536 800
rect 32984 0 33096 800
rect 33656 0 33768 800
rect 34216 0 34328 800
rect 34888 0 35000 800
rect 35448 0 35560 800
rect 36120 0 36232 800
rect 36680 0 36792 800
rect 37352 0 37464 800
rect 37912 0 38024 800
rect 38472 0 38584 800
rect 39144 0 39256 800
rect 39704 0 39816 800
rect 40376 0 40488 800
rect 40936 0 41048 800
rect 41608 0 41720 800
rect 42168 0 42280 800
rect 42840 0 42952 800
rect 43400 0 43512 800
rect 43960 0 44072 800
rect 44632 0 44744 800
rect 45192 0 45304 800
rect 45864 0 45976 800
rect 46424 0 46536 800
rect 47096 0 47208 800
rect 47656 0 47768 800
rect 48328 0 48440 800
rect 48888 0 49000 800
rect 49448 0 49560 800
rect 50120 0 50232 800
rect 50680 0 50792 800
rect 51352 0 51464 800
rect 51912 0 52024 800
rect 52584 0 52696 800
rect 53144 0 53256 800
rect 53816 0 53928 800
rect 54376 0 54488 800
rect 54936 0 55048 800
rect 55608 0 55720 800
rect 56168 0 56280 800
rect 56840 0 56952 800
rect 57400 0 57512 800
rect 58072 0 58184 800
rect 58632 0 58744 800
rect 59192 0 59304 800
rect 59864 0 59976 800
rect 60424 0 60536 800
rect 61096 0 61208 800
rect 61656 0 61768 800
rect 62328 0 62440 800
rect 62888 0 63000 800
rect 63560 0 63672 800
rect 64120 0 64232 800
rect 64680 0 64792 800
rect 65352 0 65464 800
rect 65912 0 66024 800
rect 66584 0 66696 800
rect 67144 0 67256 800
rect 67816 0 67928 800
rect 68376 0 68488 800
rect 69048 0 69160 800
rect 69608 0 69720 800
rect 70168 0 70280 800
rect 70840 0 70952 800
rect 71400 0 71512 800
rect 72072 0 72184 800
rect 72632 0 72744 800
rect 73304 0 73416 800
rect 73864 0 73976 800
rect 74536 0 74648 800
rect 75096 0 75208 800
rect 75656 0 75768 800
rect 76328 0 76440 800
rect 76888 0 77000 800
rect 77560 0 77672 800
rect 78120 0 78232 800
rect 78792 0 78904 800
rect 79352 0 79464 800
rect 80024 0 80136 800
rect 80584 0 80696 800
rect 81144 0 81256 800
rect 81816 0 81928 800
rect 82376 0 82488 800
rect 83048 0 83160 800
rect 83608 0 83720 800
rect 84280 0 84392 800
rect 84840 0 84952 800
rect 85512 0 85624 800
rect 86072 0 86184 800
rect 86632 0 86744 800
rect 87304 0 87416 800
rect 87864 0 87976 800
rect 88536 0 88648 800
rect 89096 0 89208 800
rect 89768 0 89880 800
rect 90328 0 90440 800
rect 91000 0 91112 800
rect 91560 0 91672 800
rect 92120 0 92232 800
rect 92792 0 92904 800
rect 93352 0 93464 800
rect 94024 0 94136 800
rect 94584 0 94696 800
rect 95256 0 95368 800
rect 95816 0 95928 800
rect 96488 0 96600 800
rect 97048 0 97160 800
rect 97608 0 97720 800
rect 98280 0 98392 800
rect 98840 0 98952 800
rect 99512 0 99624 800
rect 100072 0 100184 800
rect 100744 0 100856 800
rect 101304 0 101416 800
rect 101976 0 102088 800
rect 102536 0 102648 800
rect 103096 0 103208 800
rect 103768 0 103880 800
rect 104328 0 104440 800
rect 105000 0 105112 800
rect 105560 0 105672 800
rect 106232 0 106344 800
rect 106792 0 106904 800
rect 107464 0 107576 800
rect 108024 0 108136 800
rect 108584 0 108696 800
rect 109256 0 109368 800
rect 109816 0 109928 800
rect 110488 0 110600 800
rect 111048 0 111160 800
rect 111720 0 111832 800
rect 112280 0 112392 800
rect 112840 0 112952 800
rect 113512 0 113624 800
rect 114072 0 114184 800
rect 114744 0 114856 800
rect 115304 0 115416 800
rect 115976 0 116088 800
rect 116536 0 116648 800
rect 117208 0 117320 800
rect 117768 0 117880 800
rect 118328 0 118440 800
rect 119000 0 119112 800
rect 119560 0 119672 800
rect 120232 0 120344 800
rect 120792 0 120904 800
rect 121464 0 121576 800
rect 122024 0 122136 800
rect 122696 0 122808 800
rect 123256 0 123368 800
rect 123816 0 123928 800
rect 124488 0 124600 800
rect 125048 0 125160 800
rect 125720 0 125832 800
rect 126280 0 126392 800
rect 126952 0 127064 800
rect 127512 0 127624 800
rect 128184 0 128296 800
rect 128744 0 128856 800
rect 129304 0 129416 800
rect 129976 0 130088 800
rect 130536 0 130648 800
rect 131208 0 131320 800
rect 131768 0 131880 800
rect 132440 0 132552 800
rect 133000 0 133112 800
rect 133672 0 133784 800
rect 134232 0 134344 800
rect 134792 0 134904 800
rect 135464 0 135576 800
rect 136024 0 136136 800
rect 136696 0 136808 800
rect 137256 0 137368 800
rect 137928 0 138040 800
rect 138488 0 138600 800
rect 139160 0 139272 800
rect 139720 0 139832 800
rect 140280 0 140392 800
rect 140952 0 141064 800
rect 141512 0 141624 800
rect 142184 0 142296 800
rect 142744 0 142856 800
rect 143416 0 143528 800
rect 143976 0 144088 800
rect 144648 0 144760 800
rect 145208 0 145320 800
rect 145768 0 145880 800
rect 146440 0 146552 800
rect 147000 0 147112 800
rect 147672 0 147784 800
rect 148232 0 148344 800
rect 148904 0 149016 800
rect 149464 0 149576 800
rect 150136 0 150248 800
rect 150696 0 150808 800
rect 151256 0 151368 800
rect 151928 0 152040 800
rect 152488 0 152600 800
rect 153160 0 153272 800
rect 153720 0 153832 800
rect 154392 0 154504 800
rect 154952 0 155064 800
rect 155624 0 155736 800
rect 156184 0 156296 800
rect 156744 0 156856 800
rect 157416 0 157528 800
rect 157976 0 158088 800
rect 158648 0 158760 800
rect 159208 0 159320 800
rect 159880 0 159992 800
rect 160440 0 160552 800
rect 161112 0 161224 800
rect 161672 0 161784 800
rect 162232 0 162344 800
rect 162904 0 163016 800
rect 163464 0 163576 800
rect 164136 0 164248 800
rect 164696 0 164808 800
rect 165368 0 165480 800
rect 165928 0 166040 800
rect 166488 0 166600 800
rect 167160 0 167272 800
rect 167720 0 167832 800
rect 168392 0 168504 800
rect 168952 0 169064 800
rect 169624 0 169736 800
rect 170184 0 170296 800
rect 170856 0 170968 800
rect 171416 0 171528 800
rect 171976 0 172088 800
rect 172648 0 172760 800
rect 173208 0 173320 800
rect 173880 0 173992 800
rect 174440 0 174552 800
rect 175112 0 175224 800
rect 175672 0 175784 800
rect 176344 0 176456 800
rect 176904 0 177016 800
rect 177464 0 177576 800
rect 178136 0 178248 800
rect 178696 0 178808 800
rect 179368 0 179480 800
rect 179928 0 180040 800
rect 180600 0 180712 800
rect 181160 0 181272 800
rect 181832 0 181944 800
rect 182392 0 182504 800
rect 182952 0 183064 800
rect 183624 0 183736 800
rect 184184 0 184296 800
rect 184856 0 184968 800
rect 185416 0 185528 800
rect 186088 0 186200 800
rect 186648 0 186760 800
rect 187320 0 187432 800
rect 187880 0 187992 800
rect 188440 0 188552 800
rect 189112 0 189224 800
rect 189672 0 189784 800
rect 190344 0 190456 800
rect 190904 0 191016 800
rect 191576 0 191688 800
rect 192136 0 192248 800
rect 192808 0 192920 800
rect 193368 0 193480 800
rect 193928 0 194040 800
rect 194600 0 194712 800
rect 195160 0 195272 800
rect 195832 0 195944 800
rect 196392 0 196504 800
rect 197064 0 197176 800
rect 197624 0 197736 800
rect 198296 0 198408 800
rect 198856 0 198968 800
rect 199416 0 199528 800
rect 200088 0 200200 800
rect 200648 0 200760 800
rect 201320 0 201432 800
rect 201880 0 201992 800
rect 202552 0 202664 800
rect 203112 0 203224 800
rect 203784 0 203896 800
rect 204344 0 204456 800
rect 204904 0 205016 800
rect 205576 0 205688 800
rect 206136 0 206248 800
rect 206808 0 206920 800
rect 207368 0 207480 800
rect 208040 0 208152 800
rect 208600 0 208712 800
rect 209272 0 209384 800
rect 209832 0 209944 800
rect 210392 0 210504 800
rect 211064 0 211176 800
rect 211624 0 211736 800
rect 212296 0 212408 800
rect 212856 0 212968 800
rect 213528 0 213640 800
rect 214088 0 214200 800
rect 214760 0 214872 800
rect 215320 0 215432 800
rect 215880 0 215992 800
rect 216552 0 216664 800
rect 217112 0 217224 800
rect 217784 0 217896 800
rect 218344 0 218456 800
rect 219016 0 219128 800
rect 219576 0 219688 800
<< obsm2 >>
rect 84 14140 220 14934
rect 452 14140 892 14934
rect 1124 14140 1676 14934
rect 1908 14140 2348 14934
rect 2580 14140 3132 14934
rect 3364 14140 3804 14934
rect 4036 14140 4588 14934
rect 4820 14140 5260 14934
rect 5492 14140 6044 14934
rect 6276 14140 6716 14934
rect 6948 14140 7500 14934
rect 7732 14140 8172 14934
rect 8404 14140 8956 14934
rect 9188 14140 9628 14934
rect 9860 14140 10412 14934
rect 10644 14140 11084 14934
rect 11316 14140 11868 14934
rect 12100 14140 12540 14934
rect 12772 14140 13324 14934
rect 13556 14140 13996 14934
rect 14228 14140 14780 14934
rect 15012 14140 15452 14934
rect 15684 14140 16236 14934
rect 16468 14140 16908 14934
rect 17140 14140 17692 14934
rect 17924 14140 18364 14934
rect 18596 14140 19148 14934
rect 19380 14140 19820 14934
rect 20052 14140 20604 14934
rect 20836 14140 21276 14934
rect 21508 14140 22060 14934
rect 22292 14140 22732 14934
rect 22964 14140 23516 14934
rect 23748 14140 24188 14934
rect 24420 14140 24972 14934
rect 25204 14140 25644 14934
rect 25876 14140 26428 14934
rect 26660 14140 27100 14934
rect 27332 14140 27884 14934
rect 28116 14140 28556 14934
rect 28788 14140 29340 14934
rect 29572 14140 30012 14934
rect 30244 14140 30796 14934
rect 31028 14140 31468 14934
rect 31700 14140 32252 14934
rect 32484 14140 32924 14934
rect 33156 14140 33708 14934
rect 33940 14140 34380 14934
rect 34612 14140 35164 14934
rect 35396 14140 35836 14934
rect 36068 14140 36620 14934
rect 36852 14140 37292 14934
rect 37524 14140 38076 14934
rect 38308 14140 38748 14934
rect 38980 14140 39532 14934
rect 39764 14140 40204 14934
rect 40436 14140 40988 14934
rect 41220 14140 41660 14934
rect 41892 14140 42444 14934
rect 42676 14140 43116 14934
rect 43348 14140 43900 14934
rect 44132 14140 44572 14934
rect 44804 14140 45356 14934
rect 45588 14140 46028 14934
rect 46260 14140 46812 14934
rect 47044 14140 47484 14934
rect 47716 14140 48268 14934
rect 48500 14140 48940 14934
rect 49172 14140 49724 14934
rect 49956 14140 50396 14934
rect 50628 14140 51180 14934
rect 51412 14140 51852 14934
rect 52084 14140 52636 14934
rect 52868 14140 53308 14934
rect 53540 14140 54092 14934
rect 54324 14140 54764 14934
rect 54996 14140 55548 14934
rect 55780 14140 56332 14934
rect 56564 14140 57004 14934
rect 57236 14140 57788 14934
rect 58020 14140 58460 14934
rect 58692 14140 59244 14934
rect 59476 14140 59916 14934
rect 60148 14140 60700 14934
rect 60932 14140 61372 14934
rect 61604 14140 62156 14934
rect 62388 14140 62828 14934
rect 63060 14140 63612 14934
rect 63844 14140 64284 14934
rect 64516 14140 65068 14934
rect 65300 14140 65740 14934
rect 65972 14140 66524 14934
rect 66756 14140 67196 14934
rect 67428 14140 67980 14934
rect 68212 14140 68652 14934
rect 68884 14140 69436 14934
rect 69668 14140 70108 14934
rect 70340 14140 70892 14934
rect 71124 14140 71564 14934
rect 71796 14140 72348 14934
rect 72580 14140 73020 14934
rect 73252 14140 73804 14934
rect 74036 14140 74476 14934
rect 74708 14140 75260 14934
rect 75492 14140 75932 14934
rect 76164 14140 76716 14934
rect 76948 14140 77388 14934
rect 77620 14140 78172 14934
rect 78404 14140 78844 14934
rect 79076 14140 79628 14934
rect 79860 14140 80300 14934
rect 80532 14140 81084 14934
rect 81316 14140 81756 14934
rect 81988 14140 82540 14934
rect 82772 14140 83212 14934
rect 83444 14140 83996 14934
rect 84228 14140 84668 14934
rect 84900 14140 85452 14934
rect 85684 14140 86124 14934
rect 86356 14140 86908 14934
rect 87140 14140 87580 14934
rect 87812 14140 88364 14934
rect 88596 14140 89036 14934
rect 89268 14140 89820 14934
rect 90052 14140 90492 14934
rect 90724 14140 91276 14934
rect 91508 14140 91948 14934
rect 92180 14140 92732 14934
rect 92964 14140 93404 14934
rect 93636 14140 94188 14934
rect 94420 14140 94860 14934
rect 95092 14140 95644 14934
rect 95876 14140 96316 14934
rect 96548 14140 97100 14934
rect 97332 14140 97772 14934
rect 98004 14140 98556 14934
rect 98788 14140 99228 14934
rect 99460 14140 100012 14934
rect 100244 14140 100684 14934
rect 100916 14140 101468 14934
rect 101700 14140 102140 14934
rect 102372 14140 102924 14934
rect 103156 14140 103596 14934
rect 103828 14140 104380 14934
rect 104612 14140 105052 14934
rect 105284 14140 105836 14934
rect 106068 14140 106508 14934
rect 106740 14140 107292 14934
rect 107524 14140 107964 14934
rect 108196 14140 108748 14934
rect 108980 14140 109420 14934
rect 109652 14140 110204 14934
rect 110436 14140 110988 14934
rect 111220 14140 111660 14934
rect 111892 14140 112444 14934
rect 112676 14140 113116 14934
rect 113348 14140 113900 14934
rect 114132 14140 114572 14934
rect 114804 14140 115356 14934
rect 115588 14140 116028 14934
rect 116260 14140 116812 14934
rect 117044 14140 117484 14934
rect 117716 14140 118268 14934
rect 118500 14140 118940 14934
rect 119172 14140 119724 14934
rect 119956 14140 120396 14934
rect 120628 14140 121180 14934
rect 121412 14140 121852 14934
rect 122084 14140 122636 14934
rect 122868 14140 123308 14934
rect 123540 14140 124092 14934
rect 124324 14140 124764 14934
rect 124996 14140 125548 14934
rect 125780 14140 126220 14934
rect 126452 14140 127004 14934
rect 127236 14140 127676 14934
rect 127908 14140 128460 14934
rect 128692 14140 129132 14934
rect 129364 14140 129916 14934
rect 130148 14140 130588 14934
rect 130820 14140 131372 14934
rect 131604 14140 132044 14934
rect 132276 14140 132828 14934
rect 133060 14140 133500 14934
rect 133732 14140 134284 14934
rect 134516 14140 134956 14934
rect 135188 14140 135740 14934
rect 135972 14140 136412 14934
rect 136644 14140 137196 14934
rect 137428 14140 137868 14934
rect 138100 14140 138652 14934
rect 138884 14140 139324 14934
rect 139556 14140 140108 14934
rect 140340 14140 140780 14934
rect 141012 14140 141564 14934
rect 141796 14140 142236 14934
rect 142468 14140 143020 14934
rect 143252 14140 143692 14934
rect 143924 14140 144476 14934
rect 144708 14140 145148 14934
rect 145380 14140 145932 14934
rect 146164 14140 146604 14934
rect 146836 14140 147388 14934
rect 147620 14140 148060 14934
rect 148292 14140 148844 14934
rect 149076 14140 149516 14934
rect 149748 14140 150300 14934
rect 150532 14140 150972 14934
rect 151204 14140 151756 14934
rect 151988 14140 152428 14934
rect 152660 14140 153212 14934
rect 153444 14140 153884 14934
rect 154116 14140 154668 14934
rect 154900 14140 155340 14934
rect 155572 14140 156124 14934
rect 156356 14140 156796 14934
rect 157028 14140 157580 14934
rect 157812 14140 158252 14934
rect 158484 14140 159036 14934
rect 159268 14140 159708 14934
rect 159940 14140 160492 14934
rect 160724 14140 161164 14934
rect 161396 14140 161948 14934
rect 162180 14140 162620 14934
rect 162852 14140 163404 14934
rect 163636 14140 164076 14934
rect 164308 14140 164860 14934
rect 165092 14140 165644 14934
rect 165876 14140 166316 14934
rect 166548 14140 167100 14934
rect 167332 14140 167772 14934
rect 168004 14140 168556 14934
rect 168788 14140 169228 14934
rect 169460 14140 170012 14934
rect 170244 14140 170684 14934
rect 170916 14140 171468 14934
rect 171700 14140 172140 14934
rect 172372 14140 172924 14934
rect 173156 14140 173596 14934
rect 173828 14140 174380 14934
rect 174612 14140 175052 14934
rect 175284 14140 175836 14934
rect 176068 14140 176508 14934
rect 176740 14140 177292 14934
rect 177524 14140 177964 14934
rect 178196 14140 178748 14934
rect 178980 14140 179420 14934
rect 179652 14140 180204 14934
rect 180436 14140 180876 14934
rect 181108 14140 181660 14934
rect 181892 14140 182332 14934
rect 182564 14140 183116 14934
rect 183348 14140 183788 14934
rect 184020 14140 184572 14934
rect 184804 14140 185244 14934
rect 185476 14140 186028 14934
rect 186260 14140 186700 14934
rect 186932 14140 187484 14934
rect 187716 14140 188156 14934
rect 188388 14140 188940 14934
rect 189172 14140 189612 14934
rect 189844 14140 190396 14934
rect 190628 14140 191068 14934
rect 191300 14140 191852 14934
rect 192084 14140 192524 14934
rect 192756 14140 193308 14934
rect 193540 14140 193980 14934
rect 194212 14140 194764 14934
rect 194996 14140 195436 14934
rect 195668 14140 196220 14934
rect 196452 14140 196892 14934
rect 197124 14140 197676 14934
rect 197908 14140 198348 14934
rect 198580 14140 199132 14934
rect 199364 14140 199804 14934
rect 200036 14140 200588 14934
rect 200820 14140 201260 14934
rect 201492 14140 202044 14934
rect 202276 14140 202716 14934
rect 202948 14140 203500 14934
rect 203732 14140 204172 14934
rect 204404 14140 204956 14934
rect 205188 14140 205628 14934
rect 205860 14140 206412 14934
rect 206644 14140 207084 14934
rect 207316 14140 207868 14934
rect 208100 14140 208540 14934
rect 208772 14140 209324 14934
rect 209556 14140 209996 14934
rect 210228 14140 210780 14934
rect 211012 14140 211452 14934
rect 211684 14140 212236 14934
rect 212468 14140 212908 14934
rect 213140 14140 213692 14934
rect 213924 14140 214364 14934
rect 214596 14140 215148 14934
rect 215380 14140 215820 14934
rect 216052 14140 216604 14934
rect 216836 14140 217276 14934
rect 217508 14140 218060 14934
rect 218292 14140 218732 14934
rect 218964 14140 219516 14934
rect 84 860 219660 14140
rect 84 74 108 860
rect 340 74 668 860
rect 900 74 1228 860
rect 1460 74 1900 860
rect 2132 74 2460 860
rect 2692 74 3132 860
rect 3364 74 3692 860
rect 3924 74 4364 860
rect 4596 74 4924 860
rect 5156 74 5484 860
rect 5716 74 6156 860
rect 6388 74 6716 860
rect 6948 74 7388 860
rect 7620 74 7948 860
rect 8180 74 8620 860
rect 8852 74 9180 860
rect 9412 74 9852 860
rect 10084 74 10412 860
rect 10644 74 10972 860
rect 11204 74 11644 860
rect 11876 74 12204 860
rect 12436 74 12876 860
rect 13108 74 13436 860
rect 13668 74 14108 860
rect 14340 74 14668 860
rect 14900 74 15340 860
rect 15572 74 15900 860
rect 16132 74 16460 860
rect 16692 74 17132 860
rect 17364 74 17692 860
rect 17924 74 18364 860
rect 18596 74 18924 860
rect 19156 74 19596 860
rect 19828 74 20156 860
rect 20388 74 20828 860
rect 21060 74 21388 860
rect 21620 74 21948 860
rect 22180 74 22620 860
rect 22852 74 23180 860
rect 23412 74 23852 860
rect 24084 74 24412 860
rect 24644 74 25084 860
rect 25316 74 25644 860
rect 25876 74 26316 860
rect 26548 74 26876 860
rect 27108 74 27436 860
rect 27668 74 28108 860
rect 28340 74 28668 860
rect 28900 74 29340 860
rect 29572 74 29900 860
rect 30132 74 30572 860
rect 30804 74 31132 860
rect 31364 74 31804 860
rect 32036 74 32364 860
rect 32596 74 32924 860
rect 33156 74 33596 860
rect 33828 74 34156 860
rect 34388 74 34828 860
rect 35060 74 35388 860
rect 35620 74 36060 860
rect 36292 74 36620 860
rect 36852 74 37292 860
rect 37524 74 37852 860
rect 38084 74 38412 860
rect 38644 74 39084 860
rect 39316 74 39644 860
rect 39876 74 40316 860
rect 40548 74 40876 860
rect 41108 74 41548 860
rect 41780 74 42108 860
rect 42340 74 42780 860
rect 43012 74 43340 860
rect 43572 74 43900 860
rect 44132 74 44572 860
rect 44804 74 45132 860
rect 45364 74 45804 860
rect 46036 74 46364 860
rect 46596 74 47036 860
rect 47268 74 47596 860
rect 47828 74 48268 860
rect 48500 74 48828 860
rect 49060 74 49388 860
rect 49620 74 50060 860
rect 50292 74 50620 860
rect 50852 74 51292 860
rect 51524 74 51852 860
rect 52084 74 52524 860
rect 52756 74 53084 860
rect 53316 74 53756 860
rect 53988 74 54316 860
rect 54548 74 54876 860
rect 55108 74 55548 860
rect 55780 74 56108 860
rect 56340 74 56780 860
rect 57012 74 57340 860
rect 57572 74 58012 860
rect 58244 74 58572 860
rect 58804 74 59132 860
rect 59364 74 59804 860
rect 60036 74 60364 860
rect 60596 74 61036 860
rect 61268 74 61596 860
rect 61828 74 62268 860
rect 62500 74 62828 860
rect 63060 74 63500 860
rect 63732 74 64060 860
rect 64292 74 64620 860
rect 64852 74 65292 860
rect 65524 74 65852 860
rect 66084 74 66524 860
rect 66756 74 67084 860
rect 67316 74 67756 860
rect 67988 74 68316 860
rect 68548 74 68988 860
rect 69220 74 69548 860
rect 69780 74 70108 860
rect 70340 74 70780 860
rect 71012 74 71340 860
rect 71572 74 72012 860
rect 72244 74 72572 860
rect 72804 74 73244 860
rect 73476 74 73804 860
rect 74036 74 74476 860
rect 74708 74 75036 860
rect 75268 74 75596 860
rect 75828 74 76268 860
rect 76500 74 76828 860
rect 77060 74 77500 860
rect 77732 74 78060 860
rect 78292 74 78732 860
rect 78964 74 79292 860
rect 79524 74 79964 860
rect 80196 74 80524 860
rect 80756 74 81084 860
rect 81316 74 81756 860
rect 81988 74 82316 860
rect 82548 74 82988 860
rect 83220 74 83548 860
rect 83780 74 84220 860
rect 84452 74 84780 860
rect 85012 74 85452 860
rect 85684 74 86012 860
rect 86244 74 86572 860
rect 86804 74 87244 860
rect 87476 74 87804 860
rect 88036 74 88476 860
rect 88708 74 89036 860
rect 89268 74 89708 860
rect 89940 74 90268 860
rect 90500 74 90940 860
rect 91172 74 91500 860
rect 91732 74 92060 860
rect 92292 74 92732 860
rect 92964 74 93292 860
rect 93524 74 93964 860
rect 94196 74 94524 860
rect 94756 74 95196 860
rect 95428 74 95756 860
rect 95988 74 96428 860
rect 96660 74 96988 860
rect 97220 74 97548 860
rect 97780 74 98220 860
rect 98452 74 98780 860
rect 99012 74 99452 860
rect 99684 74 100012 860
rect 100244 74 100684 860
rect 100916 74 101244 860
rect 101476 74 101916 860
rect 102148 74 102476 860
rect 102708 74 103036 860
rect 103268 74 103708 860
rect 103940 74 104268 860
rect 104500 74 104940 860
rect 105172 74 105500 860
rect 105732 74 106172 860
rect 106404 74 106732 860
rect 106964 74 107404 860
rect 107636 74 107964 860
rect 108196 74 108524 860
rect 108756 74 109196 860
rect 109428 74 109756 860
rect 109988 74 110428 860
rect 110660 74 110988 860
rect 111220 74 111660 860
rect 111892 74 112220 860
rect 112452 74 112780 860
rect 113012 74 113452 860
rect 113684 74 114012 860
rect 114244 74 114684 860
rect 114916 74 115244 860
rect 115476 74 115916 860
rect 116148 74 116476 860
rect 116708 74 117148 860
rect 117380 74 117708 860
rect 117940 74 118268 860
rect 118500 74 118940 860
rect 119172 74 119500 860
rect 119732 74 120172 860
rect 120404 74 120732 860
rect 120964 74 121404 860
rect 121636 74 121964 860
rect 122196 74 122636 860
rect 122868 74 123196 860
rect 123428 74 123756 860
rect 123988 74 124428 860
rect 124660 74 124988 860
rect 125220 74 125660 860
rect 125892 74 126220 860
rect 126452 74 126892 860
rect 127124 74 127452 860
rect 127684 74 128124 860
rect 128356 74 128684 860
rect 128916 74 129244 860
rect 129476 74 129916 860
rect 130148 74 130476 860
rect 130708 74 131148 860
rect 131380 74 131708 860
rect 131940 74 132380 860
rect 132612 74 132940 860
rect 133172 74 133612 860
rect 133844 74 134172 860
rect 134404 74 134732 860
rect 134964 74 135404 860
rect 135636 74 135964 860
rect 136196 74 136636 860
rect 136868 74 137196 860
rect 137428 74 137868 860
rect 138100 74 138428 860
rect 138660 74 139100 860
rect 139332 74 139660 860
rect 139892 74 140220 860
rect 140452 74 140892 860
rect 141124 74 141452 860
rect 141684 74 142124 860
rect 142356 74 142684 860
rect 142916 74 143356 860
rect 143588 74 143916 860
rect 144148 74 144588 860
rect 144820 74 145148 860
rect 145380 74 145708 860
rect 145940 74 146380 860
rect 146612 74 146940 860
rect 147172 74 147612 860
rect 147844 74 148172 860
rect 148404 74 148844 860
rect 149076 74 149404 860
rect 149636 74 150076 860
rect 150308 74 150636 860
rect 150868 74 151196 860
rect 151428 74 151868 860
rect 152100 74 152428 860
rect 152660 74 153100 860
rect 153332 74 153660 860
rect 153892 74 154332 860
rect 154564 74 154892 860
rect 155124 74 155564 860
rect 155796 74 156124 860
rect 156356 74 156684 860
rect 156916 74 157356 860
rect 157588 74 157916 860
rect 158148 74 158588 860
rect 158820 74 159148 860
rect 159380 74 159820 860
rect 160052 74 160380 860
rect 160612 74 161052 860
rect 161284 74 161612 860
rect 161844 74 162172 860
rect 162404 74 162844 860
rect 163076 74 163404 860
rect 163636 74 164076 860
rect 164308 74 164636 860
rect 164868 74 165308 860
rect 165540 74 165868 860
rect 166100 74 166428 860
rect 166660 74 167100 860
rect 167332 74 167660 860
rect 167892 74 168332 860
rect 168564 74 168892 860
rect 169124 74 169564 860
rect 169796 74 170124 860
rect 170356 74 170796 860
rect 171028 74 171356 860
rect 171588 74 171916 860
rect 172148 74 172588 860
rect 172820 74 173148 860
rect 173380 74 173820 860
rect 174052 74 174380 860
rect 174612 74 175052 860
rect 175284 74 175612 860
rect 175844 74 176284 860
rect 176516 74 176844 860
rect 177076 74 177404 860
rect 177636 74 178076 860
rect 178308 74 178636 860
rect 178868 74 179308 860
rect 179540 74 179868 860
rect 180100 74 180540 860
rect 180772 74 181100 860
rect 181332 74 181772 860
rect 182004 74 182332 860
rect 182564 74 182892 860
rect 183124 74 183564 860
rect 183796 74 184124 860
rect 184356 74 184796 860
rect 185028 74 185356 860
rect 185588 74 186028 860
rect 186260 74 186588 860
rect 186820 74 187260 860
rect 187492 74 187820 860
rect 188052 74 188380 860
rect 188612 74 189052 860
rect 189284 74 189612 860
rect 189844 74 190284 860
rect 190516 74 190844 860
rect 191076 74 191516 860
rect 191748 74 192076 860
rect 192308 74 192748 860
rect 192980 74 193308 860
rect 193540 74 193868 860
rect 194100 74 194540 860
rect 194772 74 195100 860
rect 195332 74 195772 860
rect 196004 74 196332 860
rect 196564 74 197004 860
rect 197236 74 197564 860
rect 197796 74 198236 860
rect 198468 74 198796 860
rect 199028 74 199356 860
rect 199588 74 200028 860
rect 200260 74 200588 860
rect 200820 74 201260 860
rect 201492 74 201820 860
rect 202052 74 202492 860
rect 202724 74 203052 860
rect 203284 74 203724 860
rect 203956 74 204284 860
rect 204516 74 204844 860
rect 205076 74 205516 860
rect 205748 74 206076 860
rect 206308 74 206748 860
rect 206980 74 207308 860
rect 207540 74 207980 860
rect 208212 74 208540 860
rect 208772 74 209212 860
rect 209444 74 209772 860
rect 210004 74 210332 860
rect 210564 74 211004 860
rect 211236 74 211564 860
rect 211796 74 212236 860
rect 212468 74 212796 860
rect 213028 74 213468 860
rect 213700 74 214028 860
rect 214260 74 214700 860
rect 214932 74 215260 860
rect 215492 74 215820 860
rect 216052 74 216492 860
rect 216724 74 217052 860
rect 217284 74 217724 860
rect 217956 74 218284 860
rect 218516 74 218956 860
rect 219188 74 219516 860
<< metal3 >>
rect 219200 13608 220000 13720
rect 0 12376 800 12488
rect 219200 11144 220000 11256
rect 219200 8680 220000 8792
rect 0 7448 800 7560
rect 219200 6216 220000 6328
rect 219200 3752 220000 3864
rect 0 2520 800 2632
rect 219200 1288 220000 1400
<< obsm3 >>
rect 74 13780 219670 14924
rect 74 13548 219140 13780
rect 74 12548 219670 13548
rect 860 12316 219670 12548
rect 74 11316 219670 12316
rect 74 11084 219140 11316
rect 74 8852 219670 11084
rect 74 8620 219140 8852
rect 74 7620 219670 8620
rect 860 7388 219670 7620
rect 74 6388 219670 7388
rect 74 6156 219140 6388
rect 74 3924 219670 6156
rect 74 3692 219140 3924
rect 74 2692 219670 3692
rect 860 2460 219670 2692
rect 74 1460 219670 2460
rect 74 1228 219140 1460
rect 74 84 219670 1228
<< metal4 >>
rect 28348 4644 28668 10252
rect 55512 4644 55832 10252
rect 82676 4644 82996 10252
rect 109840 4644 110160 10252
rect 137004 4644 137324 10252
rect 164168 4644 164488 10252
rect 191332 4644 191652 10252
<< obsm4 >>
rect 1316 10312 217196 14978
rect 1316 4584 28288 10312
rect 28728 4584 55452 10312
rect 55892 4584 82616 10312
rect 83056 4584 109780 10312
rect 110220 4584 136944 10312
rect 137384 4584 164108 10312
rect 164548 4584 191272 10312
rect 191712 4584 217196 10312
rect 1316 74 217196 4584
<< metal5 >>
rect 1284 9437 218684 9757
rect 1284 8738 218684 9058
rect 1284 8039 218684 8359
rect 1284 7340 218684 7660
rect 1284 6641 218684 6961
rect 1284 5942 218684 6262
rect 1284 5243 218684 5563
<< obsm5 >>
rect 1300 9857 217212 14984
rect 1300 9158 217212 9337
rect 1300 8459 217212 8638
rect 1300 7760 217212 7939
rect 1300 7061 217212 7240
rect 1300 6362 217212 6541
rect 1300 5663 217212 5842
rect 1300 136 217212 5143
<< labels >>
rlabel metal4 s 28348 4644 28668 10252 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 82676 4644 82996 10252 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 137004 4644 137324 10252 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 191332 4644 191652 10252 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 1284 5243 218684 5563 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 1284 6641 218684 6961 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 1284 8039 218684 8359 6 VDD
port 1 nsew power bidirectional
rlabel metal5 s 1284 9437 218684 9757 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 55512 4644 55832 10252 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 109840 4644 110160 10252 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 164168 4644 164488 10252 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 1284 5942 218684 6262 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 1284 7340 218684 7660 6 VSS
port 2 nsew ground bidirectional
rlabel metal5 s 1284 8738 218684 9058 6 VSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 2520 800 2632 6 caravel_clk
port 3 nsew signal input
rlabel metal3 s 0 7448 800 7560 6 caravel_clk2
port 4 nsew signal input
rlabel metal3 s 0 12376 800 12488 6 caravel_rstn
port 5 nsew signal input
rlabel metal2 s 77448 14200 77560 15000 6 la_data_in_core[0]
port 6 nsew signal output
rlabel metal2 s 99288 14200 99400 15000 6 la_data_in_core[10]
port 7 nsew signal output
rlabel metal2 s 101528 14200 101640 15000 6 la_data_in_core[11]
port 8 nsew signal output
rlabel metal2 s 103656 14200 103768 15000 6 la_data_in_core[12]
port 9 nsew signal output
rlabel metal2 s 105896 14200 106008 15000 6 la_data_in_core[13]
port 10 nsew signal output
rlabel metal2 s 108024 14200 108136 15000 6 la_data_in_core[14]
port 11 nsew signal output
rlabel metal2 s 110264 14200 110376 15000 6 la_data_in_core[15]
port 12 nsew signal output
rlabel metal2 s 112504 14200 112616 15000 6 la_data_in_core[16]
port 13 nsew signal output
rlabel metal2 s 114632 14200 114744 15000 6 la_data_in_core[17]
port 14 nsew signal output
rlabel metal2 s 116872 14200 116984 15000 6 la_data_in_core[18]
port 15 nsew signal output
rlabel metal2 s 119000 14200 119112 15000 6 la_data_in_core[19]
port 16 nsew signal output
rlabel metal2 s 79688 14200 79800 15000 6 la_data_in_core[1]
port 17 nsew signal output
rlabel metal2 s 121240 14200 121352 15000 6 la_data_in_core[20]
port 18 nsew signal output
rlabel metal2 s 123368 14200 123480 15000 6 la_data_in_core[21]
port 19 nsew signal output
rlabel metal2 s 125608 14200 125720 15000 6 la_data_in_core[22]
port 20 nsew signal output
rlabel metal2 s 127736 14200 127848 15000 6 la_data_in_core[23]
port 21 nsew signal output
rlabel metal2 s 129976 14200 130088 15000 6 la_data_in_core[24]
port 22 nsew signal output
rlabel metal2 s 132104 14200 132216 15000 6 la_data_in_core[25]
port 23 nsew signal output
rlabel metal2 s 134344 14200 134456 15000 6 la_data_in_core[26]
port 24 nsew signal output
rlabel metal2 s 136472 14200 136584 15000 6 la_data_in_core[27]
port 25 nsew signal output
rlabel metal2 s 138712 14200 138824 15000 6 la_data_in_core[28]
port 26 nsew signal output
rlabel metal2 s 140840 14200 140952 15000 6 la_data_in_core[29]
port 27 nsew signal output
rlabel metal2 s 81816 14200 81928 15000 6 la_data_in_core[2]
port 28 nsew signal output
rlabel metal2 s 143080 14200 143192 15000 6 la_data_in_core[30]
port 29 nsew signal output
rlabel metal2 s 145208 14200 145320 15000 6 la_data_in_core[31]
port 30 nsew signal output
rlabel metal2 s 147448 14200 147560 15000 6 la_data_in_core[32]
port 31 nsew signal output
rlabel metal2 s 149576 14200 149688 15000 6 la_data_in_core[33]
port 32 nsew signal output
rlabel metal2 s 151816 14200 151928 15000 6 la_data_in_core[34]
port 33 nsew signal output
rlabel metal2 s 153944 14200 154056 15000 6 la_data_in_core[35]
port 34 nsew signal output
rlabel metal2 s 156184 14200 156296 15000 6 la_data_in_core[36]
port 35 nsew signal output
rlabel metal2 s 158312 14200 158424 15000 6 la_data_in_core[37]
port 36 nsew signal output
rlabel metal2 s 160552 14200 160664 15000 6 la_data_in_core[38]
port 37 nsew signal output
rlabel metal2 s 162680 14200 162792 15000 6 la_data_in_core[39]
port 38 nsew signal output
rlabel metal2 s 84056 14200 84168 15000 6 la_data_in_core[3]
port 39 nsew signal output
rlabel metal2 s 164920 14200 165032 15000 6 la_data_in_core[40]
port 40 nsew signal output
rlabel metal2 s 167160 14200 167272 15000 6 la_data_in_core[41]
port 41 nsew signal output
rlabel metal2 s 169288 14200 169400 15000 6 la_data_in_core[42]
port 42 nsew signal output
rlabel metal2 s 171528 14200 171640 15000 6 la_data_in_core[43]
port 43 nsew signal output
rlabel metal2 s 173656 14200 173768 15000 6 la_data_in_core[44]
port 44 nsew signal output
rlabel metal2 s 175896 14200 176008 15000 6 la_data_in_core[45]
port 45 nsew signal output
rlabel metal2 s 178024 14200 178136 15000 6 la_data_in_core[46]
port 46 nsew signal output
rlabel metal2 s 180264 14200 180376 15000 6 la_data_in_core[47]
port 47 nsew signal output
rlabel metal2 s 182392 14200 182504 15000 6 la_data_in_core[48]
port 48 nsew signal output
rlabel metal2 s 184632 14200 184744 15000 6 la_data_in_core[49]
port 49 nsew signal output
rlabel metal2 s 86184 14200 86296 15000 6 la_data_in_core[4]
port 50 nsew signal output
rlabel metal2 s 186760 14200 186872 15000 6 la_data_in_core[50]
port 51 nsew signal output
rlabel metal2 s 189000 14200 189112 15000 6 la_data_in_core[51]
port 52 nsew signal output
rlabel metal2 s 191128 14200 191240 15000 6 la_data_in_core[52]
port 53 nsew signal output
rlabel metal2 s 193368 14200 193480 15000 6 la_data_in_core[53]
port 54 nsew signal output
rlabel metal2 s 195496 14200 195608 15000 6 la_data_in_core[54]
port 55 nsew signal output
rlabel metal2 s 197736 14200 197848 15000 6 la_data_in_core[55]
port 56 nsew signal output
rlabel metal2 s 199864 14200 199976 15000 6 la_data_in_core[56]
port 57 nsew signal output
rlabel metal2 s 202104 14200 202216 15000 6 la_data_in_core[57]
port 58 nsew signal output
rlabel metal2 s 204232 14200 204344 15000 6 la_data_in_core[58]
port 59 nsew signal output
rlabel metal2 s 206472 14200 206584 15000 6 la_data_in_core[59]
port 60 nsew signal output
rlabel metal2 s 88424 14200 88536 15000 6 la_data_in_core[5]
port 61 nsew signal output
rlabel metal2 s 208600 14200 208712 15000 6 la_data_in_core[60]
port 62 nsew signal output
rlabel metal2 s 210840 14200 210952 15000 6 la_data_in_core[61]
port 63 nsew signal output
rlabel metal2 s 212968 14200 213080 15000 6 la_data_in_core[62]
port 64 nsew signal output
rlabel metal2 s 215208 14200 215320 15000 6 la_data_in_core[63]
port 65 nsew signal output
rlabel metal2 s 90552 14200 90664 15000 6 la_data_in_core[6]
port 66 nsew signal output
rlabel metal2 s 92792 14200 92904 15000 6 la_data_in_core[7]
port 67 nsew signal output
rlabel metal2 s 94920 14200 95032 15000 6 la_data_in_core[8]
port 68 nsew signal output
rlabel metal2 s 97160 14200 97272 15000 6 la_data_in_core[9]
port 69 nsew signal output
rlabel metal2 s 168 0 280 800 6 la_data_in_mprj[0]
port 70 nsew signal output
rlabel metal2 s 6216 0 6328 800 6 la_data_in_mprj[10]
port 71 nsew signal output
rlabel metal2 s 6776 0 6888 800 6 la_data_in_mprj[11]
port 72 nsew signal output
rlabel metal2 s 7448 0 7560 800 6 la_data_in_mprj[12]
port 73 nsew signal output
rlabel metal2 s 8008 0 8120 800 6 la_data_in_mprj[13]
port 74 nsew signal output
rlabel metal2 s 8680 0 8792 800 6 la_data_in_mprj[14]
port 75 nsew signal output
rlabel metal2 s 9240 0 9352 800 6 la_data_in_mprj[15]
port 76 nsew signal output
rlabel metal2 s 9912 0 10024 800 6 la_data_in_mprj[16]
port 77 nsew signal output
rlabel metal2 s 10472 0 10584 800 6 la_data_in_mprj[17]
port 78 nsew signal output
rlabel metal2 s 11032 0 11144 800 6 la_data_in_mprj[18]
port 79 nsew signal output
rlabel metal2 s 11704 0 11816 800 6 la_data_in_mprj[19]
port 80 nsew signal output
rlabel metal2 s 728 0 840 800 6 la_data_in_mprj[1]
port 81 nsew signal output
rlabel metal2 s 12264 0 12376 800 6 la_data_in_mprj[20]
port 82 nsew signal output
rlabel metal2 s 12936 0 13048 800 6 la_data_in_mprj[21]
port 83 nsew signal output
rlabel metal2 s 13496 0 13608 800 6 la_data_in_mprj[22]
port 84 nsew signal output
rlabel metal2 s 14168 0 14280 800 6 la_data_in_mprj[23]
port 85 nsew signal output
rlabel metal2 s 14728 0 14840 800 6 la_data_in_mprj[24]
port 86 nsew signal output
rlabel metal2 s 15400 0 15512 800 6 la_data_in_mprj[25]
port 87 nsew signal output
rlabel metal2 s 15960 0 16072 800 6 la_data_in_mprj[26]
port 88 nsew signal output
rlabel metal2 s 16520 0 16632 800 6 la_data_in_mprj[27]
port 89 nsew signal output
rlabel metal2 s 17192 0 17304 800 6 la_data_in_mprj[28]
port 90 nsew signal output
rlabel metal2 s 17752 0 17864 800 6 la_data_in_mprj[29]
port 91 nsew signal output
rlabel metal2 s 1288 0 1400 800 6 la_data_in_mprj[2]
port 92 nsew signal output
rlabel metal2 s 18424 0 18536 800 6 la_data_in_mprj[30]
port 93 nsew signal output
rlabel metal2 s 18984 0 19096 800 6 la_data_in_mprj[31]
port 94 nsew signal output
rlabel metal2 s 19656 0 19768 800 6 la_data_in_mprj[32]
port 95 nsew signal output
rlabel metal2 s 20216 0 20328 800 6 la_data_in_mprj[33]
port 96 nsew signal output
rlabel metal2 s 20888 0 21000 800 6 la_data_in_mprj[34]
port 97 nsew signal output
rlabel metal2 s 21448 0 21560 800 6 la_data_in_mprj[35]
port 98 nsew signal output
rlabel metal2 s 22008 0 22120 800 6 la_data_in_mprj[36]
port 99 nsew signal output
rlabel metal2 s 22680 0 22792 800 6 la_data_in_mprj[37]
port 100 nsew signal output
rlabel metal2 s 23240 0 23352 800 6 la_data_in_mprj[38]
port 101 nsew signal output
rlabel metal2 s 23912 0 24024 800 6 la_data_in_mprj[39]
port 102 nsew signal output
rlabel metal2 s 1960 0 2072 800 6 la_data_in_mprj[3]
port 103 nsew signal output
rlabel metal2 s 24472 0 24584 800 6 la_data_in_mprj[40]
port 104 nsew signal output
rlabel metal2 s 25144 0 25256 800 6 la_data_in_mprj[41]
port 105 nsew signal output
rlabel metal2 s 25704 0 25816 800 6 la_data_in_mprj[42]
port 106 nsew signal output
rlabel metal2 s 26376 0 26488 800 6 la_data_in_mprj[43]
port 107 nsew signal output
rlabel metal2 s 26936 0 27048 800 6 la_data_in_mprj[44]
port 108 nsew signal output
rlabel metal2 s 27496 0 27608 800 6 la_data_in_mprj[45]
port 109 nsew signal output
rlabel metal2 s 28168 0 28280 800 6 la_data_in_mprj[46]
port 110 nsew signal output
rlabel metal2 s 28728 0 28840 800 6 la_data_in_mprj[47]
port 111 nsew signal output
rlabel metal2 s 29400 0 29512 800 6 la_data_in_mprj[48]
port 112 nsew signal output
rlabel metal2 s 29960 0 30072 800 6 la_data_in_mprj[49]
port 113 nsew signal output
rlabel metal2 s 2520 0 2632 800 6 la_data_in_mprj[4]
port 114 nsew signal output
rlabel metal2 s 30632 0 30744 800 6 la_data_in_mprj[50]
port 115 nsew signal output
rlabel metal2 s 31192 0 31304 800 6 la_data_in_mprj[51]
port 116 nsew signal output
rlabel metal2 s 31864 0 31976 800 6 la_data_in_mprj[52]
port 117 nsew signal output
rlabel metal2 s 32424 0 32536 800 6 la_data_in_mprj[53]
port 118 nsew signal output
rlabel metal2 s 32984 0 33096 800 6 la_data_in_mprj[54]
port 119 nsew signal output
rlabel metal2 s 33656 0 33768 800 6 la_data_in_mprj[55]
port 120 nsew signal output
rlabel metal2 s 34216 0 34328 800 6 la_data_in_mprj[56]
port 121 nsew signal output
rlabel metal2 s 34888 0 35000 800 6 la_data_in_mprj[57]
port 122 nsew signal output
rlabel metal2 s 35448 0 35560 800 6 la_data_in_mprj[58]
port 123 nsew signal output
rlabel metal2 s 36120 0 36232 800 6 la_data_in_mprj[59]
port 124 nsew signal output
rlabel metal2 s 3192 0 3304 800 6 la_data_in_mprj[5]
port 125 nsew signal output
rlabel metal2 s 36680 0 36792 800 6 la_data_in_mprj[60]
port 126 nsew signal output
rlabel metal2 s 37352 0 37464 800 6 la_data_in_mprj[61]
port 127 nsew signal output
rlabel metal2 s 37912 0 38024 800 6 la_data_in_mprj[62]
port 128 nsew signal output
rlabel metal2 s 38472 0 38584 800 6 la_data_in_mprj[63]
port 129 nsew signal output
rlabel metal2 s 3752 0 3864 800 6 la_data_in_mprj[6]
port 130 nsew signal output
rlabel metal2 s 4424 0 4536 800 6 la_data_in_mprj[7]
port 131 nsew signal output
rlabel metal2 s 4984 0 5096 800 6 la_data_in_mprj[8]
port 132 nsew signal output
rlabel metal2 s 5544 0 5656 800 6 la_data_in_mprj[9]
port 133 nsew signal output
rlabel metal2 s 78232 14200 78344 15000 6 la_data_out_core[0]
port 134 nsew signal input
rlabel metal2 s 100072 14200 100184 15000 6 la_data_out_core[10]
port 135 nsew signal input
rlabel metal2 s 102200 14200 102312 15000 6 la_data_out_core[11]
port 136 nsew signal input
rlabel metal2 s 104440 14200 104552 15000 6 la_data_out_core[12]
port 137 nsew signal input
rlabel metal2 s 106568 14200 106680 15000 6 la_data_out_core[13]
port 138 nsew signal input
rlabel metal2 s 108808 14200 108920 15000 6 la_data_out_core[14]
port 139 nsew signal input
rlabel metal2 s 111048 14200 111160 15000 6 la_data_out_core[15]
port 140 nsew signal input
rlabel metal2 s 113176 14200 113288 15000 6 la_data_out_core[16]
port 141 nsew signal input
rlabel metal2 s 115416 14200 115528 15000 6 la_data_out_core[17]
port 142 nsew signal input
rlabel metal2 s 117544 14200 117656 15000 6 la_data_out_core[18]
port 143 nsew signal input
rlabel metal2 s 119784 14200 119896 15000 6 la_data_out_core[19]
port 144 nsew signal input
rlabel metal2 s 80360 14200 80472 15000 6 la_data_out_core[1]
port 145 nsew signal input
rlabel metal2 s 121912 14200 122024 15000 6 la_data_out_core[20]
port 146 nsew signal input
rlabel metal2 s 124152 14200 124264 15000 6 la_data_out_core[21]
port 147 nsew signal input
rlabel metal2 s 126280 14200 126392 15000 6 la_data_out_core[22]
port 148 nsew signal input
rlabel metal2 s 128520 14200 128632 15000 6 la_data_out_core[23]
port 149 nsew signal input
rlabel metal2 s 130648 14200 130760 15000 6 la_data_out_core[24]
port 150 nsew signal input
rlabel metal2 s 132888 14200 133000 15000 6 la_data_out_core[25]
port 151 nsew signal input
rlabel metal2 s 135016 14200 135128 15000 6 la_data_out_core[26]
port 152 nsew signal input
rlabel metal2 s 137256 14200 137368 15000 6 la_data_out_core[27]
port 153 nsew signal input
rlabel metal2 s 139384 14200 139496 15000 6 la_data_out_core[28]
port 154 nsew signal input
rlabel metal2 s 141624 14200 141736 15000 6 la_data_out_core[29]
port 155 nsew signal input
rlabel metal2 s 82600 14200 82712 15000 6 la_data_out_core[2]
port 156 nsew signal input
rlabel metal2 s 143752 14200 143864 15000 6 la_data_out_core[30]
port 157 nsew signal input
rlabel metal2 s 145992 14200 146104 15000 6 la_data_out_core[31]
port 158 nsew signal input
rlabel metal2 s 148120 14200 148232 15000 6 la_data_out_core[32]
port 159 nsew signal input
rlabel metal2 s 150360 14200 150472 15000 6 la_data_out_core[33]
port 160 nsew signal input
rlabel metal2 s 152488 14200 152600 15000 6 la_data_out_core[34]
port 161 nsew signal input
rlabel metal2 s 154728 14200 154840 15000 6 la_data_out_core[35]
port 162 nsew signal input
rlabel metal2 s 156856 14200 156968 15000 6 la_data_out_core[36]
port 163 nsew signal input
rlabel metal2 s 159096 14200 159208 15000 6 la_data_out_core[37]
port 164 nsew signal input
rlabel metal2 s 161224 14200 161336 15000 6 la_data_out_core[38]
port 165 nsew signal input
rlabel metal2 s 163464 14200 163576 15000 6 la_data_out_core[39]
port 166 nsew signal input
rlabel metal2 s 84728 14200 84840 15000 6 la_data_out_core[3]
port 167 nsew signal input
rlabel metal2 s 165704 14200 165816 15000 6 la_data_out_core[40]
port 168 nsew signal input
rlabel metal2 s 167832 14200 167944 15000 6 la_data_out_core[41]
port 169 nsew signal input
rlabel metal2 s 170072 14200 170184 15000 6 la_data_out_core[42]
port 170 nsew signal input
rlabel metal2 s 172200 14200 172312 15000 6 la_data_out_core[43]
port 171 nsew signal input
rlabel metal2 s 174440 14200 174552 15000 6 la_data_out_core[44]
port 172 nsew signal input
rlabel metal2 s 176568 14200 176680 15000 6 la_data_out_core[45]
port 173 nsew signal input
rlabel metal2 s 178808 14200 178920 15000 6 la_data_out_core[46]
port 174 nsew signal input
rlabel metal2 s 180936 14200 181048 15000 6 la_data_out_core[47]
port 175 nsew signal input
rlabel metal2 s 183176 14200 183288 15000 6 la_data_out_core[48]
port 176 nsew signal input
rlabel metal2 s 185304 14200 185416 15000 6 la_data_out_core[49]
port 177 nsew signal input
rlabel metal2 s 86968 14200 87080 15000 6 la_data_out_core[4]
port 178 nsew signal input
rlabel metal2 s 187544 14200 187656 15000 6 la_data_out_core[50]
port 179 nsew signal input
rlabel metal2 s 189672 14200 189784 15000 6 la_data_out_core[51]
port 180 nsew signal input
rlabel metal2 s 191912 14200 192024 15000 6 la_data_out_core[52]
port 181 nsew signal input
rlabel metal2 s 194040 14200 194152 15000 6 la_data_out_core[53]
port 182 nsew signal input
rlabel metal2 s 196280 14200 196392 15000 6 la_data_out_core[54]
port 183 nsew signal input
rlabel metal2 s 198408 14200 198520 15000 6 la_data_out_core[55]
port 184 nsew signal input
rlabel metal2 s 200648 14200 200760 15000 6 la_data_out_core[56]
port 185 nsew signal input
rlabel metal2 s 202776 14200 202888 15000 6 la_data_out_core[57]
port 186 nsew signal input
rlabel metal2 s 205016 14200 205128 15000 6 la_data_out_core[58]
port 187 nsew signal input
rlabel metal2 s 207144 14200 207256 15000 6 la_data_out_core[59]
port 188 nsew signal input
rlabel metal2 s 89096 14200 89208 15000 6 la_data_out_core[5]
port 189 nsew signal input
rlabel metal2 s 209384 14200 209496 15000 6 la_data_out_core[60]
port 190 nsew signal input
rlabel metal2 s 211512 14200 211624 15000 6 la_data_out_core[61]
port 191 nsew signal input
rlabel metal2 s 213752 14200 213864 15000 6 la_data_out_core[62]
port 192 nsew signal input
rlabel metal2 s 215880 14200 215992 15000 6 la_data_out_core[63]
port 193 nsew signal input
rlabel metal2 s 91336 14200 91448 15000 6 la_data_out_core[6]
port 194 nsew signal input
rlabel metal2 s 93464 14200 93576 15000 6 la_data_out_core[7]
port 195 nsew signal input
rlabel metal2 s 95704 14200 95816 15000 6 la_data_out_core[8]
port 196 nsew signal input
rlabel metal2 s 97832 14200 97944 15000 6 la_data_out_core[9]
port 197 nsew signal input
rlabel metal2 s 39144 0 39256 800 6 la_data_out_mprj[0]
port 198 nsew signal input
rlabel metal2 s 45192 0 45304 800 6 la_data_out_mprj[10]
port 199 nsew signal input
rlabel metal2 s 45864 0 45976 800 6 la_data_out_mprj[11]
port 200 nsew signal input
rlabel metal2 s 46424 0 46536 800 6 la_data_out_mprj[12]
port 201 nsew signal input
rlabel metal2 s 47096 0 47208 800 6 la_data_out_mprj[13]
port 202 nsew signal input
rlabel metal2 s 47656 0 47768 800 6 la_data_out_mprj[14]
port 203 nsew signal input
rlabel metal2 s 48328 0 48440 800 6 la_data_out_mprj[15]
port 204 nsew signal input
rlabel metal2 s 48888 0 49000 800 6 la_data_out_mprj[16]
port 205 nsew signal input
rlabel metal2 s 49448 0 49560 800 6 la_data_out_mprj[17]
port 206 nsew signal input
rlabel metal2 s 50120 0 50232 800 6 la_data_out_mprj[18]
port 207 nsew signal input
rlabel metal2 s 50680 0 50792 800 6 la_data_out_mprj[19]
port 208 nsew signal input
rlabel metal2 s 39704 0 39816 800 6 la_data_out_mprj[1]
port 209 nsew signal input
rlabel metal2 s 51352 0 51464 800 6 la_data_out_mprj[20]
port 210 nsew signal input
rlabel metal2 s 51912 0 52024 800 6 la_data_out_mprj[21]
port 211 nsew signal input
rlabel metal2 s 52584 0 52696 800 6 la_data_out_mprj[22]
port 212 nsew signal input
rlabel metal2 s 53144 0 53256 800 6 la_data_out_mprj[23]
port 213 nsew signal input
rlabel metal2 s 53816 0 53928 800 6 la_data_out_mprj[24]
port 214 nsew signal input
rlabel metal2 s 54376 0 54488 800 6 la_data_out_mprj[25]
port 215 nsew signal input
rlabel metal2 s 54936 0 55048 800 6 la_data_out_mprj[26]
port 216 nsew signal input
rlabel metal2 s 55608 0 55720 800 6 la_data_out_mprj[27]
port 217 nsew signal input
rlabel metal2 s 56168 0 56280 800 6 la_data_out_mprj[28]
port 218 nsew signal input
rlabel metal2 s 56840 0 56952 800 6 la_data_out_mprj[29]
port 219 nsew signal input
rlabel metal2 s 40376 0 40488 800 6 la_data_out_mprj[2]
port 220 nsew signal input
rlabel metal2 s 57400 0 57512 800 6 la_data_out_mprj[30]
port 221 nsew signal input
rlabel metal2 s 58072 0 58184 800 6 la_data_out_mprj[31]
port 222 nsew signal input
rlabel metal2 s 58632 0 58744 800 6 la_data_out_mprj[32]
port 223 nsew signal input
rlabel metal2 s 59192 0 59304 800 6 la_data_out_mprj[33]
port 224 nsew signal input
rlabel metal2 s 59864 0 59976 800 6 la_data_out_mprj[34]
port 225 nsew signal input
rlabel metal2 s 60424 0 60536 800 6 la_data_out_mprj[35]
port 226 nsew signal input
rlabel metal2 s 61096 0 61208 800 6 la_data_out_mprj[36]
port 227 nsew signal input
rlabel metal2 s 61656 0 61768 800 6 la_data_out_mprj[37]
port 228 nsew signal input
rlabel metal2 s 62328 0 62440 800 6 la_data_out_mprj[38]
port 229 nsew signal input
rlabel metal2 s 62888 0 63000 800 6 la_data_out_mprj[39]
port 230 nsew signal input
rlabel metal2 s 40936 0 41048 800 6 la_data_out_mprj[3]
port 231 nsew signal input
rlabel metal2 s 63560 0 63672 800 6 la_data_out_mprj[40]
port 232 nsew signal input
rlabel metal2 s 64120 0 64232 800 6 la_data_out_mprj[41]
port 233 nsew signal input
rlabel metal2 s 64680 0 64792 800 6 la_data_out_mprj[42]
port 234 nsew signal input
rlabel metal2 s 65352 0 65464 800 6 la_data_out_mprj[43]
port 235 nsew signal input
rlabel metal2 s 65912 0 66024 800 6 la_data_out_mprj[44]
port 236 nsew signal input
rlabel metal2 s 66584 0 66696 800 6 la_data_out_mprj[45]
port 237 nsew signal input
rlabel metal2 s 67144 0 67256 800 6 la_data_out_mprj[46]
port 238 nsew signal input
rlabel metal2 s 67816 0 67928 800 6 la_data_out_mprj[47]
port 239 nsew signal input
rlabel metal2 s 68376 0 68488 800 6 la_data_out_mprj[48]
port 240 nsew signal input
rlabel metal2 s 69048 0 69160 800 6 la_data_out_mprj[49]
port 241 nsew signal input
rlabel metal2 s 41608 0 41720 800 6 la_data_out_mprj[4]
port 242 nsew signal input
rlabel metal2 s 69608 0 69720 800 6 la_data_out_mprj[50]
port 243 nsew signal input
rlabel metal2 s 70168 0 70280 800 6 la_data_out_mprj[51]
port 244 nsew signal input
rlabel metal2 s 70840 0 70952 800 6 la_data_out_mprj[52]
port 245 nsew signal input
rlabel metal2 s 71400 0 71512 800 6 la_data_out_mprj[53]
port 246 nsew signal input
rlabel metal2 s 72072 0 72184 800 6 la_data_out_mprj[54]
port 247 nsew signal input
rlabel metal2 s 72632 0 72744 800 6 la_data_out_mprj[55]
port 248 nsew signal input
rlabel metal2 s 73304 0 73416 800 6 la_data_out_mprj[56]
port 249 nsew signal input
rlabel metal2 s 73864 0 73976 800 6 la_data_out_mprj[57]
port 250 nsew signal input
rlabel metal2 s 74536 0 74648 800 6 la_data_out_mprj[58]
port 251 nsew signal input
rlabel metal2 s 75096 0 75208 800 6 la_data_out_mprj[59]
port 252 nsew signal input
rlabel metal2 s 42168 0 42280 800 6 la_data_out_mprj[5]
port 253 nsew signal input
rlabel metal2 s 75656 0 75768 800 6 la_data_out_mprj[60]
port 254 nsew signal input
rlabel metal2 s 76328 0 76440 800 6 la_data_out_mprj[61]
port 255 nsew signal input
rlabel metal2 s 76888 0 77000 800 6 la_data_out_mprj[62]
port 256 nsew signal input
rlabel metal2 s 77560 0 77672 800 6 la_data_out_mprj[63]
port 257 nsew signal input
rlabel metal2 s 42840 0 42952 800 6 la_data_out_mprj[6]
port 258 nsew signal input
rlabel metal2 s 43400 0 43512 800 6 la_data_out_mprj[7]
port 259 nsew signal input
rlabel metal2 s 43960 0 44072 800 6 la_data_out_mprj[8]
port 260 nsew signal input
rlabel metal2 s 44632 0 44744 800 6 la_data_out_mprj[9]
port 261 nsew signal input
rlabel metal2 s 117208 0 117320 800 6 la_iena_mprj[0]
port 262 nsew signal input
rlabel metal2 s 123256 0 123368 800 6 la_iena_mprj[10]
port 263 nsew signal input
rlabel metal2 s 123816 0 123928 800 6 la_iena_mprj[11]
port 264 nsew signal input
rlabel metal2 s 124488 0 124600 800 6 la_iena_mprj[12]
port 265 nsew signal input
rlabel metal2 s 125048 0 125160 800 6 la_iena_mprj[13]
port 266 nsew signal input
rlabel metal2 s 125720 0 125832 800 6 la_iena_mprj[14]
port 267 nsew signal input
rlabel metal2 s 126280 0 126392 800 6 la_iena_mprj[15]
port 268 nsew signal input
rlabel metal2 s 126952 0 127064 800 6 la_iena_mprj[16]
port 269 nsew signal input
rlabel metal2 s 127512 0 127624 800 6 la_iena_mprj[17]
port 270 nsew signal input
rlabel metal2 s 128184 0 128296 800 6 la_iena_mprj[18]
port 271 nsew signal input
rlabel metal2 s 128744 0 128856 800 6 la_iena_mprj[19]
port 272 nsew signal input
rlabel metal2 s 117768 0 117880 800 6 la_iena_mprj[1]
port 273 nsew signal input
rlabel metal2 s 129304 0 129416 800 6 la_iena_mprj[20]
port 274 nsew signal input
rlabel metal2 s 129976 0 130088 800 6 la_iena_mprj[21]
port 275 nsew signal input
rlabel metal2 s 130536 0 130648 800 6 la_iena_mprj[22]
port 276 nsew signal input
rlabel metal2 s 131208 0 131320 800 6 la_iena_mprj[23]
port 277 nsew signal input
rlabel metal2 s 131768 0 131880 800 6 la_iena_mprj[24]
port 278 nsew signal input
rlabel metal2 s 132440 0 132552 800 6 la_iena_mprj[25]
port 279 nsew signal input
rlabel metal2 s 133000 0 133112 800 6 la_iena_mprj[26]
port 280 nsew signal input
rlabel metal2 s 133672 0 133784 800 6 la_iena_mprj[27]
port 281 nsew signal input
rlabel metal2 s 134232 0 134344 800 6 la_iena_mprj[28]
port 282 nsew signal input
rlabel metal2 s 134792 0 134904 800 6 la_iena_mprj[29]
port 283 nsew signal input
rlabel metal2 s 118328 0 118440 800 6 la_iena_mprj[2]
port 284 nsew signal input
rlabel metal2 s 135464 0 135576 800 6 la_iena_mprj[30]
port 285 nsew signal input
rlabel metal2 s 136024 0 136136 800 6 la_iena_mprj[31]
port 286 nsew signal input
rlabel metal2 s 136696 0 136808 800 6 la_iena_mprj[32]
port 287 nsew signal input
rlabel metal2 s 137256 0 137368 800 6 la_iena_mprj[33]
port 288 nsew signal input
rlabel metal2 s 137928 0 138040 800 6 la_iena_mprj[34]
port 289 nsew signal input
rlabel metal2 s 138488 0 138600 800 6 la_iena_mprj[35]
port 290 nsew signal input
rlabel metal2 s 139160 0 139272 800 6 la_iena_mprj[36]
port 291 nsew signal input
rlabel metal2 s 139720 0 139832 800 6 la_iena_mprj[37]
port 292 nsew signal input
rlabel metal2 s 140280 0 140392 800 6 la_iena_mprj[38]
port 293 nsew signal input
rlabel metal2 s 140952 0 141064 800 6 la_iena_mprj[39]
port 294 nsew signal input
rlabel metal2 s 119000 0 119112 800 6 la_iena_mprj[3]
port 295 nsew signal input
rlabel metal2 s 141512 0 141624 800 6 la_iena_mprj[40]
port 296 nsew signal input
rlabel metal2 s 142184 0 142296 800 6 la_iena_mprj[41]
port 297 nsew signal input
rlabel metal2 s 142744 0 142856 800 6 la_iena_mprj[42]
port 298 nsew signal input
rlabel metal2 s 143416 0 143528 800 6 la_iena_mprj[43]
port 299 nsew signal input
rlabel metal2 s 143976 0 144088 800 6 la_iena_mprj[44]
port 300 nsew signal input
rlabel metal2 s 144648 0 144760 800 6 la_iena_mprj[45]
port 301 nsew signal input
rlabel metal2 s 145208 0 145320 800 6 la_iena_mprj[46]
port 302 nsew signal input
rlabel metal2 s 145768 0 145880 800 6 la_iena_mprj[47]
port 303 nsew signal input
rlabel metal2 s 146440 0 146552 800 6 la_iena_mprj[48]
port 304 nsew signal input
rlabel metal2 s 147000 0 147112 800 6 la_iena_mprj[49]
port 305 nsew signal input
rlabel metal2 s 119560 0 119672 800 6 la_iena_mprj[4]
port 306 nsew signal input
rlabel metal2 s 147672 0 147784 800 6 la_iena_mprj[50]
port 307 nsew signal input
rlabel metal2 s 148232 0 148344 800 6 la_iena_mprj[51]
port 308 nsew signal input
rlabel metal2 s 148904 0 149016 800 6 la_iena_mprj[52]
port 309 nsew signal input
rlabel metal2 s 149464 0 149576 800 6 la_iena_mprj[53]
port 310 nsew signal input
rlabel metal2 s 150136 0 150248 800 6 la_iena_mprj[54]
port 311 nsew signal input
rlabel metal2 s 150696 0 150808 800 6 la_iena_mprj[55]
port 312 nsew signal input
rlabel metal2 s 151256 0 151368 800 6 la_iena_mprj[56]
port 313 nsew signal input
rlabel metal2 s 151928 0 152040 800 6 la_iena_mprj[57]
port 314 nsew signal input
rlabel metal2 s 152488 0 152600 800 6 la_iena_mprj[58]
port 315 nsew signal input
rlabel metal2 s 153160 0 153272 800 6 la_iena_mprj[59]
port 316 nsew signal input
rlabel metal2 s 120232 0 120344 800 6 la_iena_mprj[5]
port 317 nsew signal input
rlabel metal2 s 153720 0 153832 800 6 la_iena_mprj[60]
port 318 nsew signal input
rlabel metal2 s 154392 0 154504 800 6 la_iena_mprj[61]
port 319 nsew signal input
rlabel metal2 s 154952 0 155064 800 6 la_iena_mprj[62]
port 320 nsew signal input
rlabel metal2 s 155624 0 155736 800 6 la_iena_mprj[63]
port 321 nsew signal input
rlabel metal2 s 120792 0 120904 800 6 la_iena_mprj[6]
port 322 nsew signal input
rlabel metal2 s 121464 0 121576 800 6 la_iena_mprj[7]
port 323 nsew signal input
rlabel metal2 s 122024 0 122136 800 6 la_iena_mprj[8]
port 324 nsew signal input
rlabel metal2 s 122696 0 122808 800 6 la_iena_mprj[9]
port 325 nsew signal input
rlabel metal2 s 78904 14200 79016 15000 6 la_oenb_core[0]
port 326 nsew signal output
rlabel metal2 s 100744 14200 100856 15000 6 la_oenb_core[10]
port 327 nsew signal output
rlabel metal2 s 102984 14200 103096 15000 6 la_oenb_core[11]
port 328 nsew signal output
rlabel metal2 s 105112 14200 105224 15000 6 la_oenb_core[12]
port 329 nsew signal output
rlabel metal2 s 107352 14200 107464 15000 6 la_oenb_core[13]
port 330 nsew signal output
rlabel metal2 s 109480 14200 109592 15000 6 la_oenb_core[14]
port 331 nsew signal output
rlabel metal2 s 111720 14200 111832 15000 6 la_oenb_core[15]
port 332 nsew signal output
rlabel metal2 s 113960 14200 114072 15000 6 la_oenb_core[16]
port 333 nsew signal output
rlabel metal2 s 116088 14200 116200 15000 6 la_oenb_core[17]
port 334 nsew signal output
rlabel metal2 s 118328 14200 118440 15000 6 la_oenb_core[18]
port 335 nsew signal output
rlabel metal2 s 120456 14200 120568 15000 6 la_oenb_core[19]
port 336 nsew signal output
rlabel metal2 s 81144 14200 81256 15000 6 la_oenb_core[1]
port 337 nsew signal output
rlabel metal2 s 122696 14200 122808 15000 6 la_oenb_core[20]
port 338 nsew signal output
rlabel metal2 s 124824 14200 124936 15000 6 la_oenb_core[21]
port 339 nsew signal output
rlabel metal2 s 127064 14200 127176 15000 6 la_oenb_core[22]
port 340 nsew signal output
rlabel metal2 s 129192 14200 129304 15000 6 la_oenb_core[23]
port 341 nsew signal output
rlabel metal2 s 131432 14200 131544 15000 6 la_oenb_core[24]
port 342 nsew signal output
rlabel metal2 s 133560 14200 133672 15000 6 la_oenb_core[25]
port 343 nsew signal output
rlabel metal2 s 135800 14200 135912 15000 6 la_oenb_core[26]
port 344 nsew signal output
rlabel metal2 s 137928 14200 138040 15000 6 la_oenb_core[27]
port 345 nsew signal output
rlabel metal2 s 140168 14200 140280 15000 6 la_oenb_core[28]
port 346 nsew signal output
rlabel metal2 s 142296 14200 142408 15000 6 la_oenb_core[29]
port 347 nsew signal output
rlabel metal2 s 83272 14200 83384 15000 6 la_oenb_core[2]
port 348 nsew signal output
rlabel metal2 s 144536 14200 144648 15000 6 la_oenb_core[30]
port 349 nsew signal output
rlabel metal2 s 146664 14200 146776 15000 6 la_oenb_core[31]
port 350 nsew signal output
rlabel metal2 s 148904 14200 149016 15000 6 la_oenb_core[32]
port 351 nsew signal output
rlabel metal2 s 151032 14200 151144 15000 6 la_oenb_core[33]
port 352 nsew signal output
rlabel metal2 s 153272 14200 153384 15000 6 la_oenb_core[34]
port 353 nsew signal output
rlabel metal2 s 155400 14200 155512 15000 6 la_oenb_core[35]
port 354 nsew signal output
rlabel metal2 s 157640 14200 157752 15000 6 la_oenb_core[36]
port 355 nsew signal output
rlabel metal2 s 159768 14200 159880 15000 6 la_oenb_core[37]
port 356 nsew signal output
rlabel metal2 s 162008 14200 162120 15000 6 la_oenb_core[38]
port 357 nsew signal output
rlabel metal2 s 164136 14200 164248 15000 6 la_oenb_core[39]
port 358 nsew signal output
rlabel metal2 s 85512 14200 85624 15000 6 la_oenb_core[3]
port 359 nsew signal output
rlabel metal2 s 166376 14200 166488 15000 6 la_oenb_core[40]
port 360 nsew signal output
rlabel metal2 s 168616 14200 168728 15000 6 la_oenb_core[41]
port 361 nsew signal output
rlabel metal2 s 170744 14200 170856 15000 6 la_oenb_core[42]
port 362 nsew signal output
rlabel metal2 s 172984 14200 173096 15000 6 la_oenb_core[43]
port 363 nsew signal output
rlabel metal2 s 175112 14200 175224 15000 6 la_oenb_core[44]
port 364 nsew signal output
rlabel metal2 s 177352 14200 177464 15000 6 la_oenb_core[45]
port 365 nsew signal output
rlabel metal2 s 179480 14200 179592 15000 6 la_oenb_core[46]
port 366 nsew signal output
rlabel metal2 s 181720 14200 181832 15000 6 la_oenb_core[47]
port 367 nsew signal output
rlabel metal2 s 183848 14200 183960 15000 6 la_oenb_core[48]
port 368 nsew signal output
rlabel metal2 s 186088 14200 186200 15000 6 la_oenb_core[49]
port 369 nsew signal output
rlabel metal2 s 87640 14200 87752 15000 6 la_oenb_core[4]
port 370 nsew signal output
rlabel metal2 s 188216 14200 188328 15000 6 la_oenb_core[50]
port 371 nsew signal output
rlabel metal2 s 190456 14200 190568 15000 6 la_oenb_core[51]
port 372 nsew signal output
rlabel metal2 s 192584 14200 192696 15000 6 la_oenb_core[52]
port 373 nsew signal output
rlabel metal2 s 194824 14200 194936 15000 6 la_oenb_core[53]
port 374 nsew signal output
rlabel metal2 s 196952 14200 197064 15000 6 la_oenb_core[54]
port 375 nsew signal output
rlabel metal2 s 199192 14200 199304 15000 6 la_oenb_core[55]
port 376 nsew signal output
rlabel metal2 s 201320 14200 201432 15000 6 la_oenb_core[56]
port 377 nsew signal output
rlabel metal2 s 203560 14200 203672 15000 6 la_oenb_core[57]
port 378 nsew signal output
rlabel metal2 s 205688 14200 205800 15000 6 la_oenb_core[58]
port 379 nsew signal output
rlabel metal2 s 207928 14200 208040 15000 6 la_oenb_core[59]
port 380 nsew signal output
rlabel metal2 s 89880 14200 89992 15000 6 la_oenb_core[5]
port 381 nsew signal output
rlabel metal2 s 210056 14200 210168 15000 6 la_oenb_core[60]
port 382 nsew signal output
rlabel metal2 s 212296 14200 212408 15000 6 la_oenb_core[61]
port 383 nsew signal output
rlabel metal2 s 214424 14200 214536 15000 6 la_oenb_core[62]
port 384 nsew signal output
rlabel metal2 s 216664 14200 216776 15000 6 la_oenb_core[63]
port 385 nsew signal output
rlabel metal2 s 92008 14200 92120 15000 6 la_oenb_core[6]
port 386 nsew signal output
rlabel metal2 s 94248 14200 94360 15000 6 la_oenb_core[7]
port 387 nsew signal output
rlabel metal2 s 96376 14200 96488 15000 6 la_oenb_core[8]
port 388 nsew signal output
rlabel metal2 s 98616 14200 98728 15000 6 la_oenb_core[9]
port 389 nsew signal output
rlabel metal2 s 78120 0 78232 800 6 la_oenb_mprj[0]
port 390 nsew signal input
rlabel metal2 s 84280 0 84392 800 6 la_oenb_mprj[10]
port 391 nsew signal input
rlabel metal2 s 84840 0 84952 800 6 la_oenb_mprj[11]
port 392 nsew signal input
rlabel metal2 s 85512 0 85624 800 6 la_oenb_mprj[12]
port 393 nsew signal input
rlabel metal2 s 86072 0 86184 800 6 la_oenb_mprj[13]
port 394 nsew signal input
rlabel metal2 s 86632 0 86744 800 6 la_oenb_mprj[14]
port 395 nsew signal input
rlabel metal2 s 87304 0 87416 800 6 la_oenb_mprj[15]
port 396 nsew signal input
rlabel metal2 s 87864 0 87976 800 6 la_oenb_mprj[16]
port 397 nsew signal input
rlabel metal2 s 88536 0 88648 800 6 la_oenb_mprj[17]
port 398 nsew signal input
rlabel metal2 s 89096 0 89208 800 6 la_oenb_mprj[18]
port 399 nsew signal input
rlabel metal2 s 89768 0 89880 800 6 la_oenb_mprj[19]
port 400 nsew signal input
rlabel metal2 s 78792 0 78904 800 6 la_oenb_mprj[1]
port 401 nsew signal input
rlabel metal2 s 90328 0 90440 800 6 la_oenb_mprj[20]
port 402 nsew signal input
rlabel metal2 s 91000 0 91112 800 6 la_oenb_mprj[21]
port 403 nsew signal input
rlabel metal2 s 91560 0 91672 800 6 la_oenb_mprj[22]
port 404 nsew signal input
rlabel metal2 s 92120 0 92232 800 6 la_oenb_mprj[23]
port 405 nsew signal input
rlabel metal2 s 92792 0 92904 800 6 la_oenb_mprj[24]
port 406 nsew signal input
rlabel metal2 s 93352 0 93464 800 6 la_oenb_mprj[25]
port 407 nsew signal input
rlabel metal2 s 94024 0 94136 800 6 la_oenb_mprj[26]
port 408 nsew signal input
rlabel metal2 s 94584 0 94696 800 6 la_oenb_mprj[27]
port 409 nsew signal input
rlabel metal2 s 95256 0 95368 800 6 la_oenb_mprj[28]
port 410 nsew signal input
rlabel metal2 s 95816 0 95928 800 6 la_oenb_mprj[29]
port 411 nsew signal input
rlabel metal2 s 79352 0 79464 800 6 la_oenb_mprj[2]
port 412 nsew signal input
rlabel metal2 s 96488 0 96600 800 6 la_oenb_mprj[30]
port 413 nsew signal input
rlabel metal2 s 97048 0 97160 800 6 la_oenb_mprj[31]
port 414 nsew signal input
rlabel metal2 s 97608 0 97720 800 6 la_oenb_mprj[32]
port 415 nsew signal input
rlabel metal2 s 98280 0 98392 800 6 la_oenb_mprj[33]
port 416 nsew signal input
rlabel metal2 s 98840 0 98952 800 6 la_oenb_mprj[34]
port 417 nsew signal input
rlabel metal2 s 99512 0 99624 800 6 la_oenb_mprj[35]
port 418 nsew signal input
rlabel metal2 s 100072 0 100184 800 6 la_oenb_mprj[36]
port 419 nsew signal input
rlabel metal2 s 100744 0 100856 800 6 la_oenb_mprj[37]
port 420 nsew signal input
rlabel metal2 s 101304 0 101416 800 6 la_oenb_mprj[38]
port 421 nsew signal input
rlabel metal2 s 101976 0 102088 800 6 la_oenb_mprj[39]
port 422 nsew signal input
rlabel metal2 s 80024 0 80136 800 6 la_oenb_mprj[3]
port 423 nsew signal input
rlabel metal2 s 102536 0 102648 800 6 la_oenb_mprj[40]
port 424 nsew signal input
rlabel metal2 s 103096 0 103208 800 6 la_oenb_mprj[41]
port 425 nsew signal input
rlabel metal2 s 103768 0 103880 800 6 la_oenb_mprj[42]
port 426 nsew signal input
rlabel metal2 s 104328 0 104440 800 6 la_oenb_mprj[43]
port 427 nsew signal input
rlabel metal2 s 105000 0 105112 800 6 la_oenb_mprj[44]
port 428 nsew signal input
rlabel metal2 s 105560 0 105672 800 6 la_oenb_mprj[45]
port 429 nsew signal input
rlabel metal2 s 106232 0 106344 800 6 la_oenb_mprj[46]
port 430 nsew signal input
rlabel metal2 s 106792 0 106904 800 6 la_oenb_mprj[47]
port 431 nsew signal input
rlabel metal2 s 107464 0 107576 800 6 la_oenb_mprj[48]
port 432 nsew signal input
rlabel metal2 s 108024 0 108136 800 6 la_oenb_mprj[49]
port 433 nsew signal input
rlabel metal2 s 80584 0 80696 800 6 la_oenb_mprj[4]
port 434 nsew signal input
rlabel metal2 s 108584 0 108696 800 6 la_oenb_mprj[50]
port 435 nsew signal input
rlabel metal2 s 109256 0 109368 800 6 la_oenb_mprj[51]
port 436 nsew signal input
rlabel metal2 s 109816 0 109928 800 6 la_oenb_mprj[52]
port 437 nsew signal input
rlabel metal2 s 110488 0 110600 800 6 la_oenb_mprj[53]
port 438 nsew signal input
rlabel metal2 s 111048 0 111160 800 6 la_oenb_mprj[54]
port 439 nsew signal input
rlabel metal2 s 111720 0 111832 800 6 la_oenb_mprj[55]
port 440 nsew signal input
rlabel metal2 s 112280 0 112392 800 6 la_oenb_mprj[56]
port 441 nsew signal input
rlabel metal2 s 112840 0 112952 800 6 la_oenb_mprj[57]
port 442 nsew signal input
rlabel metal2 s 113512 0 113624 800 6 la_oenb_mprj[58]
port 443 nsew signal input
rlabel metal2 s 114072 0 114184 800 6 la_oenb_mprj[59]
port 444 nsew signal input
rlabel metal2 s 81144 0 81256 800 6 la_oenb_mprj[5]
port 445 nsew signal input
rlabel metal2 s 114744 0 114856 800 6 la_oenb_mprj[60]
port 446 nsew signal input
rlabel metal2 s 115304 0 115416 800 6 la_oenb_mprj[61]
port 447 nsew signal input
rlabel metal2 s 115976 0 116088 800 6 la_oenb_mprj[62]
port 448 nsew signal input
rlabel metal2 s 116536 0 116648 800 6 la_oenb_mprj[63]
port 449 nsew signal input
rlabel metal2 s 81816 0 81928 800 6 la_oenb_mprj[6]
port 450 nsew signal input
rlabel metal2 s 82376 0 82488 800 6 la_oenb_mprj[7]
port 451 nsew signal input
rlabel metal2 s 83048 0 83160 800 6 la_oenb_mprj[8]
port 452 nsew signal input
rlabel metal2 s 83608 0 83720 800 6 la_oenb_mprj[9]
port 453 nsew signal input
rlabel metal2 s 219016 0 219128 800 6 mprj_ack_i_core
port 454 nsew signal output
rlabel metal2 s 1736 14200 1848 15000 6 mprj_ack_i_user
port 455 nsew signal input
rlabel metal2 s 178136 0 178248 800 6 mprj_adr_o_core[0]
port 456 nsew signal input
rlabel metal2 s 184184 0 184296 800 6 mprj_adr_o_core[10]
port 457 nsew signal input
rlabel metal2 s 184856 0 184968 800 6 mprj_adr_o_core[11]
port 458 nsew signal input
rlabel metal2 s 185416 0 185528 800 6 mprj_adr_o_core[12]
port 459 nsew signal input
rlabel metal2 s 186088 0 186200 800 6 mprj_adr_o_core[13]
port 460 nsew signal input
rlabel metal2 s 186648 0 186760 800 6 mprj_adr_o_core[14]
port 461 nsew signal input
rlabel metal2 s 187320 0 187432 800 6 mprj_adr_o_core[15]
port 462 nsew signal input
rlabel metal2 s 187880 0 187992 800 6 mprj_adr_o_core[16]
port 463 nsew signal input
rlabel metal2 s 188440 0 188552 800 6 mprj_adr_o_core[17]
port 464 nsew signal input
rlabel metal2 s 189112 0 189224 800 6 mprj_adr_o_core[18]
port 465 nsew signal input
rlabel metal2 s 189672 0 189784 800 6 mprj_adr_o_core[19]
port 466 nsew signal input
rlabel metal2 s 178696 0 178808 800 6 mprj_adr_o_core[1]
port 467 nsew signal input
rlabel metal2 s 190344 0 190456 800 6 mprj_adr_o_core[20]
port 468 nsew signal input
rlabel metal2 s 190904 0 191016 800 6 mprj_adr_o_core[21]
port 469 nsew signal input
rlabel metal2 s 191576 0 191688 800 6 mprj_adr_o_core[22]
port 470 nsew signal input
rlabel metal2 s 192136 0 192248 800 6 mprj_adr_o_core[23]
port 471 nsew signal input
rlabel metal2 s 192808 0 192920 800 6 mprj_adr_o_core[24]
port 472 nsew signal input
rlabel metal2 s 193368 0 193480 800 6 mprj_adr_o_core[25]
port 473 nsew signal input
rlabel metal2 s 193928 0 194040 800 6 mprj_adr_o_core[26]
port 474 nsew signal input
rlabel metal2 s 194600 0 194712 800 6 mprj_adr_o_core[27]
port 475 nsew signal input
rlabel metal2 s 195160 0 195272 800 6 mprj_adr_o_core[28]
port 476 nsew signal input
rlabel metal2 s 195832 0 195944 800 6 mprj_adr_o_core[29]
port 477 nsew signal input
rlabel metal2 s 179368 0 179480 800 6 mprj_adr_o_core[2]
port 478 nsew signal input
rlabel metal2 s 196392 0 196504 800 6 mprj_adr_o_core[30]
port 479 nsew signal input
rlabel metal2 s 197064 0 197176 800 6 mprj_adr_o_core[31]
port 480 nsew signal input
rlabel metal2 s 179928 0 180040 800 6 mprj_adr_o_core[3]
port 481 nsew signal input
rlabel metal2 s 180600 0 180712 800 6 mprj_adr_o_core[4]
port 482 nsew signal input
rlabel metal2 s 181160 0 181272 800 6 mprj_adr_o_core[5]
port 483 nsew signal input
rlabel metal2 s 181832 0 181944 800 6 mprj_adr_o_core[6]
port 484 nsew signal input
rlabel metal2 s 182392 0 182504 800 6 mprj_adr_o_core[7]
port 485 nsew signal input
rlabel metal2 s 182952 0 183064 800 6 mprj_adr_o_core[8]
port 486 nsew signal input
rlabel metal2 s 183624 0 183736 800 6 mprj_adr_o_core[9]
port 487 nsew signal input
rlabel metal2 s 4648 14200 4760 15000 6 mprj_adr_o_user[0]
port 488 nsew signal output
rlabel metal2 s 29400 14200 29512 15000 6 mprj_adr_o_user[10]
port 489 nsew signal output
rlabel metal2 s 31528 14200 31640 15000 6 mprj_adr_o_user[11]
port 490 nsew signal output
rlabel metal2 s 33768 14200 33880 15000 6 mprj_adr_o_user[12]
port 491 nsew signal output
rlabel metal2 s 35896 14200 36008 15000 6 mprj_adr_o_user[13]
port 492 nsew signal output
rlabel metal2 s 38136 14200 38248 15000 6 mprj_adr_o_user[14]
port 493 nsew signal output
rlabel metal2 s 40264 14200 40376 15000 6 mprj_adr_o_user[15]
port 494 nsew signal output
rlabel metal2 s 42504 14200 42616 15000 6 mprj_adr_o_user[16]
port 495 nsew signal output
rlabel metal2 s 44632 14200 44744 15000 6 mprj_adr_o_user[17]
port 496 nsew signal output
rlabel metal2 s 46872 14200 46984 15000 6 mprj_adr_o_user[18]
port 497 nsew signal output
rlabel metal2 s 49000 14200 49112 15000 6 mprj_adr_o_user[19]
port 498 nsew signal output
rlabel metal2 s 7560 14200 7672 15000 6 mprj_adr_o_user[1]
port 499 nsew signal output
rlabel metal2 s 51240 14200 51352 15000 6 mprj_adr_o_user[20]
port 500 nsew signal output
rlabel metal2 s 53368 14200 53480 15000 6 mprj_adr_o_user[21]
port 501 nsew signal output
rlabel metal2 s 55608 14200 55720 15000 6 mprj_adr_o_user[22]
port 502 nsew signal output
rlabel metal2 s 57848 14200 57960 15000 6 mprj_adr_o_user[23]
port 503 nsew signal output
rlabel metal2 s 59976 14200 60088 15000 6 mprj_adr_o_user[24]
port 504 nsew signal output
rlabel metal2 s 62216 14200 62328 15000 6 mprj_adr_o_user[25]
port 505 nsew signal output
rlabel metal2 s 64344 14200 64456 15000 6 mprj_adr_o_user[26]
port 506 nsew signal output
rlabel metal2 s 66584 14200 66696 15000 6 mprj_adr_o_user[27]
port 507 nsew signal output
rlabel metal2 s 68712 14200 68824 15000 6 mprj_adr_o_user[28]
port 508 nsew signal output
rlabel metal2 s 70952 14200 71064 15000 6 mprj_adr_o_user[29]
port 509 nsew signal output
rlabel metal2 s 10472 14200 10584 15000 6 mprj_adr_o_user[2]
port 510 nsew signal output
rlabel metal2 s 73080 14200 73192 15000 6 mprj_adr_o_user[30]
port 511 nsew signal output
rlabel metal2 s 75320 14200 75432 15000 6 mprj_adr_o_user[31]
port 512 nsew signal output
rlabel metal2 s 13384 14200 13496 15000 6 mprj_adr_o_user[3]
port 513 nsew signal output
rlabel metal2 s 16296 14200 16408 15000 6 mprj_adr_o_user[4]
port 514 nsew signal output
rlabel metal2 s 18424 14200 18536 15000 6 mprj_adr_o_user[5]
port 515 nsew signal output
rlabel metal2 s 20664 14200 20776 15000 6 mprj_adr_o_user[6]
port 516 nsew signal output
rlabel metal2 s 22792 14200 22904 15000 6 mprj_adr_o_user[7]
port 517 nsew signal output
rlabel metal2 s 25032 14200 25144 15000 6 mprj_adr_o_user[8]
port 518 nsew signal output
rlabel metal2 s 27160 14200 27272 15000 6 mprj_adr_o_user[9]
port 519 nsew signal output
rlabel metal2 s 217784 0 217896 800 6 mprj_cyc_o_core
port 520 nsew signal input
rlabel metal2 s 2408 14200 2520 15000 6 mprj_cyc_o_user
port 521 nsew signal output
rlabel metal2 s 156184 0 156296 800 6 mprj_dat_i_core[0]
port 522 nsew signal output
rlabel metal2 s 162232 0 162344 800 6 mprj_dat_i_core[10]
port 523 nsew signal output
rlabel metal2 s 162904 0 163016 800 6 mprj_dat_i_core[11]
port 524 nsew signal output
rlabel metal2 s 163464 0 163576 800 6 mprj_dat_i_core[12]
port 525 nsew signal output
rlabel metal2 s 164136 0 164248 800 6 mprj_dat_i_core[13]
port 526 nsew signal output
rlabel metal2 s 164696 0 164808 800 6 mprj_dat_i_core[14]
port 527 nsew signal output
rlabel metal2 s 165368 0 165480 800 6 mprj_dat_i_core[15]
port 528 nsew signal output
rlabel metal2 s 165928 0 166040 800 6 mprj_dat_i_core[16]
port 529 nsew signal output
rlabel metal2 s 166488 0 166600 800 6 mprj_dat_i_core[17]
port 530 nsew signal output
rlabel metal2 s 167160 0 167272 800 6 mprj_dat_i_core[18]
port 531 nsew signal output
rlabel metal2 s 167720 0 167832 800 6 mprj_dat_i_core[19]
port 532 nsew signal output
rlabel metal2 s 156744 0 156856 800 6 mprj_dat_i_core[1]
port 533 nsew signal output
rlabel metal2 s 168392 0 168504 800 6 mprj_dat_i_core[20]
port 534 nsew signal output
rlabel metal2 s 168952 0 169064 800 6 mprj_dat_i_core[21]
port 535 nsew signal output
rlabel metal2 s 169624 0 169736 800 6 mprj_dat_i_core[22]
port 536 nsew signal output
rlabel metal2 s 170184 0 170296 800 6 mprj_dat_i_core[23]
port 537 nsew signal output
rlabel metal2 s 170856 0 170968 800 6 mprj_dat_i_core[24]
port 538 nsew signal output
rlabel metal2 s 171416 0 171528 800 6 mprj_dat_i_core[25]
port 539 nsew signal output
rlabel metal2 s 171976 0 172088 800 6 mprj_dat_i_core[26]
port 540 nsew signal output
rlabel metal2 s 172648 0 172760 800 6 mprj_dat_i_core[27]
port 541 nsew signal output
rlabel metal2 s 173208 0 173320 800 6 mprj_dat_i_core[28]
port 542 nsew signal output
rlabel metal2 s 173880 0 173992 800 6 mprj_dat_i_core[29]
port 543 nsew signal output
rlabel metal2 s 157416 0 157528 800 6 mprj_dat_i_core[2]
port 544 nsew signal output
rlabel metal2 s 174440 0 174552 800 6 mprj_dat_i_core[30]
port 545 nsew signal output
rlabel metal2 s 175112 0 175224 800 6 mprj_dat_i_core[31]
port 546 nsew signal output
rlabel metal2 s 157976 0 158088 800 6 mprj_dat_i_core[3]
port 547 nsew signal output
rlabel metal2 s 158648 0 158760 800 6 mprj_dat_i_core[4]
port 548 nsew signal output
rlabel metal2 s 159208 0 159320 800 6 mprj_dat_i_core[5]
port 549 nsew signal output
rlabel metal2 s 159880 0 159992 800 6 mprj_dat_i_core[6]
port 550 nsew signal output
rlabel metal2 s 160440 0 160552 800 6 mprj_dat_i_core[7]
port 551 nsew signal output
rlabel metal2 s 161112 0 161224 800 6 mprj_dat_i_core[8]
port 552 nsew signal output
rlabel metal2 s 161672 0 161784 800 6 mprj_dat_i_core[9]
port 553 nsew signal output
rlabel metal2 s 5320 14200 5432 15000 6 mprj_dat_i_user[0]
port 554 nsew signal input
rlabel metal2 s 30072 14200 30184 15000 6 mprj_dat_i_user[10]
port 555 nsew signal input
rlabel metal2 s 32312 14200 32424 15000 6 mprj_dat_i_user[11]
port 556 nsew signal input
rlabel metal2 s 34440 14200 34552 15000 6 mprj_dat_i_user[12]
port 557 nsew signal input
rlabel metal2 s 36680 14200 36792 15000 6 mprj_dat_i_user[13]
port 558 nsew signal input
rlabel metal2 s 38808 14200 38920 15000 6 mprj_dat_i_user[14]
port 559 nsew signal input
rlabel metal2 s 41048 14200 41160 15000 6 mprj_dat_i_user[15]
port 560 nsew signal input
rlabel metal2 s 43176 14200 43288 15000 6 mprj_dat_i_user[16]
port 561 nsew signal input
rlabel metal2 s 45416 14200 45528 15000 6 mprj_dat_i_user[17]
port 562 nsew signal input
rlabel metal2 s 47544 14200 47656 15000 6 mprj_dat_i_user[18]
port 563 nsew signal input
rlabel metal2 s 49784 14200 49896 15000 6 mprj_dat_i_user[19]
port 564 nsew signal input
rlabel metal2 s 8232 14200 8344 15000 6 mprj_dat_i_user[1]
port 565 nsew signal input
rlabel metal2 s 51912 14200 52024 15000 6 mprj_dat_i_user[20]
port 566 nsew signal input
rlabel metal2 s 54152 14200 54264 15000 6 mprj_dat_i_user[21]
port 567 nsew signal input
rlabel metal2 s 56392 14200 56504 15000 6 mprj_dat_i_user[22]
port 568 nsew signal input
rlabel metal2 s 58520 14200 58632 15000 6 mprj_dat_i_user[23]
port 569 nsew signal input
rlabel metal2 s 60760 14200 60872 15000 6 mprj_dat_i_user[24]
port 570 nsew signal input
rlabel metal2 s 62888 14200 63000 15000 6 mprj_dat_i_user[25]
port 571 nsew signal input
rlabel metal2 s 65128 14200 65240 15000 6 mprj_dat_i_user[26]
port 572 nsew signal input
rlabel metal2 s 67256 14200 67368 15000 6 mprj_dat_i_user[27]
port 573 nsew signal input
rlabel metal2 s 69496 14200 69608 15000 6 mprj_dat_i_user[28]
port 574 nsew signal input
rlabel metal2 s 71624 14200 71736 15000 6 mprj_dat_i_user[29]
port 575 nsew signal input
rlabel metal2 s 11144 14200 11256 15000 6 mprj_dat_i_user[2]
port 576 nsew signal input
rlabel metal2 s 73864 14200 73976 15000 6 mprj_dat_i_user[30]
port 577 nsew signal input
rlabel metal2 s 75992 14200 76104 15000 6 mprj_dat_i_user[31]
port 578 nsew signal input
rlabel metal2 s 14056 14200 14168 15000 6 mprj_dat_i_user[3]
port 579 nsew signal input
rlabel metal2 s 16968 14200 17080 15000 6 mprj_dat_i_user[4]
port 580 nsew signal input
rlabel metal2 s 19208 14200 19320 15000 6 mprj_dat_i_user[5]
port 581 nsew signal input
rlabel metal2 s 21336 14200 21448 15000 6 mprj_dat_i_user[6]
port 582 nsew signal input
rlabel metal2 s 23576 14200 23688 15000 6 mprj_dat_i_user[7]
port 583 nsew signal input
rlabel metal2 s 25704 14200 25816 15000 6 mprj_dat_i_user[8]
port 584 nsew signal input
rlabel metal2 s 27944 14200 28056 15000 6 mprj_dat_i_user[9]
port 585 nsew signal input
rlabel metal2 s 197624 0 197736 800 6 mprj_dat_o_core[0]
port 586 nsew signal input
rlabel metal2 s 203784 0 203896 800 6 mprj_dat_o_core[10]
port 587 nsew signal input
rlabel metal2 s 204344 0 204456 800 6 mprj_dat_o_core[11]
port 588 nsew signal input
rlabel metal2 s 204904 0 205016 800 6 mprj_dat_o_core[12]
port 589 nsew signal input
rlabel metal2 s 205576 0 205688 800 6 mprj_dat_o_core[13]
port 590 nsew signal input
rlabel metal2 s 206136 0 206248 800 6 mprj_dat_o_core[14]
port 591 nsew signal input
rlabel metal2 s 206808 0 206920 800 6 mprj_dat_o_core[15]
port 592 nsew signal input
rlabel metal2 s 207368 0 207480 800 6 mprj_dat_o_core[16]
port 593 nsew signal input
rlabel metal2 s 208040 0 208152 800 6 mprj_dat_o_core[17]
port 594 nsew signal input
rlabel metal2 s 208600 0 208712 800 6 mprj_dat_o_core[18]
port 595 nsew signal input
rlabel metal2 s 209272 0 209384 800 6 mprj_dat_o_core[19]
port 596 nsew signal input
rlabel metal2 s 198296 0 198408 800 6 mprj_dat_o_core[1]
port 597 nsew signal input
rlabel metal2 s 209832 0 209944 800 6 mprj_dat_o_core[20]
port 598 nsew signal input
rlabel metal2 s 210392 0 210504 800 6 mprj_dat_o_core[21]
port 599 nsew signal input
rlabel metal2 s 211064 0 211176 800 6 mprj_dat_o_core[22]
port 600 nsew signal input
rlabel metal2 s 211624 0 211736 800 6 mprj_dat_o_core[23]
port 601 nsew signal input
rlabel metal2 s 212296 0 212408 800 6 mprj_dat_o_core[24]
port 602 nsew signal input
rlabel metal2 s 212856 0 212968 800 6 mprj_dat_o_core[25]
port 603 nsew signal input
rlabel metal2 s 213528 0 213640 800 6 mprj_dat_o_core[26]
port 604 nsew signal input
rlabel metal2 s 214088 0 214200 800 6 mprj_dat_o_core[27]
port 605 nsew signal input
rlabel metal2 s 214760 0 214872 800 6 mprj_dat_o_core[28]
port 606 nsew signal input
rlabel metal2 s 215320 0 215432 800 6 mprj_dat_o_core[29]
port 607 nsew signal input
rlabel metal2 s 198856 0 198968 800 6 mprj_dat_o_core[2]
port 608 nsew signal input
rlabel metal2 s 215880 0 215992 800 6 mprj_dat_o_core[30]
port 609 nsew signal input
rlabel metal2 s 216552 0 216664 800 6 mprj_dat_o_core[31]
port 610 nsew signal input
rlabel metal2 s 199416 0 199528 800 6 mprj_dat_o_core[3]
port 611 nsew signal input
rlabel metal2 s 200088 0 200200 800 6 mprj_dat_o_core[4]
port 612 nsew signal input
rlabel metal2 s 200648 0 200760 800 6 mprj_dat_o_core[5]
port 613 nsew signal input
rlabel metal2 s 201320 0 201432 800 6 mprj_dat_o_core[6]
port 614 nsew signal input
rlabel metal2 s 201880 0 201992 800 6 mprj_dat_o_core[7]
port 615 nsew signal input
rlabel metal2 s 202552 0 202664 800 6 mprj_dat_o_core[8]
port 616 nsew signal input
rlabel metal2 s 203112 0 203224 800 6 mprj_dat_o_core[9]
port 617 nsew signal input
rlabel metal2 s 6104 14200 6216 15000 6 mprj_dat_o_user[0]
port 618 nsew signal output
rlabel metal2 s 30856 14200 30968 15000 6 mprj_dat_o_user[10]
port 619 nsew signal output
rlabel metal2 s 32984 14200 33096 15000 6 mprj_dat_o_user[11]
port 620 nsew signal output
rlabel metal2 s 35224 14200 35336 15000 6 mprj_dat_o_user[12]
port 621 nsew signal output
rlabel metal2 s 37352 14200 37464 15000 6 mprj_dat_o_user[13]
port 622 nsew signal output
rlabel metal2 s 39592 14200 39704 15000 6 mprj_dat_o_user[14]
port 623 nsew signal output
rlabel metal2 s 41720 14200 41832 15000 6 mprj_dat_o_user[15]
port 624 nsew signal output
rlabel metal2 s 43960 14200 44072 15000 6 mprj_dat_o_user[16]
port 625 nsew signal output
rlabel metal2 s 46088 14200 46200 15000 6 mprj_dat_o_user[17]
port 626 nsew signal output
rlabel metal2 s 48328 14200 48440 15000 6 mprj_dat_o_user[18]
port 627 nsew signal output
rlabel metal2 s 50456 14200 50568 15000 6 mprj_dat_o_user[19]
port 628 nsew signal output
rlabel metal2 s 9016 14200 9128 15000 6 mprj_dat_o_user[1]
port 629 nsew signal output
rlabel metal2 s 52696 14200 52808 15000 6 mprj_dat_o_user[20]
port 630 nsew signal output
rlabel metal2 s 54824 14200 54936 15000 6 mprj_dat_o_user[21]
port 631 nsew signal output
rlabel metal2 s 57064 14200 57176 15000 6 mprj_dat_o_user[22]
port 632 nsew signal output
rlabel metal2 s 59304 14200 59416 15000 6 mprj_dat_o_user[23]
port 633 nsew signal output
rlabel metal2 s 61432 14200 61544 15000 6 mprj_dat_o_user[24]
port 634 nsew signal output
rlabel metal2 s 63672 14200 63784 15000 6 mprj_dat_o_user[25]
port 635 nsew signal output
rlabel metal2 s 65800 14200 65912 15000 6 mprj_dat_o_user[26]
port 636 nsew signal output
rlabel metal2 s 68040 14200 68152 15000 6 mprj_dat_o_user[27]
port 637 nsew signal output
rlabel metal2 s 70168 14200 70280 15000 6 mprj_dat_o_user[28]
port 638 nsew signal output
rlabel metal2 s 72408 14200 72520 15000 6 mprj_dat_o_user[29]
port 639 nsew signal output
rlabel metal2 s 11928 14200 12040 15000 6 mprj_dat_o_user[2]
port 640 nsew signal output
rlabel metal2 s 74536 14200 74648 15000 6 mprj_dat_o_user[30]
port 641 nsew signal output
rlabel metal2 s 76776 14200 76888 15000 6 mprj_dat_o_user[31]
port 642 nsew signal output
rlabel metal2 s 14840 14200 14952 15000 6 mprj_dat_o_user[3]
port 643 nsew signal output
rlabel metal2 s 17752 14200 17864 15000 6 mprj_dat_o_user[4]
port 644 nsew signal output
rlabel metal2 s 19880 14200 19992 15000 6 mprj_dat_o_user[5]
port 645 nsew signal output
rlabel metal2 s 22120 14200 22232 15000 6 mprj_dat_o_user[6]
port 646 nsew signal output
rlabel metal2 s 24248 14200 24360 15000 6 mprj_dat_o_user[7]
port 647 nsew signal output
rlabel metal2 s 26488 14200 26600 15000 6 mprj_dat_o_user[8]
port 648 nsew signal output
rlabel metal2 s 28616 14200 28728 15000 6 mprj_dat_o_user[9]
port 649 nsew signal output
rlabel metal2 s 219576 0 219688 800 6 mprj_iena_wb
port 650 nsew signal input
rlabel metal2 s 175672 0 175784 800 6 mprj_sel_o_core[0]
port 651 nsew signal input
rlabel metal2 s 176344 0 176456 800 6 mprj_sel_o_core[1]
port 652 nsew signal input
rlabel metal2 s 176904 0 177016 800 6 mprj_sel_o_core[2]
port 653 nsew signal input
rlabel metal2 s 177464 0 177576 800 6 mprj_sel_o_core[3]
port 654 nsew signal input
rlabel metal2 s 6776 14200 6888 15000 6 mprj_sel_o_user[0]
port 655 nsew signal output
rlabel metal2 s 9688 14200 9800 15000 6 mprj_sel_o_user[1]
port 656 nsew signal output
rlabel metal2 s 12600 14200 12712 15000 6 mprj_sel_o_user[2]
port 657 nsew signal output
rlabel metal2 s 15512 14200 15624 15000 6 mprj_sel_o_user[3]
port 658 nsew signal output
rlabel metal2 s 218344 0 218456 800 6 mprj_stb_o_core
port 659 nsew signal input
rlabel metal2 s 3192 14200 3304 15000 6 mprj_stb_o_user
port 660 nsew signal output
rlabel metal2 s 217112 0 217224 800 6 mprj_we_o_core
port 661 nsew signal input
rlabel metal2 s 3864 14200 3976 15000 6 mprj_we_o_user
port 662 nsew signal output
rlabel metal2 s 280 14200 392 15000 6 user_clock
port 663 nsew signal output
rlabel metal2 s 217336 14200 217448 15000 6 user_clock2
port 664 nsew signal output
rlabel metal3 s 219200 8680 220000 8792 6 user_irq[0]
port 665 nsew signal output
rlabel metal3 s 219200 11144 220000 11256 6 user_irq[1]
port 666 nsew signal output
rlabel metal3 s 219200 13608 220000 13720 6 user_irq[2]
port 667 nsew signal output
rlabel metal2 s 218120 14200 218232 15000 6 user_irq_core[0]
port 668 nsew signal input
rlabel metal2 s 218792 14200 218904 15000 6 user_irq_core[1]
port 669 nsew signal input
rlabel metal2 s 219576 14200 219688 15000 6 user_irq_core[2]
port 670 nsew signal input
rlabel metal3 s 219200 1288 220000 1400 6 user_irq_ena[0]
port 671 nsew signal input
rlabel metal3 s 219200 3752 220000 3864 6 user_irq_ena[1]
port 672 nsew signal input
rlabel metal3 s 219200 6216 220000 6328 6 user_irq_ena[2]
port 673 nsew signal input
rlabel metal2 s 952 14200 1064 15000 6 user_reset
port 674 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 220000 15000
string GDS_END 2482568
string GDS_FILE ../gds/mgmt_protect.gds.gz
string GDS_START 68820
string LEFclass BLOCK
string LEFview TRUE
<< end >>
