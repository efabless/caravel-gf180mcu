VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO housekeeping
  CLASS BLOCK ;
  FOREIGN housekeeping ;
  ORIGIN 0.000 0.000 ;
  SIZE 620.000 BY 780.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT -0.880 8.080 0.720 768.080 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.880 8.080 620.800 9.680 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -0.880 766.480 620.800 768.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 619.200 8.080 620.800 768.080 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 22.240 4.780 23.840 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 99.040 4.780 100.640 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 4.780 177.440 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 4.780 254.240 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 4.780 331.040 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 4.780 407.840 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 4.780 484.640 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 4.780 561.440 771.380 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 21.290 624.100 22.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 81.290 624.100 82.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 141.290 624.100 142.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 201.290 624.100 202.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 261.290 624.100 262.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 321.290 624.100 322.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 381.290 624.100 382.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 441.290 624.100 442.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 501.290 624.100 502.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 561.290 624.100 562.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 621.290 624.100 622.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 681.290 624.100 682.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 741.290 624.100 742.890 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT -4.180 4.780 -2.580 771.380 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 4.780 624.100 6.380 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 769.780 624.100 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 622.500 4.780 624.100 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 25.540 4.780 27.140 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 102.340 4.780 103.940 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 179.140 4.780 180.740 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 255.940 4.780 257.540 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 332.740 4.780 334.340 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 409.540 4.780 411.140 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 486.340 4.780 487.940 771.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 563.140 4.780 564.740 771.380 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 51.290 624.100 52.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 111.290 624.100 112.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 171.290 624.100 172.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 231.290 624.100 232.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 291.290 624.100 292.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 351.290 624.100 352.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 411.290 624.100 412.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 471.290 624.100 472.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 531.290 624.100 532.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 591.290 624.100 592.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 651.290 624.100 652.890 ;
    END
    PORT
      LAYER Metal5 ;
        RECT -4.180 711.290 624.100 712.890 ;
    END
  END VSS
  PIN debug_in
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 22.960 4.000 23.520 ;
    END
  END debug_in
  PIN debug_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 29.120 4.000 29.680 ;
    END
  END debug_mode
  PIN debug_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 35.280 4.000 35.840 ;
    END
  END debug_oeb
  PIN debug_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 41.440 4.000 42.000 ;
    END
  END debug_out
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.760 4.000 54.320 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.920 4.000 60.480 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 66.080 4.000 66.640 ;
    END
  END irq[2]
  PIN mask_rev_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 393.680 0.000 394.240 4.000 ;
    END
  END mask_rev_in[0]
  PIN mask_rev_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 460.880 0.000 461.440 4.000 ;
    END
  END mask_rev_in[10]
  PIN mask_rev_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 467.600 0.000 468.160 4.000 ;
    END
  END mask_rev_in[11]
  PIN mask_rev_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 474.320 0.000 474.880 4.000 ;
    END
  END mask_rev_in[12]
  PIN mask_rev_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 481.040 0.000 481.600 4.000 ;
    END
  END mask_rev_in[13]
  PIN mask_rev_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 487.760 0.000 488.320 4.000 ;
    END
  END mask_rev_in[14]
  PIN mask_rev_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 494.480 0.000 495.040 4.000 ;
    END
  END mask_rev_in[15]
  PIN mask_rev_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 501.200 0.000 501.760 4.000 ;
    END
  END mask_rev_in[16]
  PIN mask_rev_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 507.920 0.000 508.480 4.000 ;
    END
  END mask_rev_in[17]
  PIN mask_rev_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 514.640 0.000 515.200 4.000 ;
    END
  END mask_rev_in[18]
  PIN mask_rev_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 521.360 0.000 521.920 4.000 ;
    END
  END mask_rev_in[19]
  PIN mask_rev_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 400.400 0.000 400.960 4.000 ;
    END
  END mask_rev_in[1]
  PIN mask_rev_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 528.080 0.000 528.640 4.000 ;
    END
  END mask_rev_in[20]
  PIN mask_rev_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 534.800 0.000 535.360 4.000 ;
    END
  END mask_rev_in[21]
  PIN mask_rev_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 541.520 0.000 542.080 4.000 ;
    END
  END mask_rev_in[22]
  PIN mask_rev_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 548.240 0.000 548.800 4.000 ;
    END
  END mask_rev_in[23]
  PIN mask_rev_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 554.960 0.000 555.520 4.000 ;
    END
  END mask_rev_in[24]
  PIN mask_rev_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 561.680 0.000 562.240 4.000 ;
    END
  END mask_rev_in[25]
  PIN mask_rev_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 568.400 0.000 568.960 4.000 ;
    END
  END mask_rev_in[26]
  PIN mask_rev_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 575.120 0.000 575.680 4.000 ;
    END
  END mask_rev_in[27]
  PIN mask_rev_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 581.840 0.000 582.400 4.000 ;
    END
  END mask_rev_in[28]
  PIN mask_rev_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 588.560 0.000 589.120 4.000 ;
    END
  END mask_rev_in[29]
  PIN mask_rev_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 407.120 0.000 407.680 4.000 ;
    END
  END mask_rev_in[2]
  PIN mask_rev_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 595.280 0.000 595.840 4.000 ;
    END
  END mask_rev_in[30]
  PIN mask_rev_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 602.000 0.000 602.560 4.000 ;
    END
  END mask_rev_in[31]
  PIN mask_rev_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.840 0.000 414.400 4.000 ;
    END
  END mask_rev_in[3]
  PIN mask_rev_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 420.560 0.000 421.120 4.000 ;
    END
  END mask_rev_in[4]
  PIN mask_rev_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 427.280 0.000 427.840 4.000 ;
    END
  END mask_rev_in[5]
  PIN mask_rev_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 434.000 0.000 434.560 4.000 ;
    END
  END mask_rev_in[6]
  PIN mask_rev_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 440.720 0.000 441.280 4.000 ;
    END
  END mask_rev_in[7]
  PIN mask_rev_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 447.440 0.000 448.000 4.000 ;
    END
  END mask_rev_in[8]
  PIN mask_rev_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 454.160 0.000 454.720 4.000 ;
    END
  END mask_rev_in[9]
  PIN mgmt_gpio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 72.240 620.000 72.800 ;
    END
  END mgmt_gpio_in[0]
  PIN mgmt_gpio_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 425.040 620.000 425.600 ;
    END
  END mgmt_gpio_in[10]
  PIN mgmt_gpio_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 460.320 620.000 460.880 ;
    END
  END mgmt_gpio_in[11]
  PIN mgmt_gpio_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 495.600 620.000 496.160 ;
    END
  END mgmt_gpio_in[12]
  PIN mgmt_gpio_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 530.880 620.000 531.440 ;
    END
  END mgmt_gpio_in[13]
  PIN mgmt_gpio_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 566.160 620.000 566.720 ;
    END
  END mgmt_gpio_in[14]
  PIN mgmt_gpio_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 601.440 620.000 602.000 ;
    END
  END mgmt_gpio_in[15]
  PIN mgmt_gpio_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 636.720 620.000 637.280 ;
    END
  END mgmt_gpio_in[16]
  PIN mgmt_gpio_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 672.000 620.000 672.560 ;
    END
  END mgmt_gpio_in[17]
  PIN mgmt_gpio_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 707.280 620.000 707.840 ;
    END
  END mgmt_gpio_in[18]
  PIN mgmt_gpio_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 742.560 620.000 743.120 ;
    END
  END mgmt_gpio_in[19]
  PIN mgmt_gpio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 107.520 620.000 108.080 ;
    END
  END mgmt_gpio_in[1]
  PIN mgmt_gpio_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 429.520 4.000 430.080 ;
    END
  END mgmt_gpio_in[20]
  PIN mgmt_gpio_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 448.000 4.000 448.560 ;
    END
  END mgmt_gpio_in[21]
  PIN mgmt_gpio_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 466.480 4.000 467.040 ;
    END
  END mgmt_gpio_in[22]
  PIN mgmt_gpio_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 484.960 4.000 485.520 ;
    END
  END mgmt_gpio_in[23]
  PIN mgmt_gpio_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 503.440 4.000 504.000 ;
    END
  END mgmt_gpio_in[24]
  PIN mgmt_gpio_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 521.920 4.000 522.480 ;
    END
  END mgmt_gpio_in[25]
  PIN mgmt_gpio_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 540.400 4.000 540.960 ;
    END
  END mgmt_gpio_in[26]
  PIN mgmt_gpio_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 558.880 4.000 559.440 ;
    END
  END mgmt_gpio_in[27]
  PIN mgmt_gpio_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 577.360 4.000 577.920 ;
    END
  END mgmt_gpio_in[28]
  PIN mgmt_gpio_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 595.840 4.000 596.400 ;
    END
  END mgmt_gpio_in[29]
  PIN mgmt_gpio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 142.800 620.000 143.360 ;
    END
  END mgmt_gpio_in[2]
  PIN mgmt_gpio_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 614.320 4.000 614.880 ;
    END
  END mgmt_gpio_in[30]
  PIN mgmt_gpio_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 632.800 4.000 633.360 ;
    END
  END mgmt_gpio_in[31]
  PIN mgmt_gpio_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 651.280 4.000 651.840 ;
    END
  END mgmt_gpio_in[32]
  PIN mgmt_gpio_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 669.760 4.000 670.320 ;
    END
  END mgmt_gpio_in[33]
  PIN mgmt_gpio_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 688.240 4.000 688.800 ;
    END
  END mgmt_gpio_in[34]
  PIN mgmt_gpio_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 706.720 4.000 707.280 ;
    END
  END mgmt_gpio_in[35]
  PIN mgmt_gpio_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 725.200 4.000 725.760 ;
    END
  END mgmt_gpio_in[36]
  PIN mgmt_gpio_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 743.680 4.000 744.240 ;
    END
  END mgmt_gpio_in[37]
  PIN mgmt_gpio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 178.080 620.000 178.640 ;
    END
  END mgmt_gpio_in[3]
  PIN mgmt_gpio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 213.360 620.000 213.920 ;
    END
  END mgmt_gpio_in[4]
  PIN mgmt_gpio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 248.640 620.000 249.200 ;
    END
  END mgmt_gpio_in[5]
  PIN mgmt_gpio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 283.920 620.000 284.480 ;
    END
  END mgmt_gpio_in[6]
  PIN mgmt_gpio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 319.200 620.000 319.760 ;
    END
  END mgmt_gpio_in[7]
  PIN mgmt_gpio_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 354.480 620.000 355.040 ;
    END
  END mgmt_gpio_in[8]
  PIN mgmt_gpio_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 389.760 620.000 390.320 ;
    END
  END mgmt_gpio_in[9]
  PIN mgmt_gpio_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 84.000 620.000 84.560 ;
    END
  END mgmt_gpio_oeb[0]
  PIN mgmt_gpio_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 436.800 620.000 437.360 ;
    END
  END mgmt_gpio_oeb[10]
  PIN mgmt_gpio_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 472.080 620.000 472.640 ;
    END
  END mgmt_gpio_oeb[11]
  PIN mgmt_gpio_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 507.360 620.000 507.920 ;
    END
  END mgmt_gpio_oeb[12]
  PIN mgmt_gpio_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 542.640 620.000 543.200 ;
    END
  END mgmt_gpio_oeb[13]
  PIN mgmt_gpio_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 577.920 620.000 578.480 ;
    END
  END mgmt_gpio_oeb[14]
  PIN mgmt_gpio_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 613.200 620.000 613.760 ;
    END
  END mgmt_gpio_oeb[15]
  PIN mgmt_gpio_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 648.480 620.000 649.040 ;
    END
  END mgmt_gpio_oeb[16]
  PIN mgmt_gpio_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 683.760 620.000 684.320 ;
    END
  END mgmt_gpio_oeb[17]
  PIN mgmt_gpio_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 719.040 620.000 719.600 ;
    END
  END mgmt_gpio_oeb[18]
  PIN mgmt_gpio_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 754.320 620.000 754.880 ;
    END
  END mgmt_gpio_oeb[19]
  PIN mgmt_gpio_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 119.280 620.000 119.840 ;
    END
  END mgmt_gpio_oeb[1]
  PIN mgmt_gpio_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 435.680 4.000 436.240 ;
    END
  END mgmt_gpio_oeb[20]
  PIN mgmt_gpio_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 454.160 4.000 454.720 ;
    END
  END mgmt_gpio_oeb[21]
  PIN mgmt_gpio_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 472.640 4.000 473.200 ;
    END
  END mgmt_gpio_oeb[22]
  PIN mgmt_gpio_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 491.120 4.000 491.680 ;
    END
  END mgmt_gpio_oeb[23]
  PIN mgmt_gpio_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 509.600 4.000 510.160 ;
    END
  END mgmt_gpio_oeb[24]
  PIN mgmt_gpio_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 528.080 4.000 528.640 ;
    END
  END mgmt_gpio_oeb[25]
  PIN mgmt_gpio_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 546.560 4.000 547.120 ;
    END
  END mgmt_gpio_oeb[26]
  PIN mgmt_gpio_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 565.040 4.000 565.600 ;
    END
  END mgmt_gpio_oeb[27]
  PIN mgmt_gpio_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 583.520 4.000 584.080 ;
    END
  END mgmt_gpio_oeb[28]
  PIN mgmt_gpio_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 602.000 4.000 602.560 ;
    END
  END mgmt_gpio_oeb[29]
  PIN mgmt_gpio_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 154.560 620.000 155.120 ;
    END
  END mgmt_gpio_oeb[2]
  PIN mgmt_gpio_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 620.480 4.000 621.040 ;
    END
  END mgmt_gpio_oeb[30]
  PIN mgmt_gpio_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 638.960 4.000 639.520 ;
    END
  END mgmt_gpio_oeb[31]
  PIN mgmt_gpio_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 657.440 4.000 658.000 ;
    END
  END mgmt_gpio_oeb[32]
  PIN mgmt_gpio_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 675.920 4.000 676.480 ;
    END
  END mgmt_gpio_oeb[33]
  PIN mgmt_gpio_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 694.400 4.000 694.960 ;
    END
  END mgmt_gpio_oeb[34]
  PIN mgmt_gpio_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 712.880 4.000 713.440 ;
    END
  END mgmt_gpio_oeb[35]
  PIN mgmt_gpio_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 731.360 4.000 731.920 ;
    END
  END mgmt_gpio_oeb[36]
  PIN mgmt_gpio_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 749.840 4.000 750.400 ;
    END
  END mgmt_gpio_oeb[37]
  PIN mgmt_gpio_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 189.840 620.000 190.400 ;
    END
  END mgmt_gpio_oeb[3]
  PIN mgmt_gpio_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 225.120 620.000 225.680 ;
    END
  END mgmt_gpio_oeb[4]
  PIN mgmt_gpio_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 260.400 620.000 260.960 ;
    END
  END mgmt_gpio_oeb[5]
  PIN mgmt_gpio_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 295.680 620.000 296.240 ;
    END
  END mgmt_gpio_oeb[6]
  PIN mgmt_gpio_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 330.960 620.000 331.520 ;
    END
  END mgmt_gpio_oeb[7]
  PIN mgmt_gpio_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 366.240 620.000 366.800 ;
    END
  END mgmt_gpio_oeb[8]
  PIN mgmt_gpio_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 401.520 620.000 402.080 ;
    END
  END mgmt_gpio_oeb[9]
  PIN mgmt_gpio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 95.760 620.000 96.320 ;
    END
  END mgmt_gpio_out[0]
  PIN mgmt_gpio_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 448.560 620.000 449.120 ;
    END
  END mgmt_gpio_out[10]
  PIN mgmt_gpio_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 483.840 620.000 484.400 ;
    END
  END mgmt_gpio_out[11]
  PIN mgmt_gpio_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 519.120 620.000 519.680 ;
    END
  END mgmt_gpio_out[12]
  PIN mgmt_gpio_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 554.400 620.000 554.960 ;
    END
  END mgmt_gpio_out[13]
  PIN mgmt_gpio_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 589.680 620.000 590.240 ;
    END
  END mgmt_gpio_out[14]
  PIN mgmt_gpio_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 624.960 620.000 625.520 ;
    END
  END mgmt_gpio_out[15]
  PIN mgmt_gpio_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 660.240 620.000 660.800 ;
    END
  END mgmt_gpio_out[16]
  PIN mgmt_gpio_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 695.520 620.000 696.080 ;
    END
  END mgmt_gpio_out[17]
  PIN mgmt_gpio_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 730.800 620.000 731.360 ;
    END
  END mgmt_gpio_out[18]
  PIN mgmt_gpio_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 766.080 620.000 766.640 ;
    END
  END mgmt_gpio_out[19]
  PIN mgmt_gpio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 131.040 620.000 131.600 ;
    END
  END mgmt_gpio_out[1]
  PIN mgmt_gpio_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 441.840 4.000 442.400 ;
    END
  END mgmt_gpio_out[20]
  PIN mgmt_gpio_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 460.320 4.000 460.880 ;
    END
  END mgmt_gpio_out[21]
  PIN mgmt_gpio_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 478.800 4.000 479.360 ;
    END
  END mgmt_gpio_out[22]
  PIN mgmt_gpio_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 497.280 4.000 497.840 ;
    END
  END mgmt_gpio_out[23]
  PIN mgmt_gpio_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 515.760 4.000 516.320 ;
    END
  END mgmt_gpio_out[24]
  PIN mgmt_gpio_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 534.240 4.000 534.800 ;
    END
  END mgmt_gpio_out[25]
  PIN mgmt_gpio_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 552.720 4.000 553.280 ;
    END
  END mgmt_gpio_out[26]
  PIN mgmt_gpio_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 571.200 4.000 571.760 ;
    END
  END mgmt_gpio_out[27]
  PIN mgmt_gpio_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 589.680 4.000 590.240 ;
    END
  END mgmt_gpio_out[28]
  PIN mgmt_gpio_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 608.160 4.000 608.720 ;
    END
  END mgmt_gpio_out[29]
  PIN mgmt_gpio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 166.320 620.000 166.880 ;
    END
  END mgmt_gpio_out[2]
  PIN mgmt_gpio_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 626.640 4.000 627.200 ;
    END
  END mgmt_gpio_out[30]
  PIN mgmt_gpio_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 645.120 4.000 645.680 ;
    END
  END mgmt_gpio_out[31]
  PIN mgmt_gpio_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 663.600 4.000 664.160 ;
    END
  END mgmt_gpio_out[32]
  PIN mgmt_gpio_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 682.080 4.000 682.640 ;
    END
  END mgmt_gpio_out[33]
  PIN mgmt_gpio_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 700.560 4.000 701.120 ;
    END
  END mgmt_gpio_out[34]
  PIN mgmt_gpio_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 719.040 4.000 719.600 ;
    END
  END mgmt_gpio_out[35]
  PIN mgmt_gpio_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 737.520 4.000 738.080 ;
    END
  END mgmt_gpio_out[36]
  PIN mgmt_gpio_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 756.000 4.000 756.560 ;
    END
  END mgmt_gpio_out[37]
  PIN mgmt_gpio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 201.600 620.000 202.160 ;
    END
  END mgmt_gpio_out[3]
  PIN mgmt_gpio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 236.880 620.000 237.440 ;
    END
  END mgmt_gpio_out[4]
  PIN mgmt_gpio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 272.160 620.000 272.720 ;
    END
  END mgmt_gpio_out[5]
  PIN mgmt_gpio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 307.440 620.000 308.000 ;
    END
  END mgmt_gpio_out[6]
  PIN mgmt_gpio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 342.720 620.000 343.280 ;
    END
  END mgmt_gpio_out[7]
  PIN mgmt_gpio_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 378.000 620.000 378.560 ;
    END
  END mgmt_gpio_out[8]
  PIN mgmt_gpio_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 413.280 620.000 413.840 ;
    END
  END mgmt_gpio_out[9]
  PIN pad_flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 17.360 0.000 17.920 4.000 ;
    END
  END pad_flash_clk
  PIN pad_flash_clk_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 24.080 0.000 24.640 4.000 ;
    END
  END pad_flash_clk_oe
  PIN pad_flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.800 0.000 31.360 4.000 ;
    END
  END pad_flash_csb
  PIN pad_flash_csb_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 37.520 0.000 38.080 4.000 ;
    END
  END pad_flash_csb_oe
  PIN pad_flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 44.240 0.000 44.800 4.000 ;
    END
  END pad_flash_io0_di
  PIN pad_flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.960 0.000 51.520 4.000 ;
    END
  END pad_flash_io0_do
  PIN pad_flash_io0_ie
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.680 0.000 58.240 4.000 ;
    END
  END pad_flash_io0_ie
  PIN pad_flash_io0_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 64.400 0.000 64.960 4.000 ;
    END
  END pad_flash_io0_oe
  PIN pad_flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 71.120 0.000 71.680 4.000 ;
    END
  END pad_flash_io1_di
  PIN pad_flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.840 0.000 78.400 4.000 ;
    END
  END pad_flash_io1_do
  PIN pad_flash_io1_ie
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.560 0.000 85.120 4.000 ;
    END
  END pad_flash_io1_ie
  PIN pad_flash_io1_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 91.280 0.000 91.840 4.000 ;
    END
  END pad_flash_io1_oe
  PIN pll90_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.640 0.000 179.200 4.000 ;
    END
  END pll90_sel[0]
  PIN pll90_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 185.360 0.000 185.920 4.000 ;
    END
  END pll90_sel[1]
  PIN pll90_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 192.080 0.000 192.640 4.000 ;
    END
  END pll90_sel[2]
  PIN pll_bypass
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 373.520 0.000 374.080 4.000 ;
    END
  END pll_bypass
  PIN pll_dco_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 118.160 0.000 118.720 4.000 ;
    END
  END pll_dco_ena
  PIN pll_div[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.880 0.000 125.440 4.000 ;
    END
  END pll_div[0]
  PIN pll_div[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.600 0.000 132.160 4.000 ;
    END
  END pll_div[1]
  PIN pll_div[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 138.320 0.000 138.880 4.000 ;
    END
  END pll_div[2]
  PIN pll_div[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 145.040 0.000 145.600 4.000 ;
    END
  END pll_div[3]
  PIN pll_div[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.760 0.000 152.320 4.000 ;
    END
  END pll_div[4]
  PIN pll_ena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 111.440 0.000 112.000 4.000 ;
    END
  END pll_ena
  PIN pll_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 158.480 0.000 159.040 4.000 ;
    END
  END pll_sel[0]
  PIN pll_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 165.200 0.000 165.760 4.000 ;
    END
  END pll_sel[1]
  PIN pll_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.920 0.000 172.480 4.000 ;
    END
  END pll_sel[2]
  PIN pll_trim[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 198.800 0.000 199.360 4.000 ;
    END
  END pll_trim[0]
  PIN pll_trim[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 266.000 0.000 266.560 4.000 ;
    END
  END pll_trim[10]
  PIN pll_trim[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.720 0.000 273.280 4.000 ;
    END
  END pll_trim[11]
  PIN pll_trim[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 279.440 0.000 280.000 4.000 ;
    END
  END pll_trim[12]
  PIN pll_trim[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 286.160 0.000 286.720 4.000 ;
    END
  END pll_trim[13]
  PIN pll_trim[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.880 0.000 293.440 4.000 ;
    END
  END pll_trim[14]
  PIN pll_trim[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.600 0.000 300.160 4.000 ;
    END
  END pll_trim[15]
  PIN pll_trim[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 306.320 0.000 306.880 4.000 ;
    END
  END pll_trim[16]
  PIN pll_trim[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 313.040 0.000 313.600 4.000 ;
    END
  END pll_trim[17]
  PIN pll_trim[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 319.760 0.000 320.320 4.000 ;
    END
  END pll_trim[18]
  PIN pll_trim[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 326.480 0.000 327.040 4.000 ;
    END
  END pll_trim[19]
  PIN pll_trim[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 205.520 0.000 206.080 4.000 ;
    END
  END pll_trim[1]
  PIN pll_trim[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 333.200 0.000 333.760 4.000 ;
    END
  END pll_trim[20]
  PIN pll_trim[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 339.920 0.000 340.480 4.000 ;
    END
  END pll_trim[21]
  PIN pll_trim[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 346.640 0.000 347.200 4.000 ;
    END
  END pll_trim[22]
  PIN pll_trim[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 353.360 0.000 353.920 4.000 ;
    END
  END pll_trim[23]
  PIN pll_trim[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 360.080 0.000 360.640 4.000 ;
    END
  END pll_trim[24]
  PIN pll_trim[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.800 0.000 367.360 4.000 ;
    END
  END pll_trim[25]
  PIN pll_trim[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 212.240 0.000 212.800 4.000 ;
    END
  END pll_trim[2]
  PIN pll_trim[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.960 0.000 219.520 4.000 ;
    END
  END pll_trim[3]
  PIN pll_trim[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.680 0.000 226.240 4.000 ;
    END
  END pll_trim[4]
  PIN pll_trim[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 232.400 0.000 232.960 4.000 ;
    END
  END pll_trim[5]
  PIN pll_trim[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 239.120 0.000 239.680 4.000 ;
    END
  END pll_trim[6]
  PIN pll_trim[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.840 0.000 246.400 4.000 ;
    END
  END pll_trim[7]
  PIN pll_trim[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.560 0.000 253.120 4.000 ;
    END
  END pll_trim[8]
  PIN pll_trim[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 259.280 0.000 259.840 4.000 ;
    END
  END pll_trim[9]
  PIN porb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 98.000 0.000 98.560 4.000 ;
    END
  END porb
  PIN pwr_ctrl_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 608.720 0.000 609.280 4.000 ;
    END
  END pwr_ctrl_out
  PIN qspi_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 115.360 4.000 115.920 ;
    END
  END qspi_enabled
  PIN reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.720 0.000 105.280 4.000 ;
    END
  END reset
  PIN ser_rx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 109.200 4.000 109.760 ;
    END
  END ser_rx
  PIN ser_tx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 103.040 4.000 103.600 ;
    END
  END ser_tx
  PIN serial_clock
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 13.440 620.000 14.000 ;
    END
  END serial_clock
  PIN serial_data_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 48.720 620.000 49.280 ;
    END
  END serial_data_1
  PIN serial_data_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 60.480 620.000 61.040 ;
    END
  END serial_data_2
  PIN serial_load
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 36.960 620.000 37.520 ;
    END
  END serial_load
  PIN serial_resetn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 616.000 25.200 620.000 25.760 ;
    END
  END serial_resetn
  PIN spi_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.720 4.000 91.280 ;
    END
  END spi_csb
  PIN spi_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END spi_enabled
  PIN spi_sck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.560 4.000 85.120 ;
    END
  END spi_sck
  PIN spi_sdi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 96.880 4.000 97.440 ;
    END
  END spi_sdi
  PIN spi_sdo
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 78.400 4.000 78.960 ;
    END
  END spi_sdo
  PIN spi_sdoenb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 72.240 4.000 72.800 ;
    END
  END spi_sdoenb
  PIN spimemio_flash_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 343.280 4.000 343.840 ;
    END
  END spimemio_flash_clk
  PIN spimemio_flash_csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 349.440 4.000 350.000 ;
    END
  END spimemio_flash_csb
  PIN spimemio_flash_io0_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 355.600 4.000 356.160 ;
    END
  END spimemio_flash_io0_di
  PIN spimemio_flash_io0_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 361.760 4.000 362.320 ;
    END
  END spimemio_flash_io0_do
  PIN spimemio_flash_io0_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 367.920 4.000 368.480 ;
    END
  END spimemio_flash_io0_oeb
  PIN spimemio_flash_io1_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 374.080 4.000 374.640 ;
    END
  END spimemio_flash_io1_di
  PIN spimemio_flash_io1_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 380.240 4.000 380.800 ;
    END
  END spimemio_flash_io1_do
  PIN spimemio_flash_io1_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 386.400 4.000 386.960 ;
    END
  END spimemio_flash_io1_oeb
  PIN spimemio_flash_io2_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 392.560 4.000 393.120 ;
    END
  END spimemio_flash_io2_di
  PIN spimemio_flash_io2_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 398.720 4.000 399.280 ;
    END
  END spimemio_flash_io2_do
  PIN spimemio_flash_io2_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 404.880 4.000 405.440 ;
    END
  END spimemio_flash_io2_oeb
  PIN spimemio_flash_io3_di
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 411.040 4.000 411.600 ;
    END
  END spimemio_flash_io3_di
  PIN spimemio_flash_io3_do
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 417.200 4.000 417.760 ;
    END
  END spimemio_flash_io3_do
  PIN spimemio_flash_io3_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 423.360 4.000 423.920 ;
    END
  END spimemio_flash_io3_oeb
  PIN trap
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 47.600 4.000 48.160 ;
    END
  END trap
  PIN uart_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 121.520 4.000 122.080 ;
    END
  END uart_enabled
  PIN user_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.640 0.000 11.200 4.000 ;
    END
  END user_clock
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 133.840 4.000 134.400 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.600 776.000 20.160 780.000 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.600 776.000 104.160 780.000 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 776.000 112.560 780.000 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.400 776.000 120.960 780.000 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 128.800 776.000 129.360 780.000 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.200 776.000 137.760 780.000 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 145.600 776.000 146.160 780.000 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.000 776.000 154.560 780.000 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 162.400 776.000 162.960 780.000 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 170.800 776.000 171.360 780.000 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 776.000 179.760 780.000 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 28.000 776.000 28.560 780.000 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.600 776.000 188.160 780.000 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 776.000 196.560 780.000 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.400 776.000 204.960 780.000 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 212.800 776.000 213.360 780.000 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.200 776.000 221.760 780.000 ;
    END
  END wb_adr_i[24]
  PIN wb_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 776.000 230.160 780.000 ;
    END
  END wb_adr_i[25]
  PIN wb_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.000 776.000 238.560 780.000 ;
    END
  END wb_adr_i[26]
  PIN wb_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 246.400 776.000 246.960 780.000 ;
    END
  END wb_adr_i[27]
  PIN wb_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 254.800 776.000 255.360 780.000 ;
    END
  END wb_adr_i[28]
  PIN wb_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 263.200 776.000 263.760 780.000 ;
    END
  END wb_adr_i[29]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.400 776.000 36.960 780.000 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 271.600 776.000 272.160 780.000 ;
    END
  END wb_adr_i[30]
  PIN wb_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 776.000 280.560 780.000 ;
    END
  END wb_adr_i[31]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 776.000 45.360 780.000 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.200 776.000 53.760 780.000 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 61.600 776.000 62.160 780.000 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.000 776.000 70.560 780.000 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 78.400 776.000 78.960 780.000 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.800 776.000 87.360 780.000 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 776.000 95.760 780.000 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 380.240 0.000 380.800 4.000 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 599.200 776.000 599.760 780.000 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.400 776.000 288.960 780.000 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.400 776.000 372.960 780.000 ;
    END
  END wb_dat_i[10]
  PIN wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 380.800 776.000 381.360 780.000 ;
    END
  END wb_dat_i[11]
  PIN wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 389.200 776.000 389.760 780.000 ;
    END
  END wb_dat_i[12]
  PIN wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 397.600 776.000 398.160 780.000 ;
    END
  END wb_dat_i[13]
  PIN wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.000 776.000 406.560 780.000 ;
    END
  END wb_dat_i[14]
  PIN wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 776.000 414.960 780.000 ;
    END
  END wb_dat_i[15]
  PIN wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 422.800 776.000 423.360 780.000 ;
    END
  END wb_dat_i[16]
  PIN wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 431.200 776.000 431.760 780.000 ;
    END
  END wb_dat_i[17]
  PIN wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 439.600 776.000 440.160 780.000 ;
    END
  END wb_dat_i[18]
  PIN wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 448.000 776.000 448.560 780.000 ;
    END
  END wb_dat_i[19]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 776.000 297.360 780.000 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.400 776.000 456.960 780.000 ;
    END
  END wb_dat_i[20]
  PIN wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 464.800 776.000 465.360 780.000 ;
    END
  END wb_dat_i[21]
  PIN wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.200 776.000 473.760 780.000 ;
    END
  END wb_dat_i[22]
  PIN wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 481.600 776.000 482.160 780.000 ;
    END
  END wb_dat_i[23]
  PIN wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 490.000 776.000 490.560 780.000 ;
    END
  END wb_dat_i[24]
  PIN wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 498.400 776.000 498.960 780.000 ;
    END
  END wb_dat_i[25]
  PIN wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 506.800 776.000 507.360 780.000 ;
    END
  END wb_dat_i[26]
  PIN wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 515.200 776.000 515.760 780.000 ;
    END
  END wb_dat_i[27]
  PIN wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 523.600 776.000 524.160 780.000 ;
    END
  END wb_dat_i[28]
  PIN wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 532.000 776.000 532.560 780.000 ;
    END
  END wb_dat_i[29]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 305.200 776.000 305.760 780.000 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 540.400 776.000 540.960 780.000 ;
    END
  END wb_dat_i[30]
  PIN wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 548.800 776.000 549.360 780.000 ;
    END
  END wb_dat_i[31]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 313.600 776.000 314.160 780.000 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.000 776.000 322.560 780.000 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 330.400 776.000 330.960 780.000 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 338.800 776.000 339.360 780.000 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 347.200 776.000 347.760 780.000 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 355.600 776.000 356.160 780.000 ;
    END
  END wb_dat_i[8]
  PIN wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 364.000 776.000 364.560 780.000 ;
    END
  END wb_dat_i[9]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 146.160 4.000 146.720 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.760 4.000 208.320 ;
    END
  END wb_dat_o[10]
  PIN wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 213.920 4.000 214.480 ;
    END
  END wb_dat_o[11]
  PIN wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 220.080 4.000 220.640 ;
    END
  END wb_dat_o[12]
  PIN wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 226.240 4.000 226.800 ;
    END
  END wb_dat_o[13]
  PIN wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 232.400 4.000 232.960 ;
    END
  END wb_dat_o[14]
  PIN wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 238.560 4.000 239.120 ;
    END
  END wb_dat_o[15]
  PIN wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 244.720 4.000 245.280 ;
    END
  END wb_dat_o[16]
  PIN wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 250.880 4.000 251.440 ;
    END
  END wb_dat_o[17]
  PIN wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 257.040 4.000 257.600 ;
    END
  END wb_dat_o[18]
  PIN wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 263.200 4.000 263.760 ;
    END
  END wb_dat_o[19]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 152.320 4.000 152.880 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 269.360 4.000 269.920 ;
    END
  END wb_dat_o[20]
  PIN wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 275.520 4.000 276.080 ;
    END
  END wb_dat_o[21]
  PIN wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 281.680 4.000 282.240 ;
    END
  END wb_dat_o[22]
  PIN wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 287.840 4.000 288.400 ;
    END
  END wb_dat_o[23]
  PIN wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.000 4.000 294.560 ;
    END
  END wb_dat_o[24]
  PIN wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 300.160 4.000 300.720 ;
    END
  END wb_dat_o[25]
  PIN wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 306.320 4.000 306.880 ;
    END
  END wb_dat_o[26]
  PIN wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 312.480 4.000 313.040 ;
    END
  END wb_dat_o[27]
  PIN wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.640 4.000 319.200 ;
    END
  END wb_dat_o[28]
  PIN wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 324.800 4.000 325.360 ;
    END
  END wb_dat_o[29]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 158.480 4.000 159.040 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 330.960 4.000 331.520 ;
    END
  END wb_dat_o[30]
  PIN wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 337.120 4.000 337.680 ;
    END
  END wb_dat_o[31]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 4.000 165.200 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 170.800 4.000 171.360 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 176.960 4.000 177.520 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 183.120 4.000 183.680 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 189.280 4.000 189.840 ;
    END
  END wb_dat_o[7]
  PIN wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 195.440 4.000 196.000 ;
    END
  END wb_dat_o[8]
  PIN wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END wb_dat_o[9]
  PIN wb_rstn_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.960 0.000 387.520 4.000 ;
    END
  END wb_rstn_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 557.200 776.000 557.760 780.000 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 565.600 776.000 566.160 780.000 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 574.000 776.000 574.560 780.000 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 582.400 776.000 582.960 780.000 ;
    END
  END wb_sel_i[3]
  PIN wb_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 140.000 4.000 140.560 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 590.800 776.000 591.360 780.000 ;
    END
  END wb_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 613.200 762.570 ;
      LAYER Metal2 ;
        RECT 4.060 775.700 19.300 776.000 ;
        RECT 20.460 775.700 27.700 776.000 ;
        RECT 28.860 775.700 36.100 776.000 ;
        RECT 37.260 775.700 44.500 776.000 ;
        RECT 45.660 775.700 52.900 776.000 ;
        RECT 54.060 775.700 61.300 776.000 ;
        RECT 62.460 775.700 69.700 776.000 ;
        RECT 70.860 775.700 78.100 776.000 ;
        RECT 79.260 775.700 86.500 776.000 ;
        RECT 87.660 775.700 94.900 776.000 ;
        RECT 96.060 775.700 103.300 776.000 ;
        RECT 104.460 775.700 111.700 776.000 ;
        RECT 112.860 775.700 120.100 776.000 ;
        RECT 121.260 775.700 128.500 776.000 ;
        RECT 129.660 775.700 136.900 776.000 ;
        RECT 138.060 775.700 145.300 776.000 ;
        RECT 146.460 775.700 153.700 776.000 ;
        RECT 154.860 775.700 162.100 776.000 ;
        RECT 163.260 775.700 170.500 776.000 ;
        RECT 171.660 775.700 178.900 776.000 ;
        RECT 180.060 775.700 187.300 776.000 ;
        RECT 188.460 775.700 195.700 776.000 ;
        RECT 196.860 775.700 204.100 776.000 ;
        RECT 205.260 775.700 212.500 776.000 ;
        RECT 213.660 775.700 220.900 776.000 ;
        RECT 222.060 775.700 229.300 776.000 ;
        RECT 230.460 775.700 237.700 776.000 ;
        RECT 238.860 775.700 246.100 776.000 ;
        RECT 247.260 775.700 254.500 776.000 ;
        RECT 255.660 775.700 262.900 776.000 ;
        RECT 264.060 775.700 271.300 776.000 ;
        RECT 272.460 775.700 279.700 776.000 ;
        RECT 280.860 775.700 288.100 776.000 ;
        RECT 289.260 775.700 296.500 776.000 ;
        RECT 297.660 775.700 304.900 776.000 ;
        RECT 306.060 775.700 313.300 776.000 ;
        RECT 314.460 775.700 321.700 776.000 ;
        RECT 322.860 775.700 330.100 776.000 ;
        RECT 331.260 775.700 338.500 776.000 ;
        RECT 339.660 775.700 346.900 776.000 ;
        RECT 348.060 775.700 355.300 776.000 ;
        RECT 356.460 775.700 363.700 776.000 ;
        RECT 364.860 775.700 372.100 776.000 ;
        RECT 373.260 775.700 380.500 776.000 ;
        RECT 381.660 775.700 388.900 776.000 ;
        RECT 390.060 775.700 397.300 776.000 ;
        RECT 398.460 775.700 405.700 776.000 ;
        RECT 406.860 775.700 414.100 776.000 ;
        RECT 415.260 775.700 422.500 776.000 ;
        RECT 423.660 775.700 430.900 776.000 ;
        RECT 432.060 775.700 439.300 776.000 ;
        RECT 440.460 775.700 447.700 776.000 ;
        RECT 448.860 775.700 456.100 776.000 ;
        RECT 457.260 775.700 464.500 776.000 ;
        RECT 465.660 775.700 472.900 776.000 ;
        RECT 474.060 775.700 481.300 776.000 ;
        RECT 482.460 775.700 489.700 776.000 ;
        RECT 490.860 775.700 498.100 776.000 ;
        RECT 499.260 775.700 506.500 776.000 ;
        RECT 507.660 775.700 514.900 776.000 ;
        RECT 516.060 775.700 523.300 776.000 ;
        RECT 524.460 775.700 531.700 776.000 ;
        RECT 532.860 775.700 540.100 776.000 ;
        RECT 541.260 775.700 548.500 776.000 ;
        RECT 549.660 775.700 556.900 776.000 ;
        RECT 558.060 775.700 565.300 776.000 ;
        RECT 566.460 775.700 573.700 776.000 ;
        RECT 574.860 775.700 582.100 776.000 ;
        RECT 583.260 775.700 590.500 776.000 ;
        RECT 591.660 775.700 598.900 776.000 ;
        RECT 600.060 775.700 615.300 776.000 ;
        RECT 4.060 4.300 615.300 775.700 ;
        RECT 4.060 3.500 10.340 4.300 ;
        RECT 11.500 3.500 17.060 4.300 ;
        RECT 18.220 3.500 23.780 4.300 ;
        RECT 24.940 3.500 30.500 4.300 ;
        RECT 31.660 3.500 37.220 4.300 ;
        RECT 38.380 3.500 43.940 4.300 ;
        RECT 45.100 3.500 50.660 4.300 ;
        RECT 51.820 3.500 57.380 4.300 ;
        RECT 58.540 3.500 64.100 4.300 ;
        RECT 65.260 3.500 70.820 4.300 ;
        RECT 71.980 3.500 77.540 4.300 ;
        RECT 78.700 3.500 84.260 4.300 ;
        RECT 85.420 3.500 90.980 4.300 ;
        RECT 92.140 3.500 97.700 4.300 ;
        RECT 98.860 3.500 104.420 4.300 ;
        RECT 105.580 3.500 111.140 4.300 ;
        RECT 112.300 3.500 117.860 4.300 ;
        RECT 119.020 3.500 124.580 4.300 ;
        RECT 125.740 3.500 131.300 4.300 ;
        RECT 132.460 3.500 138.020 4.300 ;
        RECT 139.180 3.500 144.740 4.300 ;
        RECT 145.900 3.500 151.460 4.300 ;
        RECT 152.620 3.500 158.180 4.300 ;
        RECT 159.340 3.500 164.900 4.300 ;
        RECT 166.060 3.500 171.620 4.300 ;
        RECT 172.780 3.500 178.340 4.300 ;
        RECT 179.500 3.500 185.060 4.300 ;
        RECT 186.220 3.500 191.780 4.300 ;
        RECT 192.940 3.500 198.500 4.300 ;
        RECT 199.660 3.500 205.220 4.300 ;
        RECT 206.380 3.500 211.940 4.300 ;
        RECT 213.100 3.500 218.660 4.300 ;
        RECT 219.820 3.500 225.380 4.300 ;
        RECT 226.540 3.500 232.100 4.300 ;
        RECT 233.260 3.500 238.820 4.300 ;
        RECT 239.980 3.500 245.540 4.300 ;
        RECT 246.700 3.500 252.260 4.300 ;
        RECT 253.420 3.500 258.980 4.300 ;
        RECT 260.140 3.500 265.700 4.300 ;
        RECT 266.860 3.500 272.420 4.300 ;
        RECT 273.580 3.500 279.140 4.300 ;
        RECT 280.300 3.500 285.860 4.300 ;
        RECT 287.020 3.500 292.580 4.300 ;
        RECT 293.740 3.500 299.300 4.300 ;
        RECT 300.460 3.500 306.020 4.300 ;
        RECT 307.180 3.500 312.740 4.300 ;
        RECT 313.900 3.500 319.460 4.300 ;
        RECT 320.620 3.500 326.180 4.300 ;
        RECT 327.340 3.500 332.900 4.300 ;
        RECT 334.060 3.500 339.620 4.300 ;
        RECT 340.780 3.500 346.340 4.300 ;
        RECT 347.500 3.500 353.060 4.300 ;
        RECT 354.220 3.500 359.780 4.300 ;
        RECT 360.940 3.500 366.500 4.300 ;
        RECT 367.660 3.500 373.220 4.300 ;
        RECT 374.380 3.500 379.940 4.300 ;
        RECT 381.100 3.500 386.660 4.300 ;
        RECT 387.820 3.500 393.380 4.300 ;
        RECT 394.540 3.500 400.100 4.300 ;
        RECT 401.260 3.500 406.820 4.300 ;
        RECT 407.980 3.500 413.540 4.300 ;
        RECT 414.700 3.500 420.260 4.300 ;
        RECT 421.420 3.500 426.980 4.300 ;
        RECT 428.140 3.500 433.700 4.300 ;
        RECT 434.860 3.500 440.420 4.300 ;
        RECT 441.580 3.500 447.140 4.300 ;
        RECT 448.300 3.500 453.860 4.300 ;
        RECT 455.020 3.500 460.580 4.300 ;
        RECT 461.740 3.500 467.300 4.300 ;
        RECT 468.460 3.500 474.020 4.300 ;
        RECT 475.180 3.500 480.740 4.300 ;
        RECT 481.900 3.500 487.460 4.300 ;
        RECT 488.620 3.500 494.180 4.300 ;
        RECT 495.340 3.500 500.900 4.300 ;
        RECT 502.060 3.500 507.620 4.300 ;
        RECT 508.780 3.500 514.340 4.300 ;
        RECT 515.500 3.500 521.060 4.300 ;
        RECT 522.220 3.500 527.780 4.300 ;
        RECT 528.940 3.500 534.500 4.300 ;
        RECT 535.660 3.500 541.220 4.300 ;
        RECT 542.380 3.500 547.940 4.300 ;
        RECT 549.100 3.500 554.660 4.300 ;
        RECT 555.820 3.500 561.380 4.300 ;
        RECT 562.540 3.500 568.100 4.300 ;
        RECT 569.260 3.500 574.820 4.300 ;
        RECT 575.980 3.500 581.540 4.300 ;
        RECT 582.700 3.500 588.260 4.300 ;
        RECT 589.420 3.500 594.980 4.300 ;
        RECT 596.140 3.500 601.700 4.300 ;
        RECT 602.860 3.500 608.420 4.300 ;
        RECT 609.580 3.500 615.300 4.300 ;
      LAYER Metal3 ;
        RECT 3.500 765.780 615.700 766.500 ;
        RECT 3.500 756.860 616.420 765.780 ;
        RECT 4.300 755.700 616.420 756.860 ;
        RECT 3.500 755.180 616.420 755.700 ;
        RECT 3.500 754.020 615.700 755.180 ;
        RECT 3.500 750.700 616.420 754.020 ;
        RECT 4.300 749.540 616.420 750.700 ;
        RECT 3.500 744.540 616.420 749.540 ;
        RECT 4.300 743.420 616.420 744.540 ;
        RECT 4.300 743.380 615.700 743.420 ;
        RECT 3.500 742.260 615.700 743.380 ;
        RECT 3.500 738.380 616.420 742.260 ;
        RECT 4.300 737.220 616.420 738.380 ;
        RECT 3.500 732.220 616.420 737.220 ;
        RECT 4.300 731.660 616.420 732.220 ;
        RECT 4.300 731.060 615.700 731.660 ;
        RECT 3.500 730.500 615.700 731.060 ;
        RECT 3.500 726.060 616.420 730.500 ;
        RECT 4.300 724.900 616.420 726.060 ;
        RECT 3.500 719.900 616.420 724.900 ;
        RECT 4.300 718.740 615.700 719.900 ;
        RECT 3.500 713.740 616.420 718.740 ;
        RECT 4.300 712.580 616.420 713.740 ;
        RECT 3.500 708.140 616.420 712.580 ;
        RECT 3.500 707.580 615.700 708.140 ;
        RECT 4.300 706.980 615.700 707.580 ;
        RECT 4.300 706.420 616.420 706.980 ;
        RECT 3.500 701.420 616.420 706.420 ;
        RECT 4.300 700.260 616.420 701.420 ;
        RECT 3.500 696.380 616.420 700.260 ;
        RECT 3.500 695.260 615.700 696.380 ;
        RECT 4.300 695.220 615.700 695.260 ;
        RECT 4.300 694.100 616.420 695.220 ;
        RECT 3.500 689.100 616.420 694.100 ;
        RECT 4.300 687.940 616.420 689.100 ;
        RECT 3.500 684.620 616.420 687.940 ;
        RECT 3.500 683.460 615.700 684.620 ;
        RECT 3.500 682.940 616.420 683.460 ;
        RECT 4.300 681.780 616.420 682.940 ;
        RECT 3.500 676.780 616.420 681.780 ;
        RECT 4.300 675.620 616.420 676.780 ;
        RECT 3.500 672.860 616.420 675.620 ;
        RECT 3.500 671.700 615.700 672.860 ;
        RECT 3.500 670.620 616.420 671.700 ;
        RECT 4.300 669.460 616.420 670.620 ;
        RECT 3.500 664.460 616.420 669.460 ;
        RECT 4.300 663.300 616.420 664.460 ;
        RECT 3.500 661.100 616.420 663.300 ;
        RECT 3.500 659.940 615.700 661.100 ;
        RECT 3.500 658.300 616.420 659.940 ;
        RECT 4.300 657.140 616.420 658.300 ;
        RECT 3.500 652.140 616.420 657.140 ;
        RECT 4.300 650.980 616.420 652.140 ;
        RECT 3.500 649.340 616.420 650.980 ;
        RECT 3.500 648.180 615.700 649.340 ;
        RECT 3.500 645.980 616.420 648.180 ;
        RECT 4.300 644.820 616.420 645.980 ;
        RECT 3.500 639.820 616.420 644.820 ;
        RECT 4.300 638.660 616.420 639.820 ;
        RECT 3.500 637.580 616.420 638.660 ;
        RECT 3.500 636.420 615.700 637.580 ;
        RECT 3.500 633.660 616.420 636.420 ;
        RECT 4.300 632.500 616.420 633.660 ;
        RECT 3.500 627.500 616.420 632.500 ;
        RECT 4.300 626.340 616.420 627.500 ;
        RECT 3.500 625.820 616.420 626.340 ;
        RECT 3.500 624.660 615.700 625.820 ;
        RECT 3.500 621.340 616.420 624.660 ;
        RECT 4.300 620.180 616.420 621.340 ;
        RECT 3.500 615.180 616.420 620.180 ;
        RECT 4.300 614.060 616.420 615.180 ;
        RECT 4.300 614.020 615.700 614.060 ;
        RECT 3.500 612.900 615.700 614.020 ;
        RECT 3.500 609.020 616.420 612.900 ;
        RECT 4.300 607.860 616.420 609.020 ;
        RECT 3.500 602.860 616.420 607.860 ;
        RECT 4.300 602.300 616.420 602.860 ;
        RECT 4.300 601.700 615.700 602.300 ;
        RECT 3.500 601.140 615.700 601.700 ;
        RECT 3.500 596.700 616.420 601.140 ;
        RECT 4.300 595.540 616.420 596.700 ;
        RECT 3.500 590.540 616.420 595.540 ;
        RECT 4.300 589.380 615.700 590.540 ;
        RECT 3.500 584.380 616.420 589.380 ;
        RECT 4.300 583.220 616.420 584.380 ;
        RECT 3.500 578.780 616.420 583.220 ;
        RECT 3.500 578.220 615.700 578.780 ;
        RECT 4.300 577.620 615.700 578.220 ;
        RECT 4.300 577.060 616.420 577.620 ;
        RECT 3.500 572.060 616.420 577.060 ;
        RECT 4.300 570.900 616.420 572.060 ;
        RECT 3.500 567.020 616.420 570.900 ;
        RECT 3.500 565.900 615.700 567.020 ;
        RECT 4.300 565.860 615.700 565.900 ;
        RECT 4.300 564.740 616.420 565.860 ;
        RECT 3.500 559.740 616.420 564.740 ;
        RECT 4.300 558.580 616.420 559.740 ;
        RECT 3.500 555.260 616.420 558.580 ;
        RECT 3.500 554.100 615.700 555.260 ;
        RECT 3.500 553.580 616.420 554.100 ;
        RECT 4.300 552.420 616.420 553.580 ;
        RECT 3.500 547.420 616.420 552.420 ;
        RECT 4.300 546.260 616.420 547.420 ;
        RECT 3.500 543.500 616.420 546.260 ;
        RECT 3.500 542.340 615.700 543.500 ;
        RECT 3.500 541.260 616.420 542.340 ;
        RECT 4.300 540.100 616.420 541.260 ;
        RECT 3.500 535.100 616.420 540.100 ;
        RECT 4.300 533.940 616.420 535.100 ;
        RECT 3.500 531.740 616.420 533.940 ;
        RECT 3.500 530.580 615.700 531.740 ;
        RECT 3.500 528.940 616.420 530.580 ;
        RECT 4.300 527.780 616.420 528.940 ;
        RECT 3.500 522.780 616.420 527.780 ;
        RECT 4.300 521.620 616.420 522.780 ;
        RECT 3.500 519.980 616.420 521.620 ;
        RECT 3.500 518.820 615.700 519.980 ;
        RECT 3.500 516.620 616.420 518.820 ;
        RECT 4.300 515.460 616.420 516.620 ;
        RECT 3.500 510.460 616.420 515.460 ;
        RECT 4.300 509.300 616.420 510.460 ;
        RECT 3.500 508.220 616.420 509.300 ;
        RECT 3.500 507.060 615.700 508.220 ;
        RECT 3.500 504.300 616.420 507.060 ;
        RECT 4.300 503.140 616.420 504.300 ;
        RECT 3.500 498.140 616.420 503.140 ;
        RECT 4.300 496.980 616.420 498.140 ;
        RECT 3.500 496.460 616.420 496.980 ;
        RECT 3.500 495.300 615.700 496.460 ;
        RECT 3.500 491.980 616.420 495.300 ;
        RECT 4.300 490.820 616.420 491.980 ;
        RECT 3.500 485.820 616.420 490.820 ;
        RECT 4.300 484.700 616.420 485.820 ;
        RECT 4.300 484.660 615.700 484.700 ;
        RECT 3.500 483.540 615.700 484.660 ;
        RECT 3.500 479.660 616.420 483.540 ;
        RECT 4.300 478.500 616.420 479.660 ;
        RECT 3.500 473.500 616.420 478.500 ;
        RECT 4.300 472.940 616.420 473.500 ;
        RECT 4.300 472.340 615.700 472.940 ;
        RECT 3.500 471.780 615.700 472.340 ;
        RECT 3.500 467.340 616.420 471.780 ;
        RECT 4.300 466.180 616.420 467.340 ;
        RECT 3.500 461.180 616.420 466.180 ;
        RECT 4.300 460.020 615.700 461.180 ;
        RECT 3.500 455.020 616.420 460.020 ;
        RECT 4.300 453.860 616.420 455.020 ;
        RECT 3.500 449.420 616.420 453.860 ;
        RECT 3.500 448.860 615.700 449.420 ;
        RECT 4.300 448.260 615.700 448.860 ;
        RECT 4.300 447.700 616.420 448.260 ;
        RECT 3.500 442.700 616.420 447.700 ;
        RECT 4.300 441.540 616.420 442.700 ;
        RECT 3.500 437.660 616.420 441.540 ;
        RECT 3.500 436.540 615.700 437.660 ;
        RECT 4.300 436.500 615.700 436.540 ;
        RECT 4.300 435.380 616.420 436.500 ;
        RECT 3.500 430.380 616.420 435.380 ;
        RECT 4.300 429.220 616.420 430.380 ;
        RECT 3.500 425.900 616.420 429.220 ;
        RECT 3.500 424.740 615.700 425.900 ;
        RECT 3.500 424.220 616.420 424.740 ;
        RECT 4.300 423.060 616.420 424.220 ;
        RECT 3.500 418.060 616.420 423.060 ;
        RECT 4.300 416.900 616.420 418.060 ;
        RECT 3.500 414.140 616.420 416.900 ;
        RECT 3.500 412.980 615.700 414.140 ;
        RECT 3.500 411.900 616.420 412.980 ;
        RECT 4.300 410.740 616.420 411.900 ;
        RECT 3.500 405.740 616.420 410.740 ;
        RECT 4.300 404.580 616.420 405.740 ;
        RECT 3.500 402.380 616.420 404.580 ;
        RECT 3.500 401.220 615.700 402.380 ;
        RECT 3.500 399.580 616.420 401.220 ;
        RECT 4.300 398.420 616.420 399.580 ;
        RECT 3.500 393.420 616.420 398.420 ;
        RECT 4.300 392.260 616.420 393.420 ;
        RECT 3.500 390.620 616.420 392.260 ;
        RECT 3.500 389.460 615.700 390.620 ;
        RECT 3.500 387.260 616.420 389.460 ;
        RECT 4.300 386.100 616.420 387.260 ;
        RECT 3.500 381.100 616.420 386.100 ;
        RECT 4.300 379.940 616.420 381.100 ;
        RECT 3.500 378.860 616.420 379.940 ;
        RECT 3.500 377.700 615.700 378.860 ;
        RECT 3.500 374.940 616.420 377.700 ;
        RECT 4.300 373.780 616.420 374.940 ;
        RECT 3.500 368.780 616.420 373.780 ;
        RECT 4.300 367.620 616.420 368.780 ;
        RECT 3.500 367.100 616.420 367.620 ;
        RECT 3.500 365.940 615.700 367.100 ;
        RECT 3.500 362.620 616.420 365.940 ;
        RECT 4.300 361.460 616.420 362.620 ;
        RECT 3.500 356.460 616.420 361.460 ;
        RECT 4.300 355.340 616.420 356.460 ;
        RECT 4.300 355.300 615.700 355.340 ;
        RECT 3.500 354.180 615.700 355.300 ;
        RECT 3.500 350.300 616.420 354.180 ;
        RECT 4.300 349.140 616.420 350.300 ;
        RECT 3.500 344.140 616.420 349.140 ;
        RECT 4.300 343.580 616.420 344.140 ;
        RECT 4.300 342.980 615.700 343.580 ;
        RECT 3.500 342.420 615.700 342.980 ;
        RECT 3.500 337.980 616.420 342.420 ;
        RECT 4.300 336.820 616.420 337.980 ;
        RECT 3.500 331.820 616.420 336.820 ;
        RECT 4.300 330.660 615.700 331.820 ;
        RECT 3.500 325.660 616.420 330.660 ;
        RECT 4.300 324.500 616.420 325.660 ;
        RECT 3.500 320.060 616.420 324.500 ;
        RECT 3.500 319.500 615.700 320.060 ;
        RECT 4.300 318.900 615.700 319.500 ;
        RECT 4.300 318.340 616.420 318.900 ;
        RECT 3.500 313.340 616.420 318.340 ;
        RECT 4.300 312.180 616.420 313.340 ;
        RECT 3.500 308.300 616.420 312.180 ;
        RECT 3.500 307.180 615.700 308.300 ;
        RECT 4.300 307.140 615.700 307.180 ;
        RECT 4.300 306.020 616.420 307.140 ;
        RECT 3.500 301.020 616.420 306.020 ;
        RECT 4.300 299.860 616.420 301.020 ;
        RECT 3.500 296.540 616.420 299.860 ;
        RECT 3.500 295.380 615.700 296.540 ;
        RECT 3.500 294.860 616.420 295.380 ;
        RECT 4.300 293.700 616.420 294.860 ;
        RECT 3.500 288.700 616.420 293.700 ;
        RECT 4.300 287.540 616.420 288.700 ;
        RECT 3.500 284.780 616.420 287.540 ;
        RECT 3.500 283.620 615.700 284.780 ;
        RECT 3.500 282.540 616.420 283.620 ;
        RECT 4.300 281.380 616.420 282.540 ;
        RECT 3.500 276.380 616.420 281.380 ;
        RECT 4.300 275.220 616.420 276.380 ;
        RECT 3.500 273.020 616.420 275.220 ;
        RECT 3.500 271.860 615.700 273.020 ;
        RECT 3.500 270.220 616.420 271.860 ;
        RECT 4.300 269.060 616.420 270.220 ;
        RECT 3.500 264.060 616.420 269.060 ;
        RECT 4.300 262.900 616.420 264.060 ;
        RECT 3.500 261.260 616.420 262.900 ;
        RECT 3.500 260.100 615.700 261.260 ;
        RECT 3.500 257.900 616.420 260.100 ;
        RECT 4.300 256.740 616.420 257.900 ;
        RECT 3.500 251.740 616.420 256.740 ;
        RECT 4.300 250.580 616.420 251.740 ;
        RECT 3.500 249.500 616.420 250.580 ;
        RECT 3.500 248.340 615.700 249.500 ;
        RECT 3.500 245.580 616.420 248.340 ;
        RECT 4.300 244.420 616.420 245.580 ;
        RECT 3.500 239.420 616.420 244.420 ;
        RECT 4.300 238.260 616.420 239.420 ;
        RECT 3.500 237.740 616.420 238.260 ;
        RECT 3.500 236.580 615.700 237.740 ;
        RECT 3.500 233.260 616.420 236.580 ;
        RECT 4.300 232.100 616.420 233.260 ;
        RECT 3.500 227.100 616.420 232.100 ;
        RECT 4.300 225.980 616.420 227.100 ;
        RECT 4.300 225.940 615.700 225.980 ;
        RECT 3.500 224.820 615.700 225.940 ;
        RECT 3.500 220.940 616.420 224.820 ;
        RECT 4.300 219.780 616.420 220.940 ;
        RECT 3.500 214.780 616.420 219.780 ;
        RECT 4.300 214.220 616.420 214.780 ;
        RECT 4.300 213.620 615.700 214.220 ;
        RECT 3.500 213.060 615.700 213.620 ;
        RECT 3.500 208.620 616.420 213.060 ;
        RECT 4.300 207.460 616.420 208.620 ;
        RECT 3.500 202.460 616.420 207.460 ;
        RECT 4.300 201.300 615.700 202.460 ;
        RECT 3.500 196.300 616.420 201.300 ;
        RECT 4.300 195.140 616.420 196.300 ;
        RECT 3.500 190.700 616.420 195.140 ;
        RECT 3.500 190.140 615.700 190.700 ;
        RECT 4.300 189.540 615.700 190.140 ;
        RECT 4.300 188.980 616.420 189.540 ;
        RECT 3.500 183.980 616.420 188.980 ;
        RECT 4.300 182.820 616.420 183.980 ;
        RECT 3.500 178.940 616.420 182.820 ;
        RECT 3.500 177.820 615.700 178.940 ;
        RECT 4.300 177.780 615.700 177.820 ;
        RECT 4.300 176.660 616.420 177.780 ;
        RECT 3.500 171.660 616.420 176.660 ;
        RECT 4.300 170.500 616.420 171.660 ;
        RECT 3.500 167.180 616.420 170.500 ;
        RECT 3.500 166.020 615.700 167.180 ;
        RECT 3.500 165.500 616.420 166.020 ;
        RECT 4.300 164.340 616.420 165.500 ;
        RECT 3.500 159.340 616.420 164.340 ;
        RECT 4.300 158.180 616.420 159.340 ;
        RECT 3.500 155.420 616.420 158.180 ;
        RECT 3.500 154.260 615.700 155.420 ;
        RECT 3.500 153.180 616.420 154.260 ;
        RECT 4.300 152.020 616.420 153.180 ;
        RECT 3.500 147.020 616.420 152.020 ;
        RECT 4.300 145.860 616.420 147.020 ;
        RECT 3.500 143.660 616.420 145.860 ;
        RECT 3.500 142.500 615.700 143.660 ;
        RECT 3.500 140.860 616.420 142.500 ;
        RECT 4.300 139.700 616.420 140.860 ;
        RECT 3.500 134.700 616.420 139.700 ;
        RECT 4.300 133.540 616.420 134.700 ;
        RECT 3.500 131.900 616.420 133.540 ;
        RECT 3.500 130.740 615.700 131.900 ;
        RECT 3.500 128.540 616.420 130.740 ;
        RECT 4.300 127.380 616.420 128.540 ;
        RECT 3.500 122.380 616.420 127.380 ;
        RECT 4.300 121.220 616.420 122.380 ;
        RECT 3.500 120.140 616.420 121.220 ;
        RECT 3.500 118.980 615.700 120.140 ;
        RECT 3.500 116.220 616.420 118.980 ;
        RECT 4.300 115.060 616.420 116.220 ;
        RECT 3.500 110.060 616.420 115.060 ;
        RECT 4.300 108.900 616.420 110.060 ;
        RECT 3.500 108.380 616.420 108.900 ;
        RECT 3.500 107.220 615.700 108.380 ;
        RECT 3.500 103.900 616.420 107.220 ;
        RECT 4.300 102.740 616.420 103.900 ;
        RECT 3.500 97.740 616.420 102.740 ;
        RECT 4.300 96.620 616.420 97.740 ;
        RECT 4.300 96.580 615.700 96.620 ;
        RECT 3.500 95.460 615.700 96.580 ;
        RECT 3.500 91.580 616.420 95.460 ;
        RECT 4.300 90.420 616.420 91.580 ;
        RECT 3.500 85.420 616.420 90.420 ;
        RECT 4.300 84.860 616.420 85.420 ;
        RECT 4.300 84.260 615.700 84.860 ;
        RECT 3.500 83.700 615.700 84.260 ;
        RECT 3.500 79.260 616.420 83.700 ;
        RECT 4.300 78.100 616.420 79.260 ;
        RECT 3.500 73.100 616.420 78.100 ;
        RECT 4.300 71.940 615.700 73.100 ;
        RECT 3.500 66.940 616.420 71.940 ;
        RECT 4.300 65.780 616.420 66.940 ;
        RECT 3.500 61.340 616.420 65.780 ;
        RECT 3.500 60.780 615.700 61.340 ;
        RECT 4.300 60.180 615.700 60.780 ;
        RECT 4.300 59.620 616.420 60.180 ;
        RECT 3.500 54.620 616.420 59.620 ;
        RECT 4.300 53.460 616.420 54.620 ;
        RECT 3.500 49.580 616.420 53.460 ;
        RECT 3.500 48.460 615.700 49.580 ;
        RECT 4.300 48.420 615.700 48.460 ;
        RECT 4.300 47.300 616.420 48.420 ;
        RECT 3.500 42.300 616.420 47.300 ;
        RECT 4.300 41.140 616.420 42.300 ;
        RECT 3.500 37.820 616.420 41.140 ;
        RECT 3.500 36.660 615.700 37.820 ;
        RECT 3.500 36.140 616.420 36.660 ;
        RECT 4.300 34.980 616.420 36.140 ;
        RECT 3.500 29.980 616.420 34.980 ;
        RECT 4.300 28.820 616.420 29.980 ;
        RECT 3.500 26.060 616.420 28.820 ;
        RECT 3.500 24.900 615.700 26.060 ;
        RECT 3.500 23.820 616.420 24.900 ;
        RECT 4.300 22.660 616.420 23.820 ;
        RECT 3.500 14.300 616.420 22.660 ;
        RECT 3.500 13.140 615.700 14.300 ;
        RECT 3.500 1.260 616.420 13.140 ;
      LAYER Metal4 ;
        RECT 7.420 4.480 21.940 758.710 ;
        RECT 24.140 4.480 25.240 758.710 ;
        RECT 27.440 4.480 98.740 758.710 ;
        RECT 100.940 4.480 102.040 758.710 ;
        RECT 104.240 4.480 175.540 758.710 ;
        RECT 177.740 4.480 178.840 758.710 ;
        RECT 181.040 4.480 252.340 758.710 ;
        RECT 254.540 4.480 255.640 758.710 ;
        RECT 257.840 4.480 329.140 758.710 ;
        RECT 331.340 4.480 332.440 758.710 ;
        RECT 334.640 4.480 405.940 758.710 ;
        RECT 408.140 4.480 409.240 758.710 ;
        RECT 411.440 4.480 482.740 758.710 ;
        RECT 484.940 4.480 486.040 758.710 ;
        RECT 488.240 4.480 559.540 758.710 ;
        RECT 561.740 4.480 562.840 758.710 ;
        RECT 565.040 4.480 611.380 758.710 ;
        RECT 7.420 0.090 611.380 4.480 ;
      LAYER Metal5 ;
        RECT 9.580 683.390 611.460 692.100 ;
        RECT 9.580 653.390 611.460 680.790 ;
        RECT 9.580 623.390 611.460 650.790 ;
        RECT 9.580 593.390 611.460 620.790 ;
        RECT 9.580 563.390 611.460 590.790 ;
        RECT 9.580 533.390 611.460 560.790 ;
        RECT 9.580 503.390 611.460 530.790 ;
        RECT 9.580 473.390 611.460 500.790 ;
        RECT 9.580 443.390 611.460 470.790 ;
        RECT 9.580 413.390 611.460 440.790 ;
        RECT 9.580 383.390 611.460 410.790 ;
        RECT 9.580 353.390 611.460 380.790 ;
        RECT 9.580 323.390 611.460 350.790 ;
        RECT 9.580 293.390 611.460 320.790 ;
        RECT 9.580 263.390 611.460 290.790 ;
        RECT 9.580 233.390 611.460 260.790 ;
        RECT 9.580 203.390 611.460 230.790 ;
        RECT 9.580 173.390 611.460 200.790 ;
        RECT 9.580 143.390 611.460 170.790 ;
        RECT 9.580 113.390 611.460 140.790 ;
        RECT 9.580 83.390 611.460 110.790 ;
        RECT 9.580 53.390 611.460 80.790 ;
        RECT 9.580 23.390 611.460 50.790 ;
        RECT 9.580 10.180 611.460 20.790 ;
        RECT 9.580 6.880 611.460 7.580 ;
        RECT 9.580 0.060 611.460 4.280 ;
  END
END housekeeping
END LIBRARY

